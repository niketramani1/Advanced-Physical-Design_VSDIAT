magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 111 127 157 467
rect 296 209 362 255
rect 396 209 490 255
rect 524 209 614 255
rect 652 209 719 255
rect 111 51 155 127
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 298 77 527
rect 18 17 77 181
rect 200 366 251 527
rect 291 404 357 493
rect 391 438 446 527
rect 493 404 559 493
rect 291 368 559 404
rect 651 332 717 465
rect 200 298 717 332
rect 200 175 262 298
rect 200 139 717 175
rect 189 17 359 89
rect 455 55 521 139
rect 562 17 617 105
rect 651 55 717 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 396 209 490 255 6 A1
port 1 nsew signal input
rlabel locali s 296 209 362 255 6 A2
port 2 nsew signal input
rlabel locali s 524 209 614 255 6 B1
port 3 nsew signal input
rlabel locali s 652 209 719 255 6 C1
port 4 nsew signal input
rlabel locali s 111 127 157 467 6 X
port 9 nsew signal output
rlabel locali s 111 51 155 127 6 X
port 9 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3411278
string GDS_START 3404714
<< end >>
