magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 103 299 169 493
rect 103 176 158 299
rect 355 215 431 265
rect 465 215 531 468
rect 565 215 631 468
rect 665 215 731 467
rect 765 215 903 265
rect 103 51 169 176
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 299 69 527
rect 203 367 305 527
rect 203 299 237 367
rect 339 333 429 493
rect 271 299 429 333
rect 17 17 69 177
rect 271 265 320 299
rect 192 215 320 265
rect 813 299 879 527
rect 203 17 252 177
rect 286 170 320 215
rect 286 51 357 170
rect 397 143 879 181
rect 397 51 463 143
rect 497 17 550 109
rect 591 51 657 143
rect 701 17 755 109
rect 813 51 879 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 765 215 903 265 6 A1
port 1 nsew signal input
rlabel locali s 665 215 731 467 6 A2
port 2 nsew signal input
rlabel locali s 565 215 631 468 6 A3
port 3 nsew signal input
rlabel locali s 465 215 531 468 6 A4
port 4 nsew signal input
rlabel locali s 355 215 431 265 6 B1
port 5 nsew signal input
rlabel locali s 103 299 169 493 6 X
port 10 nsew signal output
rlabel locali s 103 176 158 299 6 X
port 10 nsew signal output
rlabel locali s 103 51 169 176 6 X
port 10 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 551562
string GDS_START 542482
<< end >>
