magic
tech sky130A
magscale 1 2
timestamp 1624855595
<< checkpaint >>
rect -1298 -1308 2034 1852
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 93 109 177
rect 174 47 204 177
rect 258 47 288 177
rect 448 47 478 177
rect 543 47 573 177
rect 627 47 657 177
<< scpmoshvt >>
rect 79 297 109 381
rect 176 297 206 497
rect 260 297 290 497
rect 448 297 478 497
rect 544 297 574 497
rect 616 297 646 497
<< ndiff >>
rect 27 149 79 177
rect 27 115 35 149
rect 69 115 79 149
rect 27 93 79 115
rect 109 149 174 177
rect 109 115 119 149
rect 153 115 174 149
rect 109 93 174 115
rect 124 47 174 93
rect 204 101 258 177
rect 204 67 214 101
rect 248 67 258 101
rect 204 47 258 67
rect 288 93 340 177
rect 288 59 298 93
rect 332 59 340 93
rect 288 47 340 59
rect 396 161 448 177
rect 396 127 404 161
rect 438 127 448 161
rect 396 93 448 127
rect 396 59 404 93
rect 438 59 448 93
rect 396 47 448 59
rect 478 133 543 177
rect 478 99 499 133
rect 533 99 543 133
rect 478 47 543 99
rect 573 95 627 177
rect 573 61 583 95
rect 617 61 627 95
rect 573 47 627 61
rect 657 163 709 177
rect 657 129 667 163
rect 701 129 709 163
rect 657 95 709 129
rect 657 61 667 95
rect 701 61 709 95
rect 657 47 709 61
<< pdiff >>
rect 124 475 176 497
rect 124 441 132 475
rect 166 441 176 475
rect 124 381 176 441
rect 27 349 79 381
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 176 381
rect 206 339 260 497
rect 206 305 216 339
rect 250 305 260 339
rect 206 297 260 305
rect 290 475 448 497
rect 290 441 304 475
rect 338 441 396 475
rect 430 441 448 475
rect 290 297 448 441
rect 478 477 544 497
rect 478 443 500 477
rect 534 443 544 477
rect 478 409 544 443
rect 478 375 500 409
rect 534 375 544 409
rect 478 341 544 375
rect 478 307 500 341
rect 534 307 544 341
rect 478 297 544 307
rect 574 297 616 497
rect 646 477 702 497
rect 646 443 656 477
rect 690 443 702 477
rect 646 409 702 443
rect 646 375 656 409
rect 690 375 702 409
rect 646 297 702 375
<< ndiffc >>
rect 35 115 69 149
rect 119 115 153 149
rect 214 67 248 101
rect 298 59 332 93
rect 404 127 438 161
rect 404 59 438 93
rect 499 99 533 133
rect 583 61 617 95
rect 667 129 701 163
rect 667 61 701 95
<< pdiffc >>
rect 132 441 166 475
rect 35 315 69 349
rect 216 305 250 339
rect 304 441 338 475
rect 396 441 430 475
rect 500 443 534 477
rect 500 375 534 409
rect 500 307 534 341
rect 656 443 690 477
rect 656 375 690 409
<< poly >>
rect 176 497 206 523
rect 260 497 290 523
rect 448 497 478 523
rect 544 497 574 523
rect 616 497 646 523
rect 79 381 109 407
rect 79 265 109 297
rect 176 265 206 297
rect 260 265 290 297
rect 448 265 478 297
rect 544 265 574 297
rect 75 249 129 265
rect 75 215 85 249
rect 119 215 129 249
rect 75 199 129 215
rect 174 249 301 265
rect 174 215 257 249
rect 291 215 301 249
rect 174 199 301 215
rect 343 249 478 265
rect 343 215 353 249
rect 387 215 478 249
rect 343 199 478 215
rect 520 249 574 265
rect 520 215 530 249
rect 564 215 574 249
rect 520 199 574 215
rect 616 265 646 297
rect 616 249 686 265
rect 616 215 636 249
rect 670 215 686 249
rect 616 199 686 215
rect 79 177 109 199
rect 174 177 204 199
rect 258 177 288 199
rect 448 177 478 199
rect 543 177 573 199
rect 627 177 657 199
rect 79 67 109 93
rect 174 21 204 47
rect 258 21 288 47
rect 448 21 478 47
rect 543 21 573 47
rect 627 21 657 47
<< polycont >>
rect 85 215 119 249
rect 257 215 291 249
rect 353 215 387 249
rect 530 215 564 249
rect 636 215 670 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 104 475 182 527
rect 104 441 132 475
rect 166 441 182 475
rect 283 475 446 527
rect 283 441 304 475
rect 338 441 396 475
rect 430 441 446 475
rect 480 477 545 493
rect 480 443 500 477
rect 534 443 545 477
rect 480 409 545 443
rect 480 407 500 409
rect 17 373 387 407
rect 17 349 79 373
rect 17 315 35 349
rect 69 315 79 349
rect 17 299 79 315
rect 17 165 51 299
rect 119 265 155 339
rect 85 249 155 265
rect 119 215 155 249
rect 85 199 155 215
rect 189 305 216 339
rect 250 305 270 339
rect 189 299 270 305
rect 17 149 69 165
rect 17 115 35 149
rect 17 86 69 115
rect 119 149 155 165
rect 153 115 155 149
rect 119 17 155 115
rect 189 119 223 299
rect 257 249 291 265
rect 257 212 291 215
rect 353 249 387 373
rect 257 178 319 212
rect 353 199 387 215
rect 421 375 500 407
rect 534 375 545 409
rect 640 477 706 527
rect 640 443 656 477
rect 690 443 706 477
rect 640 409 706 443
rect 640 375 656 409
rect 690 375 706 409
rect 421 341 545 375
rect 421 307 500 341
rect 534 307 545 341
rect 421 291 545 307
rect 285 165 319 178
rect 421 165 455 291
rect 489 249 586 257
rect 489 215 530 249
rect 564 215 586 249
rect 620 249 719 325
rect 620 215 636 249
rect 670 215 719 249
rect 285 161 455 165
rect 285 131 404 161
rect 388 127 404 131
rect 438 127 455 161
rect 189 101 248 119
rect 189 67 214 101
rect 189 51 248 67
rect 282 93 354 97
rect 282 59 298 93
rect 332 59 354 93
rect 282 17 354 59
rect 388 93 455 127
rect 388 59 404 93
rect 438 59 455 93
rect 489 163 718 181
rect 489 147 667 163
rect 489 133 549 147
rect 489 99 499 133
rect 533 99 549 133
rect 651 129 667 147
rect 701 129 718 163
rect 489 73 549 99
rect 583 95 617 111
rect 388 51 455 59
rect 583 17 617 61
rect 651 95 718 129
rect 651 61 667 95
rect 701 61 718 95
rect 651 54 718 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 121 221 155 255 0 FreeSans 400 180 0 0 B1_N
port 3 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 85 247 119 0 FreeSans 400 180 0 0 X
port 8 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o21ba_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3683382
string GDS_START 3677094
string path 0.000 0.000 18.400 0.000 
<< end >>
