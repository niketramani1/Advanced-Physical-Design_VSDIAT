magic
tech sky130A
timestamp 1624855461
<< properties >>
string gencell sky130_fd_pr__rf_npn_05v5_W1p00L2p00
string parameter m=1
string library sky130
<< end >>
