magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1234 -1234 5270 4674
<< nwell >>
rect 180 180 3856 3260
<< pwell >>
rect 26 3286 4010 3414
rect 26 154 154 3286
rect 3882 154 4010 3286
rect 26 26 4010 154
<< psubdiff >>
rect 26 3390 4010 3414
rect 26 3356 154 3390
rect 188 3356 222 3390
rect 256 3356 290 3390
rect 324 3356 358 3390
rect 392 3356 426 3390
rect 460 3356 494 3390
rect 528 3356 562 3390
rect 596 3356 630 3390
rect 664 3356 698 3390
rect 732 3356 766 3390
rect 800 3356 834 3390
rect 868 3356 902 3390
rect 936 3356 970 3390
rect 1004 3356 1038 3390
rect 1072 3356 1106 3390
rect 1140 3356 1174 3390
rect 1208 3356 1242 3390
rect 1276 3356 1310 3390
rect 1344 3356 1378 3390
rect 1412 3356 1446 3390
rect 1480 3356 1514 3390
rect 1548 3356 1582 3390
rect 1616 3356 1650 3390
rect 1684 3356 1718 3390
rect 1752 3356 1786 3390
rect 1820 3356 1854 3390
rect 1888 3356 1922 3390
rect 1956 3356 1990 3390
rect 2024 3356 2058 3390
rect 2092 3356 2126 3390
rect 2160 3356 2194 3390
rect 2228 3356 2262 3390
rect 2296 3356 2330 3390
rect 2364 3356 2398 3390
rect 2432 3356 2466 3390
rect 2500 3356 2534 3390
rect 2568 3356 2602 3390
rect 2636 3356 2670 3390
rect 2704 3356 2738 3390
rect 2772 3356 2806 3390
rect 2840 3356 2874 3390
rect 2908 3356 2942 3390
rect 2976 3356 3010 3390
rect 3044 3356 3078 3390
rect 3112 3356 3146 3390
rect 3180 3356 3214 3390
rect 3248 3356 3282 3390
rect 3316 3356 3350 3390
rect 3384 3356 3418 3390
rect 3452 3356 3486 3390
rect 3520 3356 3554 3390
rect 3588 3356 3622 3390
rect 3656 3356 3690 3390
rect 3724 3356 3758 3390
rect 3792 3356 3826 3390
rect 3860 3356 3894 3390
rect 3928 3356 4010 3390
rect 26 3301 4010 3356
rect 26 3267 50 3301
rect 84 3286 3952 3301
rect 84 3267 154 3286
rect 26 3233 154 3267
rect 26 3199 50 3233
rect 84 3199 154 3233
rect 26 3165 154 3199
rect 26 3131 50 3165
rect 84 3131 154 3165
rect 26 3097 154 3131
rect 26 3063 50 3097
rect 84 3063 154 3097
rect 26 3029 154 3063
rect 26 2995 50 3029
rect 84 2995 154 3029
rect 26 2961 154 2995
rect 26 2927 50 2961
rect 84 2927 154 2961
rect 26 2893 154 2927
rect 26 2859 50 2893
rect 84 2859 154 2893
rect 26 2825 154 2859
rect 26 2791 50 2825
rect 84 2791 154 2825
rect 26 2757 154 2791
rect 26 2723 50 2757
rect 84 2723 154 2757
rect 26 2689 154 2723
rect 26 2655 50 2689
rect 84 2655 154 2689
rect 26 2621 154 2655
rect 26 2587 50 2621
rect 84 2587 154 2621
rect 26 2553 154 2587
rect 26 2519 50 2553
rect 84 2519 154 2553
rect 26 2485 154 2519
rect 26 2451 50 2485
rect 84 2451 154 2485
rect 26 2417 154 2451
rect 26 2383 50 2417
rect 84 2383 154 2417
rect 26 2349 154 2383
rect 26 2315 50 2349
rect 84 2315 154 2349
rect 26 2281 154 2315
rect 26 2247 50 2281
rect 84 2247 154 2281
rect 26 2213 154 2247
rect 26 2179 50 2213
rect 84 2179 154 2213
rect 26 2145 154 2179
rect 26 2111 50 2145
rect 84 2111 154 2145
rect 26 2077 154 2111
rect 26 2043 50 2077
rect 84 2043 154 2077
rect 26 2009 154 2043
rect 26 1975 50 2009
rect 84 1975 154 2009
rect 26 1941 154 1975
rect 26 1907 50 1941
rect 84 1907 154 1941
rect 26 1873 154 1907
rect 26 1839 50 1873
rect 84 1839 154 1873
rect 26 1805 154 1839
rect 26 1771 50 1805
rect 84 1771 154 1805
rect 26 1737 154 1771
rect 26 1703 50 1737
rect 84 1703 154 1737
rect 26 1669 154 1703
rect 26 1635 50 1669
rect 84 1635 154 1669
rect 26 1601 154 1635
rect 26 1567 50 1601
rect 84 1567 154 1601
rect 26 1533 154 1567
rect 26 1499 50 1533
rect 84 1499 154 1533
rect 26 1465 154 1499
rect 26 1431 50 1465
rect 84 1431 154 1465
rect 26 1397 154 1431
rect 26 1363 50 1397
rect 84 1363 154 1397
rect 26 1329 154 1363
rect 26 1295 50 1329
rect 84 1295 154 1329
rect 26 1261 154 1295
rect 26 1227 50 1261
rect 84 1227 154 1261
rect 26 1193 154 1227
rect 26 1159 50 1193
rect 84 1159 154 1193
rect 26 1125 154 1159
rect 26 1091 50 1125
rect 84 1091 154 1125
rect 26 1057 154 1091
rect 26 1023 50 1057
rect 84 1023 154 1057
rect 26 989 154 1023
rect 26 955 50 989
rect 84 955 154 989
rect 26 921 154 955
rect 26 887 50 921
rect 84 887 154 921
rect 26 853 154 887
rect 26 819 50 853
rect 84 819 154 853
rect 26 785 154 819
rect 26 751 50 785
rect 84 751 154 785
rect 26 717 154 751
rect 26 683 50 717
rect 84 683 154 717
rect 26 649 154 683
rect 26 615 50 649
rect 84 615 154 649
rect 26 581 154 615
rect 26 547 50 581
rect 84 547 154 581
rect 26 513 154 547
rect 26 479 50 513
rect 84 479 154 513
rect 26 445 154 479
rect 26 411 50 445
rect 84 411 154 445
rect 26 377 154 411
rect 26 343 50 377
rect 84 343 154 377
rect 26 309 154 343
rect 26 275 50 309
rect 84 275 154 309
rect 26 241 154 275
rect 26 207 50 241
rect 84 207 154 241
rect 26 173 154 207
rect 26 139 50 173
rect 84 154 154 173
rect 3882 3267 3952 3286
rect 3986 3267 4010 3301
rect 3882 3233 4010 3267
rect 3882 3199 3952 3233
rect 3986 3199 4010 3233
rect 3882 3165 4010 3199
rect 3882 3131 3952 3165
rect 3986 3131 4010 3165
rect 3882 3097 4010 3131
rect 3882 3063 3952 3097
rect 3986 3063 4010 3097
rect 3882 3029 4010 3063
rect 3882 2995 3952 3029
rect 3986 2995 4010 3029
rect 3882 2961 4010 2995
rect 3882 2927 3952 2961
rect 3986 2927 4010 2961
rect 3882 2893 4010 2927
rect 3882 2859 3952 2893
rect 3986 2859 4010 2893
rect 3882 2825 4010 2859
rect 3882 2791 3952 2825
rect 3986 2791 4010 2825
rect 3882 2757 4010 2791
rect 3882 2723 3952 2757
rect 3986 2723 4010 2757
rect 3882 2689 4010 2723
rect 3882 2655 3952 2689
rect 3986 2655 4010 2689
rect 3882 2621 4010 2655
rect 3882 2587 3952 2621
rect 3986 2587 4010 2621
rect 3882 2553 4010 2587
rect 3882 2519 3952 2553
rect 3986 2519 4010 2553
rect 3882 2485 4010 2519
rect 3882 2451 3952 2485
rect 3986 2451 4010 2485
rect 3882 2417 4010 2451
rect 3882 2383 3952 2417
rect 3986 2383 4010 2417
rect 3882 2349 4010 2383
rect 3882 2315 3952 2349
rect 3986 2315 4010 2349
rect 3882 2281 4010 2315
rect 3882 2247 3952 2281
rect 3986 2247 4010 2281
rect 3882 2213 4010 2247
rect 3882 2179 3952 2213
rect 3986 2179 4010 2213
rect 3882 2145 4010 2179
rect 3882 2111 3952 2145
rect 3986 2111 4010 2145
rect 3882 2077 4010 2111
rect 3882 2043 3952 2077
rect 3986 2043 4010 2077
rect 3882 2009 4010 2043
rect 3882 1975 3952 2009
rect 3986 1975 4010 2009
rect 3882 1941 4010 1975
rect 3882 1907 3952 1941
rect 3986 1907 4010 1941
rect 3882 1873 4010 1907
rect 3882 1839 3952 1873
rect 3986 1839 4010 1873
rect 3882 1805 4010 1839
rect 3882 1771 3952 1805
rect 3986 1771 4010 1805
rect 3882 1737 4010 1771
rect 3882 1703 3952 1737
rect 3986 1703 4010 1737
rect 3882 1669 4010 1703
rect 3882 1635 3952 1669
rect 3986 1635 4010 1669
rect 3882 1601 4010 1635
rect 3882 1567 3952 1601
rect 3986 1567 4010 1601
rect 3882 1533 4010 1567
rect 3882 1499 3952 1533
rect 3986 1499 4010 1533
rect 3882 1465 4010 1499
rect 3882 1431 3952 1465
rect 3986 1431 4010 1465
rect 3882 1397 4010 1431
rect 3882 1363 3952 1397
rect 3986 1363 4010 1397
rect 3882 1329 4010 1363
rect 3882 1295 3952 1329
rect 3986 1295 4010 1329
rect 3882 1261 4010 1295
rect 3882 1227 3952 1261
rect 3986 1227 4010 1261
rect 3882 1193 4010 1227
rect 3882 1159 3952 1193
rect 3986 1159 4010 1193
rect 3882 1125 4010 1159
rect 3882 1091 3952 1125
rect 3986 1091 4010 1125
rect 3882 1057 4010 1091
rect 3882 1023 3952 1057
rect 3986 1023 4010 1057
rect 3882 989 4010 1023
rect 3882 955 3952 989
rect 3986 955 4010 989
rect 3882 921 4010 955
rect 3882 887 3952 921
rect 3986 887 4010 921
rect 3882 853 4010 887
rect 3882 819 3952 853
rect 3986 819 4010 853
rect 3882 785 4010 819
rect 3882 751 3952 785
rect 3986 751 4010 785
rect 3882 717 4010 751
rect 3882 683 3952 717
rect 3986 683 4010 717
rect 3882 649 4010 683
rect 3882 615 3952 649
rect 3986 615 4010 649
rect 3882 581 4010 615
rect 3882 547 3952 581
rect 3986 547 4010 581
rect 3882 513 4010 547
rect 3882 479 3952 513
rect 3986 479 4010 513
rect 3882 445 4010 479
rect 3882 411 3952 445
rect 3986 411 4010 445
rect 3882 377 4010 411
rect 3882 343 3952 377
rect 3986 343 4010 377
rect 3882 309 4010 343
rect 3882 275 3952 309
rect 3986 275 4010 309
rect 3882 241 4010 275
rect 3882 207 3952 241
rect 3986 207 4010 241
rect 3882 173 4010 207
rect 3882 154 3952 173
rect 84 139 3952 154
rect 3986 139 4010 173
rect 26 84 4010 139
rect 26 50 144 84
rect 178 50 212 84
rect 246 50 280 84
rect 314 50 348 84
rect 382 50 416 84
rect 450 50 484 84
rect 518 50 552 84
rect 586 50 620 84
rect 654 50 688 84
rect 722 50 756 84
rect 790 50 824 84
rect 858 50 892 84
rect 926 50 960 84
rect 994 50 1028 84
rect 1062 50 1096 84
rect 1130 50 1164 84
rect 1198 50 1232 84
rect 1266 50 1300 84
rect 1334 50 1368 84
rect 1402 50 1436 84
rect 1470 50 1504 84
rect 1538 50 1572 84
rect 1606 50 1640 84
rect 1674 50 1708 84
rect 1742 50 1776 84
rect 1810 50 1844 84
rect 1878 50 1912 84
rect 1946 50 1980 84
rect 2014 50 2048 84
rect 2082 50 2116 84
rect 2150 50 2184 84
rect 2218 50 2252 84
rect 2286 50 2320 84
rect 2354 50 2388 84
rect 2422 50 2456 84
rect 2490 50 2524 84
rect 2558 50 2592 84
rect 2626 50 2660 84
rect 2694 50 2728 84
rect 2762 50 2796 84
rect 2830 50 2864 84
rect 2898 50 2932 84
rect 2966 50 3000 84
rect 3034 50 3068 84
rect 3102 50 3136 84
rect 3170 50 3204 84
rect 3238 50 3272 84
rect 3306 50 3340 84
rect 3374 50 3408 84
rect 3442 50 3476 84
rect 3510 50 3544 84
rect 3578 50 3612 84
rect 3646 50 3680 84
rect 3714 50 3748 84
rect 3782 50 3816 84
rect 3850 50 3884 84
rect 3918 50 4010 84
rect 26 26 4010 50
<< psubdiffcont >>
rect 154 3356 188 3390
rect 222 3356 256 3390
rect 290 3356 324 3390
rect 358 3356 392 3390
rect 426 3356 460 3390
rect 494 3356 528 3390
rect 562 3356 596 3390
rect 630 3356 664 3390
rect 698 3356 732 3390
rect 766 3356 800 3390
rect 834 3356 868 3390
rect 902 3356 936 3390
rect 970 3356 1004 3390
rect 1038 3356 1072 3390
rect 1106 3356 1140 3390
rect 1174 3356 1208 3390
rect 1242 3356 1276 3390
rect 1310 3356 1344 3390
rect 1378 3356 1412 3390
rect 1446 3356 1480 3390
rect 1514 3356 1548 3390
rect 1582 3356 1616 3390
rect 1650 3356 1684 3390
rect 1718 3356 1752 3390
rect 1786 3356 1820 3390
rect 1854 3356 1888 3390
rect 1922 3356 1956 3390
rect 1990 3356 2024 3390
rect 2058 3356 2092 3390
rect 2126 3356 2160 3390
rect 2194 3356 2228 3390
rect 2262 3356 2296 3390
rect 2330 3356 2364 3390
rect 2398 3356 2432 3390
rect 2466 3356 2500 3390
rect 2534 3356 2568 3390
rect 2602 3356 2636 3390
rect 2670 3356 2704 3390
rect 2738 3356 2772 3390
rect 2806 3356 2840 3390
rect 2874 3356 2908 3390
rect 2942 3356 2976 3390
rect 3010 3356 3044 3390
rect 3078 3356 3112 3390
rect 3146 3356 3180 3390
rect 3214 3356 3248 3390
rect 3282 3356 3316 3390
rect 3350 3356 3384 3390
rect 3418 3356 3452 3390
rect 3486 3356 3520 3390
rect 3554 3356 3588 3390
rect 3622 3356 3656 3390
rect 3690 3356 3724 3390
rect 3758 3356 3792 3390
rect 3826 3356 3860 3390
rect 3894 3356 3928 3390
rect 50 3267 84 3301
rect 50 3199 84 3233
rect 50 3131 84 3165
rect 50 3063 84 3097
rect 50 2995 84 3029
rect 50 2927 84 2961
rect 50 2859 84 2893
rect 50 2791 84 2825
rect 50 2723 84 2757
rect 50 2655 84 2689
rect 50 2587 84 2621
rect 50 2519 84 2553
rect 50 2451 84 2485
rect 50 2383 84 2417
rect 50 2315 84 2349
rect 50 2247 84 2281
rect 50 2179 84 2213
rect 50 2111 84 2145
rect 50 2043 84 2077
rect 50 1975 84 2009
rect 50 1907 84 1941
rect 50 1839 84 1873
rect 50 1771 84 1805
rect 50 1703 84 1737
rect 50 1635 84 1669
rect 50 1567 84 1601
rect 50 1499 84 1533
rect 50 1431 84 1465
rect 50 1363 84 1397
rect 50 1295 84 1329
rect 50 1227 84 1261
rect 50 1159 84 1193
rect 50 1091 84 1125
rect 50 1023 84 1057
rect 50 955 84 989
rect 50 887 84 921
rect 50 819 84 853
rect 50 751 84 785
rect 50 683 84 717
rect 50 615 84 649
rect 50 547 84 581
rect 50 479 84 513
rect 50 411 84 445
rect 50 343 84 377
rect 50 275 84 309
rect 50 207 84 241
rect 50 139 84 173
rect 3952 3267 3986 3301
rect 3952 3199 3986 3233
rect 3952 3131 3986 3165
rect 3952 3063 3986 3097
rect 3952 2995 3986 3029
rect 3952 2927 3986 2961
rect 3952 2859 3986 2893
rect 3952 2791 3986 2825
rect 3952 2723 3986 2757
rect 3952 2655 3986 2689
rect 3952 2587 3986 2621
rect 3952 2519 3986 2553
rect 3952 2451 3986 2485
rect 3952 2383 3986 2417
rect 3952 2315 3986 2349
rect 3952 2247 3986 2281
rect 3952 2179 3986 2213
rect 3952 2111 3986 2145
rect 3952 2043 3986 2077
rect 3952 1975 3986 2009
rect 3952 1907 3986 1941
rect 3952 1839 3986 1873
rect 3952 1771 3986 1805
rect 3952 1703 3986 1737
rect 3952 1635 3986 1669
rect 3952 1567 3986 1601
rect 3952 1499 3986 1533
rect 3952 1431 3986 1465
rect 3952 1363 3986 1397
rect 3952 1295 3986 1329
rect 3952 1227 3986 1261
rect 3952 1159 3986 1193
rect 3952 1091 3986 1125
rect 3952 1023 3986 1057
rect 3952 955 3986 989
rect 3952 887 3986 921
rect 3952 819 3986 853
rect 3952 751 3986 785
rect 3952 683 3986 717
rect 3952 615 3986 649
rect 3952 547 3986 581
rect 3952 479 3986 513
rect 3952 411 3986 445
rect 3952 343 3986 377
rect 3952 275 3986 309
rect 3952 207 3986 241
rect 3952 139 3986 173
rect 144 50 178 84
rect 212 50 246 84
rect 280 50 314 84
rect 348 50 382 84
rect 416 50 450 84
rect 484 50 518 84
rect 552 50 586 84
rect 620 50 654 84
rect 688 50 722 84
rect 756 50 790 84
rect 824 50 858 84
rect 892 50 926 84
rect 960 50 994 84
rect 1028 50 1062 84
rect 1096 50 1130 84
rect 1164 50 1198 84
rect 1232 50 1266 84
rect 1300 50 1334 84
rect 1368 50 1402 84
rect 1436 50 1470 84
rect 1504 50 1538 84
rect 1572 50 1606 84
rect 1640 50 1674 84
rect 1708 50 1742 84
rect 1776 50 1810 84
rect 1844 50 1878 84
rect 1912 50 1946 84
rect 1980 50 2014 84
rect 2048 50 2082 84
rect 2116 50 2150 84
rect 2184 50 2218 84
rect 2252 50 2286 84
rect 2320 50 2354 84
rect 2388 50 2422 84
rect 2456 50 2490 84
rect 2524 50 2558 84
rect 2592 50 2626 84
rect 2660 50 2694 84
rect 2728 50 2762 84
rect 2796 50 2830 84
rect 2864 50 2898 84
rect 2932 50 2966 84
rect 3000 50 3034 84
rect 3068 50 3102 84
rect 3136 50 3170 84
rect 3204 50 3238 84
rect 3272 50 3306 84
rect 3340 50 3374 84
rect 3408 50 3442 84
rect 3476 50 3510 84
rect 3544 50 3578 84
rect 3612 50 3646 84
rect 3680 50 3714 84
rect 3748 50 3782 84
rect 3816 50 3850 84
rect 3884 50 3918 84
<< locali >>
rect 26 3390 4010 3414
rect 26 3356 154 3390
rect 188 3356 222 3390
rect 256 3356 290 3390
rect 324 3356 358 3390
rect 392 3356 426 3390
rect 460 3356 494 3390
rect 528 3356 562 3390
rect 596 3356 630 3390
rect 664 3356 698 3390
rect 732 3356 766 3390
rect 800 3356 834 3390
rect 868 3356 902 3390
rect 936 3356 970 3390
rect 1004 3356 1038 3390
rect 1072 3356 1106 3390
rect 1140 3356 1174 3390
rect 1208 3356 1242 3390
rect 1276 3356 1310 3390
rect 1344 3356 1378 3390
rect 1412 3356 1446 3390
rect 1480 3356 1514 3390
rect 1548 3356 1582 3390
rect 1616 3356 1650 3390
rect 1684 3356 1718 3390
rect 1752 3356 1786 3390
rect 1820 3356 1854 3390
rect 1888 3356 1922 3390
rect 1956 3356 1990 3390
rect 2024 3356 2058 3390
rect 2092 3356 2126 3390
rect 2160 3356 2194 3390
rect 2228 3356 2262 3390
rect 2296 3356 2330 3390
rect 2364 3356 2398 3390
rect 2432 3356 2466 3390
rect 2500 3356 2534 3390
rect 2568 3356 2602 3390
rect 2636 3356 2670 3390
rect 2704 3356 2738 3390
rect 2772 3356 2806 3390
rect 2840 3356 2874 3390
rect 2908 3356 2942 3390
rect 2976 3356 3010 3390
rect 3044 3356 3078 3390
rect 3112 3356 3146 3390
rect 3180 3356 3214 3390
rect 3248 3356 3282 3390
rect 3316 3356 3350 3390
rect 3384 3356 3418 3390
rect 3452 3356 3486 3390
rect 3520 3356 3554 3390
rect 3588 3356 3622 3390
rect 3656 3356 3690 3390
rect 3724 3356 3758 3390
rect 3792 3356 3826 3390
rect 3860 3356 3894 3390
rect 3928 3356 4010 3390
rect 26 3332 4010 3356
rect 26 3301 108 3332
rect 26 3267 50 3301
rect 84 3267 108 3301
rect 26 3233 108 3267
rect 26 3199 50 3233
rect 84 3199 108 3233
rect 26 3165 108 3199
rect 26 3131 50 3165
rect 84 3131 108 3165
rect 26 3097 108 3131
rect 26 3063 50 3097
rect 84 3074 108 3097
rect 26 3040 53 3063
rect 87 3040 108 3074
rect 26 3029 108 3040
rect 26 2995 50 3029
rect 84 3002 108 3029
rect 26 2968 53 2995
rect 87 2968 108 3002
rect 26 2961 108 2968
rect 26 2927 50 2961
rect 84 2930 108 2961
rect 26 2896 53 2927
rect 87 2896 108 2930
rect 26 2893 108 2896
rect 26 2859 50 2893
rect 84 2859 108 2893
rect 26 2858 108 2859
rect 26 2825 53 2858
rect 26 2791 50 2825
rect 87 2824 108 2858
rect 84 2791 108 2824
rect 26 2786 108 2791
rect 26 2757 53 2786
rect 26 2723 50 2757
rect 87 2752 108 2786
rect 84 2723 108 2752
rect 26 2714 108 2723
rect 26 2689 53 2714
rect 26 2655 50 2689
rect 87 2680 108 2714
rect 84 2655 108 2680
rect 26 2642 108 2655
rect 26 2621 53 2642
rect 26 2587 50 2621
rect 87 2608 108 2642
rect 84 2587 108 2608
rect 26 2570 108 2587
rect 26 2553 53 2570
rect 26 2519 50 2553
rect 87 2536 108 2570
rect 84 2519 108 2536
rect 26 2498 108 2519
rect 26 2485 53 2498
rect 26 2451 50 2485
rect 87 2464 108 2498
rect 84 2451 108 2464
rect 26 2426 108 2451
rect 26 2417 53 2426
rect 26 2383 50 2417
rect 87 2392 108 2426
rect 84 2383 108 2392
rect 26 2354 108 2383
rect 26 2349 53 2354
rect 26 2315 50 2349
rect 87 2320 108 2354
rect 84 2315 108 2320
rect 26 2282 108 2315
rect 26 2281 53 2282
rect 26 2247 50 2281
rect 87 2248 108 2282
rect 84 2247 108 2248
rect 26 2213 108 2247
rect 26 2179 50 2213
rect 84 2210 108 2213
rect 26 2176 53 2179
rect 87 2176 108 2210
rect 26 2145 108 2176
rect 26 2111 50 2145
rect 84 2138 108 2145
rect 26 2104 53 2111
rect 87 2104 108 2138
rect 26 2077 108 2104
rect 26 2043 50 2077
rect 84 2066 108 2077
rect 26 2032 53 2043
rect 87 2032 108 2066
rect 26 2009 108 2032
rect 26 1975 50 2009
rect 84 1994 108 2009
rect 26 1960 53 1975
rect 87 1960 108 1994
rect 26 1941 108 1960
rect 26 1907 50 1941
rect 84 1922 108 1941
rect 26 1888 53 1907
rect 87 1888 108 1922
rect 26 1873 108 1888
rect 26 1839 50 1873
rect 84 1850 108 1873
rect 26 1816 53 1839
rect 87 1816 108 1850
rect 26 1805 108 1816
rect 26 1771 50 1805
rect 84 1778 108 1805
rect 26 1744 53 1771
rect 87 1744 108 1778
rect 26 1737 108 1744
rect 26 1703 50 1737
rect 84 1706 108 1737
rect 26 1672 53 1703
rect 87 1672 108 1706
rect 26 1669 108 1672
rect 26 1635 50 1669
rect 84 1635 108 1669
rect 26 1634 108 1635
rect 26 1601 53 1634
rect 26 1567 50 1601
rect 87 1600 108 1634
rect 84 1567 108 1600
rect 26 1562 108 1567
rect 26 1533 53 1562
rect 26 1499 50 1533
rect 87 1528 108 1562
rect 84 1499 108 1528
rect 26 1490 108 1499
rect 26 1465 53 1490
rect 26 1431 50 1465
rect 87 1456 108 1490
rect 84 1431 108 1456
rect 26 1418 108 1431
rect 26 1397 53 1418
rect 26 1363 50 1397
rect 87 1384 108 1418
rect 84 1363 108 1384
rect 26 1346 108 1363
rect 26 1329 53 1346
rect 26 1295 50 1329
rect 87 1312 108 1346
rect 84 1295 108 1312
rect 26 1274 108 1295
rect 26 1261 53 1274
rect 26 1227 50 1261
rect 87 1240 108 1274
rect 84 1227 108 1240
rect 26 1202 108 1227
rect 26 1193 53 1202
rect 26 1159 50 1193
rect 87 1168 108 1202
rect 84 1159 108 1168
rect 26 1130 108 1159
rect 26 1125 53 1130
rect 26 1091 50 1125
rect 87 1096 108 1130
rect 84 1091 108 1096
rect 26 1058 108 1091
rect 26 1057 53 1058
rect 26 1023 50 1057
rect 87 1024 108 1058
rect 84 1023 108 1024
rect 26 989 108 1023
rect 26 955 50 989
rect 84 986 108 989
rect 26 952 53 955
rect 87 952 108 986
rect 26 921 108 952
rect 26 887 50 921
rect 84 914 108 921
rect 26 880 53 887
rect 87 880 108 914
rect 26 853 108 880
rect 26 819 50 853
rect 84 842 108 853
rect 26 808 53 819
rect 87 808 108 842
rect 26 785 108 808
rect 26 751 50 785
rect 84 770 108 785
rect 26 736 53 751
rect 87 736 108 770
rect 26 717 108 736
rect 26 683 50 717
rect 84 698 108 717
rect 26 664 53 683
rect 87 664 108 698
rect 26 649 108 664
rect 26 615 50 649
rect 84 626 108 649
rect 26 592 53 615
rect 87 592 108 626
rect 26 581 108 592
rect 26 547 50 581
rect 84 554 108 581
rect 26 520 53 547
rect 87 520 108 554
rect 26 513 108 520
rect 26 479 50 513
rect 84 482 108 513
rect 26 448 53 479
rect 87 448 108 482
rect 26 445 108 448
rect 26 411 50 445
rect 84 411 108 445
rect 26 410 108 411
rect 26 377 53 410
rect 26 343 50 377
rect 87 376 108 410
rect 84 343 108 376
rect 26 338 108 343
rect 26 309 53 338
rect 26 275 50 309
rect 87 304 108 338
rect 84 275 108 304
rect 26 266 108 275
rect 26 241 53 266
rect 26 207 50 241
rect 87 232 108 266
rect 84 207 108 232
rect 26 194 108 207
rect 26 173 53 194
rect 87 180 108 194
rect 3928 3301 4010 3332
rect 3928 3267 3952 3301
rect 3986 3267 4010 3301
rect 3928 3233 4010 3267
rect 3928 3199 3952 3233
rect 3986 3199 4010 3233
rect 3928 3165 4010 3199
rect 3928 3131 3952 3165
rect 3986 3131 4010 3165
rect 3928 3097 4010 3131
rect 3928 3063 3952 3097
rect 3986 3074 4010 3097
rect 3928 3040 3955 3063
rect 3989 3040 4010 3074
rect 3928 3029 4010 3040
rect 3928 2995 3952 3029
rect 3986 3002 4010 3029
rect 3928 2968 3955 2995
rect 3989 2968 4010 3002
rect 3928 2961 4010 2968
rect 3928 2927 3952 2961
rect 3986 2930 4010 2961
rect 3928 2896 3955 2927
rect 3989 2896 4010 2930
rect 3928 2893 4010 2896
rect 3928 2859 3952 2893
rect 3986 2859 4010 2893
rect 3928 2858 4010 2859
rect 3928 2825 3955 2858
rect 3928 2791 3952 2825
rect 3989 2824 4010 2858
rect 3986 2791 4010 2824
rect 3928 2786 4010 2791
rect 3928 2757 3955 2786
rect 3928 2723 3952 2757
rect 3989 2752 4010 2786
rect 3986 2723 4010 2752
rect 3928 2714 4010 2723
rect 3928 2689 3955 2714
rect 3928 2655 3952 2689
rect 3989 2680 4010 2714
rect 3986 2655 4010 2680
rect 3928 2642 4010 2655
rect 3928 2621 3955 2642
rect 3928 2587 3952 2621
rect 3989 2608 4010 2642
rect 3986 2587 4010 2608
rect 3928 2570 4010 2587
rect 3928 2553 3955 2570
rect 3928 2519 3952 2553
rect 3989 2536 4010 2570
rect 3986 2519 4010 2536
rect 3928 2498 4010 2519
rect 3928 2485 3955 2498
rect 3928 2451 3952 2485
rect 3989 2464 4010 2498
rect 3986 2451 4010 2464
rect 3928 2426 4010 2451
rect 3928 2417 3955 2426
rect 3928 2383 3952 2417
rect 3989 2392 4010 2426
rect 3986 2383 4010 2392
rect 3928 2354 4010 2383
rect 3928 2349 3955 2354
rect 3928 2315 3952 2349
rect 3989 2320 4010 2354
rect 3986 2315 4010 2320
rect 3928 2282 4010 2315
rect 3928 2281 3955 2282
rect 3928 2247 3952 2281
rect 3989 2248 4010 2282
rect 3986 2247 4010 2248
rect 3928 2213 4010 2247
rect 3928 2179 3952 2213
rect 3986 2210 4010 2213
rect 3928 2176 3955 2179
rect 3989 2176 4010 2210
rect 3928 2145 4010 2176
rect 3928 2111 3952 2145
rect 3986 2138 4010 2145
rect 3928 2104 3955 2111
rect 3989 2104 4010 2138
rect 3928 2077 4010 2104
rect 3928 2043 3952 2077
rect 3986 2066 4010 2077
rect 3928 2032 3955 2043
rect 3989 2032 4010 2066
rect 3928 2009 4010 2032
rect 3928 1975 3952 2009
rect 3986 1994 4010 2009
rect 3928 1960 3955 1975
rect 3989 1960 4010 1994
rect 3928 1941 4010 1960
rect 3928 1907 3952 1941
rect 3986 1922 4010 1941
rect 3928 1888 3955 1907
rect 3989 1888 4010 1922
rect 3928 1873 4010 1888
rect 3928 1839 3952 1873
rect 3986 1850 4010 1873
rect 3928 1816 3955 1839
rect 3989 1816 4010 1850
rect 3928 1805 4010 1816
rect 3928 1771 3952 1805
rect 3986 1778 4010 1805
rect 3928 1744 3955 1771
rect 3989 1744 4010 1778
rect 3928 1737 4010 1744
rect 3928 1703 3952 1737
rect 3986 1706 4010 1737
rect 3928 1672 3955 1703
rect 3989 1672 4010 1706
rect 3928 1669 4010 1672
rect 3928 1635 3952 1669
rect 3986 1635 4010 1669
rect 3928 1634 4010 1635
rect 3928 1601 3955 1634
rect 3928 1567 3952 1601
rect 3989 1600 4010 1634
rect 3986 1567 4010 1600
rect 3928 1562 4010 1567
rect 3928 1533 3955 1562
rect 3928 1499 3952 1533
rect 3989 1528 4010 1562
rect 3986 1499 4010 1528
rect 3928 1490 4010 1499
rect 3928 1465 3955 1490
rect 3928 1431 3952 1465
rect 3989 1456 4010 1490
rect 3986 1431 4010 1456
rect 3928 1418 4010 1431
rect 3928 1397 3955 1418
rect 3928 1363 3952 1397
rect 3989 1384 4010 1418
rect 3986 1363 4010 1384
rect 3928 1346 4010 1363
rect 3928 1329 3955 1346
rect 3928 1295 3952 1329
rect 3989 1312 4010 1346
rect 3986 1295 4010 1312
rect 3928 1274 4010 1295
rect 3928 1261 3955 1274
rect 3928 1227 3952 1261
rect 3989 1240 4010 1274
rect 3986 1227 4010 1240
rect 3928 1202 4010 1227
rect 3928 1193 3955 1202
rect 3928 1159 3952 1193
rect 3989 1168 4010 1202
rect 3986 1159 4010 1168
rect 3928 1130 4010 1159
rect 3928 1125 3955 1130
rect 3928 1091 3952 1125
rect 3989 1096 4010 1130
rect 3986 1091 4010 1096
rect 3928 1058 4010 1091
rect 3928 1057 3955 1058
rect 3928 1023 3952 1057
rect 3989 1024 4010 1058
rect 3986 1023 4010 1024
rect 3928 989 4010 1023
rect 3928 955 3952 989
rect 3986 986 4010 989
rect 3928 952 3955 955
rect 3989 952 4010 986
rect 3928 921 4010 952
rect 3928 887 3952 921
rect 3986 914 4010 921
rect 3928 880 3955 887
rect 3989 880 4010 914
rect 3928 853 4010 880
rect 3928 819 3952 853
rect 3986 842 4010 853
rect 3928 808 3955 819
rect 3989 808 4010 842
rect 3928 785 4010 808
rect 3928 751 3952 785
rect 3986 770 4010 785
rect 3928 736 3955 751
rect 3989 736 4010 770
rect 3928 717 4010 736
rect 3928 683 3952 717
rect 3986 698 4010 717
rect 3928 664 3955 683
rect 3989 664 4010 698
rect 3928 649 4010 664
rect 3928 615 3952 649
rect 3986 626 4010 649
rect 3928 592 3955 615
rect 3989 592 4010 626
rect 3928 581 4010 592
rect 3928 547 3952 581
rect 3986 554 4010 581
rect 3928 520 3955 547
rect 3989 520 4010 554
rect 3928 513 4010 520
rect 3928 479 3952 513
rect 3986 482 4010 513
rect 3928 448 3955 479
rect 3989 448 4010 482
rect 3928 445 4010 448
rect 3928 411 3952 445
rect 3986 411 4010 445
rect 3928 410 4010 411
rect 3928 377 3955 410
rect 3928 343 3952 377
rect 3989 376 4010 410
rect 3986 343 4010 376
rect 3928 338 4010 343
rect 3928 309 3955 338
rect 3928 275 3952 309
rect 3989 304 4010 338
rect 3986 275 4010 304
rect 3928 266 4010 275
rect 3928 241 3955 266
rect 3928 207 3952 241
rect 3989 232 4010 266
rect 3986 207 4010 232
rect 3928 194 4010 207
rect 3928 180 3955 194
rect 87 173 3955 180
rect 26 139 50 173
rect 87 160 3952 173
rect 3989 160 4010 194
rect 84 139 3952 160
rect 3986 139 4010 160
rect 26 84 4010 139
rect 26 50 144 84
rect 178 50 212 84
rect 246 50 280 84
rect 314 50 348 84
rect 382 50 416 84
rect 450 50 484 84
rect 518 50 552 84
rect 586 50 620 84
rect 654 50 688 84
rect 722 50 756 84
rect 790 50 824 84
rect 858 50 892 84
rect 926 50 960 84
rect 994 50 1028 84
rect 1062 50 1096 84
rect 1130 50 1164 84
rect 1198 50 1232 84
rect 1266 50 1300 84
rect 1334 50 1368 84
rect 1402 50 1436 84
rect 1470 50 1504 84
rect 1538 50 1572 84
rect 1606 50 1640 84
rect 1674 50 1708 84
rect 1742 50 1776 84
rect 1810 50 1844 84
rect 1878 50 1912 84
rect 1946 50 1980 84
rect 2014 50 2048 84
rect 2082 50 2116 84
rect 2150 50 2184 84
rect 2218 50 2252 84
rect 2286 50 2320 84
rect 2354 50 2388 84
rect 2422 50 2456 84
rect 2490 50 2524 84
rect 2558 50 2592 84
rect 2626 50 2660 84
rect 2694 50 2728 84
rect 2762 50 2796 84
rect 2830 50 2864 84
rect 2898 50 2932 84
rect 2966 50 3000 84
rect 3034 50 3068 84
rect 3102 50 3136 84
rect 3170 50 3204 84
rect 3238 50 3272 84
rect 3306 50 3340 84
rect 3374 50 3408 84
rect 3442 50 3476 84
rect 3510 50 3544 84
rect 3578 50 3612 84
rect 3646 50 3680 84
rect 3714 50 3748 84
rect 3782 50 3816 84
rect 3850 50 3884 84
rect 3918 50 4010 84
rect 26 26 4010 50
<< viali >>
rect 53 3063 84 3074
rect 84 3063 87 3074
rect 53 3040 87 3063
rect 53 2995 84 3002
rect 84 2995 87 3002
rect 53 2968 87 2995
rect 53 2927 84 2930
rect 84 2927 87 2930
rect 53 2896 87 2927
rect 53 2825 87 2858
rect 53 2824 84 2825
rect 84 2824 87 2825
rect 53 2757 87 2786
rect 53 2752 84 2757
rect 84 2752 87 2757
rect 53 2689 87 2714
rect 53 2680 84 2689
rect 84 2680 87 2689
rect 53 2621 87 2642
rect 53 2608 84 2621
rect 84 2608 87 2621
rect 53 2553 87 2570
rect 53 2536 84 2553
rect 84 2536 87 2553
rect 53 2485 87 2498
rect 53 2464 84 2485
rect 84 2464 87 2485
rect 53 2417 87 2426
rect 53 2392 84 2417
rect 84 2392 87 2417
rect 53 2349 87 2354
rect 53 2320 84 2349
rect 84 2320 87 2349
rect 53 2281 87 2282
rect 53 2248 84 2281
rect 84 2248 87 2281
rect 53 2179 84 2210
rect 84 2179 87 2210
rect 53 2176 87 2179
rect 53 2111 84 2138
rect 84 2111 87 2138
rect 53 2104 87 2111
rect 53 2043 84 2066
rect 84 2043 87 2066
rect 53 2032 87 2043
rect 53 1975 84 1994
rect 84 1975 87 1994
rect 53 1960 87 1975
rect 53 1907 84 1922
rect 84 1907 87 1922
rect 53 1888 87 1907
rect 53 1839 84 1850
rect 84 1839 87 1850
rect 53 1816 87 1839
rect 53 1771 84 1778
rect 84 1771 87 1778
rect 53 1744 87 1771
rect 53 1703 84 1706
rect 84 1703 87 1706
rect 53 1672 87 1703
rect 53 1601 87 1634
rect 53 1600 84 1601
rect 84 1600 87 1601
rect 53 1533 87 1562
rect 53 1528 84 1533
rect 84 1528 87 1533
rect 53 1465 87 1490
rect 53 1456 84 1465
rect 84 1456 87 1465
rect 53 1397 87 1418
rect 53 1384 84 1397
rect 84 1384 87 1397
rect 53 1329 87 1346
rect 53 1312 84 1329
rect 84 1312 87 1329
rect 53 1261 87 1274
rect 53 1240 84 1261
rect 84 1240 87 1261
rect 53 1193 87 1202
rect 53 1168 84 1193
rect 84 1168 87 1193
rect 53 1125 87 1130
rect 53 1096 84 1125
rect 84 1096 87 1125
rect 53 1057 87 1058
rect 53 1024 84 1057
rect 84 1024 87 1057
rect 53 955 84 986
rect 84 955 87 986
rect 53 952 87 955
rect 53 887 84 914
rect 84 887 87 914
rect 53 880 87 887
rect 53 819 84 842
rect 84 819 87 842
rect 53 808 87 819
rect 53 751 84 770
rect 84 751 87 770
rect 53 736 87 751
rect 53 683 84 698
rect 84 683 87 698
rect 53 664 87 683
rect 53 615 84 626
rect 84 615 87 626
rect 53 592 87 615
rect 53 547 84 554
rect 84 547 87 554
rect 53 520 87 547
rect 53 479 84 482
rect 84 479 87 482
rect 53 448 87 479
rect 53 377 87 410
rect 53 376 84 377
rect 84 376 87 377
rect 53 309 87 338
rect 53 304 84 309
rect 84 304 87 309
rect 53 241 87 266
rect 53 232 84 241
rect 84 232 87 241
rect 53 173 87 194
rect 3955 3063 3986 3074
rect 3986 3063 3989 3074
rect 3955 3040 3989 3063
rect 3955 2995 3986 3002
rect 3986 2995 3989 3002
rect 3955 2968 3989 2995
rect 3955 2927 3986 2930
rect 3986 2927 3989 2930
rect 3955 2896 3989 2927
rect 3955 2825 3989 2858
rect 3955 2824 3986 2825
rect 3986 2824 3989 2825
rect 3955 2757 3989 2786
rect 3955 2752 3986 2757
rect 3986 2752 3989 2757
rect 3955 2689 3989 2714
rect 3955 2680 3986 2689
rect 3986 2680 3989 2689
rect 3955 2621 3989 2642
rect 3955 2608 3986 2621
rect 3986 2608 3989 2621
rect 3955 2553 3989 2570
rect 3955 2536 3986 2553
rect 3986 2536 3989 2553
rect 3955 2485 3989 2498
rect 3955 2464 3986 2485
rect 3986 2464 3989 2485
rect 3955 2417 3989 2426
rect 3955 2392 3986 2417
rect 3986 2392 3989 2417
rect 3955 2349 3989 2354
rect 3955 2320 3986 2349
rect 3986 2320 3989 2349
rect 3955 2281 3989 2282
rect 3955 2248 3986 2281
rect 3986 2248 3989 2281
rect 3955 2179 3986 2210
rect 3986 2179 3989 2210
rect 3955 2176 3989 2179
rect 3955 2111 3986 2138
rect 3986 2111 3989 2138
rect 3955 2104 3989 2111
rect 3955 2043 3986 2066
rect 3986 2043 3989 2066
rect 3955 2032 3989 2043
rect 3955 1975 3986 1994
rect 3986 1975 3989 1994
rect 3955 1960 3989 1975
rect 3955 1907 3986 1922
rect 3986 1907 3989 1922
rect 3955 1888 3989 1907
rect 3955 1839 3986 1850
rect 3986 1839 3989 1850
rect 3955 1816 3989 1839
rect 3955 1771 3986 1778
rect 3986 1771 3989 1778
rect 3955 1744 3989 1771
rect 3955 1703 3986 1706
rect 3986 1703 3989 1706
rect 3955 1672 3989 1703
rect 3955 1601 3989 1634
rect 3955 1600 3986 1601
rect 3986 1600 3989 1601
rect 3955 1533 3989 1562
rect 3955 1528 3986 1533
rect 3986 1528 3989 1533
rect 3955 1465 3989 1490
rect 3955 1456 3986 1465
rect 3986 1456 3989 1465
rect 3955 1397 3989 1418
rect 3955 1384 3986 1397
rect 3986 1384 3989 1397
rect 3955 1329 3989 1346
rect 3955 1312 3986 1329
rect 3986 1312 3989 1329
rect 3955 1261 3989 1274
rect 3955 1240 3986 1261
rect 3986 1240 3989 1261
rect 3955 1193 3989 1202
rect 3955 1168 3986 1193
rect 3986 1168 3989 1193
rect 3955 1125 3989 1130
rect 3955 1096 3986 1125
rect 3986 1096 3989 1125
rect 3955 1057 3989 1058
rect 3955 1024 3986 1057
rect 3986 1024 3989 1057
rect 3955 955 3986 986
rect 3986 955 3989 986
rect 3955 952 3989 955
rect 3955 887 3986 914
rect 3986 887 3989 914
rect 3955 880 3989 887
rect 3955 819 3986 842
rect 3986 819 3989 842
rect 3955 808 3989 819
rect 3955 751 3986 770
rect 3986 751 3989 770
rect 3955 736 3989 751
rect 3955 683 3986 698
rect 3986 683 3989 698
rect 3955 664 3989 683
rect 3955 615 3986 626
rect 3986 615 3989 626
rect 3955 592 3989 615
rect 3955 547 3986 554
rect 3986 547 3989 554
rect 3955 520 3989 547
rect 3955 479 3986 482
rect 3986 479 3989 482
rect 3955 448 3989 479
rect 3955 377 3989 410
rect 3955 376 3986 377
rect 3986 376 3989 377
rect 3955 309 3989 338
rect 3955 304 3986 309
rect 3986 304 3989 309
rect 3955 241 3989 266
rect 3955 232 3986 241
rect 3986 232 3989 241
rect 3955 173 3989 194
rect 53 160 84 173
rect 84 160 87 173
rect 3955 160 3986 173
rect 3986 160 3989 173
<< metal1 >>
rect 26 3074 108 3087
rect 26 3040 53 3074
rect 87 3040 108 3074
rect 26 3002 108 3040
rect 26 2968 53 3002
rect 87 2968 108 3002
rect 26 2930 108 2968
rect 26 2896 53 2930
rect 87 2896 108 2930
rect 26 2858 108 2896
rect 26 2824 53 2858
rect 87 2824 108 2858
rect 26 2786 108 2824
rect 26 2752 53 2786
rect 87 2752 108 2786
rect 26 2714 108 2752
rect 26 2680 53 2714
rect 87 2680 108 2714
rect 26 2642 108 2680
rect 26 2608 53 2642
rect 87 2608 108 2642
rect 26 2570 108 2608
rect 26 2536 53 2570
rect 87 2536 108 2570
rect 26 2498 108 2536
rect 26 2464 53 2498
rect 87 2464 108 2498
rect 26 2426 108 2464
rect 26 2392 53 2426
rect 87 2392 108 2426
rect 26 2354 108 2392
rect 26 2320 53 2354
rect 87 2320 108 2354
rect 26 2282 108 2320
rect 26 2248 53 2282
rect 87 2248 108 2282
rect 26 2210 108 2248
rect 26 2176 53 2210
rect 87 2176 108 2210
rect 26 2138 108 2176
rect 26 2104 53 2138
rect 87 2104 108 2138
rect 26 2066 108 2104
rect 26 2032 53 2066
rect 87 2032 108 2066
rect 26 1994 108 2032
rect 26 1960 53 1994
rect 87 1960 108 1994
rect 26 1922 108 1960
rect 26 1888 53 1922
rect 87 1888 108 1922
rect 26 1850 108 1888
rect 26 1816 53 1850
rect 87 1816 108 1850
rect 26 1778 108 1816
rect 26 1744 53 1778
rect 87 1744 108 1778
rect 26 1706 108 1744
rect 26 1672 53 1706
rect 87 1672 108 1706
rect 26 1634 108 1672
rect 26 1600 53 1634
rect 87 1600 108 1634
rect 26 1562 108 1600
rect 26 1528 53 1562
rect 87 1528 108 1562
rect 26 1490 108 1528
rect 26 1456 53 1490
rect 87 1456 108 1490
rect 26 1418 108 1456
rect 26 1384 53 1418
rect 87 1384 108 1418
rect 26 1346 108 1384
rect 26 1312 53 1346
rect 87 1312 108 1346
rect 26 1274 108 1312
rect 26 1240 53 1274
rect 87 1240 108 1274
rect 26 1202 108 1240
rect 26 1168 53 1202
rect 87 1168 108 1202
rect 26 1130 108 1168
rect 26 1096 53 1130
rect 87 1096 108 1130
rect 26 1058 108 1096
rect 26 1024 53 1058
rect 87 1024 108 1058
rect 26 986 108 1024
rect 26 952 53 986
rect 87 952 108 986
rect 26 914 108 952
rect 26 880 53 914
rect 87 880 108 914
rect 26 842 108 880
rect 26 808 53 842
rect 87 808 108 842
rect 26 770 108 808
rect 26 736 53 770
rect 87 736 108 770
rect 26 698 108 736
rect 26 664 53 698
rect 87 664 108 698
rect 26 626 108 664
rect 26 592 53 626
rect 87 592 108 626
rect 26 554 108 592
rect 26 520 53 554
rect 87 520 108 554
rect 26 482 108 520
rect 26 448 53 482
rect 87 448 108 482
rect 26 410 108 448
rect 26 376 53 410
rect 87 376 108 410
rect 26 338 108 376
rect 26 304 53 338
rect 87 304 108 338
rect 26 266 108 304
rect 26 232 53 266
rect 87 232 108 266
rect 26 194 108 232
rect 26 160 53 194
rect 87 160 108 194
rect 26 154 108 160
rect 3928 3074 4010 3087
rect 3928 3040 3955 3074
rect 3989 3040 4010 3074
rect 3928 3002 4010 3040
rect 3928 2968 3955 3002
rect 3989 2968 4010 3002
rect 3928 2930 4010 2968
rect 3928 2896 3955 2930
rect 3989 2896 4010 2930
rect 3928 2858 4010 2896
rect 3928 2824 3955 2858
rect 3989 2824 4010 2858
rect 3928 2786 4010 2824
rect 3928 2752 3955 2786
rect 3989 2752 4010 2786
rect 3928 2714 4010 2752
rect 3928 2680 3955 2714
rect 3989 2680 4010 2714
rect 3928 2642 4010 2680
rect 3928 2608 3955 2642
rect 3989 2608 4010 2642
rect 3928 2570 4010 2608
rect 3928 2536 3955 2570
rect 3989 2536 4010 2570
rect 3928 2498 4010 2536
rect 3928 2464 3955 2498
rect 3989 2464 4010 2498
rect 3928 2426 4010 2464
rect 3928 2392 3955 2426
rect 3989 2392 4010 2426
rect 3928 2354 4010 2392
rect 3928 2320 3955 2354
rect 3989 2320 4010 2354
rect 3928 2282 4010 2320
rect 3928 2248 3955 2282
rect 3989 2248 4010 2282
rect 3928 2210 4010 2248
rect 3928 2176 3955 2210
rect 3989 2176 4010 2210
rect 3928 2138 4010 2176
rect 3928 2104 3955 2138
rect 3989 2104 4010 2138
rect 3928 2066 4010 2104
rect 3928 2032 3955 2066
rect 3989 2032 4010 2066
rect 3928 1994 4010 2032
rect 3928 1960 3955 1994
rect 3989 1960 4010 1994
rect 3928 1922 4010 1960
rect 3928 1888 3955 1922
rect 3989 1888 4010 1922
rect 3928 1850 4010 1888
rect 3928 1816 3955 1850
rect 3989 1816 4010 1850
rect 3928 1778 4010 1816
rect 3928 1744 3955 1778
rect 3989 1744 4010 1778
rect 3928 1706 4010 1744
rect 3928 1672 3955 1706
rect 3989 1672 4010 1706
rect 3928 1634 4010 1672
rect 3928 1600 3955 1634
rect 3989 1600 4010 1634
rect 3928 1562 4010 1600
rect 3928 1528 3955 1562
rect 3989 1528 4010 1562
rect 3928 1490 4010 1528
rect 3928 1456 3955 1490
rect 3989 1456 4010 1490
rect 3928 1418 4010 1456
rect 3928 1384 3955 1418
rect 3989 1384 4010 1418
rect 3928 1346 4010 1384
rect 3928 1312 3955 1346
rect 3989 1312 4010 1346
rect 3928 1274 4010 1312
rect 3928 1240 3955 1274
rect 3989 1240 4010 1274
rect 3928 1202 4010 1240
rect 3928 1168 3955 1202
rect 3989 1168 4010 1202
rect 3928 1130 4010 1168
rect 3928 1096 3955 1130
rect 3989 1096 4010 1130
rect 3928 1058 4010 1096
rect 3928 1024 3955 1058
rect 3989 1024 4010 1058
rect 3928 986 4010 1024
rect 3928 952 3955 986
rect 3989 952 4010 986
rect 3928 914 4010 952
rect 3928 880 3955 914
rect 3989 880 4010 914
rect 3928 842 4010 880
rect 3928 808 3955 842
rect 3989 808 4010 842
rect 3928 770 4010 808
rect 3928 736 3955 770
rect 3989 736 4010 770
rect 3928 698 4010 736
rect 3928 664 3955 698
rect 3989 664 4010 698
rect 3928 626 4010 664
rect 3928 592 3955 626
rect 3989 592 4010 626
rect 3928 554 4010 592
rect 3928 520 3955 554
rect 3989 520 4010 554
rect 3928 482 4010 520
rect 3928 448 3955 482
rect 3989 448 4010 482
rect 3928 410 4010 448
rect 3928 376 3955 410
rect 3989 376 4010 410
rect 3928 338 4010 376
rect 3928 304 3955 338
rect 3989 304 4010 338
rect 3928 266 4010 304
rect 3928 232 3955 266
rect 3989 232 4010 266
rect 3928 194 4010 232
rect 3928 160 3955 194
rect 3989 160 4010 194
rect 3928 154 4010 160
use sky130_fd_pr__tpl1__example_55959141808686  sky130_fd_pr__tpl1__example_55959141808686_0
timestamp 1624855509
transform -1 0 3942 0 1 26
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808686  sky130_fd_pr__tpl1__example_55959141808686_1
timestamp 1624855509
transform -1 0 3952 0 1 3332
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808685  sky130_fd_pr__tpl1__example_55959141808685_0
timestamp 1624855509
transform 1 0 26 0 1 115
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808685  sky130_fd_pr__tpl1__example_55959141808685_1
timestamp 1624855509
transform 1 0 3928 0 1 115
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808684  sky130_fd_pr__via_l1m1__example_55959141808684_0
timestamp 1624855509
transform 1 0 3955 0 1 160
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808684  sky130_fd_pr__via_l1m1__example_55959141808684_1
timestamp 1624855509
transform 1 0 53 0 1 160
box 0 0 1 1
use sky130_fd_io__gnd2gnd_diff  sky130_fd_io__gnd2gnd_diff_0
array 0 3 824 0 0 3052
timestamp 1624855509
transform 1 0 632 0 1 220
box 0 0 300 3000
use sky130_fd_io__gnd2gnd_tap  sky130_fd_io__gnd2gnd_tap_0
array 0 4 824 0 0 3052
timestamp 1624855509
transform 1 0 220 0 1 220
box 0 0 300 3000
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 14500020
string GDS_START 14498388
<< end >>
