magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1260 -1286 1626 1652
<< scnmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
<< ndiff >>
rect 0 185 60 336
rect 0 151 8 185
rect 42 151 60 185
rect 0 0 60 151
rect 90 185 168 336
rect 90 151 112 185
rect 146 151 168 185
rect 90 0 168 151
rect 198 185 276 336
rect 198 151 220 185
rect 254 151 276 185
rect 198 0 276 151
rect 306 185 366 336
rect 306 151 324 185
rect 358 151 366 185
rect 306 0 366 151
<< ndiffc >>
rect 8 151 42 185
rect 112 151 146 185
rect 220 151 254 185
rect 324 151 358 185
<< poly >>
rect 60 362 306 392
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
<< locali >>
rect 112 235 358 269
rect 8 185 42 201
rect 8 135 42 151
rect 112 185 146 235
rect 112 135 146 151
rect 220 185 254 201
rect 220 135 254 151
rect 324 185 358 235
rect 324 135 358 151
use contact_11  contact_11_0
timestamp 1624857261
transform 1 0 316 0 1 135
box 0 0 1 1
use contact_11  contact_11_1
timestamp 1624857261
transform 1 0 212 0 1 135
box 0 0 1 1
use contact_11  contact_11_2
timestamp 1624857261
transform 1 0 104 0 1 135
box 0 0 1 1
use contact_11  contact_11_3
timestamp 1624857261
transform 1 0 0 0 1 135
box 0 0 1 1
<< labels >>
rlabel poly s 183 377 183 377 4 G
rlabel locali s 237 168 237 168 4 S
rlabel locali s 25 168 25 168 4 S
rlabel locali s 235 252 235 252 4 D
<< properties >>
string FIXED_BBOX -25 -26 391 392
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 9064806
string GDS_START 9063634
<< end >>
