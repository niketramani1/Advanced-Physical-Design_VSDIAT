magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 18 289 389 323
rect 18 215 125 289
rect 159 215 280 255
rect 323 215 389 289
rect 549 391 607 493
rect 816 391 866 425
rect 549 357 866 391
rect 549 215 643 357
rect 682 289 1087 323
rect 682 215 748 289
rect 792 215 900 255
rect 946 215 1087 289
rect 549 129 615 215
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 30 359 80 527
rect 115 393 165 493
rect 199 427 249 527
rect 367 427 515 527
rect 283 393 333 425
rect 115 357 457 393
rect 423 265 457 357
rect 641 425 698 527
rect 732 459 950 493
rect 732 425 782 459
rect 900 357 950 459
rect 993 359 1034 527
rect 423 199 515 265
rect 423 181 457 199
rect 39 17 73 179
rect 107 95 157 179
rect 191 145 457 181
rect 191 129 257 145
rect 649 147 1042 181
rect 107 61 341 95
rect 375 17 409 111
rect 465 95 515 111
rect 649 95 706 147
rect 808 145 1042 147
rect 465 51 706 95
rect 740 17 774 111
rect 808 51 874 145
rect 908 17 942 111
rect 976 51 1042 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 323 215 389 289 6 A1_N
port 1 nsew signal input
rlabel locali s 18 289 389 323 6 A1_N
port 1 nsew signal input
rlabel locali s 18 215 125 289 6 A1_N
port 1 nsew signal input
rlabel locali s 159 215 280 255 6 A2_N
port 2 nsew signal input
rlabel locali s 946 215 1087 289 6 B1
port 3 nsew signal input
rlabel locali s 682 289 1087 323 6 B1
port 3 nsew signal input
rlabel locali s 682 215 748 289 6 B1
port 3 nsew signal input
rlabel locali s 792 215 900 255 6 B2
port 4 nsew signal input
rlabel locali s 816 391 866 425 6 Y
port 9 nsew signal output
rlabel locali s 549 391 607 493 6 Y
port 9 nsew signal output
rlabel locali s 549 357 866 391 6 Y
port 9 nsew signal output
rlabel locali s 549 215 643 357 6 Y
port 9 nsew signal output
rlabel locali s 549 129 615 215 6 Y
port 9 nsew signal output
rlabel metal1 s 0 -48 1104 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1137096
string GDS_START 1128598
<< end >>
