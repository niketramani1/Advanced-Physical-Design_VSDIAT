magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1302 -1260 1405 1560
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_0
timestamp 1624855509
transform -1 0 -14 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 145 300 145 300 0 FreeSans 300 0 0 0 D
flabel comment s -42 267 -42 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 1886714
string GDS_START 1885730
<< end >>
