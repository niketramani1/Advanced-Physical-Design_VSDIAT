magic
tech sky130A
magscale 1 2
timestamp 1624855514
<< obsli1 >>
rect 0 46 16000 39941
<< metal1 >>
rect 12486 0 12538 261
<< obsm1 >>
rect 0 317 16000 40000
rect 0 52 12430 317
rect 12594 52 16000 317
<< metal2 >>
rect 675 0 721 895
rect 1084 0 1130 895
rect 1226 0 1278 310
rect 2551 0 2603 1070
rect 3262 0 3314 464
rect 4471 0 4523 1285
rect 5320 0 5372 541
rect 5698 0 5750 814
rect 6150 0 6202 453
rect 6363 0 6415 668
rect 7092 0 7144 310
rect 7678 0 7730 618
rect 9049 0 9101 1018
rect 9971 0 10023 109
rect 13367 0 13419 239
rect 13655 0 13785 454
rect 15256 0 15384 411
rect 15522 0 15574 237
rect 15741 0 15781 243
rect 15943 0 15983 35574
<< obsm2 >>
rect 42 35630 15983 40000
rect 42 1341 15887 35630
rect 42 1126 4415 1341
rect 42 951 2495 1126
rect 42 50 619 951
rect 777 50 1028 951
rect 1186 366 2495 951
rect 1334 50 2495 366
rect 2659 520 4415 1126
rect 2659 50 3206 520
rect 3370 50 4415 520
rect 4579 1074 15887 1341
rect 4579 870 8993 1074
rect 4579 597 5642 870
rect 4579 50 5264 597
rect 5428 50 5642 597
rect 5806 724 8993 870
rect 5806 509 6307 724
rect 6471 674 8993 724
rect 5806 50 6094 509
rect 6258 50 6307 509
rect 6471 366 7622 674
rect 6471 50 7036 366
rect 7200 50 7622 366
rect 7786 50 8993 674
rect 9157 510 15887 1074
rect 9157 295 13599 510
rect 13841 467 15887 510
rect 9157 165 13311 295
rect 9157 50 9915 165
rect 10079 50 13311 165
rect 13475 50 13599 295
rect 13841 50 15200 467
rect 15440 299 15887 467
rect 15440 293 15685 299
rect 15440 50 15466 293
rect 15630 50 15685 293
rect 15837 50 15887 299
<< metal3 >>
rect 80 0 204 35697
rect 9173 0 9239 7361
rect 15716 0 15782 36955
rect 15848 0 15914 37912
<< obsm3 >>
rect 80 37992 15914 40000
rect 80 37035 15768 37992
rect 80 35777 15636 37035
rect 284 7441 15636 35777
rect 284 0 9093 7441
rect 9319 0 15636 7441
<< metal4 >>
rect 1714 24211 1960 24248
rect 1962 24241 2500 24250
rect 1714 24002 2500 24211
rect 1503 23971 1714 24002
rect 1743 24001 2500 24002
rect 1503 23791 2500 23971
rect 400 21317 2500 23791
rect 1566 21283 2500 21317
rect 1566 21242 1641 21283
rect 1660 21242 2500 21253
rect 1641 21043 2500 21242
rect 1641 21006 1877 21043
rect 1900 21006 2500 21013
rect 1877 20953 2500 21006
rect 1877 20879 2004 20953
rect 13606 14007 16000 19000
rect 12189 12817 16000 13707
rect 14315 11647 16000 12537
rect 9418 11281 16000 11347
rect 7752 10625 16000 11221
rect 10893 9673 16000 10269
rect 11141 8317 16000 9247
rect 4770 6377 16000 7067
rect 4306 5167 16000 6097
rect 10314 2987 16000 3677
rect 14053 1777 16000 2707
rect 15362 407 16000 1497
<< obsm4 >>
rect 0 24330 16000 40000
rect 0 24328 1882 24330
rect 0 24082 1634 24328
rect 0 23871 1423 24082
rect 0 21237 320 23871
rect 0 21162 1486 21237
rect 0 20926 1561 21162
rect 0 20799 1797 20926
rect 2580 20873 16000 24330
rect 2084 20799 16000 20873
rect 0 19080 16000 20799
rect 0 13927 13526 19080
rect 0 13787 16000 13927
rect 0 12737 12109 13787
rect 0 12617 16000 12737
rect 0 11567 14235 12617
rect 0 11427 16000 11567
rect 0 11301 9338 11427
rect 0 10545 7672 11301
rect 0 10349 16000 10545
rect 0 9593 10813 10349
rect 0 9327 16000 9593
rect 0 8237 11061 9327
rect 0 7147 16000 8237
rect 0 6297 4690 7147
rect 0 6177 16000 6297
rect 0 5087 4226 6177
rect 0 3757 16000 5087
rect 0 2907 10234 3757
rect 0 2787 16000 2907
rect 0 1697 13973 2787
rect 0 1577 16000 1697
rect 0 327 15282 1577
rect 0 107 16000 327
<< metal5 >>
rect 2220 20879 14760 33402
<< obsm5 >>
rect 1960 33722 15040 34697
rect 1960 19617 15040 20559
<< labels >>
rlabel metal4 s 7752 10625 16000 11221 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 10893 9673 16000 10269 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal1 s 12486 0 12538 261 6 ANALOG_EN
port 3 nsew signal input
rlabel metal3 s 9173 0 9239 7361 6 ANALOG_POL
port 4 nsew signal input
rlabel metal2 s 6150 0 6202 453 6 ANALOG_SEL
port 5 nsew signal input
rlabel metal2 s 9971 0 10023 109 6 DM[0]
port 6 nsew signal input
rlabel metal2 s 13367 0 13419 239 6 DM[1]
port 7 nsew signal input
rlabel metal2 s 5698 0 5750 814 6 DM[2]
port 8 nsew signal input
rlabel metal2 s 7092 0 7144 310 6 ENABLE_H
port 9 nsew signal input
rlabel metal2 s 7678 0 7730 618 6 ENABLE_INP_H
port 10 nsew signal input
rlabel metal2 s 2551 0 2603 1070 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel metal3 s 15716 0 15782 36955 6 ENABLE_VDDIO
port 12 nsew signal input
rlabel metal2 s 3262 0 3314 464 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel metal2 s 6363 0 6415 668 6 HLD_H_N
port 14 nsew signal input
rlabel metal2 s 5320 0 5372 541 6 HLD_OVR
port 15 nsew signal input
rlabel metal2 s 1084 0 1130 895 6 IB_MODE_SEL
port 16 nsew signal input
rlabel metal3 s 15848 0 15914 37912 6 IN
port 17 nsew signal output
rlabel metal2 s 9049 0 9101 1018 6 INP_DIS
port 18 nsew signal input
rlabel metal3 s 80 0 204 35697 6 IN_H
port 19 nsew signal output
rlabel metal2 s 675 0 721 895 6 OE_N
port 20 nsew signal input
rlabel metal2 s 4471 0 4523 1285 6 OUT
port 21 nsew signal input
rlabel metal5 s 2220 20879 14760 33402 6 PAD
port 22 nsew signal bidirectional
rlabel metal2 s 15256 0 15384 411 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel metal2 s 13655 0 13785 454 6 PAD_A_ESD_1_H
port 24 nsew signal bidirectional
rlabel metal2 s 13682 21 13684 23 6 PAD_A_ESD_1_H
port 24 nsew signal bidirectional
rlabel metal4 s 400 21317 2500 23791 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1503 23791 1714 24002 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1533 23791 2500 23821 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1563 23821 2500 23851 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1566 21242 1641 21317 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1570 21313 2500 21317 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1593 23851 2500 23881 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1600 21283 2500 21313 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1623 23881 2500 23911 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1641 21006 1877 21242 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1653 23911 2500 23941 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1660 21223 2500 21253 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1683 23941 2500 23971 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1690 21193 2500 21223 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1714 24002 1960 24248 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1720 21163 2500 21193 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1743 24001 2500 24031 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1750 21133 2500 21163 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1773 24031 2500 24061 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1780 21103 2500 21133 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1803 24061 2500 24091 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1810 21073 2500 21103 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1833 24091 2500 24121 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1840 21043 2500 21073 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1863 24121 2500 24151 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1877 20879 2004 21006 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1893 24151 2500 24181 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1900 20983 2500 21013 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1923 24181 2500 24211 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1930 20953 2500 20983 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal4 s 1962 24241 2500 24250 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel metal2 s 15522 0 15574 237 6 SLOW
port 26 nsew signal input
rlabel metal2 s 15741 0 15781 243 6 TIE_HI_ESD
port 27 nsew signal output
rlabel metal2 s 15760 21 15762 23 6 TIE_HI_ESD
port 27 nsew signal output
rlabel metal2 s 15943 0 15983 35574 6 TIE_LO_ESD
port 28 nsew signal output
rlabel metal2 s 1226 0 1278 310 6 VTRIP_SEL
port 29 nsew signal input
rlabel metal4 s 14053 1777 16000 2707 6 VCCD
port 30 nsew power bidirectional
rlabel metal4 s 15362 407 16000 1497 6 VCCHIB
port 31 nsew power bidirectional
rlabel metal4 s 10314 2987 16000 3677 6 VDDA
port 32 nsew power bidirectional
rlabel metal4 s 13606 14007 16000 19000 6 VDDIO
port 33 nsew power bidirectional
rlabel metal4 s 12189 12817 16000 13707 6 VDDIO_Q
port 34 nsew power bidirectional
rlabel metal4 s 9418 11281 16000 11347 6 VSSA
port 35 nsew ground bidirectional
rlabel metal4 s 11141 8317 16000 9247 6 VSSD
port 36 nsew ground bidirectional
rlabel metal4 s 4306 5167 16000 6097 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 14315 11647 16000 12537 6 VSSIO_Q
port 38 nsew ground bidirectional
rlabel metal4 s 4770 6377 16000 7067 6 VSWITCH
port 39 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 16000 40000
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 8058748
string GDS_START 6287582
<< end >>
