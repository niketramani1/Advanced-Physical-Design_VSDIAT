magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1310 -3204 4201 1261
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_1
timestamp 1624855509
transform 1 0 2940 0 1 -1944
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_0
timestamp 1624855509
transform 1 0 -50 0 1 0
box 0 0 1 1
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 14463290
string GDS_START 14459626
<< end >>
