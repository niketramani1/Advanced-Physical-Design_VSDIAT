magic
tech sky130A
magscale 1 2
timestamp 1624855514
<< obsm3 >>
rect 100 4768 14940 39600
<< metal4 >>
rect 111 39529 175 39593
rect 191 39529 255 39593
rect 271 39529 335 39593
rect 351 39529 415 39593
rect 431 39529 495 39593
rect 511 39529 575 39593
rect 591 39529 655 39593
rect 671 39529 735 39593
rect 751 39529 815 39593
rect 831 39529 895 39593
rect 911 39529 975 39593
rect 991 39529 1055 39593
rect 1071 39529 1135 39593
rect 1151 39529 1215 39593
rect 1231 39529 1295 39593
rect 1311 39529 1375 39593
rect 1391 39529 1455 39593
rect 1471 39529 1535 39593
rect 1551 39529 1615 39593
rect 1631 39529 1695 39593
rect 1711 39529 1775 39593
rect 1791 39529 1855 39593
rect 1871 39529 1935 39593
rect 1951 39529 2015 39593
rect 2031 39529 2095 39593
rect 2111 39529 2175 39593
rect 2191 39529 2255 39593
rect 2271 39529 2335 39593
rect 2351 39529 2415 39593
rect 2431 39529 2495 39593
rect 2511 39529 2575 39593
rect 12416 39529 12480 39593
rect 12498 39529 12562 39593
rect 12580 39529 12644 39593
rect 12662 39529 12726 39593
rect 12744 39529 12808 39593
rect 12826 39529 12890 39593
rect 12908 39529 12972 39593
rect 12990 39529 13054 39593
rect 13072 39529 13136 39593
rect 13154 39529 13218 39593
rect 13236 39529 13300 39593
rect 13318 39529 13382 39593
rect 13400 39529 13464 39593
rect 13482 39529 13546 39593
rect 13564 39529 13628 39593
rect 13646 39529 13710 39593
rect 13728 39529 13792 39593
rect 13810 39529 13874 39593
rect 13892 39529 13956 39593
rect 13974 39529 14038 39593
rect 14056 39529 14120 39593
rect 14138 39529 14202 39593
rect 14220 39529 14284 39593
rect 14302 39529 14366 39593
rect 14384 39529 14448 39593
rect 14466 39529 14530 39593
rect 14548 39529 14612 39593
rect 14630 39529 14694 39593
rect 14712 39529 14776 39593
rect 14794 39529 14858 39593
rect 14876 39529 14940 39593
rect 111 39448 175 39512
rect 191 39448 255 39512
rect 271 39448 335 39512
rect 351 39448 415 39512
rect 431 39448 495 39512
rect 511 39448 575 39512
rect 591 39448 655 39512
rect 671 39448 735 39512
rect 751 39448 815 39512
rect 831 39448 895 39512
rect 911 39448 975 39512
rect 991 39448 1055 39512
rect 1071 39448 1135 39512
rect 1151 39448 1215 39512
rect 1231 39448 1295 39512
rect 1311 39448 1375 39512
rect 1391 39448 1455 39512
rect 1471 39448 1535 39512
rect 1551 39448 1615 39512
rect 1631 39448 1695 39512
rect 1711 39448 1775 39512
rect 1791 39448 1855 39512
rect 1871 39448 1935 39512
rect 1951 39448 2015 39512
rect 2031 39448 2095 39512
rect 2111 39448 2175 39512
rect 2191 39448 2255 39512
rect 2271 39448 2335 39512
rect 2351 39448 2415 39512
rect 2431 39448 2495 39512
rect 2511 39448 2575 39512
rect 12416 39448 12480 39512
rect 12498 39448 12562 39512
rect 12580 39448 12644 39512
rect 12662 39448 12726 39512
rect 12744 39448 12808 39512
rect 12826 39448 12890 39512
rect 12908 39448 12972 39512
rect 12990 39448 13054 39512
rect 13072 39448 13136 39512
rect 13154 39448 13218 39512
rect 13236 39448 13300 39512
rect 13318 39448 13382 39512
rect 13400 39448 13464 39512
rect 13482 39448 13546 39512
rect 13564 39448 13628 39512
rect 13646 39448 13710 39512
rect 13728 39448 13792 39512
rect 13810 39448 13874 39512
rect 13892 39448 13956 39512
rect 13974 39448 14038 39512
rect 14056 39448 14120 39512
rect 14138 39448 14202 39512
rect 14220 39448 14284 39512
rect 14302 39448 14366 39512
rect 14384 39448 14448 39512
rect 14466 39448 14530 39512
rect 14548 39448 14612 39512
rect 14630 39448 14694 39512
rect 14712 39448 14776 39512
rect 14794 39448 14858 39512
rect 14876 39448 14940 39512
rect 111 39367 175 39431
rect 191 39367 255 39431
rect 271 39367 335 39431
rect 351 39367 415 39431
rect 431 39367 495 39431
rect 511 39367 575 39431
rect 591 39367 655 39431
rect 671 39367 735 39431
rect 751 39367 815 39431
rect 831 39367 895 39431
rect 911 39367 975 39431
rect 991 39367 1055 39431
rect 1071 39367 1135 39431
rect 1151 39367 1215 39431
rect 1231 39367 1295 39431
rect 1311 39367 1375 39431
rect 1391 39367 1455 39431
rect 1471 39367 1535 39431
rect 1551 39367 1615 39431
rect 1631 39367 1695 39431
rect 1711 39367 1775 39431
rect 1791 39367 1855 39431
rect 1871 39367 1935 39431
rect 1951 39367 2015 39431
rect 2031 39367 2095 39431
rect 2111 39367 2175 39431
rect 2191 39367 2255 39431
rect 2271 39367 2335 39431
rect 2351 39367 2415 39431
rect 2431 39367 2495 39431
rect 2511 39367 2575 39431
rect 12416 39367 12480 39431
rect 12498 39367 12562 39431
rect 12580 39367 12644 39431
rect 12662 39367 12726 39431
rect 12744 39367 12808 39431
rect 12826 39367 12890 39431
rect 12908 39367 12972 39431
rect 12990 39367 13054 39431
rect 13072 39367 13136 39431
rect 13154 39367 13218 39431
rect 13236 39367 13300 39431
rect 13318 39367 13382 39431
rect 13400 39367 13464 39431
rect 13482 39367 13546 39431
rect 13564 39367 13628 39431
rect 13646 39367 13710 39431
rect 13728 39367 13792 39431
rect 13810 39367 13874 39431
rect 13892 39367 13956 39431
rect 13974 39367 14038 39431
rect 14056 39367 14120 39431
rect 14138 39367 14202 39431
rect 14220 39367 14284 39431
rect 14302 39367 14366 39431
rect 14384 39367 14448 39431
rect 14466 39367 14530 39431
rect 14548 39367 14612 39431
rect 14630 39367 14694 39431
rect 14712 39367 14776 39431
rect 14794 39367 14858 39431
rect 14876 39367 14940 39431
rect 111 39286 175 39350
rect 191 39286 255 39350
rect 271 39286 335 39350
rect 351 39286 415 39350
rect 431 39286 495 39350
rect 511 39286 575 39350
rect 591 39286 655 39350
rect 671 39286 735 39350
rect 751 39286 815 39350
rect 831 39286 895 39350
rect 911 39286 975 39350
rect 991 39286 1055 39350
rect 1071 39286 1135 39350
rect 1151 39286 1215 39350
rect 1231 39286 1295 39350
rect 1311 39286 1375 39350
rect 1391 39286 1455 39350
rect 1471 39286 1535 39350
rect 1551 39286 1615 39350
rect 1631 39286 1695 39350
rect 1711 39286 1775 39350
rect 1791 39286 1855 39350
rect 1871 39286 1935 39350
rect 1951 39286 2015 39350
rect 2031 39286 2095 39350
rect 2111 39286 2175 39350
rect 2191 39286 2255 39350
rect 2271 39286 2335 39350
rect 2351 39286 2415 39350
rect 2431 39286 2495 39350
rect 2511 39286 2575 39350
rect 12416 39286 12480 39350
rect 12498 39286 12562 39350
rect 12580 39286 12644 39350
rect 12662 39286 12726 39350
rect 12744 39286 12808 39350
rect 12826 39286 12890 39350
rect 12908 39286 12972 39350
rect 12990 39286 13054 39350
rect 13072 39286 13136 39350
rect 13154 39286 13218 39350
rect 13236 39286 13300 39350
rect 13318 39286 13382 39350
rect 13400 39286 13464 39350
rect 13482 39286 13546 39350
rect 13564 39286 13628 39350
rect 13646 39286 13710 39350
rect 13728 39286 13792 39350
rect 13810 39286 13874 39350
rect 13892 39286 13956 39350
rect 13974 39286 14038 39350
rect 14056 39286 14120 39350
rect 14138 39286 14202 39350
rect 14220 39286 14284 39350
rect 14302 39286 14366 39350
rect 14384 39286 14448 39350
rect 14466 39286 14530 39350
rect 14548 39286 14612 39350
rect 14630 39286 14694 39350
rect 14712 39286 14776 39350
rect 14794 39286 14858 39350
rect 14876 39286 14940 39350
rect 111 39205 175 39269
rect 191 39205 255 39269
rect 271 39205 335 39269
rect 351 39205 415 39269
rect 431 39205 495 39269
rect 511 39205 575 39269
rect 591 39205 655 39269
rect 671 39205 735 39269
rect 751 39205 815 39269
rect 831 39205 895 39269
rect 911 39205 975 39269
rect 991 39205 1055 39269
rect 1071 39205 1135 39269
rect 1151 39205 1215 39269
rect 1231 39205 1295 39269
rect 1311 39205 1375 39269
rect 1391 39205 1455 39269
rect 1471 39205 1535 39269
rect 1551 39205 1615 39269
rect 1631 39205 1695 39269
rect 1711 39205 1775 39269
rect 1791 39205 1855 39269
rect 1871 39205 1935 39269
rect 1951 39205 2015 39269
rect 2031 39205 2095 39269
rect 2111 39205 2175 39269
rect 2191 39205 2255 39269
rect 2271 39205 2335 39269
rect 2351 39205 2415 39269
rect 2431 39205 2495 39269
rect 2511 39205 2575 39269
rect 12416 39205 12480 39269
rect 12498 39205 12562 39269
rect 12580 39205 12644 39269
rect 12662 39205 12726 39269
rect 12744 39205 12808 39269
rect 12826 39205 12890 39269
rect 12908 39205 12972 39269
rect 12990 39205 13054 39269
rect 13072 39205 13136 39269
rect 13154 39205 13218 39269
rect 13236 39205 13300 39269
rect 13318 39205 13382 39269
rect 13400 39205 13464 39269
rect 13482 39205 13546 39269
rect 13564 39205 13628 39269
rect 13646 39205 13710 39269
rect 13728 39205 13792 39269
rect 13810 39205 13874 39269
rect 13892 39205 13956 39269
rect 13974 39205 14038 39269
rect 14056 39205 14120 39269
rect 14138 39205 14202 39269
rect 14220 39205 14284 39269
rect 14302 39205 14366 39269
rect 14384 39205 14448 39269
rect 14466 39205 14530 39269
rect 14548 39205 14612 39269
rect 14630 39205 14694 39269
rect 14712 39205 14776 39269
rect 14794 39205 14858 39269
rect 14876 39205 14940 39269
rect 111 39124 175 39188
rect 191 39124 255 39188
rect 271 39124 335 39188
rect 351 39124 415 39188
rect 431 39124 495 39188
rect 511 39124 575 39188
rect 591 39124 655 39188
rect 671 39124 735 39188
rect 751 39124 815 39188
rect 831 39124 895 39188
rect 911 39124 975 39188
rect 991 39124 1055 39188
rect 1071 39124 1135 39188
rect 1151 39124 1215 39188
rect 1231 39124 1295 39188
rect 1311 39124 1375 39188
rect 1391 39124 1455 39188
rect 1471 39124 1535 39188
rect 1551 39124 1615 39188
rect 1631 39124 1695 39188
rect 1711 39124 1775 39188
rect 1791 39124 1855 39188
rect 1871 39124 1935 39188
rect 1951 39124 2015 39188
rect 2031 39124 2095 39188
rect 2111 39124 2175 39188
rect 2191 39124 2255 39188
rect 2271 39124 2335 39188
rect 2351 39124 2415 39188
rect 2431 39124 2495 39188
rect 2511 39124 2575 39188
rect 12416 39124 12480 39188
rect 12498 39124 12562 39188
rect 12580 39124 12644 39188
rect 12662 39124 12726 39188
rect 12744 39124 12808 39188
rect 12826 39124 12890 39188
rect 12908 39124 12972 39188
rect 12990 39124 13054 39188
rect 13072 39124 13136 39188
rect 13154 39124 13218 39188
rect 13236 39124 13300 39188
rect 13318 39124 13382 39188
rect 13400 39124 13464 39188
rect 13482 39124 13546 39188
rect 13564 39124 13628 39188
rect 13646 39124 13710 39188
rect 13728 39124 13792 39188
rect 13810 39124 13874 39188
rect 13892 39124 13956 39188
rect 13974 39124 14038 39188
rect 14056 39124 14120 39188
rect 14138 39124 14202 39188
rect 14220 39124 14284 39188
rect 14302 39124 14366 39188
rect 14384 39124 14448 39188
rect 14466 39124 14530 39188
rect 14548 39124 14612 39188
rect 14630 39124 14694 39188
rect 14712 39124 14776 39188
rect 14794 39124 14858 39188
rect 14876 39124 14940 39188
rect 111 39043 175 39107
rect 191 39043 255 39107
rect 271 39043 335 39107
rect 351 39043 415 39107
rect 431 39043 495 39107
rect 511 39043 575 39107
rect 591 39043 655 39107
rect 671 39043 735 39107
rect 751 39043 815 39107
rect 831 39043 895 39107
rect 911 39043 975 39107
rect 991 39043 1055 39107
rect 1071 39043 1135 39107
rect 1151 39043 1215 39107
rect 1231 39043 1295 39107
rect 1311 39043 1375 39107
rect 1391 39043 1455 39107
rect 1471 39043 1535 39107
rect 1551 39043 1615 39107
rect 1631 39043 1695 39107
rect 1711 39043 1775 39107
rect 1791 39043 1855 39107
rect 1871 39043 1935 39107
rect 1951 39043 2015 39107
rect 2031 39043 2095 39107
rect 2111 39043 2175 39107
rect 2191 39043 2255 39107
rect 2271 39043 2335 39107
rect 2351 39043 2415 39107
rect 2431 39043 2495 39107
rect 2511 39043 2575 39107
rect 12416 39043 12480 39107
rect 12498 39043 12562 39107
rect 12580 39043 12644 39107
rect 12662 39043 12726 39107
rect 12744 39043 12808 39107
rect 12826 39043 12890 39107
rect 12908 39043 12972 39107
rect 12990 39043 13054 39107
rect 13072 39043 13136 39107
rect 13154 39043 13218 39107
rect 13236 39043 13300 39107
rect 13318 39043 13382 39107
rect 13400 39043 13464 39107
rect 13482 39043 13546 39107
rect 13564 39043 13628 39107
rect 13646 39043 13710 39107
rect 13728 39043 13792 39107
rect 13810 39043 13874 39107
rect 13892 39043 13956 39107
rect 13974 39043 14038 39107
rect 14056 39043 14120 39107
rect 14138 39043 14202 39107
rect 14220 39043 14284 39107
rect 14302 39043 14366 39107
rect 14384 39043 14448 39107
rect 14466 39043 14530 39107
rect 14548 39043 14612 39107
rect 14630 39043 14694 39107
rect 14712 39043 14776 39107
rect 14794 39043 14858 39107
rect 14876 39043 14940 39107
rect 111 38962 175 39026
rect 191 38962 255 39026
rect 271 38962 335 39026
rect 351 38962 415 39026
rect 431 38962 495 39026
rect 511 38962 575 39026
rect 591 38962 655 39026
rect 671 38962 735 39026
rect 751 38962 815 39026
rect 831 38962 895 39026
rect 911 38962 975 39026
rect 991 38962 1055 39026
rect 1071 38962 1135 39026
rect 1151 38962 1215 39026
rect 1231 38962 1295 39026
rect 1311 38962 1375 39026
rect 1391 38962 1455 39026
rect 1471 38962 1535 39026
rect 1551 38962 1615 39026
rect 1631 38962 1695 39026
rect 1711 38962 1775 39026
rect 1791 38962 1855 39026
rect 1871 38962 1935 39026
rect 1951 38962 2015 39026
rect 2031 38962 2095 39026
rect 2111 38962 2175 39026
rect 2191 38962 2255 39026
rect 2271 38962 2335 39026
rect 2351 38962 2415 39026
rect 2431 38962 2495 39026
rect 2511 38962 2575 39026
rect 12416 38962 12480 39026
rect 12498 38962 12562 39026
rect 12580 38962 12644 39026
rect 12662 38962 12726 39026
rect 12744 38962 12808 39026
rect 12826 38962 12890 39026
rect 12908 38962 12972 39026
rect 12990 38962 13054 39026
rect 13072 38962 13136 39026
rect 13154 38962 13218 39026
rect 13236 38962 13300 39026
rect 13318 38962 13382 39026
rect 13400 38962 13464 39026
rect 13482 38962 13546 39026
rect 13564 38962 13628 39026
rect 13646 38962 13710 39026
rect 13728 38962 13792 39026
rect 13810 38962 13874 39026
rect 13892 38962 13956 39026
rect 13974 38962 14038 39026
rect 14056 38962 14120 39026
rect 14138 38962 14202 39026
rect 14220 38962 14284 39026
rect 14302 38962 14366 39026
rect 14384 38962 14448 39026
rect 14466 38962 14530 39026
rect 14548 38962 14612 39026
rect 14630 38962 14694 39026
rect 14712 38962 14776 39026
rect 14794 38962 14858 39026
rect 14876 38962 14940 39026
rect 111 38881 175 38945
rect 191 38881 255 38945
rect 271 38881 335 38945
rect 351 38881 415 38945
rect 431 38881 495 38945
rect 511 38881 575 38945
rect 591 38881 655 38945
rect 671 38881 735 38945
rect 751 38881 815 38945
rect 831 38881 895 38945
rect 911 38881 975 38945
rect 991 38881 1055 38945
rect 1071 38881 1135 38945
rect 1151 38881 1215 38945
rect 1231 38881 1295 38945
rect 1311 38881 1375 38945
rect 1391 38881 1455 38945
rect 1471 38881 1535 38945
rect 1551 38881 1615 38945
rect 1631 38881 1695 38945
rect 1711 38881 1775 38945
rect 1791 38881 1855 38945
rect 1871 38881 1935 38945
rect 1951 38881 2015 38945
rect 2031 38881 2095 38945
rect 2111 38881 2175 38945
rect 2191 38881 2255 38945
rect 2271 38881 2335 38945
rect 2351 38881 2415 38945
rect 2431 38881 2495 38945
rect 2511 38881 2575 38945
rect 12416 38881 12480 38945
rect 12498 38881 12562 38945
rect 12580 38881 12644 38945
rect 12662 38881 12726 38945
rect 12744 38881 12808 38945
rect 12826 38881 12890 38945
rect 12908 38881 12972 38945
rect 12990 38881 13054 38945
rect 13072 38881 13136 38945
rect 13154 38881 13218 38945
rect 13236 38881 13300 38945
rect 13318 38881 13382 38945
rect 13400 38881 13464 38945
rect 13482 38881 13546 38945
rect 13564 38881 13628 38945
rect 13646 38881 13710 38945
rect 13728 38881 13792 38945
rect 13810 38881 13874 38945
rect 13892 38881 13956 38945
rect 13974 38881 14038 38945
rect 14056 38881 14120 38945
rect 14138 38881 14202 38945
rect 14220 38881 14284 38945
rect 14302 38881 14366 38945
rect 14384 38881 14448 38945
rect 14466 38881 14530 38945
rect 14548 38881 14612 38945
rect 14630 38881 14694 38945
rect 14712 38881 14776 38945
rect 14794 38881 14858 38945
rect 14876 38881 14940 38945
rect 111 38800 175 38864
rect 191 38800 255 38864
rect 271 38800 335 38864
rect 351 38800 415 38864
rect 431 38800 495 38864
rect 511 38800 575 38864
rect 591 38800 655 38864
rect 671 38800 735 38864
rect 751 38800 815 38864
rect 831 38800 895 38864
rect 911 38800 975 38864
rect 991 38800 1055 38864
rect 1071 38800 1135 38864
rect 1151 38800 1215 38864
rect 1231 38800 1295 38864
rect 1311 38800 1375 38864
rect 1391 38800 1455 38864
rect 1471 38800 1535 38864
rect 1551 38800 1615 38864
rect 1631 38800 1695 38864
rect 1711 38800 1775 38864
rect 1791 38800 1855 38864
rect 1871 38800 1935 38864
rect 1951 38800 2015 38864
rect 2031 38800 2095 38864
rect 2111 38800 2175 38864
rect 2191 38800 2255 38864
rect 2271 38800 2335 38864
rect 2351 38800 2415 38864
rect 2431 38800 2495 38864
rect 2511 38800 2575 38864
rect 12416 38800 12480 38864
rect 12498 38800 12562 38864
rect 12580 38800 12644 38864
rect 12662 38800 12726 38864
rect 12744 38800 12808 38864
rect 12826 38800 12890 38864
rect 12908 38800 12972 38864
rect 12990 38800 13054 38864
rect 13072 38800 13136 38864
rect 13154 38800 13218 38864
rect 13236 38800 13300 38864
rect 13318 38800 13382 38864
rect 13400 38800 13464 38864
rect 13482 38800 13546 38864
rect 13564 38800 13628 38864
rect 13646 38800 13710 38864
rect 13728 38800 13792 38864
rect 13810 38800 13874 38864
rect 13892 38800 13956 38864
rect 13974 38800 14038 38864
rect 14056 38800 14120 38864
rect 14138 38800 14202 38864
rect 14220 38800 14284 38864
rect 14302 38800 14366 38864
rect 14384 38800 14448 38864
rect 14466 38800 14530 38864
rect 14548 38800 14612 38864
rect 14630 38800 14694 38864
rect 14712 38800 14776 38864
rect 14794 38800 14858 38864
rect 14876 38800 14940 38864
rect 111 38719 175 38783
rect 191 38719 255 38783
rect 271 38719 335 38783
rect 351 38719 415 38783
rect 431 38719 495 38783
rect 511 38719 575 38783
rect 591 38719 655 38783
rect 671 38719 735 38783
rect 751 38719 815 38783
rect 831 38719 895 38783
rect 911 38719 975 38783
rect 991 38719 1055 38783
rect 1071 38719 1135 38783
rect 1151 38719 1215 38783
rect 1231 38719 1295 38783
rect 1311 38719 1375 38783
rect 1391 38719 1455 38783
rect 1471 38719 1535 38783
rect 1551 38719 1615 38783
rect 1631 38719 1695 38783
rect 1711 38719 1775 38783
rect 1791 38719 1855 38783
rect 1871 38719 1935 38783
rect 1951 38719 2015 38783
rect 2031 38719 2095 38783
rect 2111 38719 2175 38783
rect 2191 38719 2255 38783
rect 2271 38719 2335 38783
rect 2351 38719 2415 38783
rect 2431 38719 2495 38783
rect 2511 38719 2575 38783
rect 12416 38719 12480 38783
rect 12498 38719 12562 38783
rect 12580 38719 12644 38783
rect 12662 38719 12726 38783
rect 12744 38719 12808 38783
rect 12826 38719 12890 38783
rect 12908 38719 12972 38783
rect 12990 38719 13054 38783
rect 13072 38719 13136 38783
rect 13154 38719 13218 38783
rect 13236 38719 13300 38783
rect 13318 38719 13382 38783
rect 13400 38719 13464 38783
rect 13482 38719 13546 38783
rect 13564 38719 13628 38783
rect 13646 38719 13710 38783
rect 13728 38719 13792 38783
rect 13810 38719 13874 38783
rect 13892 38719 13956 38783
rect 13974 38719 14038 38783
rect 14056 38719 14120 38783
rect 14138 38719 14202 38783
rect 14220 38719 14284 38783
rect 14302 38719 14366 38783
rect 14384 38719 14448 38783
rect 14466 38719 14530 38783
rect 14548 38719 14612 38783
rect 14630 38719 14694 38783
rect 14712 38719 14776 38783
rect 14794 38719 14858 38783
rect 14876 38719 14940 38783
rect 111 38638 175 38702
rect 191 38638 255 38702
rect 271 38638 335 38702
rect 351 38638 415 38702
rect 431 38638 495 38702
rect 511 38638 575 38702
rect 591 38638 655 38702
rect 671 38638 735 38702
rect 751 38638 815 38702
rect 831 38638 895 38702
rect 911 38638 975 38702
rect 991 38638 1055 38702
rect 1071 38638 1135 38702
rect 1151 38638 1215 38702
rect 1231 38638 1295 38702
rect 1311 38638 1375 38702
rect 1391 38638 1455 38702
rect 1471 38638 1535 38702
rect 1551 38638 1615 38702
rect 1631 38638 1695 38702
rect 1711 38638 1775 38702
rect 1791 38638 1855 38702
rect 1871 38638 1935 38702
rect 1951 38638 2015 38702
rect 2031 38638 2095 38702
rect 2111 38638 2175 38702
rect 2191 38638 2255 38702
rect 2271 38638 2335 38702
rect 2351 38638 2415 38702
rect 2431 38638 2495 38702
rect 2511 38638 2575 38702
rect 12416 38638 12480 38702
rect 12498 38638 12562 38702
rect 12580 38638 12644 38702
rect 12662 38638 12726 38702
rect 12744 38638 12808 38702
rect 12826 38638 12890 38702
rect 12908 38638 12972 38702
rect 12990 38638 13054 38702
rect 13072 38638 13136 38702
rect 13154 38638 13218 38702
rect 13236 38638 13300 38702
rect 13318 38638 13382 38702
rect 13400 38638 13464 38702
rect 13482 38638 13546 38702
rect 13564 38638 13628 38702
rect 13646 38638 13710 38702
rect 13728 38638 13792 38702
rect 13810 38638 13874 38702
rect 13892 38638 13956 38702
rect 13974 38638 14038 38702
rect 14056 38638 14120 38702
rect 14138 38638 14202 38702
rect 14220 38638 14284 38702
rect 14302 38638 14366 38702
rect 14384 38638 14448 38702
rect 14466 38638 14530 38702
rect 14548 38638 14612 38702
rect 14630 38638 14694 38702
rect 14712 38638 14776 38702
rect 14794 38638 14858 38702
rect 14876 38638 14940 38702
rect 111 38557 175 38621
rect 191 38557 255 38621
rect 271 38557 335 38621
rect 351 38557 415 38621
rect 431 38557 495 38621
rect 511 38557 575 38621
rect 591 38557 655 38621
rect 671 38557 735 38621
rect 751 38557 815 38621
rect 831 38557 895 38621
rect 911 38557 975 38621
rect 991 38557 1055 38621
rect 1071 38557 1135 38621
rect 1151 38557 1215 38621
rect 1231 38557 1295 38621
rect 1311 38557 1375 38621
rect 1391 38557 1455 38621
rect 1471 38557 1535 38621
rect 1551 38557 1615 38621
rect 1631 38557 1695 38621
rect 1711 38557 1775 38621
rect 1791 38557 1855 38621
rect 1871 38557 1935 38621
rect 1951 38557 2015 38621
rect 2031 38557 2095 38621
rect 2111 38557 2175 38621
rect 2191 38557 2255 38621
rect 2271 38557 2335 38621
rect 2351 38557 2415 38621
rect 2431 38557 2495 38621
rect 2511 38557 2575 38621
rect 12416 38557 12480 38621
rect 12498 38557 12562 38621
rect 12580 38557 12644 38621
rect 12662 38557 12726 38621
rect 12744 38557 12808 38621
rect 12826 38557 12890 38621
rect 12908 38557 12972 38621
rect 12990 38557 13054 38621
rect 13072 38557 13136 38621
rect 13154 38557 13218 38621
rect 13236 38557 13300 38621
rect 13318 38557 13382 38621
rect 13400 38557 13464 38621
rect 13482 38557 13546 38621
rect 13564 38557 13628 38621
rect 13646 38557 13710 38621
rect 13728 38557 13792 38621
rect 13810 38557 13874 38621
rect 13892 38557 13956 38621
rect 13974 38557 14038 38621
rect 14056 38557 14120 38621
rect 14138 38557 14202 38621
rect 14220 38557 14284 38621
rect 14302 38557 14366 38621
rect 14384 38557 14448 38621
rect 14466 38557 14530 38621
rect 14548 38557 14612 38621
rect 14630 38557 14694 38621
rect 14712 38557 14776 38621
rect 14794 38557 14858 38621
rect 14876 38557 14940 38621
rect 111 38476 175 38540
rect 191 38476 255 38540
rect 271 38476 335 38540
rect 351 38476 415 38540
rect 431 38476 495 38540
rect 511 38476 575 38540
rect 591 38476 655 38540
rect 671 38476 735 38540
rect 751 38476 815 38540
rect 831 38476 895 38540
rect 911 38476 975 38540
rect 991 38476 1055 38540
rect 1071 38476 1135 38540
rect 1151 38476 1215 38540
rect 1231 38476 1295 38540
rect 1311 38476 1375 38540
rect 1391 38476 1455 38540
rect 1471 38476 1535 38540
rect 1551 38476 1615 38540
rect 1631 38476 1695 38540
rect 1711 38476 1775 38540
rect 1791 38476 1855 38540
rect 1871 38476 1935 38540
rect 1951 38476 2015 38540
rect 2031 38476 2095 38540
rect 2111 38476 2175 38540
rect 2191 38476 2255 38540
rect 2271 38476 2335 38540
rect 2351 38476 2415 38540
rect 2431 38476 2495 38540
rect 2511 38476 2575 38540
rect 12416 38476 12480 38540
rect 12498 38476 12562 38540
rect 12580 38476 12644 38540
rect 12662 38476 12726 38540
rect 12744 38476 12808 38540
rect 12826 38476 12890 38540
rect 12908 38476 12972 38540
rect 12990 38476 13054 38540
rect 13072 38476 13136 38540
rect 13154 38476 13218 38540
rect 13236 38476 13300 38540
rect 13318 38476 13382 38540
rect 13400 38476 13464 38540
rect 13482 38476 13546 38540
rect 13564 38476 13628 38540
rect 13646 38476 13710 38540
rect 13728 38476 13792 38540
rect 13810 38476 13874 38540
rect 13892 38476 13956 38540
rect 13974 38476 14038 38540
rect 14056 38476 14120 38540
rect 14138 38476 14202 38540
rect 14220 38476 14284 38540
rect 14302 38476 14366 38540
rect 14384 38476 14448 38540
rect 14466 38476 14530 38540
rect 14548 38476 14612 38540
rect 14630 38476 14694 38540
rect 14712 38476 14776 38540
rect 14794 38476 14858 38540
rect 14876 38476 14940 38540
rect 111 38395 175 38459
rect 191 38395 255 38459
rect 271 38395 335 38459
rect 351 38395 415 38459
rect 431 38395 495 38459
rect 511 38395 575 38459
rect 591 38395 655 38459
rect 671 38395 735 38459
rect 751 38395 815 38459
rect 831 38395 895 38459
rect 911 38395 975 38459
rect 991 38395 1055 38459
rect 1071 38395 1135 38459
rect 1151 38395 1215 38459
rect 1231 38395 1295 38459
rect 1311 38395 1375 38459
rect 1391 38395 1455 38459
rect 1471 38395 1535 38459
rect 1551 38395 1615 38459
rect 1631 38395 1695 38459
rect 1711 38395 1775 38459
rect 1791 38395 1855 38459
rect 1871 38395 1935 38459
rect 1951 38395 2015 38459
rect 2031 38395 2095 38459
rect 2111 38395 2175 38459
rect 2191 38395 2255 38459
rect 2271 38395 2335 38459
rect 2351 38395 2415 38459
rect 2431 38395 2495 38459
rect 2511 38395 2575 38459
rect 12416 38395 12480 38459
rect 12498 38395 12562 38459
rect 12580 38395 12644 38459
rect 12662 38395 12726 38459
rect 12744 38395 12808 38459
rect 12826 38395 12890 38459
rect 12908 38395 12972 38459
rect 12990 38395 13054 38459
rect 13072 38395 13136 38459
rect 13154 38395 13218 38459
rect 13236 38395 13300 38459
rect 13318 38395 13382 38459
rect 13400 38395 13464 38459
rect 13482 38395 13546 38459
rect 13564 38395 13628 38459
rect 13646 38395 13710 38459
rect 13728 38395 13792 38459
rect 13810 38395 13874 38459
rect 13892 38395 13956 38459
rect 13974 38395 14038 38459
rect 14056 38395 14120 38459
rect 14138 38395 14202 38459
rect 14220 38395 14284 38459
rect 14302 38395 14366 38459
rect 14384 38395 14448 38459
rect 14466 38395 14530 38459
rect 14548 38395 14612 38459
rect 14630 38395 14694 38459
rect 14712 38395 14776 38459
rect 14794 38395 14858 38459
rect 14876 38395 14940 38459
rect 111 38314 175 38378
rect 191 38314 255 38378
rect 271 38314 335 38378
rect 351 38314 415 38378
rect 431 38314 495 38378
rect 511 38314 575 38378
rect 591 38314 655 38378
rect 671 38314 735 38378
rect 751 38314 815 38378
rect 831 38314 895 38378
rect 911 38314 975 38378
rect 991 38314 1055 38378
rect 1071 38314 1135 38378
rect 1151 38314 1215 38378
rect 1231 38314 1295 38378
rect 1311 38314 1375 38378
rect 1391 38314 1455 38378
rect 1471 38314 1535 38378
rect 1551 38314 1615 38378
rect 1631 38314 1695 38378
rect 1711 38314 1775 38378
rect 1791 38314 1855 38378
rect 1871 38314 1935 38378
rect 1951 38314 2015 38378
rect 2031 38314 2095 38378
rect 2111 38314 2175 38378
rect 2191 38314 2255 38378
rect 2271 38314 2335 38378
rect 2351 38314 2415 38378
rect 2431 38314 2495 38378
rect 2511 38314 2575 38378
rect 12416 38314 12480 38378
rect 12498 38314 12562 38378
rect 12580 38314 12644 38378
rect 12662 38314 12726 38378
rect 12744 38314 12808 38378
rect 12826 38314 12890 38378
rect 12908 38314 12972 38378
rect 12990 38314 13054 38378
rect 13072 38314 13136 38378
rect 13154 38314 13218 38378
rect 13236 38314 13300 38378
rect 13318 38314 13382 38378
rect 13400 38314 13464 38378
rect 13482 38314 13546 38378
rect 13564 38314 13628 38378
rect 13646 38314 13710 38378
rect 13728 38314 13792 38378
rect 13810 38314 13874 38378
rect 13892 38314 13956 38378
rect 13974 38314 14038 38378
rect 14056 38314 14120 38378
rect 14138 38314 14202 38378
rect 14220 38314 14284 38378
rect 14302 38314 14366 38378
rect 14384 38314 14448 38378
rect 14466 38314 14530 38378
rect 14548 38314 14612 38378
rect 14630 38314 14694 38378
rect 14712 38314 14776 38378
rect 14794 38314 14858 38378
rect 14876 38314 14940 38378
rect 111 38233 175 38297
rect 191 38233 255 38297
rect 271 38233 335 38297
rect 351 38233 415 38297
rect 431 38233 495 38297
rect 511 38233 575 38297
rect 591 38233 655 38297
rect 671 38233 735 38297
rect 751 38233 815 38297
rect 831 38233 895 38297
rect 911 38233 975 38297
rect 991 38233 1055 38297
rect 1071 38233 1135 38297
rect 1151 38233 1215 38297
rect 1231 38233 1295 38297
rect 1311 38233 1375 38297
rect 1391 38233 1455 38297
rect 1471 38233 1535 38297
rect 1551 38233 1615 38297
rect 1631 38233 1695 38297
rect 1711 38233 1775 38297
rect 1791 38233 1855 38297
rect 1871 38233 1935 38297
rect 1951 38233 2015 38297
rect 2031 38233 2095 38297
rect 2111 38233 2175 38297
rect 2191 38233 2255 38297
rect 2271 38233 2335 38297
rect 2351 38233 2415 38297
rect 2431 38233 2495 38297
rect 2511 38233 2575 38297
rect 12416 38233 12480 38297
rect 12498 38233 12562 38297
rect 12580 38233 12644 38297
rect 12662 38233 12726 38297
rect 12744 38233 12808 38297
rect 12826 38233 12890 38297
rect 12908 38233 12972 38297
rect 12990 38233 13054 38297
rect 13072 38233 13136 38297
rect 13154 38233 13218 38297
rect 13236 38233 13300 38297
rect 13318 38233 13382 38297
rect 13400 38233 13464 38297
rect 13482 38233 13546 38297
rect 13564 38233 13628 38297
rect 13646 38233 13710 38297
rect 13728 38233 13792 38297
rect 13810 38233 13874 38297
rect 13892 38233 13956 38297
rect 13974 38233 14038 38297
rect 14056 38233 14120 38297
rect 14138 38233 14202 38297
rect 14220 38233 14284 38297
rect 14302 38233 14366 38297
rect 14384 38233 14448 38297
rect 14466 38233 14530 38297
rect 14548 38233 14612 38297
rect 14630 38233 14694 38297
rect 14712 38233 14776 38297
rect 14794 38233 14858 38297
rect 14876 38233 14940 38297
rect 111 38152 175 38216
rect 191 38152 255 38216
rect 271 38152 335 38216
rect 351 38152 415 38216
rect 431 38152 495 38216
rect 511 38152 575 38216
rect 591 38152 655 38216
rect 671 38152 735 38216
rect 751 38152 815 38216
rect 831 38152 895 38216
rect 911 38152 975 38216
rect 991 38152 1055 38216
rect 1071 38152 1135 38216
rect 1151 38152 1215 38216
rect 1231 38152 1295 38216
rect 1311 38152 1375 38216
rect 1391 38152 1455 38216
rect 1471 38152 1535 38216
rect 1551 38152 1615 38216
rect 1631 38152 1695 38216
rect 1711 38152 1775 38216
rect 1791 38152 1855 38216
rect 1871 38152 1935 38216
rect 1951 38152 2015 38216
rect 2031 38152 2095 38216
rect 2111 38152 2175 38216
rect 2191 38152 2255 38216
rect 2271 38152 2335 38216
rect 2351 38152 2415 38216
rect 2431 38152 2495 38216
rect 2511 38152 2575 38216
rect 12416 38152 12480 38216
rect 12498 38152 12562 38216
rect 12580 38152 12644 38216
rect 12662 38152 12726 38216
rect 12744 38152 12808 38216
rect 12826 38152 12890 38216
rect 12908 38152 12972 38216
rect 12990 38152 13054 38216
rect 13072 38152 13136 38216
rect 13154 38152 13218 38216
rect 13236 38152 13300 38216
rect 13318 38152 13382 38216
rect 13400 38152 13464 38216
rect 13482 38152 13546 38216
rect 13564 38152 13628 38216
rect 13646 38152 13710 38216
rect 13728 38152 13792 38216
rect 13810 38152 13874 38216
rect 13892 38152 13956 38216
rect 13974 38152 14038 38216
rect 14056 38152 14120 38216
rect 14138 38152 14202 38216
rect 14220 38152 14284 38216
rect 14302 38152 14366 38216
rect 14384 38152 14448 38216
rect 14466 38152 14530 38216
rect 14548 38152 14612 38216
rect 14630 38152 14694 38216
rect 14712 38152 14776 38216
rect 14794 38152 14858 38216
rect 14876 38152 14940 38216
rect 111 38071 175 38135
rect 191 38071 255 38135
rect 271 38071 335 38135
rect 351 38071 415 38135
rect 431 38071 495 38135
rect 511 38071 575 38135
rect 591 38071 655 38135
rect 671 38071 735 38135
rect 751 38071 815 38135
rect 831 38071 895 38135
rect 911 38071 975 38135
rect 991 38071 1055 38135
rect 1071 38071 1135 38135
rect 1151 38071 1215 38135
rect 1231 38071 1295 38135
rect 1311 38071 1375 38135
rect 1391 38071 1455 38135
rect 1471 38071 1535 38135
rect 1551 38071 1615 38135
rect 1631 38071 1695 38135
rect 1711 38071 1775 38135
rect 1791 38071 1855 38135
rect 1871 38071 1935 38135
rect 1951 38071 2015 38135
rect 2031 38071 2095 38135
rect 2111 38071 2175 38135
rect 2191 38071 2255 38135
rect 2271 38071 2335 38135
rect 2351 38071 2415 38135
rect 2431 38071 2495 38135
rect 2511 38071 2575 38135
rect 12416 38071 12480 38135
rect 12498 38071 12562 38135
rect 12580 38071 12644 38135
rect 12662 38071 12726 38135
rect 12744 38071 12808 38135
rect 12826 38071 12890 38135
rect 12908 38071 12972 38135
rect 12990 38071 13054 38135
rect 13072 38071 13136 38135
rect 13154 38071 13218 38135
rect 13236 38071 13300 38135
rect 13318 38071 13382 38135
rect 13400 38071 13464 38135
rect 13482 38071 13546 38135
rect 13564 38071 13628 38135
rect 13646 38071 13710 38135
rect 13728 38071 13792 38135
rect 13810 38071 13874 38135
rect 13892 38071 13956 38135
rect 13974 38071 14038 38135
rect 14056 38071 14120 38135
rect 14138 38071 14202 38135
rect 14220 38071 14284 38135
rect 14302 38071 14366 38135
rect 14384 38071 14448 38135
rect 14466 38071 14530 38135
rect 14548 38071 14612 38135
rect 14630 38071 14694 38135
rect 14712 38071 14776 38135
rect 14794 38071 14858 38135
rect 14876 38071 14940 38135
rect 111 37990 175 38054
rect 191 37990 255 38054
rect 271 37990 335 38054
rect 351 37990 415 38054
rect 431 37990 495 38054
rect 511 37990 575 38054
rect 591 37990 655 38054
rect 671 37990 735 38054
rect 751 37990 815 38054
rect 831 37990 895 38054
rect 911 37990 975 38054
rect 991 37990 1055 38054
rect 1071 37990 1135 38054
rect 1151 37990 1215 38054
rect 1231 37990 1295 38054
rect 1311 37990 1375 38054
rect 1391 37990 1455 38054
rect 1471 37990 1535 38054
rect 1551 37990 1615 38054
rect 1631 37990 1695 38054
rect 1711 37990 1775 38054
rect 1791 37990 1855 38054
rect 1871 37990 1935 38054
rect 1951 37990 2015 38054
rect 2031 37990 2095 38054
rect 2111 37990 2175 38054
rect 2191 37990 2255 38054
rect 2271 37990 2335 38054
rect 2351 37990 2415 38054
rect 2431 37990 2495 38054
rect 2511 37990 2575 38054
rect 12416 37990 12480 38054
rect 12498 37990 12562 38054
rect 12580 37990 12644 38054
rect 12662 37990 12726 38054
rect 12744 37990 12808 38054
rect 12826 37990 12890 38054
rect 12908 37990 12972 38054
rect 12990 37990 13054 38054
rect 13072 37990 13136 38054
rect 13154 37990 13218 38054
rect 13236 37990 13300 38054
rect 13318 37990 13382 38054
rect 13400 37990 13464 38054
rect 13482 37990 13546 38054
rect 13564 37990 13628 38054
rect 13646 37990 13710 38054
rect 13728 37990 13792 38054
rect 13810 37990 13874 38054
rect 13892 37990 13956 38054
rect 13974 37990 14038 38054
rect 14056 37990 14120 38054
rect 14138 37990 14202 38054
rect 14220 37990 14284 38054
rect 14302 37990 14366 38054
rect 14384 37990 14448 38054
rect 14466 37990 14530 38054
rect 14548 37990 14612 38054
rect 14630 37990 14694 38054
rect 14712 37990 14776 38054
rect 14794 37990 14858 38054
rect 14876 37990 14940 38054
rect 111 37909 175 37973
rect 191 37909 255 37973
rect 271 37909 335 37973
rect 351 37909 415 37973
rect 431 37909 495 37973
rect 511 37909 575 37973
rect 591 37909 655 37973
rect 671 37909 735 37973
rect 751 37909 815 37973
rect 831 37909 895 37973
rect 911 37909 975 37973
rect 991 37909 1055 37973
rect 1071 37909 1135 37973
rect 1151 37909 1215 37973
rect 1231 37909 1295 37973
rect 1311 37909 1375 37973
rect 1391 37909 1455 37973
rect 1471 37909 1535 37973
rect 1551 37909 1615 37973
rect 1631 37909 1695 37973
rect 1711 37909 1775 37973
rect 1791 37909 1855 37973
rect 1871 37909 1935 37973
rect 1951 37909 2015 37973
rect 2031 37909 2095 37973
rect 2111 37909 2175 37973
rect 2191 37909 2255 37973
rect 2271 37909 2335 37973
rect 2351 37909 2415 37973
rect 2431 37909 2495 37973
rect 2511 37909 2575 37973
rect 12416 37909 12480 37973
rect 12498 37909 12562 37973
rect 12580 37909 12644 37973
rect 12662 37909 12726 37973
rect 12744 37909 12808 37973
rect 12826 37909 12890 37973
rect 12908 37909 12972 37973
rect 12990 37909 13054 37973
rect 13072 37909 13136 37973
rect 13154 37909 13218 37973
rect 13236 37909 13300 37973
rect 13318 37909 13382 37973
rect 13400 37909 13464 37973
rect 13482 37909 13546 37973
rect 13564 37909 13628 37973
rect 13646 37909 13710 37973
rect 13728 37909 13792 37973
rect 13810 37909 13874 37973
rect 13892 37909 13956 37973
rect 13974 37909 14038 37973
rect 14056 37909 14120 37973
rect 14138 37909 14202 37973
rect 14220 37909 14284 37973
rect 14302 37909 14366 37973
rect 14384 37909 14448 37973
rect 14466 37909 14530 37973
rect 14548 37909 14612 37973
rect 14630 37909 14694 37973
rect 14712 37909 14776 37973
rect 14794 37909 14858 37973
rect 14876 37909 14940 37973
rect 111 37828 175 37892
rect 191 37828 255 37892
rect 271 37828 335 37892
rect 351 37828 415 37892
rect 431 37828 495 37892
rect 511 37828 575 37892
rect 591 37828 655 37892
rect 671 37828 735 37892
rect 751 37828 815 37892
rect 831 37828 895 37892
rect 911 37828 975 37892
rect 991 37828 1055 37892
rect 1071 37828 1135 37892
rect 1151 37828 1215 37892
rect 1231 37828 1295 37892
rect 1311 37828 1375 37892
rect 1391 37828 1455 37892
rect 1471 37828 1535 37892
rect 1551 37828 1615 37892
rect 1631 37828 1695 37892
rect 1711 37828 1775 37892
rect 1791 37828 1855 37892
rect 1871 37828 1935 37892
rect 1951 37828 2015 37892
rect 2031 37828 2095 37892
rect 2111 37828 2175 37892
rect 2191 37828 2255 37892
rect 2271 37828 2335 37892
rect 2351 37828 2415 37892
rect 2431 37828 2495 37892
rect 2511 37828 2575 37892
rect 12416 37828 12480 37892
rect 12498 37828 12562 37892
rect 12580 37828 12644 37892
rect 12662 37828 12726 37892
rect 12744 37828 12808 37892
rect 12826 37828 12890 37892
rect 12908 37828 12972 37892
rect 12990 37828 13054 37892
rect 13072 37828 13136 37892
rect 13154 37828 13218 37892
rect 13236 37828 13300 37892
rect 13318 37828 13382 37892
rect 13400 37828 13464 37892
rect 13482 37828 13546 37892
rect 13564 37828 13628 37892
rect 13646 37828 13710 37892
rect 13728 37828 13792 37892
rect 13810 37828 13874 37892
rect 13892 37828 13956 37892
rect 13974 37828 14038 37892
rect 14056 37828 14120 37892
rect 14138 37828 14202 37892
rect 14220 37828 14284 37892
rect 14302 37828 14366 37892
rect 14384 37828 14448 37892
rect 14466 37828 14530 37892
rect 14548 37828 14612 37892
rect 14630 37828 14694 37892
rect 14712 37828 14776 37892
rect 14794 37828 14858 37892
rect 14876 37828 14940 37892
rect 111 37747 175 37811
rect 191 37747 255 37811
rect 271 37747 335 37811
rect 351 37747 415 37811
rect 431 37747 495 37811
rect 511 37747 575 37811
rect 591 37747 655 37811
rect 671 37747 735 37811
rect 751 37747 815 37811
rect 831 37747 895 37811
rect 911 37747 975 37811
rect 991 37747 1055 37811
rect 1071 37747 1135 37811
rect 1151 37747 1215 37811
rect 1231 37747 1295 37811
rect 1311 37747 1375 37811
rect 1391 37747 1455 37811
rect 1471 37747 1535 37811
rect 1551 37747 1615 37811
rect 1631 37747 1695 37811
rect 1711 37747 1775 37811
rect 1791 37747 1855 37811
rect 1871 37747 1935 37811
rect 1951 37747 2015 37811
rect 2031 37747 2095 37811
rect 2111 37747 2175 37811
rect 2191 37747 2255 37811
rect 2271 37747 2335 37811
rect 2351 37747 2415 37811
rect 2431 37747 2495 37811
rect 2511 37747 2575 37811
rect 12416 37747 12480 37811
rect 12498 37747 12562 37811
rect 12580 37747 12644 37811
rect 12662 37747 12726 37811
rect 12744 37747 12808 37811
rect 12826 37747 12890 37811
rect 12908 37747 12972 37811
rect 12990 37747 13054 37811
rect 13072 37747 13136 37811
rect 13154 37747 13218 37811
rect 13236 37747 13300 37811
rect 13318 37747 13382 37811
rect 13400 37747 13464 37811
rect 13482 37747 13546 37811
rect 13564 37747 13628 37811
rect 13646 37747 13710 37811
rect 13728 37747 13792 37811
rect 13810 37747 13874 37811
rect 13892 37747 13956 37811
rect 13974 37747 14038 37811
rect 14056 37747 14120 37811
rect 14138 37747 14202 37811
rect 14220 37747 14284 37811
rect 14302 37747 14366 37811
rect 14384 37747 14448 37811
rect 14466 37747 14530 37811
rect 14548 37747 14612 37811
rect 14630 37747 14694 37811
rect 14712 37747 14776 37811
rect 14794 37747 14858 37811
rect 14876 37747 14940 37811
rect 111 37666 175 37730
rect 191 37666 255 37730
rect 271 37666 335 37730
rect 351 37666 415 37730
rect 431 37666 495 37730
rect 511 37666 575 37730
rect 591 37666 655 37730
rect 671 37666 735 37730
rect 751 37666 815 37730
rect 831 37666 895 37730
rect 911 37666 975 37730
rect 991 37666 1055 37730
rect 1071 37666 1135 37730
rect 1151 37666 1215 37730
rect 1231 37666 1295 37730
rect 1311 37666 1375 37730
rect 1391 37666 1455 37730
rect 1471 37666 1535 37730
rect 1551 37666 1615 37730
rect 1631 37666 1695 37730
rect 1711 37666 1775 37730
rect 1791 37666 1855 37730
rect 1871 37666 1935 37730
rect 1951 37666 2015 37730
rect 2031 37666 2095 37730
rect 2111 37666 2175 37730
rect 2191 37666 2255 37730
rect 2271 37666 2335 37730
rect 2351 37666 2415 37730
rect 2431 37666 2495 37730
rect 2511 37666 2575 37730
rect 12416 37666 12480 37730
rect 12498 37666 12562 37730
rect 12580 37666 12644 37730
rect 12662 37666 12726 37730
rect 12744 37666 12808 37730
rect 12826 37666 12890 37730
rect 12908 37666 12972 37730
rect 12990 37666 13054 37730
rect 13072 37666 13136 37730
rect 13154 37666 13218 37730
rect 13236 37666 13300 37730
rect 13318 37666 13382 37730
rect 13400 37666 13464 37730
rect 13482 37666 13546 37730
rect 13564 37666 13628 37730
rect 13646 37666 13710 37730
rect 13728 37666 13792 37730
rect 13810 37666 13874 37730
rect 13892 37666 13956 37730
rect 13974 37666 14038 37730
rect 14056 37666 14120 37730
rect 14138 37666 14202 37730
rect 14220 37666 14284 37730
rect 14302 37666 14366 37730
rect 14384 37666 14448 37730
rect 14466 37666 14530 37730
rect 14548 37666 14612 37730
rect 14630 37666 14694 37730
rect 14712 37666 14776 37730
rect 14794 37666 14858 37730
rect 14876 37666 14940 37730
rect 111 37585 175 37649
rect 191 37585 255 37649
rect 271 37585 335 37649
rect 351 37585 415 37649
rect 431 37585 495 37649
rect 511 37585 575 37649
rect 591 37585 655 37649
rect 671 37585 735 37649
rect 751 37585 815 37649
rect 831 37585 895 37649
rect 911 37585 975 37649
rect 991 37585 1055 37649
rect 1071 37585 1135 37649
rect 1151 37585 1215 37649
rect 1231 37585 1295 37649
rect 1311 37585 1375 37649
rect 1391 37585 1455 37649
rect 1471 37585 1535 37649
rect 1551 37585 1615 37649
rect 1631 37585 1695 37649
rect 1711 37585 1775 37649
rect 1791 37585 1855 37649
rect 1871 37585 1935 37649
rect 1951 37585 2015 37649
rect 2031 37585 2095 37649
rect 2111 37585 2175 37649
rect 2191 37585 2255 37649
rect 2271 37585 2335 37649
rect 2351 37585 2415 37649
rect 2431 37585 2495 37649
rect 2511 37585 2575 37649
rect 12416 37585 12480 37649
rect 12498 37585 12562 37649
rect 12580 37585 12644 37649
rect 12662 37585 12726 37649
rect 12744 37585 12808 37649
rect 12826 37585 12890 37649
rect 12908 37585 12972 37649
rect 12990 37585 13054 37649
rect 13072 37585 13136 37649
rect 13154 37585 13218 37649
rect 13236 37585 13300 37649
rect 13318 37585 13382 37649
rect 13400 37585 13464 37649
rect 13482 37585 13546 37649
rect 13564 37585 13628 37649
rect 13646 37585 13710 37649
rect 13728 37585 13792 37649
rect 13810 37585 13874 37649
rect 13892 37585 13956 37649
rect 13974 37585 14038 37649
rect 14056 37585 14120 37649
rect 14138 37585 14202 37649
rect 14220 37585 14284 37649
rect 14302 37585 14366 37649
rect 14384 37585 14448 37649
rect 14466 37585 14530 37649
rect 14548 37585 14612 37649
rect 14630 37585 14694 37649
rect 14712 37585 14776 37649
rect 14794 37585 14858 37649
rect 14876 37585 14940 37649
rect 111 37504 175 37568
rect 191 37504 255 37568
rect 271 37504 335 37568
rect 351 37504 415 37568
rect 431 37504 495 37568
rect 511 37504 575 37568
rect 591 37504 655 37568
rect 671 37504 735 37568
rect 751 37504 815 37568
rect 831 37504 895 37568
rect 911 37504 975 37568
rect 991 37504 1055 37568
rect 1071 37504 1135 37568
rect 1151 37504 1215 37568
rect 1231 37504 1295 37568
rect 1311 37504 1375 37568
rect 1391 37504 1455 37568
rect 1471 37504 1535 37568
rect 1551 37504 1615 37568
rect 1631 37504 1695 37568
rect 1711 37504 1775 37568
rect 1791 37504 1855 37568
rect 1871 37504 1935 37568
rect 1951 37504 2015 37568
rect 2031 37504 2095 37568
rect 2111 37504 2175 37568
rect 2191 37504 2255 37568
rect 2271 37504 2335 37568
rect 2351 37504 2415 37568
rect 2431 37504 2495 37568
rect 2511 37504 2575 37568
rect 12416 37504 12480 37568
rect 12498 37504 12562 37568
rect 12580 37504 12644 37568
rect 12662 37504 12726 37568
rect 12744 37504 12808 37568
rect 12826 37504 12890 37568
rect 12908 37504 12972 37568
rect 12990 37504 13054 37568
rect 13072 37504 13136 37568
rect 13154 37504 13218 37568
rect 13236 37504 13300 37568
rect 13318 37504 13382 37568
rect 13400 37504 13464 37568
rect 13482 37504 13546 37568
rect 13564 37504 13628 37568
rect 13646 37504 13710 37568
rect 13728 37504 13792 37568
rect 13810 37504 13874 37568
rect 13892 37504 13956 37568
rect 13974 37504 14038 37568
rect 14056 37504 14120 37568
rect 14138 37504 14202 37568
rect 14220 37504 14284 37568
rect 14302 37504 14366 37568
rect 14384 37504 14448 37568
rect 14466 37504 14530 37568
rect 14548 37504 14612 37568
rect 14630 37504 14694 37568
rect 14712 37504 14776 37568
rect 14794 37504 14858 37568
rect 14876 37504 14940 37568
rect 111 37423 175 37487
rect 191 37423 255 37487
rect 271 37423 335 37487
rect 351 37423 415 37487
rect 431 37423 495 37487
rect 511 37423 575 37487
rect 591 37423 655 37487
rect 671 37423 735 37487
rect 751 37423 815 37487
rect 831 37423 895 37487
rect 911 37423 975 37487
rect 991 37423 1055 37487
rect 1071 37423 1135 37487
rect 1151 37423 1215 37487
rect 1231 37423 1295 37487
rect 1311 37423 1375 37487
rect 1391 37423 1455 37487
rect 1471 37423 1535 37487
rect 1551 37423 1615 37487
rect 1631 37423 1695 37487
rect 1711 37423 1775 37487
rect 1791 37423 1855 37487
rect 1871 37423 1935 37487
rect 1951 37423 2015 37487
rect 2031 37423 2095 37487
rect 2111 37423 2175 37487
rect 2191 37423 2255 37487
rect 2271 37423 2335 37487
rect 2351 37423 2415 37487
rect 2431 37423 2495 37487
rect 2511 37423 2575 37487
rect 12416 37423 12480 37487
rect 12498 37423 12562 37487
rect 12580 37423 12644 37487
rect 12662 37423 12726 37487
rect 12744 37423 12808 37487
rect 12826 37423 12890 37487
rect 12908 37423 12972 37487
rect 12990 37423 13054 37487
rect 13072 37423 13136 37487
rect 13154 37423 13218 37487
rect 13236 37423 13300 37487
rect 13318 37423 13382 37487
rect 13400 37423 13464 37487
rect 13482 37423 13546 37487
rect 13564 37423 13628 37487
rect 13646 37423 13710 37487
rect 13728 37423 13792 37487
rect 13810 37423 13874 37487
rect 13892 37423 13956 37487
rect 13974 37423 14038 37487
rect 14056 37423 14120 37487
rect 14138 37423 14202 37487
rect 14220 37423 14284 37487
rect 14302 37423 14366 37487
rect 14384 37423 14448 37487
rect 14466 37423 14530 37487
rect 14548 37423 14612 37487
rect 14630 37423 14694 37487
rect 14712 37423 14776 37487
rect 14794 37423 14858 37487
rect 14876 37423 14940 37487
rect 111 37342 175 37406
rect 191 37342 255 37406
rect 271 37342 335 37406
rect 351 37342 415 37406
rect 431 37342 495 37406
rect 511 37342 575 37406
rect 591 37342 655 37406
rect 671 37342 735 37406
rect 751 37342 815 37406
rect 831 37342 895 37406
rect 911 37342 975 37406
rect 991 37342 1055 37406
rect 1071 37342 1135 37406
rect 1151 37342 1215 37406
rect 1231 37342 1295 37406
rect 1311 37342 1375 37406
rect 1391 37342 1455 37406
rect 1471 37342 1535 37406
rect 1551 37342 1615 37406
rect 1631 37342 1695 37406
rect 1711 37342 1775 37406
rect 1791 37342 1855 37406
rect 1871 37342 1935 37406
rect 1951 37342 2015 37406
rect 2031 37342 2095 37406
rect 2111 37342 2175 37406
rect 2191 37342 2255 37406
rect 2271 37342 2335 37406
rect 2351 37342 2415 37406
rect 2431 37342 2495 37406
rect 2511 37342 2575 37406
rect 12416 37342 12480 37406
rect 12498 37342 12562 37406
rect 12580 37342 12644 37406
rect 12662 37342 12726 37406
rect 12744 37342 12808 37406
rect 12826 37342 12890 37406
rect 12908 37342 12972 37406
rect 12990 37342 13054 37406
rect 13072 37342 13136 37406
rect 13154 37342 13218 37406
rect 13236 37342 13300 37406
rect 13318 37342 13382 37406
rect 13400 37342 13464 37406
rect 13482 37342 13546 37406
rect 13564 37342 13628 37406
rect 13646 37342 13710 37406
rect 13728 37342 13792 37406
rect 13810 37342 13874 37406
rect 13892 37342 13956 37406
rect 13974 37342 14038 37406
rect 14056 37342 14120 37406
rect 14138 37342 14202 37406
rect 14220 37342 14284 37406
rect 14302 37342 14366 37406
rect 14384 37342 14448 37406
rect 14466 37342 14530 37406
rect 14548 37342 14612 37406
rect 14630 37342 14694 37406
rect 14712 37342 14776 37406
rect 14794 37342 14858 37406
rect 14876 37342 14940 37406
rect 111 37261 175 37325
rect 191 37261 255 37325
rect 271 37261 335 37325
rect 351 37261 415 37325
rect 431 37261 495 37325
rect 511 37261 575 37325
rect 591 37261 655 37325
rect 671 37261 735 37325
rect 751 37261 815 37325
rect 831 37261 895 37325
rect 911 37261 975 37325
rect 991 37261 1055 37325
rect 1071 37261 1135 37325
rect 1151 37261 1215 37325
rect 1231 37261 1295 37325
rect 1311 37261 1375 37325
rect 1391 37261 1455 37325
rect 1471 37261 1535 37325
rect 1551 37261 1615 37325
rect 1631 37261 1695 37325
rect 1711 37261 1775 37325
rect 1791 37261 1855 37325
rect 1871 37261 1935 37325
rect 1951 37261 2015 37325
rect 2031 37261 2095 37325
rect 2111 37261 2175 37325
rect 2191 37261 2255 37325
rect 2271 37261 2335 37325
rect 2351 37261 2415 37325
rect 2431 37261 2495 37325
rect 2511 37261 2575 37325
rect 12416 37261 12480 37325
rect 12498 37261 12562 37325
rect 12580 37261 12644 37325
rect 12662 37261 12726 37325
rect 12744 37261 12808 37325
rect 12826 37261 12890 37325
rect 12908 37261 12972 37325
rect 12990 37261 13054 37325
rect 13072 37261 13136 37325
rect 13154 37261 13218 37325
rect 13236 37261 13300 37325
rect 13318 37261 13382 37325
rect 13400 37261 13464 37325
rect 13482 37261 13546 37325
rect 13564 37261 13628 37325
rect 13646 37261 13710 37325
rect 13728 37261 13792 37325
rect 13810 37261 13874 37325
rect 13892 37261 13956 37325
rect 13974 37261 14038 37325
rect 14056 37261 14120 37325
rect 14138 37261 14202 37325
rect 14220 37261 14284 37325
rect 14302 37261 14366 37325
rect 14384 37261 14448 37325
rect 14466 37261 14530 37325
rect 14548 37261 14612 37325
rect 14630 37261 14694 37325
rect 14712 37261 14776 37325
rect 14794 37261 14858 37325
rect 14876 37261 14940 37325
rect 111 37180 175 37244
rect 191 37180 255 37244
rect 271 37180 335 37244
rect 351 37180 415 37244
rect 431 37180 495 37244
rect 511 37180 575 37244
rect 591 37180 655 37244
rect 671 37180 735 37244
rect 751 37180 815 37244
rect 831 37180 895 37244
rect 911 37180 975 37244
rect 991 37180 1055 37244
rect 1071 37180 1135 37244
rect 1151 37180 1215 37244
rect 1231 37180 1295 37244
rect 1311 37180 1375 37244
rect 1391 37180 1455 37244
rect 1471 37180 1535 37244
rect 1551 37180 1615 37244
rect 1631 37180 1695 37244
rect 1711 37180 1775 37244
rect 1791 37180 1855 37244
rect 1871 37180 1935 37244
rect 1951 37180 2015 37244
rect 2031 37180 2095 37244
rect 2111 37180 2175 37244
rect 2191 37180 2255 37244
rect 2271 37180 2335 37244
rect 2351 37180 2415 37244
rect 2431 37180 2495 37244
rect 2511 37180 2575 37244
rect 12416 37180 12480 37244
rect 12498 37180 12562 37244
rect 12580 37180 12644 37244
rect 12662 37180 12726 37244
rect 12744 37180 12808 37244
rect 12826 37180 12890 37244
rect 12908 37180 12972 37244
rect 12990 37180 13054 37244
rect 13072 37180 13136 37244
rect 13154 37180 13218 37244
rect 13236 37180 13300 37244
rect 13318 37180 13382 37244
rect 13400 37180 13464 37244
rect 13482 37180 13546 37244
rect 13564 37180 13628 37244
rect 13646 37180 13710 37244
rect 13728 37180 13792 37244
rect 13810 37180 13874 37244
rect 13892 37180 13956 37244
rect 13974 37180 14038 37244
rect 14056 37180 14120 37244
rect 14138 37180 14202 37244
rect 14220 37180 14284 37244
rect 14302 37180 14366 37244
rect 14384 37180 14448 37244
rect 14466 37180 14530 37244
rect 14548 37180 14612 37244
rect 14630 37180 14694 37244
rect 14712 37180 14776 37244
rect 14794 37180 14858 37244
rect 14876 37180 14940 37244
rect 111 37099 175 37163
rect 191 37099 255 37163
rect 271 37099 335 37163
rect 351 37099 415 37163
rect 431 37099 495 37163
rect 511 37099 575 37163
rect 591 37099 655 37163
rect 671 37099 735 37163
rect 751 37099 815 37163
rect 831 37099 895 37163
rect 911 37099 975 37163
rect 991 37099 1055 37163
rect 1071 37099 1135 37163
rect 1151 37099 1215 37163
rect 1231 37099 1295 37163
rect 1311 37099 1375 37163
rect 1391 37099 1455 37163
rect 1471 37099 1535 37163
rect 1551 37099 1615 37163
rect 1631 37099 1695 37163
rect 1711 37099 1775 37163
rect 1791 37099 1855 37163
rect 1871 37099 1935 37163
rect 1951 37099 2015 37163
rect 2031 37099 2095 37163
rect 2111 37099 2175 37163
rect 2191 37099 2255 37163
rect 2271 37099 2335 37163
rect 2351 37099 2415 37163
rect 2431 37099 2495 37163
rect 2511 37099 2575 37163
rect 12416 37099 12480 37163
rect 12498 37099 12562 37163
rect 12580 37099 12644 37163
rect 12662 37099 12726 37163
rect 12744 37099 12808 37163
rect 12826 37099 12890 37163
rect 12908 37099 12972 37163
rect 12990 37099 13054 37163
rect 13072 37099 13136 37163
rect 13154 37099 13218 37163
rect 13236 37099 13300 37163
rect 13318 37099 13382 37163
rect 13400 37099 13464 37163
rect 13482 37099 13546 37163
rect 13564 37099 13628 37163
rect 13646 37099 13710 37163
rect 13728 37099 13792 37163
rect 13810 37099 13874 37163
rect 13892 37099 13956 37163
rect 13974 37099 14038 37163
rect 14056 37099 14120 37163
rect 14138 37099 14202 37163
rect 14220 37099 14284 37163
rect 14302 37099 14366 37163
rect 14384 37099 14448 37163
rect 14466 37099 14530 37163
rect 14548 37099 14612 37163
rect 14630 37099 14694 37163
rect 14712 37099 14776 37163
rect 14794 37099 14858 37163
rect 14876 37099 14940 37163
rect 111 37018 175 37082
rect 191 37018 255 37082
rect 271 37018 335 37082
rect 351 37018 415 37082
rect 431 37018 495 37082
rect 511 37018 575 37082
rect 591 37018 655 37082
rect 671 37018 735 37082
rect 751 37018 815 37082
rect 831 37018 895 37082
rect 911 37018 975 37082
rect 991 37018 1055 37082
rect 1071 37018 1135 37082
rect 1151 37018 1215 37082
rect 1231 37018 1295 37082
rect 1311 37018 1375 37082
rect 1391 37018 1455 37082
rect 1471 37018 1535 37082
rect 1551 37018 1615 37082
rect 1631 37018 1695 37082
rect 1711 37018 1775 37082
rect 1791 37018 1855 37082
rect 1871 37018 1935 37082
rect 1951 37018 2015 37082
rect 2031 37018 2095 37082
rect 2111 37018 2175 37082
rect 2191 37018 2255 37082
rect 2271 37018 2335 37082
rect 2351 37018 2415 37082
rect 2431 37018 2495 37082
rect 2511 37018 2575 37082
rect 12416 37018 12480 37082
rect 12498 37018 12562 37082
rect 12580 37018 12644 37082
rect 12662 37018 12726 37082
rect 12744 37018 12808 37082
rect 12826 37018 12890 37082
rect 12908 37018 12972 37082
rect 12990 37018 13054 37082
rect 13072 37018 13136 37082
rect 13154 37018 13218 37082
rect 13236 37018 13300 37082
rect 13318 37018 13382 37082
rect 13400 37018 13464 37082
rect 13482 37018 13546 37082
rect 13564 37018 13628 37082
rect 13646 37018 13710 37082
rect 13728 37018 13792 37082
rect 13810 37018 13874 37082
rect 13892 37018 13956 37082
rect 13974 37018 14038 37082
rect 14056 37018 14120 37082
rect 14138 37018 14202 37082
rect 14220 37018 14284 37082
rect 14302 37018 14366 37082
rect 14384 37018 14448 37082
rect 14466 37018 14530 37082
rect 14548 37018 14612 37082
rect 14630 37018 14694 37082
rect 14712 37018 14776 37082
rect 14794 37018 14858 37082
rect 14876 37018 14940 37082
rect 111 36937 175 37001
rect 191 36937 255 37001
rect 271 36937 335 37001
rect 351 36937 415 37001
rect 431 36937 495 37001
rect 511 36937 575 37001
rect 591 36937 655 37001
rect 671 36937 735 37001
rect 751 36937 815 37001
rect 831 36937 895 37001
rect 911 36937 975 37001
rect 991 36937 1055 37001
rect 1071 36937 1135 37001
rect 1151 36937 1215 37001
rect 1231 36937 1295 37001
rect 1311 36937 1375 37001
rect 1391 36937 1455 37001
rect 1471 36937 1535 37001
rect 1551 36937 1615 37001
rect 1631 36937 1695 37001
rect 1711 36937 1775 37001
rect 1791 36937 1855 37001
rect 1871 36937 1935 37001
rect 1951 36937 2015 37001
rect 2031 36937 2095 37001
rect 2111 36937 2175 37001
rect 2191 36937 2255 37001
rect 2271 36937 2335 37001
rect 2351 36937 2415 37001
rect 2431 36937 2495 37001
rect 2511 36937 2575 37001
rect 12416 36937 12480 37001
rect 12498 36937 12562 37001
rect 12580 36937 12644 37001
rect 12662 36937 12726 37001
rect 12744 36937 12808 37001
rect 12826 36937 12890 37001
rect 12908 36937 12972 37001
rect 12990 36937 13054 37001
rect 13072 36937 13136 37001
rect 13154 36937 13218 37001
rect 13236 36937 13300 37001
rect 13318 36937 13382 37001
rect 13400 36937 13464 37001
rect 13482 36937 13546 37001
rect 13564 36937 13628 37001
rect 13646 36937 13710 37001
rect 13728 36937 13792 37001
rect 13810 36937 13874 37001
rect 13892 36937 13956 37001
rect 13974 36937 14038 37001
rect 14056 36937 14120 37001
rect 14138 36937 14202 37001
rect 14220 36937 14284 37001
rect 14302 36937 14366 37001
rect 14384 36937 14448 37001
rect 14466 36937 14530 37001
rect 14548 36937 14612 37001
rect 14630 36937 14694 37001
rect 14712 36937 14776 37001
rect 14794 36937 14858 37001
rect 14876 36937 14940 37001
rect 111 36856 175 36920
rect 191 36856 255 36920
rect 271 36856 335 36920
rect 351 36856 415 36920
rect 431 36856 495 36920
rect 511 36856 575 36920
rect 591 36856 655 36920
rect 671 36856 735 36920
rect 751 36856 815 36920
rect 831 36856 895 36920
rect 911 36856 975 36920
rect 991 36856 1055 36920
rect 1071 36856 1135 36920
rect 1151 36856 1215 36920
rect 1231 36856 1295 36920
rect 1311 36856 1375 36920
rect 1391 36856 1455 36920
rect 1471 36856 1535 36920
rect 1551 36856 1615 36920
rect 1631 36856 1695 36920
rect 1711 36856 1775 36920
rect 1791 36856 1855 36920
rect 1871 36856 1935 36920
rect 1951 36856 2015 36920
rect 2031 36856 2095 36920
rect 2111 36856 2175 36920
rect 2191 36856 2255 36920
rect 2271 36856 2335 36920
rect 2351 36856 2415 36920
rect 2431 36856 2495 36920
rect 2511 36856 2575 36920
rect 12416 36856 12480 36920
rect 12498 36856 12562 36920
rect 12580 36856 12644 36920
rect 12662 36856 12726 36920
rect 12744 36856 12808 36920
rect 12826 36856 12890 36920
rect 12908 36856 12972 36920
rect 12990 36856 13054 36920
rect 13072 36856 13136 36920
rect 13154 36856 13218 36920
rect 13236 36856 13300 36920
rect 13318 36856 13382 36920
rect 13400 36856 13464 36920
rect 13482 36856 13546 36920
rect 13564 36856 13628 36920
rect 13646 36856 13710 36920
rect 13728 36856 13792 36920
rect 13810 36856 13874 36920
rect 13892 36856 13956 36920
rect 13974 36856 14038 36920
rect 14056 36856 14120 36920
rect 14138 36856 14202 36920
rect 14220 36856 14284 36920
rect 14302 36856 14366 36920
rect 14384 36856 14448 36920
rect 14466 36856 14530 36920
rect 14548 36856 14612 36920
rect 14630 36856 14694 36920
rect 14712 36856 14776 36920
rect 14794 36856 14858 36920
rect 14876 36856 14940 36920
rect 111 36775 175 36839
rect 191 36775 255 36839
rect 271 36775 335 36839
rect 351 36775 415 36839
rect 431 36775 495 36839
rect 511 36775 575 36839
rect 591 36775 655 36839
rect 671 36775 735 36839
rect 751 36775 815 36839
rect 831 36775 895 36839
rect 911 36775 975 36839
rect 991 36775 1055 36839
rect 1071 36775 1135 36839
rect 1151 36775 1215 36839
rect 1231 36775 1295 36839
rect 1311 36775 1375 36839
rect 1391 36775 1455 36839
rect 1471 36775 1535 36839
rect 1551 36775 1615 36839
rect 1631 36775 1695 36839
rect 1711 36775 1775 36839
rect 1791 36775 1855 36839
rect 1871 36775 1935 36839
rect 1951 36775 2015 36839
rect 2031 36775 2095 36839
rect 2111 36775 2175 36839
rect 2191 36775 2255 36839
rect 2271 36775 2335 36839
rect 2351 36775 2415 36839
rect 2431 36775 2495 36839
rect 2511 36775 2575 36839
rect 12416 36775 12480 36839
rect 12498 36775 12562 36839
rect 12580 36775 12644 36839
rect 12662 36775 12726 36839
rect 12744 36775 12808 36839
rect 12826 36775 12890 36839
rect 12908 36775 12972 36839
rect 12990 36775 13054 36839
rect 13072 36775 13136 36839
rect 13154 36775 13218 36839
rect 13236 36775 13300 36839
rect 13318 36775 13382 36839
rect 13400 36775 13464 36839
rect 13482 36775 13546 36839
rect 13564 36775 13628 36839
rect 13646 36775 13710 36839
rect 13728 36775 13792 36839
rect 13810 36775 13874 36839
rect 13892 36775 13956 36839
rect 13974 36775 14038 36839
rect 14056 36775 14120 36839
rect 14138 36775 14202 36839
rect 14220 36775 14284 36839
rect 14302 36775 14366 36839
rect 14384 36775 14448 36839
rect 14466 36775 14530 36839
rect 14548 36775 14612 36839
rect 14630 36775 14694 36839
rect 14712 36775 14776 36839
rect 14794 36775 14858 36839
rect 14876 36775 14940 36839
rect 111 36694 175 36758
rect 191 36694 255 36758
rect 271 36694 335 36758
rect 351 36694 415 36758
rect 431 36694 495 36758
rect 511 36694 575 36758
rect 591 36694 655 36758
rect 671 36694 735 36758
rect 751 36694 815 36758
rect 831 36694 895 36758
rect 911 36694 975 36758
rect 991 36694 1055 36758
rect 1071 36694 1135 36758
rect 1151 36694 1215 36758
rect 1231 36694 1295 36758
rect 1311 36694 1375 36758
rect 1391 36694 1455 36758
rect 1471 36694 1535 36758
rect 1551 36694 1615 36758
rect 1631 36694 1695 36758
rect 1711 36694 1775 36758
rect 1791 36694 1855 36758
rect 1871 36694 1935 36758
rect 1951 36694 2015 36758
rect 2031 36694 2095 36758
rect 2111 36694 2175 36758
rect 2191 36694 2255 36758
rect 2271 36694 2335 36758
rect 2351 36694 2415 36758
rect 2431 36694 2495 36758
rect 2511 36694 2575 36758
rect 12416 36694 12480 36758
rect 12498 36694 12562 36758
rect 12580 36694 12644 36758
rect 12662 36694 12726 36758
rect 12744 36694 12808 36758
rect 12826 36694 12890 36758
rect 12908 36694 12972 36758
rect 12990 36694 13054 36758
rect 13072 36694 13136 36758
rect 13154 36694 13218 36758
rect 13236 36694 13300 36758
rect 13318 36694 13382 36758
rect 13400 36694 13464 36758
rect 13482 36694 13546 36758
rect 13564 36694 13628 36758
rect 13646 36694 13710 36758
rect 13728 36694 13792 36758
rect 13810 36694 13874 36758
rect 13892 36694 13956 36758
rect 13974 36694 14038 36758
rect 14056 36694 14120 36758
rect 14138 36694 14202 36758
rect 14220 36694 14284 36758
rect 14302 36694 14366 36758
rect 14384 36694 14448 36758
rect 14466 36694 14530 36758
rect 14548 36694 14612 36758
rect 14630 36694 14694 36758
rect 14712 36694 14776 36758
rect 14794 36694 14858 36758
rect 14876 36694 14940 36758
rect 111 36613 175 36677
rect 191 36613 255 36677
rect 271 36613 335 36677
rect 351 36613 415 36677
rect 431 36613 495 36677
rect 511 36613 575 36677
rect 591 36613 655 36677
rect 671 36613 735 36677
rect 751 36613 815 36677
rect 831 36613 895 36677
rect 911 36613 975 36677
rect 991 36613 1055 36677
rect 1071 36613 1135 36677
rect 1151 36613 1215 36677
rect 1231 36613 1295 36677
rect 1311 36613 1375 36677
rect 1391 36613 1455 36677
rect 1471 36613 1535 36677
rect 1551 36613 1615 36677
rect 1631 36613 1695 36677
rect 1711 36613 1775 36677
rect 1791 36613 1855 36677
rect 1871 36613 1935 36677
rect 1951 36613 2015 36677
rect 2031 36613 2095 36677
rect 2111 36613 2175 36677
rect 2191 36613 2255 36677
rect 2271 36613 2335 36677
rect 2351 36613 2415 36677
rect 2431 36613 2495 36677
rect 2511 36613 2575 36677
rect 12416 36613 12480 36677
rect 12498 36613 12562 36677
rect 12580 36613 12644 36677
rect 12662 36613 12726 36677
rect 12744 36613 12808 36677
rect 12826 36613 12890 36677
rect 12908 36613 12972 36677
rect 12990 36613 13054 36677
rect 13072 36613 13136 36677
rect 13154 36613 13218 36677
rect 13236 36613 13300 36677
rect 13318 36613 13382 36677
rect 13400 36613 13464 36677
rect 13482 36613 13546 36677
rect 13564 36613 13628 36677
rect 13646 36613 13710 36677
rect 13728 36613 13792 36677
rect 13810 36613 13874 36677
rect 13892 36613 13956 36677
rect 13974 36613 14038 36677
rect 14056 36613 14120 36677
rect 14138 36613 14202 36677
rect 14220 36613 14284 36677
rect 14302 36613 14366 36677
rect 14384 36613 14448 36677
rect 14466 36613 14530 36677
rect 14548 36613 14612 36677
rect 14630 36613 14694 36677
rect 14712 36613 14776 36677
rect 14794 36613 14858 36677
rect 14876 36613 14940 36677
rect 111 36532 175 36596
rect 191 36532 255 36596
rect 271 36532 335 36596
rect 351 36532 415 36596
rect 431 36532 495 36596
rect 511 36532 575 36596
rect 591 36532 655 36596
rect 671 36532 735 36596
rect 751 36532 815 36596
rect 831 36532 895 36596
rect 911 36532 975 36596
rect 991 36532 1055 36596
rect 1071 36532 1135 36596
rect 1151 36532 1215 36596
rect 1231 36532 1295 36596
rect 1311 36532 1375 36596
rect 1391 36532 1455 36596
rect 1471 36532 1535 36596
rect 1551 36532 1615 36596
rect 1631 36532 1695 36596
rect 1711 36532 1775 36596
rect 1791 36532 1855 36596
rect 1871 36532 1935 36596
rect 1951 36532 2015 36596
rect 2031 36532 2095 36596
rect 2111 36532 2175 36596
rect 2191 36532 2255 36596
rect 2271 36532 2335 36596
rect 2351 36532 2415 36596
rect 2431 36532 2495 36596
rect 2511 36532 2575 36596
rect 12416 36532 12480 36596
rect 12498 36532 12562 36596
rect 12580 36532 12644 36596
rect 12662 36532 12726 36596
rect 12744 36532 12808 36596
rect 12826 36532 12890 36596
rect 12908 36532 12972 36596
rect 12990 36532 13054 36596
rect 13072 36532 13136 36596
rect 13154 36532 13218 36596
rect 13236 36532 13300 36596
rect 13318 36532 13382 36596
rect 13400 36532 13464 36596
rect 13482 36532 13546 36596
rect 13564 36532 13628 36596
rect 13646 36532 13710 36596
rect 13728 36532 13792 36596
rect 13810 36532 13874 36596
rect 13892 36532 13956 36596
rect 13974 36532 14038 36596
rect 14056 36532 14120 36596
rect 14138 36532 14202 36596
rect 14220 36532 14284 36596
rect 14302 36532 14366 36596
rect 14384 36532 14448 36596
rect 14466 36532 14530 36596
rect 14548 36532 14612 36596
rect 14630 36532 14694 36596
rect 14712 36532 14776 36596
rect 14794 36532 14858 36596
rect 14876 36532 14940 36596
rect 111 36451 175 36515
rect 191 36451 255 36515
rect 271 36451 335 36515
rect 351 36451 415 36515
rect 431 36451 495 36515
rect 511 36451 575 36515
rect 591 36451 655 36515
rect 671 36451 735 36515
rect 751 36451 815 36515
rect 831 36451 895 36515
rect 911 36451 975 36515
rect 991 36451 1055 36515
rect 1071 36451 1135 36515
rect 1151 36451 1215 36515
rect 1231 36451 1295 36515
rect 1311 36451 1375 36515
rect 1391 36451 1455 36515
rect 1471 36451 1535 36515
rect 1551 36451 1615 36515
rect 1631 36451 1695 36515
rect 1711 36451 1775 36515
rect 1791 36451 1855 36515
rect 1871 36451 1935 36515
rect 1951 36451 2015 36515
rect 2031 36451 2095 36515
rect 2111 36451 2175 36515
rect 2191 36451 2255 36515
rect 2271 36451 2335 36515
rect 2351 36451 2415 36515
rect 2431 36451 2495 36515
rect 2511 36451 2575 36515
rect 12416 36451 12480 36515
rect 12498 36451 12562 36515
rect 12580 36451 12644 36515
rect 12662 36451 12726 36515
rect 12744 36451 12808 36515
rect 12826 36451 12890 36515
rect 12908 36451 12972 36515
rect 12990 36451 13054 36515
rect 13072 36451 13136 36515
rect 13154 36451 13218 36515
rect 13236 36451 13300 36515
rect 13318 36451 13382 36515
rect 13400 36451 13464 36515
rect 13482 36451 13546 36515
rect 13564 36451 13628 36515
rect 13646 36451 13710 36515
rect 13728 36451 13792 36515
rect 13810 36451 13874 36515
rect 13892 36451 13956 36515
rect 13974 36451 14038 36515
rect 14056 36451 14120 36515
rect 14138 36451 14202 36515
rect 14220 36451 14284 36515
rect 14302 36451 14366 36515
rect 14384 36451 14448 36515
rect 14466 36451 14530 36515
rect 14548 36451 14612 36515
rect 14630 36451 14694 36515
rect 14712 36451 14776 36515
rect 14794 36451 14858 36515
rect 14876 36451 14940 36515
rect 111 36370 175 36434
rect 191 36370 255 36434
rect 271 36370 335 36434
rect 351 36370 415 36434
rect 431 36370 495 36434
rect 511 36370 575 36434
rect 591 36370 655 36434
rect 671 36370 735 36434
rect 751 36370 815 36434
rect 831 36370 895 36434
rect 911 36370 975 36434
rect 991 36370 1055 36434
rect 1071 36370 1135 36434
rect 1151 36370 1215 36434
rect 1231 36370 1295 36434
rect 1311 36370 1375 36434
rect 1391 36370 1455 36434
rect 1471 36370 1535 36434
rect 1551 36370 1615 36434
rect 1631 36370 1695 36434
rect 1711 36370 1775 36434
rect 1791 36370 1855 36434
rect 1871 36370 1935 36434
rect 1951 36370 2015 36434
rect 2031 36370 2095 36434
rect 2111 36370 2175 36434
rect 2191 36370 2255 36434
rect 2271 36370 2335 36434
rect 2351 36370 2415 36434
rect 2431 36370 2495 36434
rect 2511 36370 2575 36434
rect 12416 36370 12480 36434
rect 12498 36370 12562 36434
rect 12580 36370 12644 36434
rect 12662 36370 12726 36434
rect 12744 36370 12808 36434
rect 12826 36370 12890 36434
rect 12908 36370 12972 36434
rect 12990 36370 13054 36434
rect 13072 36370 13136 36434
rect 13154 36370 13218 36434
rect 13236 36370 13300 36434
rect 13318 36370 13382 36434
rect 13400 36370 13464 36434
rect 13482 36370 13546 36434
rect 13564 36370 13628 36434
rect 13646 36370 13710 36434
rect 13728 36370 13792 36434
rect 13810 36370 13874 36434
rect 13892 36370 13956 36434
rect 13974 36370 14038 36434
rect 14056 36370 14120 36434
rect 14138 36370 14202 36434
rect 14220 36370 14284 36434
rect 14302 36370 14366 36434
rect 14384 36370 14448 36434
rect 14466 36370 14530 36434
rect 14548 36370 14612 36434
rect 14630 36370 14694 36434
rect 14712 36370 14776 36434
rect 14794 36370 14858 36434
rect 14876 36370 14940 36434
rect 111 36289 175 36353
rect 191 36289 255 36353
rect 271 36289 335 36353
rect 351 36289 415 36353
rect 431 36289 495 36353
rect 511 36289 575 36353
rect 591 36289 655 36353
rect 671 36289 735 36353
rect 751 36289 815 36353
rect 831 36289 895 36353
rect 911 36289 975 36353
rect 991 36289 1055 36353
rect 1071 36289 1135 36353
rect 1151 36289 1215 36353
rect 1231 36289 1295 36353
rect 1311 36289 1375 36353
rect 1391 36289 1455 36353
rect 1471 36289 1535 36353
rect 1551 36289 1615 36353
rect 1631 36289 1695 36353
rect 1711 36289 1775 36353
rect 1791 36289 1855 36353
rect 1871 36289 1935 36353
rect 1951 36289 2015 36353
rect 2031 36289 2095 36353
rect 2111 36289 2175 36353
rect 2191 36289 2255 36353
rect 2271 36289 2335 36353
rect 2351 36289 2415 36353
rect 2431 36289 2495 36353
rect 2511 36289 2575 36353
rect 12416 36289 12480 36353
rect 12498 36289 12562 36353
rect 12580 36289 12644 36353
rect 12662 36289 12726 36353
rect 12744 36289 12808 36353
rect 12826 36289 12890 36353
rect 12908 36289 12972 36353
rect 12990 36289 13054 36353
rect 13072 36289 13136 36353
rect 13154 36289 13218 36353
rect 13236 36289 13300 36353
rect 13318 36289 13382 36353
rect 13400 36289 13464 36353
rect 13482 36289 13546 36353
rect 13564 36289 13628 36353
rect 13646 36289 13710 36353
rect 13728 36289 13792 36353
rect 13810 36289 13874 36353
rect 13892 36289 13956 36353
rect 13974 36289 14038 36353
rect 14056 36289 14120 36353
rect 14138 36289 14202 36353
rect 14220 36289 14284 36353
rect 14302 36289 14366 36353
rect 14384 36289 14448 36353
rect 14466 36289 14530 36353
rect 14548 36289 14612 36353
rect 14630 36289 14694 36353
rect 14712 36289 14776 36353
rect 14794 36289 14858 36353
rect 14876 36289 14940 36353
rect 111 34768 2575 36272
rect 12416 36208 12480 36272
rect 12498 36208 12562 36272
rect 12580 36208 12644 36272
rect 12662 36208 12726 36272
rect 12744 36208 12808 36272
rect 12826 36208 12890 36272
rect 12908 36208 12972 36272
rect 12990 36208 13054 36272
rect 13072 36208 13136 36272
rect 13154 36208 13218 36272
rect 13236 36208 13300 36272
rect 13318 36208 13382 36272
rect 13400 36208 13464 36272
rect 13482 36208 13546 36272
rect 13564 36208 13628 36272
rect 13646 36208 13710 36272
rect 13728 36208 13792 36272
rect 13810 36208 13874 36272
rect 13892 36208 13956 36272
rect 13974 36208 14038 36272
rect 14056 36208 14120 36272
rect 14138 36208 14202 36272
rect 14220 36208 14284 36272
rect 14302 36208 14366 36272
rect 14384 36208 14448 36272
rect 14466 36208 14530 36272
rect 14548 36208 14612 36272
rect 14630 36208 14694 36272
rect 14712 36208 14776 36272
rect 14794 36208 14858 36272
rect 14876 36208 14940 36272
rect 12416 36128 12480 36192
rect 12498 36128 12562 36192
rect 12580 36128 12644 36192
rect 12662 36128 12726 36192
rect 12744 36128 12808 36192
rect 12826 36128 12890 36192
rect 12908 36128 12972 36192
rect 12990 36128 13054 36192
rect 13072 36128 13136 36192
rect 13154 36128 13218 36192
rect 13236 36128 13300 36192
rect 13318 36128 13382 36192
rect 13400 36128 13464 36192
rect 13482 36128 13546 36192
rect 13564 36128 13628 36192
rect 13646 36128 13710 36192
rect 13728 36128 13792 36192
rect 13810 36128 13874 36192
rect 13892 36128 13956 36192
rect 13974 36128 14038 36192
rect 14056 36128 14120 36192
rect 14138 36128 14202 36192
rect 14220 36128 14284 36192
rect 14302 36128 14366 36192
rect 14384 36128 14448 36192
rect 14466 36128 14530 36192
rect 14548 36128 14612 36192
rect 14630 36128 14694 36192
rect 14712 36128 14776 36192
rect 14794 36128 14858 36192
rect 14876 36128 14940 36192
rect 12416 36048 12480 36112
rect 12498 36048 12562 36112
rect 12580 36048 12644 36112
rect 12662 36048 12726 36112
rect 12744 36048 12808 36112
rect 12826 36048 12890 36112
rect 12908 36048 12972 36112
rect 12990 36048 13054 36112
rect 13072 36048 13136 36112
rect 13154 36048 13218 36112
rect 13236 36048 13300 36112
rect 13318 36048 13382 36112
rect 13400 36048 13464 36112
rect 13482 36048 13546 36112
rect 13564 36048 13628 36112
rect 13646 36048 13710 36112
rect 13728 36048 13792 36112
rect 13810 36048 13874 36112
rect 13892 36048 13956 36112
rect 13974 36048 14038 36112
rect 14056 36048 14120 36112
rect 14138 36048 14202 36112
rect 14220 36048 14284 36112
rect 14302 36048 14366 36112
rect 14384 36048 14448 36112
rect 14466 36048 14530 36112
rect 14548 36048 14612 36112
rect 14630 36048 14694 36112
rect 14712 36048 14776 36112
rect 14794 36048 14858 36112
rect 14876 36048 14940 36112
rect 12416 35968 12480 36032
rect 12498 35968 12562 36032
rect 12580 35968 12644 36032
rect 12662 35968 12726 36032
rect 12744 35968 12808 36032
rect 12826 35968 12890 36032
rect 12908 35968 12972 36032
rect 12990 35968 13054 36032
rect 13072 35968 13136 36032
rect 13154 35968 13218 36032
rect 13236 35968 13300 36032
rect 13318 35968 13382 36032
rect 13400 35968 13464 36032
rect 13482 35968 13546 36032
rect 13564 35968 13628 36032
rect 13646 35968 13710 36032
rect 13728 35968 13792 36032
rect 13810 35968 13874 36032
rect 13892 35968 13956 36032
rect 13974 35968 14038 36032
rect 14056 35968 14120 36032
rect 14138 35968 14202 36032
rect 14220 35968 14284 36032
rect 14302 35968 14366 36032
rect 14384 35968 14448 36032
rect 14466 35968 14530 36032
rect 14548 35968 14612 36032
rect 14630 35968 14694 36032
rect 14712 35968 14776 36032
rect 14794 35968 14858 36032
rect 14876 35968 14940 36032
rect 12416 35888 12480 35952
rect 12498 35888 12562 35952
rect 12580 35888 12644 35952
rect 12662 35888 12726 35952
rect 12744 35888 12808 35952
rect 12826 35888 12890 35952
rect 12908 35888 12972 35952
rect 12990 35888 13054 35952
rect 13072 35888 13136 35952
rect 13154 35888 13218 35952
rect 13236 35888 13300 35952
rect 13318 35888 13382 35952
rect 13400 35888 13464 35952
rect 13482 35888 13546 35952
rect 13564 35888 13628 35952
rect 13646 35888 13710 35952
rect 13728 35888 13792 35952
rect 13810 35888 13874 35952
rect 13892 35888 13956 35952
rect 13974 35888 14038 35952
rect 14056 35888 14120 35952
rect 14138 35888 14202 35952
rect 14220 35888 14284 35952
rect 14302 35888 14366 35952
rect 14384 35888 14448 35952
rect 14466 35888 14530 35952
rect 14548 35888 14612 35952
rect 14630 35888 14694 35952
rect 14712 35888 14776 35952
rect 14794 35888 14858 35952
rect 14876 35888 14940 35952
rect 12416 35808 12480 35872
rect 12498 35808 12562 35872
rect 12580 35808 12644 35872
rect 12662 35808 12726 35872
rect 12744 35808 12808 35872
rect 12826 35808 12890 35872
rect 12908 35808 12972 35872
rect 12990 35808 13054 35872
rect 13072 35808 13136 35872
rect 13154 35808 13218 35872
rect 13236 35808 13300 35872
rect 13318 35808 13382 35872
rect 13400 35808 13464 35872
rect 13482 35808 13546 35872
rect 13564 35808 13628 35872
rect 13646 35808 13710 35872
rect 13728 35808 13792 35872
rect 13810 35808 13874 35872
rect 13892 35808 13956 35872
rect 13974 35808 14038 35872
rect 14056 35808 14120 35872
rect 14138 35808 14202 35872
rect 14220 35808 14284 35872
rect 14302 35808 14366 35872
rect 14384 35808 14448 35872
rect 14466 35808 14530 35872
rect 14548 35808 14612 35872
rect 14630 35808 14694 35872
rect 14712 35808 14776 35872
rect 14794 35808 14858 35872
rect 14876 35808 14940 35872
rect 12416 35728 12480 35792
rect 12498 35728 12562 35792
rect 12580 35728 12644 35792
rect 12662 35728 12726 35792
rect 12744 35728 12808 35792
rect 12826 35728 12890 35792
rect 12908 35728 12972 35792
rect 12990 35728 13054 35792
rect 13072 35728 13136 35792
rect 13154 35728 13218 35792
rect 13236 35728 13300 35792
rect 13318 35728 13382 35792
rect 13400 35728 13464 35792
rect 13482 35728 13546 35792
rect 13564 35728 13628 35792
rect 13646 35728 13710 35792
rect 13728 35728 13792 35792
rect 13810 35728 13874 35792
rect 13892 35728 13956 35792
rect 13974 35728 14038 35792
rect 14056 35728 14120 35792
rect 14138 35728 14202 35792
rect 14220 35728 14284 35792
rect 14302 35728 14366 35792
rect 14384 35728 14448 35792
rect 14466 35728 14530 35792
rect 14548 35728 14612 35792
rect 14630 35728 14694 35792
rect 14712 35728 14776 35792
rect 14794 35728 14858 35792
rect 14876 35728 14940 35792
rect 12416 35648 12480 35712
rect 12498 35648 12562 35712
rect 12580 35648 12644 35712
rect 12662 35648 12726 35712
rect 12744 35648 12808 35712
rect 12826 35648 12890 35712
rect 12908 35648 12972 35712
rect 12990 35648 13054 35712
rect 13072 35648 13136 35712
rect 13154 35648 13218 35712
rect 13236 35648 13300 35712
rect 13318 35648 13382 35712
rect 13400 35648 13464 35712
rect 13482 35648 13546 35712
rect 13564 35648 13628 35712
rect 13646 35648 13710 35712
rect 13728 35648 13792 35712
rect 13810 35648 13874 35712
rect 13892 35648 13956 35712
rect 13974 35648 14038 35712
rect 14056 35648 14120 35712
rect 14138 35648 14202 35712
rect 14220 35648 14284 35712
rect 14302 35648 14366 35712
rect 14384 35648 14448 35712
rect 14466 35648 14530 35712
rect 14548 35648 14612 35712
rect 14630 35648 14694 35712
rect 14712 35648 14776 35712
rect 14794 35648 14858 35712
rect 14876 35648 14940 35712
rect 12416 35568 12480 35632
rect 12498 35568 12562 35632
rect 12580 35568 12644 35632
rect 12662 35568 12726 35632
rect 12744 35568 12808 35632
rect 12826 35568 12890 35632
rect 12908 35568 12972 35632
rect 12990 35568 13054 35632
rect 13072 35568 13136 35632
rect 13154 35568 13218 35632
rect 13236 35568 13300 35632
rect 13318 35568 13382 35632
rect 13400 35568 13464 35632
rect 13482 35568 13546 35632
rect 13564 35568 13628 35632
rect 13646 35568 13710 35632
rect 13728 35568 13792 35632
rect 13810 35568 13874 35632
rect 13892 35568 13956 35632
rect 13974 35568 14038 35632
rect 14056 35568 14120 35632
rect 14138 35568 14202 35632
rect 14220 35568 14284 35632
rect 14302 35568 14366 35632
rect 14384 35568 14448 35632
rect 14466 35568 14530 35632
rect 14548 35568 14612 35632
rect 14630 35568 14694 35632
rect 14712 35568 14776 35632
rect 14794 35568 14858 35632
rect 14876 35568 14940 35632
rect 12416 35488 12480 35552
rect 12498 35488 12562 35552
rect 12580 35488 12644 35552
rect 12662 35488 12726 35552
rect 12744 35488 12808 35552
rect 12826 35488 12890 35552
rect 12908 35488 12972 35552
rect 12990 35488 13054 35552
rect 13072 35488 13136 35552
rect 13154 35488 13218 35552
rect 13236 35488 13300 35552
rect 13318 35488 13382 35552
rect 13400 35488 13464 35552
rect 13482 35488 13546 35552
rect 13564 35488 13628 35552
rect 13646 35488 13710 35552
rect 13728 35488 13792 35552
rect 13810 35488 13874 35552
rect 13892 35488 13956 35552
rect 13974 35488 14038 35552
rect 14056 35488 14120 35552
rect 14138 35488 14202 35552
rect 14220 35488 14284 35552
rect 14302 35488 14366 35552
rect 14384 35488 14448 35552
rect 14466 35488 14530 35552
rect 14548 35488 14612 35552
rect 14630 35488 14694 35552
rect 14712 35488 14776 35552
rect 14794 35488 14858 35552
rect 14876 35488 14940 35552
rect 12416 35408 12480 35472
rect 12498 35408 12562 35472
rect 12580 35408 12644 35472
rect 12662 35408 12726 35472
rect 12744 35408 12808 35472
rect 12826 35408 12890 35472
rect 12908 35408 12972 35472
rect 12990 35408 13054 35472
rect 13072 35408 13136 35472
rect 13154 35408 13218 35472
rect 13236 35408 13300 35472
rect 13318 35408 13382 35472
rect 13400 35408 13464 35472
rect 13482 35408 13546 35472
rect 13564 35408 13628 35472
rect 13646 35408 13710 35472
rect 13728 35408 13792 35472
rect 13810 35408 13874 35472
rect 13892 35408 13956 35472
rect 13974 35408 14038 35472
rect 14056 35408 14120 35472
rect 14138 35408 14202 35472
rect 14220 35408 14284 35472
rect 14302 35408 14366 35472
rect 14384 35408 14448 35472
rect 14466 35408 14530 35472
rect 14548 35408 14612 35472
rect 14630 35408 14694 35472
rect 14712 35408 14776 35472
rect 14794 35408 14858 35472
rect 14876 35408 14940 35472
rect 12416 35328 12480 35392
rect 12498 35328 12562 35392
rect 12580 35328 12644 35392
rect 12662 35328 12726 35392
rect 12744 35328 12808 35392
rect 12826 35328 12890 35392
rect 12908 35328 12972 35392
rect 12990 35328 13054 35392
rect 13072 35328 13136 35392
rect 13154 35328 13218 35392
rect 13236 35328 13300 35392
rect 13318 35328 13382 35392
rect 13400 35328 13464 35392
rect 13482 35328 13546 35392
rect 13564 35328 13628 35392
rect 13646 35328 13710 35392
rect 13728 35328 13792 35392
rect 13810 35328 13874 35392
rect 13892 35328 13956 35392
rect 13974 35328 14038 35392
rect 14056 35328 14120 35392
rect 14138 35328 14202 35392
rect 14220 35328 14284 35392
rect 14302 35328 14366 35392
rect 14384 35328 14448 35392
rect 14466 35328 14530 35392
rect 14548 35328 14612 35392
rect 14630 35328 14694 35392
rect 14712 35328 14776 35392
rect 14794 35328 14858 35392
rect 14876 35328 14940 35392
rect 12416 35248 12480 35312
rect 12498 35248 12562 35312
rect 12580 35248 12644 35312
rect 12662 35248 12726 35312
rect 12744 35248 12808 35312
rect 12826 35248 12890 35312
rect 12908 35248 12972 35312
rect 12990 35248 13054 35312
rect 13072 35248 13136 35312
rect 13154 35248 13218 35312
rect 13236 35248 13300 35312
rect 13318 35248 13382 35312
rect 13400 35248 13464 35312
rect 13482 35248 13546 35312
rect 13564 35248 13628 35312
rect 13646 35248 13710 35312
rect 13728 35248 13792 35312
rect 13810 35248 13874 35312
rect 13892 35248 13956 35312
rect 13974 35248 14038 35312
rect 14056 35248 14120 35312
rect 14138 35248 14202 35312
rect 14220 35248 14284 35312
rect 14302 35248 14366 35312
rect 14384 35248 14448 35312
rect 14466 35248 14530 35312
rect 14548 35248 14612 35312
rect 14630 35248 14694 35312
rect 14712 35248 14776 35312
rect 14794 35248 14858 35312
rect 14876 35248 14940 35312
rect 12416 35168 12480 35232
rect 12498 35168 12562 35232
rect 12580 35168 12644 35232
rect 12662 35168 12726 35232
rect 12744 35168 12808 35232
rect 12826 35168 12890 35232
rect 12908 35168 12972 35232
rect 12990 35168 13054 35232
rect 13072 35168 13136 35232
rect 13154 35168 13218 35232
rect 13236 35168 13300 35232
rect 13318 35168 13382 35232
rect 13400 35168 13464 35232
rect 13482 35168 13546 35232
rect 13564 35168 13628 35232
rect 13646 35168 13710 35232
rect 13728 35168 13792 35232
rect 13810 35168 13874 35232
rect 13892 35168 13956 35232
rect 13974 35168 14038 35232
rect 14056 35168 14120 35232
rect 14138 35168 14202 35232
rect 14220 35168 14284 35232
rect 14302 35168 14366 35232
rect 14384 35168 14448 35232
rect 14466 35168 14530 35232
rect 14548 35168 14612 35232
rect 14630 35168 14694 35232
rect 14712 35168 14776 35232
rect 14794 35168 14858 35232
rect 14876 35168 14940 35232
rect 12416 35088 12480 35152
rect 12498 35088 12562 35152
rect 12580 35088 12644 35152
rect 12662 35088 12726 35152
rect 12744 35088 12808 35152
rect 12826 35088 12890 35152
rect 12908 35088 12972 35152
rect 12990 35088 13054 35152
rect 13072 35088 13136 35152
rect 13154 35088 13218 35152
rect 13236 35088 13300 35152
rect 13318 35088 13382 35152
rect 13400 35088 13464 35152
rect 13482 35088 13546 35152
rect 13564 35088 13628 35152
rect 13646 35088 13710 35152
rect 13728 35088 13792 35152
rect 13810 35088 13874 35152
rect 13892 35088 13956 35152
rect 13974 35088 14038 35152
rect 14056 35088 14120 35152
rect 14138 35088 14202 35152
rect 14220 35088 14284 35152
rect 14302 35088 14366 35152
rect 14384 35088 14448 35152
rect 14466 35088 14530 35152
rect 14548 35088 14612 35152
rect 14630 35088 14694 35152
rect 14712 35088 14776 35152
rect 14794 35088 14858 35152
rect 14876 35088 14940 35152
rect 12416 35008 12480 35072
rect 12498 35008 12562 35072
rect 12580 35008 12644 35072
rect 12662 35008 12726 35072
rect 12744 35008 12808 35072
rect 12826 35008 12890 35072
rect 12908 35008 12972 35072
rect 12990 35008 13054 35072
rect 13072 35008 13136 35072
rect 13154 35008 13218 35072
rect 13236 35008 13300 35072
rect 13318 35008 13382 35072
rect 13400 35008 13464 35072
rect 13482 35008 13546 35072
rect 13564 35008 13628 35072
rect 13646 35008 13710 35072
rect 13728 35008 13792 35072
rect 13810 35008 13874 35072
rect 13892 35008 13956 35072
rect 13974 35008 14038 35072
rect 14056 35008 14120 35072
rect 14138 35008 14202 35072
rect 14220 35008 14284 35072
rect 14302 35008 14366 35072
rect 14384 35008 14448 35072
rect 14466 35008 14530 35072
rect 14548 35008 14612 35072
rect 14630 35008 14694 35072
rect 14712 35008 14776 35072
rect 14794 35008 14858 35072
rect 14876 35008 14940 35072
rect 12416 34928 12480 34992
rect 12498 34928 12562 34992
rect 12580 34928 12644 34992
rect 12662 34928 12726 34992
rect 12744 34928 12808 34992
rect 12826 34928 12890 34992
rect 12908 34928 12972 34992
rect 12990 34928 13054 34992
rect 13072 34928 13136 34992
rect 13154 34928 13218 34992
rect 13236 34928 13300 34992
rect 13318 34928 13382 34992
rect 13400 34928 13464 34992
rect 13482 34928 13546 34992
rect 13564 34928 13628 34992
rect 13646 34928 13710 34992
rect 13728 34928 13792 34992
rect 13810 34928 13874 34992
rect 13892 34928 13956 34992
rect 13974 34928 14038 34992
rect 14056 34928 14120 34992
rect 14138 34928 14202 34992
rect 14220 34928 14284 34992
rect 14302 34928 14366 34992
rect 14384 34928 14448 34992
rect 14466 34928 14530 34992
rect 14548 34928 14612 34992
rect 14630 34928 14694 34992
rect 14712 34928 14776 34992
rect 14794 34928 14858 34992
rect 14876 34928 14940 34992
rect 12416 34848 12480 34912
rect 12498 34848 12562 34912
rect 12580 34848 12644 34912
rect 12662 34848 12726 34912
rect 12744 34848 12808 34912
rect 12826 34848 12890 34912
rect 12908 34848 12972 34912
rect 12990 34848 13054 34912
rect 13072 34848 13136 34912
rect 13154 34848 13218 34912
rect 13236 34848 13300 34912
rect 13318 34848 13382 34912
rect 13400 34848 13464 34912
rect 13482 34848 13546 34912
rect 13564 34848 13628 34912
rect 13646 34848 13710 34912
rect 13728 34848 13792 34912
rect 13810 34848 13874 34912
rect 13892 34848 13956 34912
rect 13974 34848 14038 34912
rect 14056 34848 14120 34912
rect 14138 34848 14202 34912
rect 14220 34848 14284 34912
rect 14302 34848 14366 34912
rect 14384 34848 14448 34912
rect 14466 34848 14530 34912
rect 14548 34848 14612 34912
rect 14630 34848 14694 34912
rect 14712 34848 14776 34912
rect 14794 34848 14858 34912
rect 14876 34848 14940 34912
rect 12416 34768 12480 34832
rect 12498 34768 12562 34832
rect 12580 34768 12644 34832
rect 12662 34768 12726 34832
rect 12744 34768 12808 34832
rect 12826 34768 12890 34832
rect 12908 34768 12972 34832
rect 12990 34768 13054 34832
rect 13072 34768 13136 34832
rect 13154 34768 13218 34832
rect 13236 34768 13300 34832
rect 13318 34768 13382 34832
rect 13400 34768 13464 34832
rect 13482 34768 13546 34832
rect 13564 34768 13628 34832
rect 13646 34768 13710 34832
rect 13728 34768 13792 34832
rect 13810 34768 13874 34832
rect 13892 34768 13956 34832
rect 13974 34768 14038 34832
rect 14056 34768 14120 34832
rect 14138 34768 14202 34832
rect 14220 34768 14284 34832
rect 14302 34768 14366 34832
rect 14384 34768 14448 34832
rect 14466 34768 14530 34832
rect 14548 34768 14612 34832
rect 14630 34768 14694 34832
rect 14712 34768 14776 34832
rect 14794 34768 14858 34832
rect 14876 34768 14940 34832
rect 106 12070 170 12134
rect 188 12070 252 12134
rect 270 12070 334 12134
rect 352 12070 416 12134
rect 434 12070 498 12134
rect 516 12070 580 12134
rect 598 12070 662 12134
rect 679 12070 743 12134
rect 760 12070 824 12134
rect 841 12070 905 12134
rect 922 12070 986 12134
rect 1003 12070 1067 12134
rect 1084 12070 1148 12134
rect 1165 12070 1229 12134
rect 1246 12070 1310 12134
rect 1327 12070 1391 12134
rect 1408 12070 1472 12134
rect 1489 12070 1553 12134
rect 1570 12070 1634 12134
rect 1651 12070 1715 12134
rect 1732 12070 1796 12134
rect 1813 12070 1877 12134
rect 1894 12070 1958 12134
rect 1975 12070 2039 12134
rect 2056 12070 2120 12134
rect 2137 12070 2201 12134
rect 2218 12070 2282 12134
rect 2299 12070 2363 12134
rect 2380 12070 2444 12134
rect 2461 12070 2525 12134
rect 2542 12070 2606 12134
rect 2623 12070 2687 12134
rect 2704 12070 2768 12134
rect 2785 12070 2849 12134
rect 2866 12070 2930 12134
rect 2947 12070 3011 12134
rect 3028 12070 3092 12134
rect 3109 12070 3173 12134
rect 3190 12070 3254 12134
rect 3271 12070 3335 12134
rect 3352 12070 3416 12134
rect 3433 12070 3497 12134
rect 3514 12070 3578 12134
rect 3595 12070 3659 12134
rect 3676 12070 3740 12134
rect 3757 12070 3821 12134
rect 3838 12070 3902 12134
rect 3919 12070 3983 12134
rect 4000 12070 4064 12134
rect 4081 12070 4145 12134
rect 4162 12070 4226 12134
rect 4243 12070 4307 12134
rect 4324 12070 4388 12134
rect 4405 12070 4469 12134
rect 4486 12070 4550 12134
rect 4567 12070 4631 12134
rect 4648 12070 4712 12134
rect 4729 12070 4793 12134
rect 4810 12070 4874 12134
rect 10157 12070 10221 12134
rect 10239 12070 10303 12134
rect 10321 12070 10385 12134
rect 10403 12070 10467 12134
rect 10485 12070 10549 12134
rect 10567 12070 10631 12134
rect 10649 12070 10713 12134
rect 10731 12070 10795 12134
rect 10813 12070 10877 12134
rect 10895 12070 10959 12134
rect 10977 12070 11041 12134
rect 11059 12070 11123 12134
rect 11141 12070 11205 12134
rect 11223 12070 11287 12134
rect 11305 12070 11369 12134
rect 11386 12070 11450 12134
rect 11467 12070 11531 12134
rect 11548 12070 11612 12134
rect 11629 12070 11693 12134
rect 11710 12070 11774 12134
rect 11791 12070 11855 12134
rect 11872 12070 11936 12134
rect 11953 12070 12017 12134
rect 12034 12070 12098 12134
rect 12115 12070 12179 12134
rect 12196 12070 12260 12134
rect 12277 12070 12341 12134
rect 12358 12070 12422 12134
rect 12439 12070 12503 12134
rect 12520 12070 12584 12134
rect 12601 12070 12665 12134
rect 12682 12070 12746 12134
rect 12763 12070 12827 12134
rect 12844 12070 12908 12134
rect 12925 12070 12989 12134
rect 13006 12070 13070 12134
rect 13087 12070 13151 12134
rect 13168 12070 13232 12134
rect 13249 12070 13313 12134
rect 13330 12070 13394 12134
rect 13411 12070 13475 12134
rect 13492 12070 13556 12134
rect 13573 12070 13637 12134
rect 13654 12070 13718 12134
rect 13735 12070 13799 12134
rect 13816 12070 13880 12134
rect 13897 12070 13961 12134
rect 13978 12070 14042 12134
rect 14059 12070 14123 12134
rect 14140 12070 14204 12134
rect 14221 12070 14285 12134
rect 14302 12070 14366 12134
rect 14383 12070 14447 12134
rect 14464 12070 14528 12134
rect 14545 12070 14609 12134
rect 14626 12070 14690 12134
rect 14707 12070 14771 12134
rect 14788 12070 14852 12134
rect 106 11988 170 12052
rect 188 11988 252 12052
rect 270 11988 334 12052
rect 352 11988 416 12052
rect 434 11988 498 12052
rect 516 11988 580 12052
rect 598 11988 662 12052
rect 679 11988 743 12052
rect 760 11988 824 12052
rect 841 11988 905 12052
rect 922 11988 986 12052
rect 1003 11988 1067 12052
rect 1084 11988 1148 12052
rect 1165 11988 1229 12052
rect 1246 11988 1310 12052
rect 1327 11988 1391 12052
rect 1408 11988 1472 12052
rect 1489 11988 1553 12052
rect 1570 11988 1634 12052
rect 1651 11988 1715 12052
rect 1732 11988 1796 12052
rect 1813 11988 1877 12052
rect 1894 11988 1958 12052
rect 1975 11988 2039 12052
rect 2056 11988 2120 12052
rect 2137 11988 2201 12052
rect 2218 11988 2282 12052
rect 2299 11988 2363 12052
rect 2380 11988 2444 12052
rect 2461 11988 2525 12052
rect 2542 11988 2606 12052
rect 2623 11988 2687 12052
rect 2704 11988 2768 12052
rect 2785 11988 2849 12052
rect 2866 11988 2930 12052
rect 2947 11988 3011 12052
rect 3028 11988 3092 12052
rect 3109 11988 3173 12052
rect 3190 11988 3254 12052
rect 3271 11988 3335 12052
rect 3352 11988 3416 12052
rect 3433 11988 3497 12052
rect 3514 11988 3578 12052
rect 3595 11988 3659 12052
rect 3676 11988 3740 12052
rect 3757 11988 3821 12052
rect 3838 11988 3902 12052
rect 3919 11988 3983 12052
rect 4000 11988 4064 12052
rect 4081 11988 4145 12052
rect 4162 11988 4226 12052
rect 4243 11988 4307 12052
rect 4324 11988 4388 12052
rect 4405 11988 4469 12052
rect 4486 11988 4550 12052
rect 4567 11988 4631 12052
rect 4648 11988 4712 12052
rect 4729 11988 4793 12052
rect 4810 11988 4874 12052
rect 10157 11988 10221 12052
rect 10239 11988 10303 12052
rect 10321 11988 10385 12052
rect 10403 11988 10467 12052
rect 10485 11988 10549 12052
rect 10567 11988 10631 12052
rect 10649 11988 10713 12052
rect 10731 11988 10795 12052
rect 10813 11988 10877 12052
rect 10895 11988 10959 12052
rect 10977 11988 11041 12052
rect 11059 11988 11123 12052
rect 11141 11988 11205 12052
rect 11223 11988 11287 12052
rect 11305 11988 11369 12052
rect 11386 11988 11450 12052
rect 11467 11988 11531 12052
rect 11548 11988 11612 12052
rect 11629 11988 11693 12052
rect 11710 11988 11774 12052
rect 11791 11988 11855 12052
rect 11872 11988 11936 12052
rect 11953 11988 12017 12052
rect 12034 11988 12098 12052
rect 12115 11988 12179 12052
rect 12196 11988 12260 12052
rect 12277 11988 12341 12052
rect 12358 11988 12422 12052
rect 12439 11988 12503 12052
rect 12520 11988 12584 12052
rect 12601 11988 12665 12052
rect 12682 11988 12746 12052
rect 12763 11988 12827 12052
rect 12844 11988 12908 12052
rect 12925 11988 12989 12052
rect 13006 11988 13070 12052
rect 13087 11988 13151 12052
rect 13168 11988 13232 12052
rect 13249 11988 13313 12052
rect 13330 11988 13394 12052
rect 13411 11988 13475 12052
rect 13492 11988 13556 12052
rect 13573 11988 13637 12052
rect 13654 11988 13718 12052
rect 13735 11988 13799 12052
rect 13816 11988 13880 12052
rect 13897 11988 13961 12052
rect 13978 11988 14042 12052
rect 14059 11988 14123 12052
rect 14140 11988 14204 12052
rect 14221 11988 14285 12052
rect 14302 11988 14366 12052
rect 14383 11988 14447 12052
rect 14464 11988 14528 12052
rect 14545 11988 14609 12052
rect 14626 11988 14690 12052
rect 14707 11988 14771 12052
rect 14788 11988 14852 12052
rect 106 11906 170 11970
rect 188 11906 252 11970
rect 270 11906 334 11970
rect 352 11906 416 11970
rect 434 11906 498 11970
rect 516 11906 580 11970
rect 598 11906 662 11970
rect 679 11906 743 11970
rect 760 11906 824 11970
rect 841 11906 905 11970
rect 922 11906 986 11970
rect 1003 11906 1067 11970
rect 1084 11906 1148 11970
rect 1165 11906 1229 11970
rect 1246 11906 1310 11970
rect 1327 11906 1391 11970
rect 1408 11906 1472 11970
rect 1489 11906 1553 11970
rect 1570 11906 1634 11970
rect 1651 11906 1715 11970
rect 1732 11906 1796 11970
rect 1813 11906 1877 11970
rect 1894 11906 1958 11970
rect 1975 11906 2039 11970
rect 2056 11906 2120 11970
rect 2137 11906 2201 11970
rect 2218 11906 2282 11970
rect 2299 11906 2363 11970
rect 2380 11906 2444 11970
rect 2461 11906 2525 11970
rect 2542 11906 2606 11970
rect 2623 11906 2687 11970
rect 2704 11906 2768 11970
rect 2785 11906 2849 11970
rect 2866 11906 2930 11970
rect 2947 11906 3011 11970
rect 3028 11906 3092 11970
rect 3109 11906 3173 11970
rect 3190 11906 3254 11970
rect 3271 11906 3335 11970
rect 3352 11906 3416 11970
rect 3433 11906 3497 11970
rect 3514 11906 3578 11970
rect 3595 11906 3659 11970
rect 3676 11906 3740 11970
rect 3757 11906 3821 11970
rect 3838 11906 3902 11970
rect 3919 11906 3983 11970
rect 4000 11906 4064 11970
rect 4081 11906 4145 11970
rect 4162 11906 4226 11970
rect 4243 11906 4307 11970
rect 4324 11906 4388 11970
rect 4405 11906 4469 11970
rect 4486 11906 4550 11970
rect 4567 11906 4631 11970
rect 4648 11906 4712 11970
rect 4729 11906 4793 11970
rect 4810 11906 4874 11970
rect 10157 11906 10221 11970
rect 10239 11906 10303 11970
rect 10321 11906 10385 11970
rect 10403 11906 10467 11970
rect 10485 11906 10549 11970
rect 10567 11906 10631 11970
rect 10649 11906 10713 11970
rect 10731 11906 10795 11970
rect 10813 11906 10877 11970
rect 10895 11906 10959 11970
rect 10977 11906 11041 11970
rect 11059 11906 11123 11970
rect 11141 11906 11205 11970
rect 11223 11906 11287 11970
rect 11305 11906 11369 11970
rect 11386 11906 11450 11970
rect 11467 11906 11531 11970
rect 11548 11906 11612 11970
rect 11629 11906 11693 11970
rect 11710 11906 11774 11970
rect 11791 11906 11855 11970
rect 11872 11906 11936 11970
rect 11953 11906 12017 11970
rect 12034 11906 12098 11970
rect 12115 11906 12179 11970
rect 12196 11906 12260 11970
rect 12277 11906 12341 11970
rect 12358 11906 12422 11970
rect 12439 11906 12503 11970
rect 12520 11906 12584 11970
rect 12601 11906 12665 11970
rect 12682 11906 12746 11970
rect 12763 11906 12827 11970
rect 12844 11906 12908 11970
rect 12925 11906 12989 11970
rect 13006 11906 13070 11970
rect 13087 11906 13151 11970
rect 13168 11906 13232 11970
rect 13249 11906 13313 11970
rect 13330 11906 13394 11970
rect 13411 11906 13475 11970
rect 13492 11906 13556 11970
rect 13573 11906 13637 11970
rect 13654 11906 13718 11970
rect 13735 11906 13799 11970
rect 13816 11906 13880 11970
rect 13897 11906 13961 11970
rect 13978 11906 14042 11970
rect 14059 11906 14123 11970
rect 14140 11906 14204 11970
rect 14221 11906 14285 11970
rect 14302 11906 14366 11970
rect 14383 11906 14447 11970
rect 14464 11906 14528 11970
rect 14545 11906 14609 11970
rect 14626 11906 14690 11970
rect 14707 11906 14771 11970
rect 14788 11906 14852 11970
rect 106 11824 170 11888
rect 188 11824 252 11888
rect 270 11824 334 11888
rect 352 11824 416 11888
rect 434 11824 498 11888
rect 516 11824 580 11888
rect 598 11824 662 11888
rect 679 11824 743 11888
rect 760 11824 824 11888
rect 841 11824 905 11888
rect 922 11824 986 11888
rect 1003 11824 1067 11888
rect 1084 11824 1148 11888
rect 1165 11824 1229 11888
rect 1246 11824 1310 11888
rect 1327 11824 1391 11888
rect 1408 11824 1472 11888
rect 1489 11824 1553 11888
rect 1570 11824 1634 11888
rect 1651 11824 1715 11888
rect 1732 11824 1796 11888
rect 1813 11824 1877 11888
rect 1894 11824 1958 11888
rect 1975 11824 2039 11888
rect 2056 11824 2120 11888
rect 2137 11824 2201 11888
rect 2218 11824 2282 11888
rect 2299 11824 2363 11888
rect 2380 11824 2444 11888
rect 2461 11824 2525 11888
rect 2542 11824 2606 11888
rect 2623 11824 2687 11888
rect 2704 11824 2768 11888
rect 2785 11824 2849 11888
rect 2866 11824 2930 11888
rect 2947 11824 3011 11888
rect 3028 11824 3092 11888
rect 3109 11824 3173 11888
rect 3190 11824 3254 11888
rect 3271 11824 3335 11888
rect 3352 11824 3416 11888
rect 3433 11824 3497 11888
rect 3514 11824 3578 11888
rect 3595 11824 3659 11888
rect 3676 11824 3740 11888
rect 3757 11824 3821 11888
rect 3838 11824 3902 11888
rect 3919 11824 3983 11888
rect 4000 11824 4064 11888
rect 4081 11824 4145 11888
rect 4162 11824 4226 11888
rect 4243 11824 4307 11888
rect 4324 11824 4388 11888
rect 4405 11824 4469 11888
rect 4486 11824 4550 11888
rect 4567 11824 4631 11888
rect 4648 11824 4712 11888
rect 4729 11824 4793 11888
rect 4810 11824 4874 11888
rect 10157 11824 10221 11888
rect 10239 11824 10303 11888
rect 10321 11824 10385 11888
rect 10403 11824 10467 11888
rect 10485 11824 10549 11888
rect 10567 11824 10631 11888
rect 10649 11824 10713 11888
rect 10731 11824 10795 11888
rect 10813 11824 10877 11888
rect 10895 11824 10959 11888
rect 10977 11824 11041 11888
rect 11059 11824 11123 11888
rect 11141 11824 11205 11888
rect 11223 11824 11287 11888
rect 11305 11824 11369 11888
rect 11386 11824 11450 11888
rect 11467 11824 11531 11888
rect 11548 11824 11612 11888
rect 11629 11824 11693 11888
rect 11710 11824 11774 11888
rect 11791 11824 11855 11888
rect 11872 11824 11936 11888
rect 11953 11824 12017 11888
rect 12034 11824 12098 11888
rect 12115 11824 12179 11888
rect 12196 11824 12260 11888
rect 12277 11824 12341 11888
rect 12358 11824 12422 11888
rect 12439 11824 12503 11888
rect 12520 11824 12584 11888
rect 12601 11824 12665 11888
rect 12682 11824 12746 11888
rect 12763 11824 12827 11888
rect 12844 11824 12908 11888
rect 12925 11824 12989 11888
rect 13006 11824 13070 11888
rect 13087 11824 13151 11888
rect 13168 11824 13232 11888
rect 13249 11824 13313 11888
rect 13330 11824 13394 11888
rect 13411 11824 13475 11888
rect 13492 11824 13556 11888
rect 13573 11824 13637 11888
rect 13654 11824 13718 11888
rect 13735 11824 13799 11888
rect 13816 11824 13880 11888
rect 13897 11824 13961 11888
rect 13978 11824 14042 11888
rect 14059 11824 14123 11888
rect 14140 11824 14204 11888
rect 14221 11824 14285 11888
rect 14302 11824 14366 11888
rect 14383 11824 14447 11888
rect 14464 11824 14528 11888
rect 14545 11824 14609 11888
rect 14626 11824 14690 11888
rect 14707 11824 14771 11888
rect 14788 11824 14852 11888
rect 106 11742 170 11806
rect 188 11742 252 11806
rect 270 11742 334 11806
rect 352 11742 416 11806
rect 434 11742 498 11806
rect 516 11742 580 11806
rect 598 11742 662 11806
rect 679 11742 743 11806
rect 760 11742 824 11806
rect 841 11742 905 11806
rect 922 11742 986 11806
rect 1003 11742 1067 11806
rect 1084 11742 1148 11806
rect 1165 11742 1229 11806
rect 1246 11742 1310 11806
rect 1327 11742 1391 11806
rect 1408 11742 1472 11806
rect 1489 11742 1553 11806
rect 1570 11742 1634 11806
rect 1651 11742 1715 11806
rect 1732 11742 1796 11806
rect 1813 11742 1877 11806
rect 1894 11742 1958 11806
rect 1975 11742 2039 11806
rect 2056 11742 2120 11806
rect 2137 11742 2201 11806
rect 2218 11742 2282 11806
rect 2299 11742 2363 11806
rect 2380 11742 2444 11806
rect 2461 11742 2525 11806
rect 2542 11742 2606 11806
rect 2623 11742 2687 11806
rect 2704 11742 2768 11806
rect 2785 11742 2849 11806
rect 2866 11742 2930 11806
rect 2947 11742 3011 11806
rect 3028 11742 3092 11806
rect 3109 11742 3173 11806
rect 3190 11742 3254 11806
rect 3271 11742 3335 11806
rect 3352 11742 3416 11806
rect 3433 11742 3497 11806
rect 3514 11742 3578 11806
rect 3595 11742 3659 11806
rect 3676 11742 3740 11806
rect 3757 11742 3821 11806
rect 3838 11742 3902 11806
rect 3919 11742 3983 11806
rect 4000 11742 4064 11806
rect 4081 11742 4145 11806
rect 4162 11742 4226 11806
rect 4243 11742 4307 11806
rect 4324 11742 4388 11806
rect 4405 11742 4469 11806
rect 4486 11742 4550 11806
rect 4567 11742 4631 11806
rect 4648 11742 4712 11806
rect 4729 11742 4793 11806
rect 4810 11742 4874 11806
rect 10157 11742 10221 11806
rect 10239 11742 10303 11806
rect 10321 11742 10385 11806
rect 10403 11742 10467 11806
rect 10485 11742 10549 11806
rect 10567 11742 10631 11806
rect 10649 11742 10713 11806
rect 10731 11742 10795 11806
rect 10813 11742 10877 11806
rect 10895 11742 10959 11806
rect 10977 11742 11041 11806
rect 11059 11742 11123 11806
rect 11141 11742 11205 11806
rect 11223 11742 11287 11806
rect 11305 11742 11369 11806
rect 11386 11742 11450 11806
rect 11467 11742 11531 11806
rect 11548 11742 11612 11806
rect 11629 11742 11693 11806
rect 11710 11742 11774 11806
rect 11791 11742 11855 11806
rect 11872 11742 11936 11806
rect 11953 11742 12017 11806
rect 12034 11742 12098 11806
rect 12115 11742 12179 11806
rect 12196 11742 12260 11806
rect 12277 11742 12341 11806
rect 12358 11742 12422 11806
rect 12439 11742 12503 11806
rect 12520 11742 12584 11806
rect 12601 11742 12665 11806
rect 12682 11742 12746 11806
rect 12763 11742 12827 11806
rect 12844 11742 12908 11806
rect 12925 11742 12989 11806
rect 13006 11742 13070 11806
rect 13087 11742 13151 11806
rect 13168 11742 13232 11806
rect 13249 11742 13313 11806
rect 13330 11742 13394 11806
rect 13411 11742 13475 11806
rect 13492 11742 13556 11806
rect 13573 11742 13637 11806
rect 13654 11742 13718 11806
rect 13735 11742 13799 11806
rect 13816 11742 13880 11806
rect 13897 11742 13961 11806
rect 13978 11742 14042 11806
rect 14059 11742 14123 11806
rect 14140 11742 14204 11806
rect 14221 11742 14285 11806
rect 14302 11742 14366 11806
rect 14383 11742 14447 11806
rect 14464 11742 14528 11806
rect 14545 11742 14609 11806
rect 14626 11742 14690 11806
rect 14707 11742 14771 11806
rect 14788 11742 14852 11806
rect 106 11660 170 11724
rect 188 11660 252 11724
rect 270 11660 334 11724
rect 352 11660 416 11724
rect 434 11660 498 11724
rect 516 11660 580 11724
rect 598 11660 662 11724
rect 679 11660 743 11724
rect 760 11660 824 11724
rect 841 11660 905 11724
rect 922 11660 986 11724
rect 1003 11660 1067 11724
rect 1084 11660 1148 11724
rect 1165 11660 1229 11724
rect 1246 11660 1310 11724
rect 1327 11660 1391 11724
rect 1408 11660 1472 11724
rect 1489 11660 1553 11724
rect 1570 11660 1634 11724
rect 1651 11660 1715 11724
rect 1732 11660 1796 11724
rect 1813 11660 1877 11724
rect 1894 11660 1958 11724
rect 1975 11660 2039 11724
rect 2056 11660 2120 11724
rect 2137 11660 2201 11724
rect 2218 11660 2282 11724
rect 2299 11660 2363 11724
rect 2380 11660 2444 11724
rect 2461 11660 2525 11724
rect 2542 11660 2606 11724
rect 2623 11660 2687 11724
rect 2704 11660 2768 11724
rect 2785 11660 2849 11724
rect 2866 11660 2930 11724
rect 2947 11660 3011 11724
rect 3028 11660 3092 11724
rect 3109 11660 3173 11724
rect 3190 11660 3254 11724
rect 3271 11660 3335 11724
rect 3352 11660 3416 11724
rect 3433 11660 3497 11724
rect 3514 11660 3578 11724
rect 3595 11660 3659 11724
rect 3676 11660 3740 11724
rect 3757 11660 3821 11724
rect 3838 11660 3902 11724
rect 3919 11660 3983 11724
rect 4000 11660 4064 11724
rect 4081 11660 4145 11724
rect 4162 11660 4226 11724
rect 4243 11660 4307 11724
rect 4324 11660 4388 11724
rect 4405 11660 4469 11724
rect 4486 11660 4550 11724
rect 4567 11660 4631 11724
rect 4648 11660 4712 11724
rect 4729 11660 4793 11724
rect 4810 11660 4874 11724
rect 10157 11660 10221 11724
rect 10239 11660 10303 11724
rect 10321 11660 10385 11724
rect 10403 11660 10467 11724
rect 10485 11660 10549 11724
rect 10567 11660 10631 11724
rect 10649 11660 10713 11724
rect 10731 11660 10795 11724
rect 10813 11660 10877 11724
rect 10895 11660 10959 11724
rect 10977 11660 11041 11724
rect 11059 11660 11123 11724
rect 11141 11660 11205 11724
rect 11223 11660 11287 11724
rect 11305 11660 11369 11724
rect 11386 11660 11450 11724
rect 11467 11660 11531 11724
rect 11548 11660 11612 11724
rect 11629 11660 11693 11724
rect 11710 11660 11774 11724
rect 11791 11660 11855 11724
rect 11872 11660 11936 11724
rect 11953 11660 12017 11724
rect 12034 11660 12098 11724
rect 12115 11660 12179 11724
rect 12196 11660 12260 11724
rect 12277 11660 12341 11724
rect 12358 11660 12422 11724
rect 12439 11660 12503 11724
rect 12520 11660 12584 11724
rect 12601 11660 12665 11724
rect 12682 11660 12746 11724
rect 12763 11660 12827 11724
rect 12844 11660 12908 11724
rect 12925 11660 12989 11724
rect 13006 11660 13070 11724
rect 13087 11660 13151 11724
rect 13168 11660 13232 11724
rect 13249 11660 13313 11724
rect 13330 11660 13394 11724
rect 13411 11660 13475 11724
rect 13492 11660 13556 11724
rect 13573 11660 13637 11724
rect 13654 11660 13718 11724
rect 13735 11660 13799 11724
rect 13816 11660 13880 11724
rect 13897 11660 13961 11724
rect 13978 11660 14042 11724
rect 14059 11660 14123 11724
rect 14140 11660 14204 11724
rect 14221 11660 14285 11724
rect 14302 11660 14366 11724
rect 14383 11660 14447 11724
rect 14464 11660 14528 11724
rect 14545 11660 14609 11724
rect 14626 11660 14690 11724
rect 14707 11660 14771 11724
rect 14788 11660 14852 11724
rect 106 11578 170 11642
rect 188 11578 252 11642
rect 270 11578 334 11642
rect 352 11578 416 11642
rect 434 11578 498 11642
rect 516 11578 580 11642
rect 598 11578 662 11642
rect 679 11578 743 11642
rect 760 11578 824 11642
rect 841 11578 905 11642
rect 922 11578 986 11642
rect 1003 11578 1067 11642
rect 1084 11578 1148 11642
rect 1165 11578 1229 11642
rect 1246 11578 1310 11642
rect 1327 11578 1391 11642
rect 1408 11578 1472 11642
rect 1489 11578 1553 11642
rect 1570 11578 1634 11642
rect 1651 11578 1715 11642
rect 1732 11578 1796 11642
rect 1813 11578 1877 11642
rect 1894 11578 1958 11642
rect 1975 11578 2039 11642
rect 2056 11578 2120 11642
rect 2137 11578 2201 11642
rect 2218 11578 2282 11642
rect 2299 11578 2363 11642
rect 2380 11578 2444 11642
rect 2461 11578 2525 11642
rect 2542 11578 2606 11642
rect 2623 11578 2687 11642
rect 2704 11578 2768 11642
rect 2785 11578 2849 11642
rect 2866 11578 2930 11642
rect 2947 11578 3011 11642
rect 3028 11578 3092 11642
rect 3109 11578 3173 11642
rect 3190 11578 3254 11642
rect 3271 11578 3335 11642
rect 3352 11578 3416 11642
rect 3433 11578 3497 11642
rect 3514 11578 3578 11642
rect 3595 11578 3659 11642
rect 3676 11578 3740 11642
rect 3757 11578 3821 11642
rect 3838 11578 3902 11642
rect 3919 11578 3983 11642
rect 4000 11578 4064 11642
rect 4081 11578 4145 11642
rect 4162 11578 4226 11642
rect 4243 11578 4307 11642
rect 4324 11578 4388 11642
rect 4405 11578 4469 11642
rect 4486 11578 4550 11642
rect 4567 11578 4631 11642
rect 4648 11578 4712 11642
rect 4729 11578 4793 11642
rect 4810 11578 4874 11642
rect 10157 11578 10221 11642
rect 10239 11578 10303 11642
rect 10321 11578 10385 11642
rect 10403 11578 10467 11642
rect 10485 11578 10549 11642
rect 10567 11578 10631 11642
rect 10649 11578 10713 11642
rect 10731 11578 10795 11642
rect 10813 11578 10877 11642
rect 10895 11578 10959 11642
rect 10977 11578 11041 11642
rect 11059 11578 11123 11642
rect 11141 11578 11205 11642
rect 11223 11578 11287 11642
rect 11305 11578 11369 11642
rect 11386 11578 11450 11642
rect 11467 11578 11531 11642
rect 11548 11578 11612 11642
rect 11629 11578 11693 11642
rect 11710 11578 11774 11642
rect 11791 11578 11855 11642
rect 11872 11578 11936 11642
rect 11953 11578 12017 11642
rect 12034 11578 12098 11642
rect 12115 11578 12179 11642
rect 12196 11578 12260 11642
rect 12277 11578 12341 11642
rect 12358 11578 12422 11642
rect 12439 11578 12503 11642
rect 12520 11578 12584 11642
rect 12601 11578 12665 11642
rect 12682 11578 12746 11642
rect 12763 11578 12827 11642
rect 12844 11578 12908 11642
rect 12925 11578 12989 11642
rect 13006 11578 13070 11642
rect 13087 11578 13151 11642
rect 13168 11578 13232 11642
rect 13249 11578 13313 11642
rect 13330 11578 13394 11642
rect 13411 11578 13475 11642
rect 13492 11578 13556 11642
rect 13573 11578 13637 11642
rect 13654 11578 13718 11642
rect 13735 11578 13799 11642
rect 13816 11578 13880 11642
rect 13897 11578 13961 11642
rect 13978 11578 14042 11642
rect 14059 11578 14123 11642
rect 14140 11578 14204 11642
rect 14221 11578 14285 11642
rect 14302 11578 14366 11642
rect 14383 11578 14447 11642
rect 14464 11578 14528 11642
rect 14545 11578 14609 11642
rect 14626 11578 14690 11642
rect 14707 11578 14771 11642
rect 14788 11578 14852 11642
rect 106 11496 170 11560
rect 188 11496 252 11560
rect 270 11496 334 11560
rect 352 11496 416 11560
rect 434 11496 498 11560
rect 516 11496 580 11560
rect 598 11496 662 11560
rect 679 11496 743 11560
rect 760 11496 824 11560
rect 841 11496 905 11560
rect 922 11496 986 11560
rect 1003 11496 1067 11560
rect 1084 11496 1148 11560
rect 1165 11496 1229 11560
rect 1246 11496 1310 11560
rect 1327 11496 1391 11560
rect 1408 11496 1472 11560
rect 1489 11496 1553 11560
rect 1570 11496 1634 11560
rect 1651 11496 1715 11560
rect 1732 11496 1796 11560
rect 1813 11496 1877 11560
rect 1894 11496 1958 11560
rect 1975 11496 2039 11560
rect 2056 11496 2120 11560
rect 2137 11496 2201 11560
rect 2218 11496 2282 11560
rect 2299 11496 2363 11560
rect 2380 11496 2444 11560
rect 2461 11496 2525 11560
rect 2542 11496 2606 11560
rect 2623 11496 2687 11560
rect 2704 11496 2768 11560
rect 2785 11496 2849 11560
rect 2866 11496 2930 11560
rect 2947 11496 3011 11560
rect 3028 11496 3092 11560
rect 3109 11496 3173 11560
rect 3190 11496 3254 11560
rect 3271 11496 3335 11560
rect 3352 11496 3416 11560
rect 3433 11496 3497 11560
rect 3514 11496 3578 11560
rect 3595 11496 3659 11560
rect 3676 11496 3740 11560
rect 3757 11496 3821 11560
rect 3838 11496 3902 11560
rect 3919 11496 3983 11560
rect 4000 11496 4064 11560
rect 4081 11496 4145 11560
rect 4162 11496 4226 11560
rect 4243 11496 4307 11560
rect 4324 11496 4388 11560
rect 4405 11496 4469 11560
rect 4486 11496 4550 11560
rect 4567 11496 4631 11560
rect 4648 11496 4712 11560
rect 4729 11496 4793 11560
rect 4810 11496 4874 11560
rect 10157 11496 10221 11560
rect 10239 11496 10303 11560
rect 10321 11496 10385 11560
rect 10403 11496 10467 11560
rect 10485 11496 10549 11560
rect 10567 11496 10631 11560
rect 10649 11496 10713 11560
rect 10731 11496 10795 11560
rect 10813 11496 10877 11560
rect 10895 11496 10959 11560
rect 10977 11496 11041 11560
rect 11059 11496 11123 11560
rect 11141 11496 11205 11560
rect 11223 11496 11287 11560
rect 11305 11496 11369 11560
rect 11386 11496 11450 11560
rect 11467 11496 11531 11560
rect 11548 11496 11612 11560
rect 11629 11496 11693 11560
rect 11710 11496 11774 11560
rect 11791 11496 11855 11560
rect 11872 11496 11936 11560
rect 11953 11496 12017 11560
rect 12034 11496 12098 11560
rect 12115 11496 12179 11560
rect 12196 11496 12260 11560
rect 12277 11496 12341 11560
rect 12358 11496 12422 11560
rect 12439 11496 12503 11560
rect 12520 11496 12584 11560
rect 12601 11496 12665 11560
rect 12682 11496 12746 11560
rect 12763 11496 12827 11560
rect 12844 11496 12908 11560
rect 12925 11496 12989 11560
rect 13006 11496 13070 11560
rect 13087 11496 13151 11560
rect 13168 11496 13232 11560
rect 13249 11496 13313 11560
rect 13330 11496 13394 11560
rect 13411 11496 13475 11560
rect 13492 11496 13556 11560
rect 13573 11496 13637 11560
rect 13654 11496 13718 11560
rect 13735 11496 13799 11560
rect 13816 11496 13880 11560
rect 13897 11496 13961 11560
rect 13978 11496 14042 11560
rect 14059 11496 14123 11560
rect 14140 11496 14204 11560
rect 14221 11496 14285 11560
rect 14302 11496 14366 11560
rect 14383 11496 14447 11560
rect 14464 11496 14528 11560
rect 14545 11496 14609 11560
rect 14626 11496 14690 11560
rect 14707 11496 14771 11560
rect 14788 11496 14852 11560
rect 106 11414 170 11478
rect 188 11414 252 11478
rect 270 11414 334 11478
rect 352 11414 416 11478
rect 434 11414 498 11478
rect 516 11414 580 11478
rect 598 11414 662 11478
rect 679 11414 743 11478
rect 760 11414 824 11478
rect 841 11414 905 11478
rect 922 11414 986 11478
rect 1003 11414 1067 11478
rect 1084 11414 1148 11478
rect 1165 11414 1229 11478
rect 1246 11414 1310 11478
rect 1327 11414 1391 11478
rect 1408 11414 1472 11478
rect 1489 11414 1553 11478
rect 1570 11414 1634 11478
rect 1651 11414 1715 11478
rect 1732 11414 1796 11478
rect 1813 11414 1877 11478
rect 1894 11414 1958 11478
rect 1975 11414 2039 11478
rect 2056 11414 2120 11478
rect 2137 11414 2201 11478
rect 2218 11414 2282 11478
rect 2299 11414 2363 11478
rect 2380 11414 2444 11478
rect 2461 11414 2525 11478
rect 2542 11414 2606 11478
rect 2623 11414 2687 11478
rect 2704 11414 2768 11478
rect 2785 11414 2849 11478
rect 2866 11414 2930 11478
rect 2947 11414 3011 11478
rect 3028 11414 3092 11478
rect 3109 11414 3173 11478
rect 3190 11414 3254 11478
rect 3271 11414 3335 11478
rect 3352 11414 3416 11478
rect 3433 11414 3497 11478
rect 3514 11414 3578 11478
rect 3595 11414 3659 11478
rect 3676 11414 3740 11478
rect 3757 11414 3821 11478
rect 3838 11414 3902 11478
rect 3919 11414 3983 11478
rect 4000 11414 4064 11478
rect 4081 11414 4145 11478
rect 4162 11414 4226 11478
rect 4243 11414 4307 11478
rect 4324 11414 4388 11478
rect 4405 11414 4469 11478
rect 4486 11414 4550 11478
rect 4567 11414 4631 11478
rect 4648 11414 4712 11478
rect 4729 11414 4793 11478
rect 4810 11414 4874 11478
rect 10157 11414 10221 11478
rect 10239 11414 10303 11478
rect 10321 11414 10385 11478
rect 10403 11414 10467 11478
rect 10485 11414 10549 11478
rect 10567 11414 10631 11478
rect 10649 11414 10713 11478
rect 10731 11414 10795 11478
rect 10813 11414 10877 11478
rect 10895 11414 10959 11478
rect 10977 11414 11041 11478
rect 11059 11414 11123 11478
rect 11141 11414 11205 11478
rect 11223 11414 11287 11478
rect 11305 11414 11369 11478
rect 11386 11414 11450 11478
rect 11467 11414 11531 11478
rect 11548 11414 11612 11478
rect 11629 11414 11693 11478
rect 11710 11414 11774 11478
rect 11791 11414 11855 11478
rect 11872 11414 11936 11478
rect 11953 11414 12017 11478
rect 12034 11414 12098 11478
rect 12115 11414 12179 11478
rect 12196 11414 12260 11478
rect 12277 11414 12341 11478
rect 12358 11414 12422 11478
rect 12439 11414 12503 11478
rect 12520 11414 12584 11478
rect 12601 11414 12665 11478
rect 12682 11414 12746 11478
rect 12763 11414 12827 11478
rect 12844 11414 12908 11478
rect 12925 11414 12989 11478
rect 13006 11414 13070 11478
rect 13087 11414 13151 11478
rect 13168 11414 13232 11478
rect 13249 11414 13313 11478
rect 13330 11414 13394 11478
rect 13411 11414 13475 11478
rect 13492 11414 13556 11478
rect 13573 11414 13637 11478
rect 13654 11414 13718 11478
rect 13735 11414 13799 11478
rect 13816 11414 13880 11478
rect 13897 11414 13961 11478
rect 13978 11414 14042 11478
rect 14059 11414 14123 11478
rect 14140 11414 14204 11478
rect 14221 11414 14285 11478
rect 14302 11414 14366 11478
rect 14383 11414 14447 11478
rect 14464 11414 14528 11478
rect 14545 11414 14609 11478
rect 14626 11414 14690 11478
rect 14707 11414 14771 11478
rect 14788 11414 14852 11478
rect 106 11332 170 11396
rect 188 11332 252 11396
rect 270 11332 334 11396
rect 352 11332 416 11396
rect 434 11332 498 11396
rect 516 11332 580 11396
rect 598 11332 662 11396
rect 679 11332 743 11396
rect 760 11332 824 11396
rect 841 11332 905 11396
rect 922 11332 986 11396
rect 1003 11332 1067 11396
rect 1084 11332 1148 11396
rect 1165 11332 1229 11396
rect 1246 11332 1310 11396
rect 1327 11332 1391 11396
rect 1408 11332 1472 11396
rect 1489 11332 1553 11396
rect 1570 11332 1634 11396
rect 1651 11332 1715 11396
rect 1732 11332 1796 11396
rect 1813 11332 1877 11396
rect 1894 11332 1958 11396
rect 1975 11332 2039 11396
rect 2056 11332 2120 11396
rect 2137 11332 2201 11396
rect 2218 11332 2282 11396
rect 2299 11332 2363 11396
rect 2380 11332 2444 11396
rect 2461 11332 2525 11396
rect 2542 11332 2606 11396
rect 2623 11332 2687 11396
rect 2704 11332 2768 11396
rect 2785 11332 2849 11396
rect 2866 11332 2930 11396
rect 2947 11332 3011 11396
rect 3028 11332 3092 11396
rect 3109 11332 3173 11396
rect 3190 11332 3254 11396
rect 3271 11332 3335 11396
rect 3352 11332 3416 11396
rect 3433 11332 3497 11396
rect 3514 11332 3578 11396
rect 3595 11332 3659 11396
rect 3676 11332 3740 11396
rect 3757 11332 3821 11396
rect 3838 11332 3902 11396
rect 3919 11332 3983 11396
rect 4000 11332 4064 11396
rect 4081 11332 4145 11396
rect 4162 11332 4226 11396
rect 4243 11332 4307 11396
rect 4324 11332 4388 11396
rect 4405 11332 4469 11396
rect 4486 11332 4550 11396
rect 4567 11332 4631 11396
rect 4648 11332 4712 11396
rect 4729 11332 4793 11396
rect 4810 11332 4874 11396
rect 10157 11332 10221 11396
rect 10239 11332 10303 11396
rect 10321 11332 10385 11396
rect 10403 11332 10467 11396
rect 10485 11332 10549 11396
rect 10567 11332 10631 11396
rect 10649 11332 10713 11396
rect 10731 11332 10795 11396
rect 10813 11332 10877 11396
rect 10895 11332 10959 11396
rect 10977 11332 11041 11396
rect 11059 11332 11123 11396
rect 11141 11332 11205 11396
rect 11223 11332 11287 11396
rect 11305 11332 11369 11396
rect 11386 11332 11450 11396
rect 11467 11332 11531 11396
rect 11548 11332 11612 11396
rect 11629 11332 11693 11396
rect 11710 11332 11774 11396
rect 11791 11332 11855 11396
rect 11872 11332 11936 11396
rect 11953 11332 12017 11396
rect 12034 11332 12098 11396
rect 12115 11332 12179 11396
rect 12196 11332 12260 11396
rect 12277 11332 12341 11396
rect 12358 11332 12422 11396
rect 12439 11332 12503 11396
rect 12520 11332 12584 11396
rect 12601 11332 12665 11396
rect 12682 11332 12746 11396
rect 12763 11332 12827 11396
rect 12844 11332 12908 11396
rect 12925 11332 12989 11396
rect 13006 11332 13070 11396
rect 13087 11332 13151 11396
rect 13168 11332 13232 11396
rect 13249 11332 13313 11396
rect 13330 11332 13394 11396
rect 13411 11332 13475 11396
rect 13492 11332 13556 11396
rect 13573 11332 13637 11396
rect 13654 11332 13718 11396
rect 13735 11332 13799 11396
rect 13816 11332 13880 11396
rect 13897 11332 13961 11396
rect 13978 11332 14042 11396
rect 14059 11332 14123 11396
rect 14140 11332 14204 11396
rect 14221 11332 14285 11396
rect 14302 11332 14366 11396
rect 14383 11332 14447 11396
rect 14464 11332 14528 11396
rect 14545 11332 14609 11396
rect 14626 11332 14690 11396
rect 14707 11332 14771 11396
rect 14788 11332 14852 11396
rect 106 11250 170 11314
rect 188 11250 252 11314
rect 270 11250 334 11314
rect 352 11250 416 11314
rect 434 11250 498 11314
rect 516 11250 580 11314
rect 598 11250 662 11314
rect 679 11250 743 11314
rect 760 11250 824 11314
rect 841 11250 905 11314
rect 922 11250 986 11314
rect 1003 11250 1067 11314
rect 1084 11250 1148 11314
rect 1165 11250 1229 11314
rect 1246 11250 1310 11314
rect 1327 11250 1391 11314
rect 1408 11250 1472 11314
rect 1489 11250 1553 11314
rect 1570 11250 1634 11314
rect 1651 11250 1715 11314
rect 1732 11250 1796 11314
rect 1813 11250 1877 11314
rect 1894 11250 1958 11314
rect 1975 11250 2039 11314
rect 2056 11250 2120 11314
rect 2137 11250 2201 11314
rect 2218 11250 2282 11314
rect 2299 11250 2363 11314
rect 2380 11250 2444 11314
rect 2461 11250 2525 11314
rect 2542 11250 2606 11314
rect 2623 11250 2687 11314
rect 2704 11250 2768 11314
rect 2785 11250 2849 11314
rect 2866 11250 2930 11314
rect 2947 11250 3011 11314
rect 3028 11250 3092 11314
rect 3109 11250 3173 11314
rect 3190 11250 3254 11314
rect 3271 11250 3335 11314
rect 3352 11250 3416 11314
rect 3433 11250 3497 11314
rect 3514 11250 3578 11314
rect 3595 11250 3659 11314
rect 3676 11250 3740 11314
rect 3757 11250 3821 11314
rect 3838 11250 3902 11314
rect 3919 11250 3983 11314
rect 4000 11250 4064 11314
rect 4081 11250 4145 11314
rect 4162 11250 4226 11314
rect 4243 11250 4307 11314
rect 4324 11250 4388 11314
rect 4405 11250 4469 11314
rect 4486 11250 4550 11314
rect 4567 11250 4631 11314
rect 4648 11250 4712 11314
rect 4729 11250 4793 11314
rect 4810 11250 4874 11314
rect 10157 11250 10221 11314
rect 10239 11250 10303 11314
rect 10321 11250 10385 11314
rect 10403 11250 10467 11314
rect 10485 11250 10549 11314
rect 10567 11250 10631 11314
rect 10649 11250 10713 11314
rect 10731 11250 10795 11314
rect 10813 11250 10877 11314
rect 10895 11250 10959 11314
rect 10977 11250 11041 11314
rect 11059 11250 11123 11314
rect 11141 11250 11205 11314
rect 11223 11250 11287 11314
rect 11305 11250 11369 11314
rect 11386 11250 11450 11314
rect 11467 11250 11531 11314
rect 11548 11250 11612 11314
rect 11629 11250 11693 11314
rect 11710 11250 11774 11314
rect 11791 11250 11855 11314
rect 11872 11250 11936 11314
rect 11953 11250 12017 11314
rect 12034 11250 12098 11314
rect 12115 11250 12179 11314
rect 12196 11250 12260 11314
rect 12277 11250 12341 11314
rect 12358 11250 12422 11314
rect 12439 11250 12503 11314
rect 12520 11250 12584 11314
rect 12601 11250 12665 11314
rect 12682 11250 12746 11314
rect 12763 11250 12827 11314
rect 12844 11250 12908 11314
rect 12925 11250 12989 11314
rect 13006 11250 13070 11314
rect 13087 11250 13151 11314
rect 13168 11250 13232 11314
rect 13249 11250 13313 11314
rect 13330 11250 13394 11314
rect 13411 11250 13475 11314
rect 13492 11250 13556 11314
rect 13573 11250 13637 11314
rect 13654 11250 13718 11314
rect 13735 11250 13799 11314
rect 13816 11250 13880 11314
rect 13897 11250 13961 11314
rect 13978 11250 14042 11314
rect 14059 11250 14123 11314
rect 14140 11250 14204 11314
rect 14221 11250 14285 11314
rect 14302 11250 14366 11314
rect 14383 11250 14447 11314
rect 14464 11250 14528 11314
rect 14545 11250 14609 11314
rect 14626 11250 14690 11314
rect 14707 11250 14771 11314
rect 14788 11250 14852 11314
rect 0 10225 15000 10821
rect 0 9273 15000 9869
rect 106 5630 170 5694
rect 188 5630 252 5694
rect 270 5630 334 5694
rect 352 5630 416 5694
rect 434 5630 498 5694
rect 516 5630 580 5694
rect 598 5630 662 5694
rect 679 5630 743 5694
rect 760 5630 824 5694
rect 841 5630 905 5694
rect 922 5630 986 5694
rect 1003 5630 1067 5694
rect 1084 5630 1148 5694
rect 1165 5630 1229 5694
rect 1246 5630 1310 5694
rect 1327 5630 1391 5694
rect 1408 5630 1472 5694
rect 1489 5630 1553 5694
rect 1570 5630 1634 5694
rect 1651 5630 1715 5694
rect 1732 5630 1796 5694
rect 1813 5630 1877 5694
rect 1894 5630 1958 5694
rect 1975 5630 2039 5694
rect 2056 5630 2120 5694
rect 2137 5630 2201 5694
rect 2218 5630 2282 5694
rect 2299 5630 2363 5694
rect 2380 5630 2444 5694
rect 2461 5630 2525 5694
rect 2542 5630 2606 5694
rect 2623 5630 2687 5694
rect 2704 5630 2768 5694
rect 2785 5630 2849 5694
rect 2866 5630 2930 5694
rect 2947 5630 3011 5694
rect 3028 5630 3092 5694
rect 3109 5630 3173 5694
rect 3190 5630 3254 5694
rect 3271 5630 3335 5694
rect 3352 5630 3416 5694
rect 3433 5630 3497 5694
rect 3514 5630 3578 5694
rect 3595 5630 3659 5694
rect 3676 5630 3740 5694
rect 3757 5630 3821 5694
rect 3838 5630 3902 5694
rect 3919 5630 3983 5694
rect 4000 5630 4064 5694
rect 4081 5630 4145 5694
rect 4162 5630 4226 5694
rect 4243 5630 4307 5694
rect 4324 5630 4388 5694
rect 4405 5630 4469 5694
rect 4486 5630 4550 5694
rect 4567 5630 4631 5694
rect 4648 5630 4712 5694
rect 4729 5630 4793 5694
rect 4810 5630 4874 5694
rect 10157 5630 10221 5694
rect 10239 5630 10303 5694
rect 10321 5630 10385 5694
rect 10403 5630 10467 5694
rect 10485 5630 10549 5694
rect 10567 5630 10631 5694
rect 10649 5630 10713 5694
rect 10731 5630 10795 5694
rect 10813 5630 10877 5694
rect 10895 5630 10959 5694
rect 10977 5630 11041 5694
rect 11059 5630 11123 5694
rect 11141 5630 11205 5694
rect 11223 5630 11287 5694
rect 11305 5630 11369 5694
rect 11386 5630 11450 5694
rect 11467 5630 11531 5694
rect 11548 5630 11612 5694
rect 11629 5630 11693 5694
rect 11710 5630 11774 5694
rect 11791 5630 11855 5694
rect 11872 5630 11936 5694
rect 11953 5630 12017 5694
rect 12034 5630 12098 5694
rect 12115 5630 12179 5694
rect 12196 5630 12260 5694
rect 12277 5630 12341 5694
rect 12358 5630 12422 5694
rect 12439 5630 12503 5694
rect 12520 5630 12584 5694
rect 12601 5630 12665 5694
rect 12682 5630 12746 5694
rect 12763 5630 12827 5694
rect 12844 5630 12908 5694
rect 12925 5630 12989 5694
rect 13006 5630 13070 5694
rect 13087 5630 13151 5694
rect 13168 5630 13232 5694
rect 13249 5630 13313 5694
rect 13330 5630 13394 5694
rect 13411 5630 13475 5694
rect 13492 5630 13556 5694
rect 13573 5630 13637 5694
rect 13654 5630 13718 5694
rect 13735 5630 13799 5694
rect 13816 5630 13880 5694
rect 13897 5630 13961 5694
rect 13978 5630 14042 5694
rect 14059 5630 14123 5694
rect 14140 5630 14204 5694
rect 14221 5630 14285 5694
rect 14302 5630 14366 5694
rect 14383 5630 14447 5694
rect 14464 5630 14528 5694
rect 14545 5630 14609 5694
rect 14626 5630 14690 5694
rect 14707 5630 14771 5694
rect 14788 5630 14852 5694
rect 106 5544 170 5608
rect 188 5544 252 5608
rect 270 5544 334 5608
rect 352 5544 416 5608
rect 434 5544 498 5608
rect 516 5544 580 5608
rect 598 5544 662 5608
rect 679 5544 743 5608
rect 760 5544 824 5608
rect 841 5544 905 5608
rect 922 5544 986 5608
rect 1003 5544 1067 5608
rect 1084 5544 1148 5608
rect 1165 5544 1229 5608
rect 1246 5544 1310 5608
rect 1327 5544 1391 5608
rect 1408 5544 1472 5608
rect 1489 5544 1553 5608
rect 1570 5544 1634 5608
rect 1651 5544 1715 5608
rect 1732 5544 1796 5608
rect 1813 5544 1877 5608
rect 1894 5544 1958 5608
rect 1975 5544 2039 5608
rect 2056 5544 2120 5608
rect 2137 5544 2201 5608
rect 2218 5544 2282 5608
rect 2299 5544 2363 5608
rect 2380 5544 2444 5608
rect 2461 5544 2525 5608
rect 2542 5544 2606 5608
rect 2623 5544 2687 5608
rect 2704 5544 2768 5608
rect 2785 5544 2849 5608
rect 2866 5544 2930 5608
rect 2947 5544 3011 5608
rect 3028 5544 3092 5608
rect 3109 5544 3173 5608
rect 3190 5544 3254 5608
rect 3271 5544 3335 5608
rect 3352 5544 3416 5608
rect 3433 5544 3497 5608
rect 3514 5544 3578 5608
rect 3595 5544 3659 5608
rect 3676 5544 3740 5608
rect 3757 5544 3821 5608
rect 3838 5544 3902 5608
rect 3919 5544 3983 5608
rect 4000 5544 4064 5608
rect 4081 5544 4145 5608
rect 4162 5544 4226 5608
rect 4243 5544 4307 5608
rect 4324 5544 4388 5608
rect 4405 5544 4469 5608
rect 4486 5544 4550 5608
rect 4567 5544 4631 5608
rect 4648 5544 4712 5608
rect 4729 5544 4793 5608
rect 4810 5544 4874 5608
rect 10157 5544 10221 5608
rect 10239 5544 10303 5608
rect 10321 5544 10385 5608
rect 10403 5544 10467 5608
rect 10485 5544 10549 5608
rect 10567 5544 10631 5608
rect 10649 5544 10713 5608
rect 10731 5544 10795 5608
rect 10813 5544 10877 5608
rect 10895 5544 10959 5608
rect 10977 5544 11041 5608
rect 11059 5544 11123 5608
rect 11141 5544 11205 5608
rect 11223 5544 11287 5608
rect 11305 5544 11369 5608
rect 11386 5544 11450 5608
rect 11467 5544 11531 5608
rect 11548 5544 11612 5608
rect 11629 5544 11693 5608
rect 11710 5544 11774 5608
rect 11791 5544 11855 5608
rect 11872 5544 11936 5608
rect 11953 5544 12017 5608
rect 12034 5544 12098 5608
rect 12115 5544 12179 5608
rect 12196 5544 12260 5608
rect 12277 5544 12341 5608
rect 12358 5544 12422 5608
rect 12439 5544 12503 5608
rect 12520 5544 12584 5608
rect 12601 5544 12665 5608
rect 12682 5544 12746 5608
rect 12763 5544 12827 5608
rect 12844 5544 12908 5608
rect 12925 5544 12989 5608
rect 13006 5544 13070 5608
rect 13087 5544 13151 5608
rect 13168 5544 13232 5608
rect 13249 5544 13313 5608
rect 13330 5544 13394 5608
rect 13411 5544 13475 5608
rect 13492 5544 13556 5608
rect 13573 5544 13637 5608
rect 13654 5544 13718 5608
rect 13735 5544 13799 5608
rect 13816 5544 13880 5608
rect 13897 5544 13961 5608
rect 13978 5544 14042 5608
rect 14059 5544 14123 5608
rect 14140 5544 14204 5608
rect 14221 5544 14285 5608
rect 14302 5544 14366 5608
rect 14383 5544 14447 5608
rect 14464 5544 14528 5608
rect 14545 5544 14609 5608
rect 14626 5544 14690 5608
rect 14707 5544 14771 5608
rect 14788 5544 14852 5608
rect 106 5458 170 5522
rect 188 5458 252 5522
rect 270 5458 334 5522
rect 352 5458 416 5522
rect 434 5458 498 5522
rect 516 5458 580 5522
rect 598 5458 662 5522
rect 679 5458 743 5522
rect 760 5458 824 5522
rect 841 5458 905 5522
rect 922 5458 986 5522
rect 1003 5458 1067 5522
rect 1084 5458 1148 5522
rect 1165 5458 1229 5522
rect 1246 5458 1310 5522
rect 1327 5458 1391 5522
rect 1408 5458 1472 5522
rect 1489 5458 1553 5522
rect 1570 5458 1634 5522
rect 1651 5458 1715 5522
rect 1732 5458 1796 5522
rect 1813 5458 1877 5522
rect 1894 5458 1958 5522
rect 1975 5458 2039 5522
rect 2056 5458 2120 5522
rect 2137 5458 2201 5522
rect 2218 5458 2282 5522
rect 2299 5458 2363 5522
rect 2380 5458 2444 5522
rect 2461 5458 2525 5522
rect 2542 5458 2606 5522
rect 2623 5458 2687 5522
rect 2704 5458 2768 5522
rect 2785 5458 2849 5522
rect 2866 5458 2930 5522
rect 2947 5458 3011 5522
rect 3028 5458 3092 5522
rect 3109 5458 3173 5522
rect 3190 5458 3254 5522
rect 3271 5458 3335 5522
rect 3352 5458 3416 5522
rect 3433 5458 3497 5522
rect 3514 5458 3578 5522
rect 3595 5458 3659 5522
rect 3676 5458 3740 5522
rect 3757 5458 3821 5522
rect 3838 5458 3902 5522
rect 3919 5458 3983 5522
rect 4000 5458 4064 5522
rect 4081 5458 4145 5522
rect 4162 5458 4226 5522
rect 4243 5458 4307 5522
rect 4324 5458 4388 5522
rect 4405 5458 4469 5522
rect 4486 5458 4550 5522
rect 4567 5458 4631 5522
rect 4648 5458 4712 5522
rect 4729 5458 4793 5522
rect 4810 5458 4874 5522
rect 10157 5458 10221 5522
rect 10239 5458 10303 5522
rect 10321 5458 10385 5522
rect 10403 5458 10467 5522
rect 10485 5458 10549 5522
rect 10567 5458 10631 5522
rect 10649 5458 10713 5522
rect 10731 5458 10795 5522
rect 10813 5458 10877 5522
rect 10895 5458 10959 5522
rect 10977 5458 11041 5522
rect 11059 5458 11123 5522
rect 11141 5458 11205 5522
rect 11223 5458 11287 5522
rect 11305 5458 11369 5522
rect 11386 5458 11450 5522
rect 11467 5458 11531 5522
rect 11548 5458 11612 5522
rect 11629 5458 11693 5522
rect 11710 5458 11774 5522
rect 11791 5458 11855 5522
rect 11872 5458 11936 5522
rect 11953 5458 12017 5522
rect 12034 5458 12098 5522
rect 12115 5458 12179 5522
rect 12196 5458 12260 5522
rect 12277 5458 12341 5522
rect 12358 5458 12422 5522
rect 12439 5458 12503 5522
rect 12520 5458 12584 5522
rect 12601 5458 12665 5522
rect 12682 5458 12746 5522
rect 12763 5458 12827 5522
rect 12844 5458 12908 5522
rect 12925 5458 12989 5522
rect 13006 5458 13070 5522
rect 13087 5458 13151 5522
rect 13168 5458 13232 5522
rect 13249 5458 13313 5522
rect 13330 5458 13394 5522
rect 13411 5458 13475 5522
rect 13492 5458 13556 5522
rect 13573 5458 13637 5522
rect 13654 5458 13718 5522
rect 13735 5458 13799 5522
rect 13816 5458 13880 5522
rect 13897 5458 13961 5522
rect 13978 5458 14042 5522
rect 14059 5458 14123 5522
rect 14140 5458 14204 5522
rect 14221 5458 14285 5522
rect 14302 5458 14366 5522
rect 14383 5458 14447 5522
rect 14464 5458 14528 5522
rect 14545 5458 14609 5522
rect 14626 5458 14690 5522
rect 14707 5458 14771 5522
rect 14788 5458 14852 5522
rect 106 5372 170 5436
rect 188 5372 252 5436
rect 270 5372 334 5436
rect 352 5372 416 5436
rect 434 5372 498 5436
rect 516 5372 580 5436
rect 598 5372 662 5436
rect 679 5372 743 5436
rect 760 5372 824 5436
rect 841 5372 905 5436
rect 922 5372 986 5436
rect 1003 5372 1067 5436
rect 1084 5372 1148 5436
rect 1165 5372 1229 5436
rect 1246 5372 1310 5436
rect 1327 5372 1391 5436
rect 1408 5372 1472 5436
rect 1489 5372 1553 5436
rect 1570 5372 1634 5436
rect 1651 5372 1715 5436
rect 1732 5372 1796 5436
rect 1813 5372 1877 5436
rect 1894 5372 1958 5436
rect 1975 5372 2039 5436
rect 2056 5372 2120 5436
rect 2137 5372 2201 5436
rect 2218 5372 2282 5436
rect 2299 5372 2363 5436
rect 2380 5372 2444 5436
rect 2461 5372 2525 5436
rect 2542 5372 2606 5436
rect 2623 5372 2687 5436
rect 2704 5372 2768 5436
rect 2785 5372 2849 5436
rect 2866 5372 2930 5436
rect 2947 5372 3011 5436
rect 3028 5372 3092 5436
rect 3109 5372 3173 5436
rect 3190 5372 3254 5436
rect 3271 5372 3335 5436
rect 3352 5372 3416 5436
rect 3433 5372 3497 5436
rect 3514 5372 3578 5436
rect 3595 5372 3659 5436
rect 3676 5372 3740 5436
rect 3757 5372 3821 5436
rect 3838 5372 3902 5436
rect 3919 5372 3983 5436
rect 4000 5372 4064 5436
rect 4081 5372 4145 5436
rect 4162 5372 4226 5436
rect 4243 5372 4307 5436
rect 4324 5372 4388 5436
rect 4405 5372 4469 5436
rect 4486 5372 4550 5436
rect 4567 5372 4631 5436
rect 4648 5372 4712 5436
rect 4729 5372 4793 5436
rect 4810 5372 4874 5436
rect 10157 5372 10221 5436
rect 10239 5372 10303 5436
rect 10321 5372 10385 5436
rect 10403 5372 10467 5436
rect 10485 5372 10549 5436
rect 10567 5372 10631 5436
rect 10649 5372 10713 5436
rect 10731 5372 10795 5436
rect 10813 5372 10877 5436
rect 10895 5372 10959 5436
rect 10977 5372 11041 5436
rect 11059 5372 11123 5436
rect 11141 5372 11205 5436
rect 11223 5372 11287 5436
rect 11305 5372 11369 5436
rect 11386 5372 11450 5436
rect 11467 5372 11531 5436
rect 11548 5372 11612 5436
rect 11629 5372 11693 5436
rect 11710 5372 11774 5436
rect 11791 5372 11855 5436
rect 11872 5372 11936 5436
rect 11953 5372 12017 5436
rect 12034 5372 12098 5436
rect 12115 5372 12179 5436
rect 12196 5372 12260 5436
rect 12277 5372 12341 5436
rect 12358 5372 12422 5436
rect 12439 5372 12503 5436
rect 12520 5372 12584 5436
rect 12601 5372 12665 5436
rect 12682 5372 12746 5436
rect 12763 5372 12827 5436
rect 12844 5372 12908 5436
rect 12925 5372 12989 5436
rect 13006 5372 13070 5436
rect 13087 5372 13151 5436
rect 13168 5372 13232 5436
rect 13249 5372 13313 5436
rect 13330 5372 13394 5436
rect 13411 5372 13475 5436
rect 13492 5372 13556 5436
rect 13573 5372 13637 5436
rect 13654 5372 13718 5436
rect 13735 5372 13799 5436
rect 13816 5372 13880 5436
rect 13897 5372 13961 5436
rect 13978 5372 14042 5436
rect 14059 5372 14123 5436
rect 14140 5372 14204 5436
rect 14221 5372 14285 5436
rect 14302 5372 14366 5436
rect 14383 5372 14447 5436
rect 14464 5372 14528 5436
rect 14545 5372 14609 5436
rect 14626 5372 14690 5436
rect 14707 5372 14771 5436
rect 14788 5372 14852 5436
rect 106 5286 170 5350
rect 188 5286 252 5350
rect 270 5286 334 5350
rect 352 5286 416 5350
rect 434 5286 498 5350
rect 516 5286 580 5350
rect 598 5286 662 5350
rect 679 5286 743 5350
rect 760 5286 824 5350
rect 841 5286 905 5350
rect 922 5286 986 5350
rect 1003 5286 1067 5350
rect 1084 5286 1148 5350
rect 1165 5286 1229 5350
rect 1246 5286 1310 5350
rect 1327 5286 1391 5350
rect 1408 5286 1472 5350
rect 1489 5286 1553 5350
rect 1570 5286 1634 5350
rect 1651 5286 1715 5350
rect 1732 5286 1796 5350
rect 1813 5286 1877 5350
rect 1894 5286 1958 5350
rect 1975 5286 2039 5350
rect 2056 5286 2120 5350
rect 2137 5286 2201 5350
rect 2218 5286 2282 5350
rect 2299 5286 2363 5350
rect 2380 5286 2444 5350
rect 2461 5286 2525 5350
rect 2542 5286 2606 5350
rect 2623 5286 2687 5350
rect 2704 5286 2768 5350
rect 2785 5286 2849 5350
rect 2866 5286 2930 5350
rect 2947 5286 3011 5350
rect 3028 5286 3092 5350
rect 3109 5286 3173 5350
rect 3190 5286 3254 5350
rect 3271 5286 3335 5350
rect 3352 5286 3416 5350
rect 3433 5286 3497 5350
rect 3514 5286 3578 5350
rect 3595 5286 3659 5350
rect 3676 5286 3740 5350
rect 3757 5286 3821 5350
rect 3838 5286 3902 5350
rect 3919 5286 3983 5350
rect 4000 5286 4064 5350
rect 4081 5286 4145 5350
rect 4162 5286 4226 5350
rect 4243 5286 4307 5350
rect 4324 5286 4388 5350
rect 4405 5286 4469 5350
rect 4486 5286 4550 5350
rect 4567 5286 4631 5350
rect 4648 5286 4712 5350
rect 4729 5286 4793 5350
rect 4810 5286 4874 5350
rect 10157 5286 10221 5350
rect 10239 5286 10303 5350
rect 10321 5286 10385 5350
rect 10403 5286 10467 5350
rect 10485 5286 10549 5350
rect 10567 5286 10631 5350
rect 10649 5286 10713 5350
rect 10731 5286 10795 5350
rect 10813 5286 10877 5350
rect 10895 5286 10959 5350
rect 10977 5286 11041 5350
rect 11059 5286 11123 5350
rect 11141 5286 11205 5350
rect 11223 5286 11287 5350
rect 11305 5286 11369 5350
rect 11386 5286 11450 5350
rect 11467 5286 11531 5350
rect 11548 5286 11612 5350
rect 11629 5286 11693 5350
rect 11710 5286 11774 5350
rect 11791 5286 11855 5350
rect 11872 5286 11936 5350
rect 11953 5286 12017 5350
rect 12034 5286 12098 5350
rect 12115 5286 12179 5350
rect 12196 5286 12260 5350
rect 12277 5286 12341 5350
rect 12358 5286 12422 5350
rect 12439 5286 12503 5350
rect 12520 5286 12584 5350
rect 12601 5286 12665 5350
rect 12682 5286 12746 5350
rect 12763 5286 12827 5350
rect 12844 5286 12908 5350
rect 12925 5286 12989 5350
rect 13006 5286 13070 5350
rect 13087 5286 13151 5350
rect 13168 5286 13232 5350
rect 13249 5286 13313 5350
rect 13330 5286 13394 5350
rect 13411 5286 13475 5350
rect 13492 5286 13556 5350
rect 13573 5286 13637 5350
rect 13654 5286 13718 5350
rect 13735 5286 13799 5350
rect 13816 5286 13880 5350
rect 13897 5286 13961 5350
rect 13978 5286 14042 5350
rect 14059 5286 14123 5350
rect 14140 5286 14204 5350
rect 14221 5286 14285 5350
rect 14302 5286 14366 5350
rect 14383 5286 14447 5350
rect 14464 5286 14528 5350
rect 14545 5286 14609 5350
rect 14626 5286 14690 5350
rect 14707 5286 14771 5350
rect 14788 5286 14852 5350
rect 106 5200 170 5264
rect 188 5200 252 5264
rect 270 5200 334 5264
rect 352 5200 416 5264
rect 434 5200 498 5264
rect 516 5200 580 5264
rect 598 5200 662 5264
rect 679 5200 743 5264
rect 760 5200 824 5264
rect 841 5200 905 5264
rect 922 5200 986 5264
rect 1003 5200 1067 5264
rect 1084 5200 1148 5264
rect 1165 5200 1229 5264
rect 1246 5200 1310 5264
rect 1327 5200 1391 5264
rect 1408 5200 1472 5264
rect 1489 5200 1553 5264
rect 1570 5200 1634 5264
rect 1651 5200 1715 5264
rect 1732 5200 1796 5264
rect 1813 5200 1877 5264
rect 1894 5200 1958 5264
rect 1975 5200 2039 5264
rect 2056 5200 2120 5264
rect 2137 5200 2201 5264
rect 2218 5200 2282 5264
rect 2299 5200 2363 5264
rect 2380 5200 2444 5264
rect 2461 5200 2525 5264
rect 2542 5200 2606 5264
rect 2623 5200 2687 5264
rect 2704 5200 2768 5264
rect 2785 5200 2849 5264
rect 2866 5200 2930 5264
rect 2947 5200 3011 5264
rect 3028 5200 3092 5264
rect 3109 5200 3173 5264
rect 3190 5200 3254 5264
rect 3271 5200 3335 5264
rect 3352 5200 3416 5264
rect 3433 5200 3497 5264
rect 3514 5200 3578 5264
rect 3595 5200 3659 5264
rect 3676 5200 3740 5264
rect 3757 5200 3821 5264
rect 3838 5200 3902 5264
rect 3919 5200 3983 5264
rect 4000 5200 4064 5264
rect 4081 5200 4145 5264
rect 4162 5200 4226 5264
rect 4243 5200 4307 5264
rect 4324 5200 4388 5264
rect 4405 5200 4469 5264
rect 4486 5200 4550 5264
rect 4567 5200 4631 5264
rect 4648 5200 4712 5264
rect 4729 5200 4793 5264
rect 4810 5200 4874 5264
rect 10157 5200 10221 5264
rect 10239 5200 10303 5264
rect 10321 5200 10385 5264
rect 10403 5200 10467 5264
rect 10485 5200 10549 5264
rect 10567 5200 10631 5264
rect 10649 5200 10713 5264
rect 10731 5200 10795 5264
rect 10813 5200 10877 5264
rect 10895 5200 10959 5264
rect 10977 5200 11041 5264
rect 11059 5200 11123 5264
rect 11141 5200 11205 5264
rect 11223 5200 11287 5264
rect 11305 5200 11369 5264
rect 11386 5200 11450 5264
rect 11467 5200 11531 5264
rect 11548 5200 11612 5264
rect 11629 5200 11693 5264
rect 11710 5200 11774 5264
rect 11791 5200 11855 5264
rect 11872 5200 11936 5264
rect 11953 5200 12017 5264
rect 12034 5200 12098 5264
rect 12115 5200 12179 5264
rect 12196 5200 12260 5264
rect 12277 5200 12341 5264
rect 12358 5200 12422 5264
rect 12439 5200 12503 5264
rect 12520 5200 12584 5264
rect 12601 5200 12665 5264
rect 12682 5200 12746 5264
rect 12763 5200 12827 5264
rect 12844 5200 12908 5264
rect 12925 5200 12989 5264
rect 13006 5200 13070 5264
rect 13087 5200 13151 5264
rect 13168 5200 13232 5264
rect 13249 5200 13313 5264
rect 13330 5200 13394 5264
rect 13411 5200 13475 5264
rect 13492 5200 13556 5264
rect 13573 5200 13637 5264
rect 13654 5200 13718 5264
rect 13735 5200 13799 5264
rect 13816 5200 13880 5264
rect 13897 5200 13961 5264
rect 13978 5200 14042 5264
rect 14059 5200 14123 5264
rect 14140 5200 14204 5264
rect 14221 5200 14285 5264
rect 14302 5200 14366 5264
rect 14383 5200 14447 5264
rect 14464 5200 14528 5264
rect 14545 5200 14609 5264
rect 14626 5200 14690 5264
rect 14707 5200 14771 5264
rect 14788 5200 14852 5264
rect 106 5114 170 5178
rect 188 5114 252 5178
rect 270 5114 334 5178
rect 352 5114 416 5178
rect 434 5114 498 5178
rect 516 5114 580 5178
rect 598 5114 662 5178
rect 679 5114 743 5178
rect 760 5114 824 5178
rect 841 5114 905 5178
rect 922 5114 986 5178
rect 1003 5114 1067 5178
rect 1084 5114 1148 5178
rect 1165 5114 1229 5178
rect 1246 5114 1310 5178
rect 1327 5114 1391 5178
rect 1408 5114 1472 5178
rect 1489 5114 1553 5178
rect 1570 5114 1634 5178
rect 1651 5114 1715 5178
rect 1732 5114 1796 5178
rect 1813 5114 1877 5178
rect 1894 5114 1958 5178
rect 1975 5114 2039 5178
rect 2056 5114 2120 5178
rect 2137 5114 2201 5178
rect 2218 5114 2282 5178
rect 2299 5114 2363 5178
rect 2380 5114 2444 5178
rect 2461 5114 2525 5178
rect 2542 5114 2606 5178
rect 2623 5114 2687 5178
rect 2704 5114 2768 5178
rect 2785 5114 2849 5178
rect 2866 5114 2930 5178
rect 2947 5114 3011 5178
rect 3028 5114 3092 5178
rect 3109 5114 3173 5178
rect 3190 5114 3254 5178
rect 3271 5114 3335 5178
rect 3352 5114 3416 5178
rect 3433 5114 3497 5178
rect 3514 5114 3578 5178
rect 3595 5114 3659 5178
rect 3676 5114 3740 5178
rect 3757 5114 3821 5178
rect 3838 5114 3902 5178
rect 3919 5114 3983 5178
rect 4000 5114 4064 5178
rect 4081 5114 4145 5178
rect 4162 5114 4226 5178
rect 4243 5114 4307 5178
rect 4324 5114 4388 5178
rect 4405 5114 4469 5178
rect 4486 5114 4550 5178
rect 4567 5114 4631 5178
rect 4648 5114 4712 5178
rect 4729 5114 4793 5178
rect 4810 5114 4874 5178
rect 10157 5114 10221 5178
rect 10239 5114 10303 5178
rect 10321 5114 10385 5178
rect 10403 5114 10467 5178
rect 10485 5114 10549 5178
rect 10567 5114 10631 5178
rect 10649 5114 10713 5178
rect 10731 5114 10795 5178
rect 10813 5114 10877 5178
rect 10895 5114 10959 5178
rect 10977 5114 11041 5178
rect 11059 5114 11123 5178
rect 11141 5114 11205 5178
rect 11223 5114 11287 5178
rect 11305 5114 11369 5178
rect 11386 5114 11450 5178
rect 11467 5114 11531 5178
rect 11548 5114 11612 5178
rect 11629 5114 11693 5178
rect 11710 5114 11774 5178
rect 11791 5114 11855 5178
rect 11872 5114 11936 5178
rect 11953 5114 12017 5178
rect 12034 5114 12098 5178
rect 12115 5114 12179 5178
rect 12196 5114 12260 5178
rect 12277 5114 12341 5178
rect 12358 5114 12422 5178
rect 12439 5114 12503 5178
rect 12520 5114 12584 5178
rect 12601 5114 12665 5178
rect 12682 5114 12746 5178
rect 12763 5114 12827 5178
rect 12844 5114 12908 5178
rect 12925 5114 12989 5178
rect 13006 5114 13070 5178
rect 13087 5114 13151 5178
rect 13168 5114 13232 5178
rect 13249 5114 13313 5178
rect 13330 5114 13394 5178
rect 13411 5114 13475 5178
rect 13492 5114 13556 5178
rect 13573 5114 13637 5178
rect 13654 5114 13718 5178
rect 13735 5114 13799 5178
rect 13816 5114 13880 5178
rect 13897 5114 13961 5178
rect 13978 5114 14042 5178
rect 14059 5114 14123 5178
rect 14140 5114 14204 5178
rect 14221 5114 14285 5178
rect 14302 5114 14366 5178
rect 14383 5114 14447 5178
rect 14464 5114 14528 5178
rect 14545 5114 14609 5178
rect 14626 5114 14690 5178
rect 14707 5114 14771 5178
rect 14788 5114 14852 5178
rect 106 5028 170 5092
rect 188 5028 252 5092
rect 270 5028 334 5092
rect 352 5028 416 5092
rect 434 5028 498 5092
rect 516 5028 580 5092
rect 598 5028 662 5092
rect 679 5028 743 5092
rect 760 5028 824 5092
rect 841 5028 905 5092
rect 922 5028 986 5092
rect 1003 5028 1067 5092
rect 1084 5028 1148 5092
rect 1165 5028 1229 5092
rect 1246 5028 1310 5092
rect 1327 5028 1391 5092
rect 1408 5028 1472 5092
rect 1489 5028 1553 5092
rect 1570 5028 1634 5092
rect 1651 5028 1715 5092
rect 1732 5028 1796 5092
rect 1813 5028 1877 5092
rect 1894 5028 1958 5092
rect 1975 5028 2039 5092
rect 2056 5028 2120 5092
rect 2137 5028 2201 5092
rect 2218 5028 2282 5092
rect 2299 5028 2363 5092
rect 2380 5028 2444 5092
rect 2461 5028 2525 5092
rect 2542 5028 2606 5092
rect 2623 5028 2687 5092
rect 2704 5028 2768 5092
rect 2785 5028 2849 5092
rect 2866 5028 2930 5092
rect 2947 5028 3011 5092
rect 3028 5028 3092 5092
rect 3109 5028 3173 5092
rect 3190 5028 3254 5092
rect 3271 5028 3335 5092
rect 3352 5028 3416 5092
rect 3433 5028 3497 5092
rect 3514 5028 3578 5092
rect 3595 5028 3659 5092
rect 3676 5028 3740 5092
rect 3757 5028 3821 5092
rect 3838 5028 3902 5092
rect 3919 5028 3983 5092
rect 4000 5028 4064 5092
rect 4081 5028 4145 5092
rect 4162 5028 4226 5092
rect 4243 5028 4307 5092
rect 4324 5028 4388 5092
rect 4405 5028 4469 5092
rect 4486 5028 4550 5092
rect 4567 5028 4631 5092
rect 4648 5028 4712 5092
rect 4729 5028 4793 5092
rect 4810 5028 4874 5092
rect 10157 5028 10221 5092
rect 10239 5028 10303 5092
rect 10321 5028 10385 5092
rect 10403 5028 10467 5092
rect 10485 5028 10549 5092
rect 10567 5028 10631 5092
rect 10649 5028 10713 5092
rect 10731 5028 10795 5092
rect 10813 5028 10877 5092
rect 10895 5028 10959 5092
rect 10977 5028 11041 5092
rect 11059 5028 11123 5092
rect 11141 5028 11205 5092
rect 11223 5028 11287 5092
rect 11305 5028 11369 5092
rect 11386 5028 11450 5092
rect 11467 5028 11531 5092
rect 11548 5028 11612 5092
rect 11629 5028 11693 5092
rect 11710 5028 11774 5092
rect 11791 5028 11855 5092
rect 11872 5028 11936 5092
rect 11953 5028 12017 5092
rect 12034 5028 12098 5092
rect 12115 5028 12179 5092
rect 12196 5028 12260 5092
rect 12277 5028 12341 5092
rect 12358 5028 12422 5092
rect 12439 5028 12503 5092
rect 12520 5028 12584 5092
rect 12601 5028 12665 5092
rect 12682 5028 12746 5092
rect 12763 5028 12827 5092
rect 12844 5028 12908 5092
rect 12925 5028 12989 5092
rect 13006 5028 13070 5092
rect 13087 5028 13151 5092
rect 13168 5028 13232 5092
rect 13249 5028 13313 5092
rect 13330 5028 13394 5092
rect 13411 5028 13475 5092
rect 13492 5028 13556 5092
rect 13573 5028 13637 5092
rect 13654 5028 13718 5092
rect 13735 5028 13799 5092
rect 13816 5028 13880 5092
rect 13897 5028 13961 5092
rect 13978 5028 14042 5092
rect 14059 5028 14123 5092
rect 14140 5028 14204 5092
rect 14221 5028 14285 5092
rect 14302 5028 14366 5092
rect 14383 5028 14447 5092
rect 14464 5028 14528 5092
rect 14545 5028 14609 5092
rect 14626 5028 14690 5092
rect 14707 5028 14771 5092
rect 14788 5028 14852 5092
rect 106 4942 170 5006
rect 188 4942 252 5006
rect 270 4942 334 5006
rect 352 4942 416 5006
rect 434 4942 498 5006
rect 516 4942 580 5006
rect 598 4942 662 5006
rect 679 4942 743 5006
rect 760 4942 824 5006
rect 841 4942 905 5006
rect 922 4942 986 5006
rect 1003 4942 1067 5006
rect 1084 4942 1148 5006
rect 1165 4942 1229 5006
rect 1246 4942 1310 5006
rect 1327 4942 1391 5006
rect 1408 4942 1472 5006
rect 1489 4942 1553 5006
rect 1570 4942 1634 5006
rect 1651 4942 1715 5006
rect 1732 4942 1796 5006
rect 1813 4942 1877 5006
rect 1894 4942 1958 5006
rect 1975 4942 2039 5006
rect 2056 4942 2120 5006
rect 2137 4942 2201 5006
rect 2218 4942 2282 5006
rect 2299 4942 2363 5006
rect 2380 4942 2444 5006
rect 2461 4942 2525 5006
rect 2542 4942 2606 5006
rect 2623 4942 2687 5006
rect 2704 4942 2768 5006
rect 2785 4942 2849 5006
rect 2866 4942 2930 5006
rect 2947 4942 3011 5006
rect 3028 4942 3092 5006
rect 3109 4942 3173 5006
rect 3190 4942 3254 5006
rect 3271 4942 3335 5006
rect 3352 4942 3416 5006
rect 3433 4942 3497 5006
rect 3514 4942 3578 5006
rect 3595 4942 3659 5006
rect 3676 4942 3740 5006
rect 3757 4942 3821 5006
rect 3838 4942 3902 5006
rect 3919 4942 3983 5006
rect 4000 4942 4064 5006
rect 4081 4942 4145 5006
rect 4162 4942 4226 5006
rect 4243 4942 4307 5006
rect 4324 4942 4388 5006
rect 4405 4942 4469 5006
rect 4486 4942 4550 5006
rect 4567 4942 4631 5006
rect 4648 4942 4712 5006
rect 4729 4942 4793 5006
rect 4810 4942 4874 5006
rect 10157 4942 10221 5006
rect 10239 4942 10303 5006
rect 10321 4942 10385 5006
rect 10403 4942 10467 5006
rect 10485 4942 10549 5006
rect 10567 4942 10631 5006
rect 10649 4942 10713 5006
rect 10731 4942 10795 5006
rect 10813 4942 10877 5006
rect 10895 4942 10959 5006
rect 10977 4942 11041 5006
rect 11059 4942 11123 5006
rect 11141 4942 11205 5006
rect 11223 4942 11287 5006
rect 11305 4942 11369 5006
rect 11386 4942 11450 5006
rect 11467 4942 11531 5006
rect 11548 4942 11612 5006
rect 11629 4942 11693 5006
rect 11710 4942 11774 5006
rect 11791 4942 11855 5006
rect 11872 4942 11936 5006
rect 11953 4942 12017 5006
rect 12034 4942 12098 5006
rect 12115 4942 12179 5006
rect 12196 4942 12260 5006
rect 12277 4942 12341 5006
rect 12358 4942 12422 5006
rect 12439 4942 12503 5006
rect 12520 4942 12584 5006
rect 12601 4942 12665 5006
rect 12682 4942 12746 5006
rect 12763 4942 12827 5006
rect 12844 4942 12908 5006
rect 12925 4942 12989 5006
rect 13006 4942 13070 5006
rect 13087 4942 13151 5006
rect 13168 4942 13232 5006
rect 13249 4942 13313 5006
rect 13330 4942 13394 5006
rect 13411 4942 13475 5006
rect 13492 4942 13556 5006
rect 13573 4942 13637 5006
rect 13654 4942 13718 5006
rect 13735 4942 13799 5006
rect 13816 4942 13880 5006
rect 13897 4942 13961 5006
rect 13978 4942 14042 5006
rect 14059 4942 14123 5006
rect 14140 4942 14204 5006
rect 14221 4942 14285 5006
rect 14302 4942 14366 5006
rect 14383 4942 14447 5006
rect 14464 4942 14528 5006
rect 14545 4942 14609 5006
rect 14626 4942 14690 5006
rect 14707 4942 14771 5006
rect 14788 4942 14852 5006
rect 106 4856 170 4920
rect 188 4856 252 4920
rect 270 4856 334 4920
rect 352 4856 416 4920
rect 434 4856 498 4920
rect 516 4856 580 4920
rect 598 4856 662 4920
rect 679 4856 743 4920
rect 760 4856 824 4920
rect 841 4856 905 4920
rect 922 4856 986 4920
rect 1003 4856 1067 4920
rect 1084 4856 1148 4920
rect 1165 4856 1229 4920
rect 1246 4856 1310 4920
rect 1327 4856 1391 4920
rect 1408 4856 1472 4920
rect 1489 4856 1553 4920
rect 1570 4856 1634 4920
rect 1651 4856 1715 4920
rect 1732 4856 1796 4920
rect 1813 4856 1877 4920
rect 1894 4856 1958 4920
rect 1975 4856 2039 4920
rect 2056 4856 2120 4920
rect 2137 4856 2201 4920
rect 2218 4856 2282 4920
rect 2299 4856 2363 4920
rect 2380 4856 2444 4920
rect 2461 4856 2525 4920
rect 2542 4856 2606 4920
rect 2623 4856 2687 4920
rect 2704 4856 2768 4920
rect 2785 4856 2849 4920
rect 2866 4856 2930 4920
rect 2947 4856 3011 4920
rect 3028 4856 3092 4920
rect 3109 4856 3173 4920
rect 3190 4856 3254 4920
rect 3271 4856 3335 4920
rect 3352 4856 3416 4920
rect 3433 4856 3497 4920
rect 3514 4856 3578 4920
rect 3595 4856 3659 4920
rect 3676 4856 3740 4920
rect 3757 4856 3821 4920
rect 3838 4856 3902 4920
rect 3919 4856 3983 4920
rect 4000 4856 4064 4920
rect 4081 4856 4145 4920
rect 4162 4856 4226 4920
rect 4243 4856 4307 4920
rect 4324 4856 4388 4920
rect 4405 4856 4469 4920
rect 4486 4856 4550 4920
rect 4567 4856 4631 4920
rect 4648 4856 4712 4920
rect 4729 4856 4793 4920
rect 4810 4856 4874 4920
rect 10157 4856 10221 4920
rect 10239 4856 10303 4920
rect 10321 4856 10385 4920
rect 10403 4856 10467 4920
rect 10485 4856 10549 4920
rect 10567 4856 10631 4920
rect 10649 4856 10713 4920
rect 10731 4856 10795 4920
rect 10813 4856 10877 4920
rect 10895 4856 10959 4920
rect 10977 4856 11041 4920
rect 11059 4856 11123 4920
rect 11141 4856 11205 4920
rect 11223 4856 11287 4920
rect 11305 4856 11369 4920
rect 11386 4856 11450 4920
rect 11467 4856 11531 4920
rect 11548 4856 11612 4920
rect 11629 4856 11693 4920
rect 11710 4856 11774 4920
rect 11791 4856 11855 4920
rect 11872 4856 11936 4920
rect 11953 4856 12017 4920
rect 12034 4856 12098 4920
rect 12115 4856 12179 4920
rect 12196 4856 12260 4920
rect 12277 4856 12341 4920
rect 12358 4856 12422 4920
rect 12439 4856 12503 4920
rect 12520 4856 12584 4920
rect 12601 4856 12665 4920
rect 12682 4856 12746 4920
rect 12763 4856 12827 4920
rect 12844 4856 12908 4920
rect 12925 4856 12989 4920
rect 13006 4856 13070 4920
rect 13087 4856 13151 4920
rect 13168 4856 13232 4920
rect 13249 4856 13313 4920
rect 13330 4856 13394 4920
rect 13411 4856 13475 4920
rect 13492 4856 13556 4920
rect 13573 4856 13637 4920
rect 13654 4856 13718 4920
rect 13735 4856 13799 4920
rect 13816 4856 13880 4920
rect 13897 4856 13961 4920
rect 13978 4856 14042 4920
rect 14059 4856 14123 4920
rect 14140 4856 14204 4920
rect 14221 4856 14285 4920
rect 14302 4856 14366 4920
rect 14383 4856 14447 4920
rect 14464 4856 14528 4920
rect 14545 4856 14609 4920
rect 14626 4856 14690 4920
rect 14707 4856 14771 4920
rect 14788 4856 14852 4920
rect 106 4770 170 4834
rect 188 4770 252 4834
rect 270 4770 334 4834
rect 352 4770 416 4834
rect 434 4770 498 4834
rect 516 4770 580 4834
rect 598 4770 662 4834
rect 679 4770 743 4834
rect 760 4770 824 4834
rect 841 4770 905 4834
rect 922 4770 986 4834
rect 1003 4770 1067 4834
rect 1084 4770 1148 4834
rect 1165 4770 1229 4834
rect 1246 4770 1310 4834
rect 1327 4770 1391 4834
rect 1408 4770 1472 4834
rect 1489 4770 1553 4834
rect 1570 4770 1634 4834
rect 1651 4770 1715 4834
rect 1732 4770 1796 4834
rect 1813 4770 1877 4834
rect 1894 4770 1958 4834
rect 1975 4770 2039 4834
rect 2056 4770 2120 4834
rect 2137 4770 2201 4834
rect 2218 4770 2282 4834
rect 2299 4770 2363 4834
rect 2380 4770 2444 4834
rect 2461 4770 2525 4834
rect 2542 4770 2606 4834
rect 2623 4770 2687 4834
rect 2704 4770 2768 4834
rect 2785 4770 2849 4834
rect 2866 4770 2930 4834
rect 2947 4770 3011 4834
rect 3028 4770 3092 4834
rect 3109 4770 3173 4834
rect 3190 4770 3254 4834
rect 3271 4770 3335 4834
rect 3352 4770 3416 4834
rect 3433 4770 3497 4834
rect 3514 4770 3578 4834
rect 3595 4770 3659 4834
rect 3676 4770 3740 4834
rect 3757 4770 3821 4834
rect 3838 4770 3902 4834
rect 3919 4770 3983 4834
rect 4000 4770 4064 4834
rect 4081 4770 4145 4834
rect 4162 4770 4226 4834
rect 4243 4770 4307 4834
rect 4324 4770 4388 4834
rect 4405 4770 4469 4834
rect 4486 4770 4550 4834
rect 4567 4770 4631 4834
rect 4648 4770 4712 4834
rect 4729 4770 4793 4834
rect 4810 4770 4874 4834
rect 10157 4770 10221 4834
rect 10239 4770 10303 4834
rect 10321 4770 10385 4834
rect 10403 4770 10467 4834
rect 10485 4770 10549 4834
rect 10567 4770 10631 4834
rect 10649 4770 10713 4834
rect 10731 4770 10795 4834
rect 10813 4770 10877 4834
rect 10895 4770 10959 4834
rect 10977 4770 11041 4834
rect 11059 4770 11123 4834
rect 11141 4770 11205 4834
rect 11223 4770 11287 4834
rect 11305 4770 11369 4834
rect 11386 4770 11450 4834
rect 11467 4770 11531 4834
rect 11548 4770 11612 4834
rect 11629 4770 11693 4834
rect 11710 4770 11774 4834
rect 11791 4770 11855 4834
rect 11872 4770 11936 4834
rect 11953 4770 12017 4834
rect 12034 4770 12098 4834
rect 12115 4770 12179 4834
rect 12196 4770 12260 4834
rect 12277 4770 12341 4834
rect 12358 4770 12422 4834
rect 12439 4770 12503 4834
rect 12520 4770 12584 4834
rect 12601 4770 12665 4834
rect 12682 4770 12746 4834
rect 12763 4770 12827 4834
rect 12844 4770 12908 4834
rect 12925 4770 12989 4834
rect 13006 4770 13070 4834
rect 13087 4770 13151 4834
rect 13168 4770 13232 4834
rect 13249 4770 13313 4834
rect 13330 4770 13394 4834
rect 13411 4770 13475 4834
rect 13492 4770 13556 4834
rect 13573 4770 13637 4834
rect 13654 4770 13718 4834
rect 13735 4770 13799 4834
rect 13816 4770 13880 4834
rect 13897 4770 13961 4834
rect 13978 4770 14042 4834
rect 14059 4770 14123 4834
rect 14140 4770 14204 4834
rect 14221 4770 14285 4834
rect 14302 4770 14366 4834
rect 14383 4770 14447 4834
rect 14464 4770 14528 4834
rect 14545 4770 14609 4834
rect 14626 4770 14690 4834
rect 14707 4770 14771 4834
rect 14788 4770 14852 4834
<< obsm4 >>
rect 0 39593 15000 39600
rect 0 39529 111 39593
rect 175 39529 191 39593
rect 255 39529 271 39593
rect 335 39529 351 39593
rect 415 39529 431 39593
rect 495 39529 511 39593
rect 575 39529 591 39593
rect 655 39529 671 39593
rect 735 39529 751 39593
rect 815 39529 831 39593
rect 895 39529 911 39593
rect 975 39529 991 39593
rect 1055 39529 1071 39593
rect 1135 39529 1151 39593
rect 1215 39529 1231 39593
rect 1295 39529 1311 39593
rect 1375 39529 1391 39593
rect 1455 39529 1471 39593
rect 1535 39529 1551 39593
rect 1615 39529 1631 39593
rect 1695 39529 1711 39593
rect 1775 39529 1791 39593
rect 1855 39529 1871 39593
rect 1935 39529 1951 39593
rect 2015 39529 2031 39593
rect 2095 39529 2111 39593
rect 2175 39529 2191 39593
rect 2255 39529 2271 39593
rect 2335 39529 2351 39593
rect 2415 39529 2431 39593
rect 2495 39529 2511 39593
rect 2575 39529 12416 39593
rect 12480 39529 12498 39593
rect 12562 39529 12580 39593
rect 12644 39529 12662 39593
rect 12726 39529 12744 39593
rect 12808 39529 12826 39593
rect 12890 39529 12908 39593
rect 12972 39529 12990 39593
rect 13054 39529 13072 39593
rect 13136 39529 13154 39593
rect 13218 39529 13236 39593
rect 13300 39529 13318 39593
rect 13382 39529 13400 39593
rect 13464 39529 13482 39593
rect 13546 39529 13564 39593
rect 13628 39529 13646 39593
rect 13710 39529 13728 39593
rect 13792 39529 13810 39593
rect 13874 39529 13892 39593
rect 13956 39529 13974 39593
rect 14038 39529 14056 39593
rect 14120 39529 14138 39593
rect 14202 39529 14220 39593
rect 14284 39529 14302 39593
rect 14366 39529 14384 39593
rect 14448 39529 14466 39593
rect 14530 39529 14548 39593
rect 14612 39529 14630 39593
rect 14694 39529 14712 39593
rect 14776 39529 14794 39593
rect 14858 39529 14876 39593
rect 14940 39529 15000 39593
rect 0 39512 15000 39529
rect 0 39448 111 39512
rect 175 39448 191 39512
rect 255 39448 271 39512
rect 335 39448 351 39512
rect 415 39448 431 39512
rect 495 39448 511 39512
rect 575 39448 591 39512
rect 655 39448 671 39512
rect 735 39448 751 39512
rect 815 39448 831 39512
rect 895 39448 911 39512
rect 975 39448 991 39512
rect 1055 39448 1071 39512
rect 1135 39448 1151 39512
rect 1215 39448 1231 39512
rect 1295 39448 1311 39512
rect 1375 39448 1391 39512
rect 1455 39448 1471 39512
rect 1535 39448 1551 39512
rect 1615 39448 1631 39512
rect 1695 39448 1711 39512
rect 1775 39448 1791 39512
rect 1855 39448 1871 39512
rect 1935 39448 1951 39512
rect 2015 39448 2031 39512
rect 2095 39448 2111 39512
rect 2175 39448 2191 39512
rect 2255 39448 2271 39512
rect 2335 39448 2351 39512
rect 2415 39448 2431 39512
rect 2495 39448 2511 39512
rect 2575 39448 12416 39512
rect 12480 39448 12498 39512
rect 12562 39448 12580 39512
rect 12644 39448 12662 39512
rect 12726 39448 12744 39512
rect 12808 39448 12826 39512
rect 12890 39448 12908 39512
rect 12972 39448 12990 39512
rect 13054 39448 13072 39512
rect 13136 39448 13154 39512
rect 13218 39448 13236 39512
rect 13300 39448 13318 39512
rect 13382 39448 13400 39512
rect 13464 39448 13482 39512
rect 13546 39448 13564 39512
rect 13628 39448 13646 39512
rect 13710 39448 13728 39512
rect 13792 39448 13810 39512
rect 13874 39448 13892 39512
rect 13956 39448 13974 39512
rect 14038 39448 14056 39512
rect 14120 39448 14138 39512
rect 14202 39448 14220 39512
rect 14284 39448 14302 39512
rect 14366 39448 14384 39512
rect 14448 39448 14466 39512
rect 14530 39448 14548 39512
rect 14612 39448 14630 39512
rect 14694 39448 14712 39512
rect 14776 39448 14794 39512
rect 14858 39448 14876 39512
rect 14940 39448 15000 39512
rect 0 39431 15000 39448
rect 0 39367 111 39431
rect 175 39367 191 39431
rect 255 39367 271 39431
rect 335 39367 351 39431
rect 415 39367 431 39431
rect 495 39367 511 39431
rect 575 39367 591 39431
rect 655 39367 671 39431
rect 735 39367 751 39431
rect 815 39367 831 39431
rect 895 39367 911 39431
rect 975 39367 991 39431
rect 1055 39367 1071 39431
rect 1135 39367 1151 39431
rect 1215 39367 1231 39431
rect 1295 39367 1311 39431
rect 1375 39367 1391 39431
rect 1455 39367 1471 39431
rect 1535 39367 1551 39431
rect 1615 39367 1631 39431
rect 1695 39367 1711 39431
rect 1775 39367 1791 39431
rect 1855 39367 1871 39431
rect 1935 39367 1951 39431
rect 2015 39367 2031 39431
rect 2095 39367 2111 39431
rect 2175 39367 2191 39431
rect 2255 39367 2271 39431
rect 2335 39367 2351 39431
rect 2415 39367 2431 39431
rect 2495 39367 2511 39431
rect 2575 39367 12416 39431
rect 12480 39367 12498 39431
rect 12562 39367 12580 39431
rect 12644 39367 12662 39431
rect 12726 39367 12744 39431
rect 12808 39367 12826 39431
rect 12890 39367 12908 39431
rect 12972 39367 12990 39431
rect 13054 39367 13072 39431
rect 13136 39367 13154 39431
rect 13218 39367 13236 39431
rect 13300 39367 13318 39431
rect 13382 39367 13400 39431
rect 13464 39367 13482 39431
rect 13546 39367 13564 39431
rect 13628 39367 13646 39431
rect 13710 39367 13728 39431
rect 13792 39367 13810 39431
rect 13874 39367 13892 39431
rect 13956 39367 13974 39431
rect 14038 39367 14056 39431
rect 14120 39367 14138 39431
rect 14202 39367 14220 39431
rect 14284 39367 14302 39431
rect 14366 39367 14384 39431
rect 14448 39367 14466 39431
rect 14530 39367 14548 39431
rect 14612 39367 14630 39431
rect 14694 39367 14712 39431
rect 14776 39367 14794 39431
rect 14858 39367 14876 39431
rect 14940 39367 15000 39431
rect 0 39350 15000 39367
rect 0 39286 111 39350
rect 175 39286 191 39350
rect 255 39286 271 39350
rect 335 39286 351 39350
rect 415 39286 431 39350
rect 495 39286 511 39350
rect 575 39286 591 39350
rect 655 39286 671 39350
rect 735 39286 751 39350
rect 815 39286 831 39350
rect 895 39286 911 39350
rect 975 39286 991 39350
rect 1055 39286 1071 39350
rect 1135 39286 1151 39350
rect 1215 39286 1231 39350
rect 1295 39286 1311 39350
rect 1375 39286 1391 39350
rect 1455 39286 1471 39350
rect 1535 39286 1551 39350
rect 1615 39286 1631 39350
rect 1695 39286 1711 39350
rect 1775 39286 1791 39350
rect 1855 39286 1871 39350
rect 1935 39286 1951 39350
rect 2015 39286 2031 39350
rect 2095 39286 2111 39350
rect 2175 39286 2191 39350
rect 2255 39286 2271 39350
rect 2335 39286 2351 39350
rect 2415 39286 2431 39350
rect 2495 39286 2511 39350
rect 2575 39286 12416 39350
rect 12480 39286 12498 39350
rect 12562 39286 12580 39350
rect 12644 39286 12662 39350
rect 12726 39286 12744 39350
rect 12808 39286 12826 39350
rect 12890 39286 12908 39350
rect 12972 39286 12990 39350
rect 13054 39286 13072 39350
rect 13136 39286 13154 39350
rect 13218 39286 13236 39350
rect 13300 39286 13318 39350
rect 13382 39286 13400 39350
rect 13464 39286 13482 39350
rect 13546 39286 13564 39350
rect 13628 39286 13646 39350
rect 13710 39286 13728 39350
rect 13792 39286 13810 39350
rect 13874 39286 13892 39350
rect 13956 39286 13974 39350
rect 14038 39286 14056 39350
rect 14120 39286 14138 39350
rect 14202 39286 14220 39350
rect 14284 39286 14302 39350
rect 14366 39286 14384 39350
rect 14448 39286 14466 39350
rect 14530 39286 14548 39350
rect 14612 39286 14630 39350
rect 14694 39286 14712 39350
rect 14776 39286 14794 39350
rect 14858 39286 14876 39350
rect 14940 39286 15000 39350
rect 0 39269 15000 39286
rect 0 39205 111 39269
rect 175 39205 191 39269
rect 255 39205 271 39269
rect 335 39205 351 39269
rect 415 39205 431 39269
rect 495 39205 511 39269
rect 575 39205 591 39269
rect 655 39205 671 39269
rect 735 39205 751 39269
rect 815 39205 831 39269
rect 895 39205 911 39269
rect 975 39205 991 39269
rect 1055 39205 1071 39269
rect 1135 39205 1151 39269
rect 1215 39205 1231 39269
rect 1295 39205 1311 39269
rect 1375 39205 1391 39269
rect 1455 39205 1471 39269
rect 1535 39205 1551 39269
rect 1615 39205 1631 39269
rect 1695 39205 1711 39269
rect 1775 39205 1791 39269
rect 1855 39205 1871 39269
rect 1935 39205 1951 39269
rect 2015 39205 2031 39269
rect 2095 39205 2111 39269
rect 2175 39205 2191 39269
rect 2255 39205 2271 39269
rect 2335 39205 2351 39269
rect 2415 39205 2431 39269
rect 2495 39205 2511 39269
rect 2575 39205 12416 39269
rect 12480 39205 12498 39269
rect 12562 39205 12580 39269
rect 12644 39205 12662 39269
rect 12726 39205 12744 39269
rect 12808 39205 12826 39269
rect 12890 39205 12908 39269
rect 12972 39205 12990 39269
rect 13054 39205 13072 39269
rect 13136 39205 13154 39269
rect 13218 39205 13236 39269
rect 13300 39205 13318 39269
rect 13382 39205 13400 39269
rect 13464 39205 13482 39269
rect 13546 39205 13564 39269
rect 13628 39205 13646 39269
rect 13710 39205 13728 39269
rect 13792 39205 13810 39269
rect 13874 39205 13892 39269
rect 13956 39205 13974 39269
rect 14038 39205 14056 39269
rect 14120 39205 14138 39269
rect 14202 39205 14220 39269
rect 14284 39205 14302 39269
rect 14366 39205 14384 39269
rect 14448 39205 14466 39269
rect 14530 39205 14548 39269
rect 14612 39205 14630 39269
rect 14694 39205 14712 39269
rect 14776 39205 14794 39269
rect 14858 39205 14876 39269
rect 14940 39205 15000 39269
rect 0 39188 15000 39205
rect 0 39124 111 39188
rect 175 39124 191 39188
rect 255 39124 271 39188
rect 335 39124 351 39188
rect 415 39124 431 39188
rect 495 39124 511 39188
rect 575 39124 591 39188
rect 655 39124 671 39188
rect 735 39124 751 39188
rect 815 39124 831 39188
rect 895 39124 911 39188
rect 975 39124 991 39188
rect 1055 39124 1071 39188
rect 1135 39124 1151 39188
rect 1215 39124 1231 39188
rect 1295 39124 1311 39188
rect 1375 39124 1391 39188
rect 1455 39124 1471 39188
rect 1535 39124 1551 39188
rect 1615 39124 1631 39188
rect 1695 39124 1711 39188
rect 1775 39124 1791 39188
rect 1855 39124 1871 39188
rect 1935 39124 1951 39188
rect 2015 39124 2031 39188
rect 2095 39124 2111 39188
rect 2175 39124 2191 39188
rect 2255 39124 2271 39188
rect 2335 39124 2351 39188
rect 2415 39124 2431 39188
rect 2495 39124 2511 39188
rect 2575 39124 12416 39188
rect 12480 39124 12498 39188
rect 12562 39124 12580 39188
rect 12644 39124 12662 39188
rect 12726 39124 12744 39188
rect 12808 39124 12826 39188
rect 12890 39124 12908 39188
rect 12972 39124 12990 39188
rect 13054 39124 13072 39188
rect 13136 39124 13154 39188
rect 13218 39124 13236 39188
rect 13300 39124 13318 39188
rect 13382 39124 13400 39188
rect 13464 39124 13482 39188
rect 13546 39124 13564 39188
rect 13628 39124 13646 39188
rect 13710 39124 13728 39188
rect 13792 39124 13810 39188
rect 13874 39124 13892 39188
rect 13956 39124 13974 39188
rect 14038 39124 14056 39188
rect 14120 39124 14138 39188
rect 14202 39124 14220 39188
rect 14284 39124 14302 39188
rect 14366 39124 14384 39188
rect 14448 39124 14466 39188
rect 14530 39124 14548 39188
rect 14612 39124 14630 39188
rect 14694 39124 14712 39188
rect 14776 39124 14794 39188
rect 14858 39124 14876 39188
rect 14940 39124 15000 39188
rect 0 39107 15000 39124
rect 0 39043 111 39107
rect 175 39043 191 39107
rect 255 39043 271 39107
rect 335 39043 351 39107
rect 415 39043 431 39107
rect 495 39043 511 39107
rect 575 39043 591 39107
rect 655 39043 671 39107
rect 735 39043 751 39107
rect 815 39043 831 39107
rect 895 39043 911 39107
rect 975 39043 991 39107
rect 1055 39043 1071 39107
rect 1135 39043 1151 39107
rect 1215 39043 1231 39107
rect 1295 39043 1311 39107
rect 1375 39043 1391 39107
rect 1455 39043 1471 39107
rect 1535 39043 1551 39107
rect 1615 39043 1631 39107
rect 1695 39043 1711 39107
rect 1775 39043 1791 39107
rect 1855 39043 1871 39107
rect 1935 39043 1951 39107
rect 2015 39043 2031 39107
rect 2095 39043 2111 39107
rect 2175 39043 2191 39107
rect 2255 39043 2271 39107
rect 2335 39043 2351 39107
rect 2415 39043 2431 39107
rect 2495 39043 2511 39107
rect 2575 39043 12416 39107
rect 12480 39043 12498 39107
rect 12562 39043 12580 39107
rect 12644 39043 12662 39107
rect 12726 39043 12744 39107
rect 12808 39043 12826 39107
rect 12890 39043 12908 39107
rect 12972 39043 12990 39107
rect 13054 39043 13072 39107
rect 13136 39043 13154 39107
rect 13218 39043 13236 39107
rect 13300 39043 13318 39107
rect 13382 39043 13400 39107
rect 13464 39043 13482 39107
rect 13546 39043 13564 39107
rect 13628 39043 13646 39107
rect 13710 39043 13728 39107
rect 13792 39043 13810 39107
rect 13874 39043 13892 39107
rect 13956 39043 13974 39107
rect 14038 39043 14056 39107
rect 14120 39043 14138 39107
rect 14202 39043 14220 39107
rect 14284 39043 14302 39107
rect 14366 39043 14384 39107
rect 14448 39043 14466 39107
rect 14530 39043 14548 39107
rect 14612 39043 14630 39107
rect 14694 39043 14712 39107
rect 14776 39043 14794 39107
rect 14858 39043 14876 39107
rect 14940 39043 15000 39107
rect 0 39026 15000 39043
rect 0 38962 111 39026
rect 175 38962 191 39026
rect 255 38962 271 39026
rect 335 38962 351 39026
rect 415 38962 431 39026
rect 495 38962 511 39026
rect 575 38962 591 39026
rect 655 38962 671 39026
rect 735 38962 751 39026
rect 815 38962 831 39026
rect 895 38962 911 39026
rect 975 38962 991 39026
rect 1055 38962 1071 39026
rect 1135 38962 1151 39026
rect 1215 38962 1231 39026
rect 1295 38962 1311 39026
rect 1375 38962 1391 39026
rect 1455 38962 1471 39026
rect 1535 38962 1551 39026
rect 1615 38962 1631 39026
rect 1695 38962 1711 39026
rect 1775 38962 1791 39026
rect 1855 38962 1871 39026
rect 1935 38962 1951 39026
rect 2015 38962 2031 39026
rect 2095 38962 2111 39026
rect 2175 38962 2191 39026
rect 2255 38962 2271 39026
rect 2335 38962 2351 39026
rect 2415 38962 2431 39026
rect 2495 38962 2511 39026
rect 2575 38962 12416 39026
rect 12480 38962 12498 39026
rect 12562 38962 12580 39026
rect 12644 38962 12662 39026
rect 12726 38962 12744 39026
rect 12808 38962 12826 39026
rect 12890 38962 12908 39026
rect 12972 38962 12990 39026
rect 13054 38962 13072 39026
rect 13136 38962 13154 39026
rect 13218 38962 13236 39026
rect 13300 38962 13318 39026
rect 13382 38962 13400 39026
rect 13464 38962 13482 39026
rect 13546 38962 13564 39026
rect 13628 38962 13646 39026
rect 13710 38962 13728 39026
rect 13792 38962 13810 39026
rect 13874 38962 13892 39026
rect 13956 38962 13974 39026
rect 14038 38962 14056 39026
rect 14120 38962 14138 39026
rect 14202 38962 14220 39026
rect 14284 38962 14302 39026
rect 14366 38962 14384 39026
rect 14448 38962 14466 39026
rect 14530 38962 14548 39026
rect 14612 38962 14630 39026
rect 14694 38962 14712 39026
rect 14776 38962 14794 39026
rect 14858 38962 14876 39026
rect 14940 38962 15000 39026
rect 0 38945 15000 38962
rect 0 38881 111 38945
rect 175 38881 191 38945
rect 255 38881 271 38945
rect 335 38881 351 38945
rect 415 38881 431 38945
rect 495 38881 511 38945
rect 575 38881 591 38945
rect 655 38881 671 38945
rect 735 38881 751 38945
rect 815 38881 831 38945
rect 895 38881 911 38945
rect 975 38881 991 38945
rect 1055 38881 1071 38945
rect 1135 38881 1151 38945
rect 1215 38881 1231 38945
rect 1295 38881 1311 38945
rect 1375 38881 1391 38945
rect 1455 38881 1471 38945
rect 1535 38881 1551 38945
rect 1615 38881 1631 38945
rect 1695 38881 1711 38945
rect 1775 38881 1791 38945
rect 1855 38881 1871 38945
rect 1935 38881 1951 38945
rect 2015 38881 2031 38945
rect 2095 38881 2111 38945
rect 2175 38881 2191 38945
rect 2255 38881 2271 38945
rect 2335 38881 2351 38945
rect 2415 38881 2431 38945
rect 2495 38881 2511 38945
rect 2575 38881 12416 38945
rect 12480 38881 12498 38945
rect 12562 38881 12580 38945
rect 12644 38881 12662 38945
rect 12726 38881 12744 38945
rect 12808 38881 12826 38945
rect 12890 38881 12908 38945
rect 12972 38881 12990 38945
rect 13054 38881 13072 38945
rect 13136 38881 13154 38945
rect 13218 38881 13236 38945
rect 13300 38881 13318 38945
rect 13382 38881 13400 38945
rect 13464 38881 13482 38945
rect 13546 38881 13564 38945
rect 13628 38881 13646 38945
rect 13710 38881 13728 38945
rect 13792 38881 13810 38945
rect 13874 38881 13892 38945
rect 13956 38881 13974 38945
rect 14038 38881 14056 38945
rect 14120 38881 14138 38945
rect 14202 38881 14220 38945
rect 14284 38881 14302 38945
rect 14366 38881 14384 38945
rect 14448 38881 14466 38945
rect 14530 38881 14548 38945
rect 14612 38881 14630 38945
rect 14694 38881 14712 38945
rect 14776 38881 14794 38945
rect 14858 38881 14876 38945
rect 14940 38881 15000 38945
rect 0 38864 15000 38881
rect 0 38800 111 38864
rect 175 38800 191 38864
rect 255 38800 271 38864
rect 335 38800 351 38864
rect 415 38800 431 38864
rect 495 38800 511 38864
rect 575 38800 591 38864
rect 655 38800 671 38864
rect 735 38800 751 38864
rect 815 38800 831 38864
rect 895 38800 911 38864
rect 975 38800 991 38864
rect 1055 38800 1071 38864
rect 1135 38800 1151 38864
rect 1215 38800 1231 38864
rect 1295 38800 1311 38864
rect 1375 38800 1391 38864
rect 1455 38800 1471 38864
rect 1535 38800 1551 38864
rect 1615 38800 1631 38864
rect 1695 38800 1711 38864
rect 1775 38800 1791 38864
rect 1855 38800 1871 38864
rect 1935 38800 1951 38864
rect 2015 38800 2031 38864
rect 2095 38800 2111 38864
rect 2175 38800 2191 38864
rect 2255 38800 2271 38864
rect 2335 38800 2351 38864
rect 2415 38800 2431 38864
rect 2495 38800 2511 38864
rect 2575 38800 12416 38864
rect 12480 38800 12498 38864
rect 12562 38800 12580 38864
rect 12644 38800 12662 38864
rect 12726 38800 12744 38864
rect 12808 38800 12826 38864
rect 12890 38800 12908 38864
rect 12972 38800 12990 38864
rect 13054 38800 13072 38864
rect 13136 38800 13154 38864
rect 13218 38800 13236 38864
rect 13300 38800 13318 38864
rect 13382 38800 13400 38864
rect 13464 38800 13482 38864
rect 13546 38800 13564 38864
rect 13628 38800 13646 38864
rect 13710 38800 13728 38864
rect 13792 38800 13810 38864
rect 13874 38800 13892 38864
rect 13956 38800 13974 38864
rect 14038 38800 14056 38864
rect 14120 38800 14138 38864
rect 14202 38800 14220 38864
rect 14284 38800 14302 38864
rect 14366 38800 14384 38864
rect 14448 38800 14466 38864
rect 14530 38800 14548 38864
rect 14612 38800 14630 38864
rect 14694 38800 14712 38864
rect 14776 38800 14794 38864
rect 14858 38800 14876 38864
rect 14940 38800 15000 38864
rect 0 38783 15000 38800
rect 0 38719 111 38783
rect 175 38719 191 38783
rect 255 38719 271 38783
rect 335 38719 351 38783
rect 415 38719 431 38783
rect 495 38719 511 38783
rect 575 38719 591 38783
rect 655 38719 671 38783
rect 735 38719 751 38783
rect 815 38719 831 38783
rect 895 38719 911 38783
rect 975 38719 991 38783
rect 1055 38719 1071 38783
rect 1135 38719 1151 38783
rect 1215 38719 1231 38783
rect 1295 38719 1311 38783
rect 1375 38719 1391 38783
rect 1455 38719 1471 38783
rect 1535 38719 1551 38783
rect 1615 38719 1631 38783
rect 1695 38719 1711 38783
rect 1775 38719 1791 38783
rect 1855 38719 1871 38783
rect 1935 38719 1951 38783
rect 2015 38719 2031 38783
rect 2095 38719 2111 38783
rect 2175 38719 2191 38783
rect 2255 38719 2271 38783
rect 2335 38719 2351 38783
rect 2415 38719 2431 38783
rect 2495 38719 2511 38783
rect 2575 38719 12416 38783
rect 12480 38719 12498 38783
rect 12562 38719 12580 38783
rect 12644 38719 12662 38783
rect 12726 38719 12744 38783
rect 12808 38719 12826 38783
rect 12890 38719 12908 38783
rect 12972 38719 12990 38783
rect 13054 38719 13072 38783
rect 13136 38719 13154 38783
rect 13218 38719 13236 38783
rect 13300 38719 13318 38783
rect 13382 38719 13400 38783
rect 13464 38719 13482 38783
rect 13546 38719 13564 38783
rect 13628 38719 13646 38783
rect 13710 38719 13728 38783
rect 13792 38719 13810 38783
rect 13874 38719 13892 38783
rect 13956 38719 13974 38783
rect 14038 38719 14056 38783
rect 14120 38719 14138 38783
rect 14202 38719 14220 38783
rect 14284 38719 14302 38783
rect 14366 38719 14384 38783
rect 14448 38719 14466 38783
rect 14530 38719 14548 38783
rect 14612 38719 14630 38783
rect 14694 38719 14712 38783
rect 14776 38719 14794 38783
rect 14858 38719 14876 38783
rect 14940 38719 15000 38783
rect 0 38702 15000 38719
rect 0 38638 111 38702
rect 175 38638 191 38702
rect 255 38638 271 38702
rect 335 38638 351 38702
rect 415 38638 431 38702
rect 495 38638 511 38702
rect 575 38638 591 38702
rect 655 38638 671 38702
rect 735 38638 751 38702
rect 815 38638 831 38702
rect 895 38638 911 38702
rect 975 38638 991 38702
rect 1055 38638 1071 38702
rect 1135 38638 1151 38702
rect 1215 38638 1231 38702
rect 1295 38638 1311 38702
rect 1375 38638 1391 38702
rect 1455 38638 1471 38702
rect 1535 38638 1551 38702
rect 1615 38638 1631 38702
rect 1695 38638 1711 38702
rect 1775 38638 1791 38702
rect 1855 38638 1871 38702
rect 1935 38638 1951 38702
rect 2015 38638 2031 38702
rect 2095 38638 2111 38702
rect 2175 38638 2191 38702
rect 2255 38638 2271 38702
rect 2335 38638 2351 38702
rect 2415 38638 2431 38702
rect 2495 38638 2511 38702
rect 2575 38638 12416 38702
rect 12480 38638 12498 38702
rect 12562 38638 12580 38702
rect 12644 38638 12662 38702
rect 12726 38638 12744 38702
rect 12808 38638 12826 38702
rect 12890 38638 12908 38702
rect 12972 38638 12990 38702
rect 13054 38638 13072 38702
rect 13136 38638 13154 38702
rect 13218 38638 13236 38702
rect 13300 38638 13318 38702
rect 13382 38638 13400 38702
rect 13464 38638 13482 38702
rect 13546 38638 13564 38702
rect 13628 38638 13646 38702
rect 13710 38638 13728 38702
rect 13792 38638 13810 38702
rect 13874 38638 13892 38702
rect 13956 38638 13974 38702
rect 14038 38638 14056 38702
rect 14120 38638 14138 38702
rect 14202 38638 14220 38702
rect 14284 38638 14302 38702
rect 14366 38638 14384 38702
rect 14448 38638 14466 38702
rect 14530 38638 14548 38702
rect 14612 38638 14630 38702
rect 14694 38638 14712 38702
rect 14776 38638 14794 38702
rect 14858 38638 14876 38702
rect 14940 38638 15000 38702
rect 0 38621 15000 38638
rect 0 38557 111 38621
rect 175 38557 191 38621
rect 255 38557 271 38621
rect 335 38557 351 38621
rect 415 38557 431 38621
rect 495 38557 511 38621
rect 575 38557 591 38621
rect 655 38557 671 38621
rect 735 38557 751 38621
rect 815 38557 831 38621
rect 895 38557 911 38621
rect 975 38557 991 38621
rect 1055 38557 1071 38621
rect 1135 38557 1151 38621
rect 1215 38557 1231 38621
rect 1295 38557 1311 38621
rect 1375 38557 1391 38621
rect 1455 38557 1471 38621
rect 1535 38557 1551 38621
rect 1615 38557 1631 38621
rect 1695 38557 1711 38621
rect 1775 38557 1791 38621
rect 1855 38557 1871 38621
rect 1935 38557 1951 38621
rect 2015 38557 2031 38621
rect 2095 38557 2111 38621
rect 2175 38557 2191 38621
rect 2255 38557 2271 38621
rect 2335 38557 2351 38621
rect 2415 38557 2431 38621
rect 2495 38557 2511 38621
rect 2575 38557 12416 38621
rect 12480 38557 12498 38621
rect 12562 38557 12580 38621
rect 12644 38557 12662 38621
rect 12726 38557 12744 38621
rect 12808 38557 12826 38621
rect 12890 38557 12908 38621
rect 12972 38557 12990 38621
rect 13054 38557 13072 38621
rect 13136 38557 13154 38621
rect 13218 38557 13236 38621
rect 13300 38557 13318 38621
rect 13382 38557 13400 38621
rect 13464 38557 13482 38621
rect 13546 38557 13564 38621
rect 13628 38557 13646 38621
rect 13710 38557 13728 38621
rect 13792 38557 13810 38621
rect 13874 38557 13892 38621
rect 13956 38557 13974 38621
rect 14038 38557 14056 38621
rect 14120 38557 14138 38621
rect 14202 38557 14220 38621
rect 14284 38557 14302 38621
rect 14366 38557 14384 38621
rect 14448 38557 14466 38621
rect 14530 38557 14548 38621
rect 14612 38557 14630 38621
rect 14694 38557 14712 38621
rect 14776 38557 14794 38621
rect 14858 38557 14876 38621
rect 14940 38557 15000 38621
rect 0 38540 15000 38557
rect 0 38476 111 38540
rect 175 38476 191 38540
rect 255 38476 271 38540
rect 335 38476 351 38540
rect 415 38476 431 38540
rect 495 38476 511 38540
rect 575 38476 591 38540
rect 655 38476 671 38540
rect 735 38476 751 38540
rect 815 38476 831 38540
rect 895 38476 911 38540
rect 975 38476 991 38540
rect 1055 38476 1071 38540
rect 1135 38476 1151 38540
rect 1215 38476 1231 38540
rect 1295 38476 1311 38540
rect 1375 38476 1391 38540
rect 1455 38476 1471 38540
rect 1535 38476 1551 38540
rect 1615 38476 1631 38540
rect 1695 38476 1711 38540
rect 1775 38476 1791 38540
rect 1855 38476 1871 38540
rect 1935 38476 1951 38540
rect 2015 38476 2031 38540
rect 2095 38476 2111 38540
rect 2175 38476 2191 38540
rect 2255 38476 2271 38540
rect 2335 38476 2351 38540
rect 2415 38476 2431 38540
rect 2495 38476 2511 38540
rect 2575 38476 12416 38540
rect 12480 38476 12498 38540
rect 12562 38476 12580 38540
rect 12644 38476 12662 38540
rect 12726 38476 12744 38540
rect 12808 38476 12826 38540
rect 12890 38476 12908 38540
rect 12972 38476 12990 38540
rect 13054 38476 13072 38540
rect 13136 38476 13154 38540
rect 13218 38476 13236 38540
rect 13300 38476 13318 38540
rect 13382 38476 13400 38540
rect 13464 38476 13482 38540
rect 13546 38476 13564 38540
rect 13628 38476 13646 38540
rect 13710 38476 13728 38540
rect 13792 38476 13810 38540
rect 13874 38476 13892 38540
rect 13956 38476 13974 38540
rect 14038 38476 14056 38540
rect 14120 38476 14138 38540
rect 14202 38476 14220 38540
rect 14284 38476 14302 38540
rect 14366 38476 14384 38540
rect 14448 38476 14466 38540
rect 14530 38476 14548 38540
rect 14612 38476 14630 38540
rect 14694 38476 14712 38540
rect 14776 38476 14794 38540
rect 14858 38476 14876 38540
rect 14940 38476 15000 38540
rect 0 38459 15000 38476
rect 0 38395 111 38459
rect 175 38395 191 38459
rect 255 38395 271 38459
rect 335 38395 351 38459
rect 415 38395 431 38459
rect 495 38395 511 38459
rect 575 38395 591 38459
rect 655 38395 671 38459
rect 735 38395 751 38459
rect 815 38395 831 38459
rect 895 38395 911 38459
rect 975 38395 991 38459
rect 1055 38395 1071 38459
rect 1135 38395 1151 38459
rect 1215 38395 1231 38459
rect 1295 38395 1311 38459
rect 1375 38395 1391 38459
rect 1455 38395 1471 38459
rect 1535 38395 1551 38459
rect 1615 38395 1631 38459
rect 1695 38395 1711 38459
rect 1775 38395 1791 38459
rect 1855 38395 1871 38459
rect 1935 38395 1951 38459
rect 2015 38395 2031 38459
rect 2095 38395 2111 38459
rect 2175 38395 2191 38459
rect 2255 38395 2271 38459
rect 2335 38395 2351 38459
rect 2415 38395 2431 38459
rect 2495 38395 2511 38459
rect 2575 38395 12416 38459
rect 12480 38395 12498 38459
rect 12562 38395 12580 38459
rect 12644 38395 12662 38459
rect 12726 38395 12744 38459
rect 12808 38395 12826 38459
rect 12890 38395 12908 38459
rect 12972 38395 12990 38459
rect 13054 38395 13072 38459
rect 13136 38395 13154 38459
rect 13218 38395 13236 38459
rect 13300 38395 13318 38459
rect 13382 38395 13400 38459
rect 13464 38395 13482 38459
rect 13546 38395 13564 38459
rect 13628 38395 13646 38459
rect 13710 38395 13728 38459
rect 13792 38395 13810 38459
rect 13874 38395 13892 38459
rect 13956 38395 13974 38459
rect 14038 38395 14056 38459
rect 14120 38395 14138 38459
rect 14202 38395 14220 38459
rect 14284 38395 14302 38459
rect 14366 38395 14384 38459
rect 14448 38395 14466 38459
rect 14530 38395 14548 38459
rect 14612 38395 14630 38459
rect 14694 38395 14712 38459
rect 14776 38395 14794 38459
rect 14858 38395 14876 38459
rect 14940 38395 15000 38459
rect 0 38378 15000 38395
rect 0 38314 111 38378
rect 175 38314 191 38378
rect 255 38314 271 38378
rect 335 38314 351 38378
rect 415 38314 431 38378
rect 495 38314 511 38378
rect 575 38314 591 38378
rect 655 38314 671 38378
rect 735 38314 751 38378
rect 815 38314 831 38378
rect 895 38314 911 38378
rect 975 38314 991 38378
rect 1055 38314 1071 38378
rect 1135 38314 1151 38378
rect 1215 38314 1231 38378
rect 1295 38314 1311 38378
rect 1375 38314 1391 38378
rect 1455 38314 1471 38378
rect 1535 38314 1551 38378
rect 1615 38314 1631 38378
rect 1695 38314 1711 38378
rect 1775 38314 1791 38378
rect 1855 38314 1871 38378
rect 1935 38314 1951 38378
rect 2015 38314 2031 38378
rect 2095 38314 2111 38378
rect 2175 38314 2191 38378
rect 2255 38314 2271 38378
rect 2335 38314 2351 38378
rect 2415 38314 2431 38378
rect 2495 38314 2511 38378
rect 2575 38314 12416 38378
rect 12480 38314 12498 38378
rect 12562 38314 12580 38378
rect 12644 38314 12662 38378
rect 12726 38314 12744 38378
rect 12808 38314 12826 38378
rect 12890 38314 12908 38378
rect 12972 38314 12990 38378
rect 13054 38314 13072 38378
rect 13136 38314 13154 38378
rect 13218 38314 13236 38378
rect 13300 38314 13318 38378
rect 13382 38314 13400 38378
rect 13464 38314 13482 38378
rect 13546 38314 13564 38378
rect 13628 38314 13646 38378
rect 13710 38314 13728 38378
rect 13792 38314 13810 38378
rect 13874 38314 13892 38378
rect 13956 38314 13974 38378
rect 14038 38314 14056 38378
rect 14120 38314 14138 38378
rect 14202 38314 14220 38378
rect 14284 38314 14302 38378
rect 14366 38314 14384 38378
rect 14448 38314 14466 38378
rect 14530 38314 14548 38378
rect 14612 38314 14630 38378
rect 14694 38314 14712 38378
rect 14776 38314 14794 38378
rect 14858 38314 14876 38378
rect 14940 38314 15000 38378
rect 0 38297 15000 38314
rect 0 38233 111 38297
rect 175 38233 191 38297
rect 255 38233 271 38297
rect 335 38233 351 38297
rect 415 38233 431 38297
rect 495 38233 511 38297
rect 575 38233 591 38297
rect 655 38233 671 38297
rect 735 38233 751 38297
rect 815 38233 831 38297
rect 895 38233 911 38297
rect 975 38233 991 38297
rect 1055 38233 1071 38297
rect 1135 38233 1151 38297
rect 1215 38233 1231 38297
rect 1295 38233 1311 38297
rect 1375 38233 1391 38297
rect 1455 38233 1471 38297
rect 1535 38233 1551 38297
rect 1615 38233 1631 38297
rect 1695 38233 1711 38297
rect 1775 38233 1791 38297
rect 1855 38233 1871 38297
rect 1935 38233 1951 38297
rect 2015 38233 2031 38297
rect 2095 38233 2111 38297
rect 2175 38233 2191 38297
rect 2255 38233 2271 38297
rect 2335 38233 2351 38297
rect 2415 38233 2431 38297
rect 2495 38233 2511 38297
rect 2575 38233 12416 38297
rect 12480 38233 12498 38297
rect 12562 38233 12580 38297
rect 12644 38233 12662 38297
rect 12726 38233 12744 38297
rect 12808 38233 12826 38297
rect 12890 38233 12908 38297
rect 12972 38233 12990 38297
rect 13054 38233 13072 38297
rect 13136 38233 13154 38297
rect 13218 38233 13236 38297
rect 13300 38233 13318 38297
rect 13382 38233 13400 38297
rect 13464 38233 13482 38297
rect 13546 38233 13564 38297
rect 13628 38233 13646 38297
rect 13710 38233 13728 38297
rect 13792 38233 13810 38297
rect 13874 38233 13892 38297
rect 13956 38233 13974 38297
rect 14038 38233 14056 38297
rect 14120 38233 14138 38297
rect 14202 38233 14220 38297
rect 14284 38233 14302 38297
rect 14366 38233 14384 38297
rect 14448 38233 14466 38297
rect 14530 38233 14548 38297
rect 14612 38233 14630 38297
rect 14694 38233 14712 38297
rect 14776 38233 14794 38297
rect 14858 38233 14876 38297
rect 14940 38233 15000 38297
rect 0 38216 15000 38233
rect 0 38152 111 38216
rect 175 38152 191 38216
rect 255 38152 271 38216
rect 335 38152 351 38216
rect 415 38152 431 38216
rect 495 38152 511 38216
rect 575 38152 591 38216
rect 655 38152 671 38216
rect 735 38152 751 38216
rect 815 38152 831 38216
rect 895 38152 911 38216
rect 975 38152 991 38216
rect 1055 38152 1071 38216
rect 1135 38152 1151 38216
rect 1215 38152 1231 38216
rect 1295 38152 1311 38216
rect 1375 38152 1391 38216
rect 1455 38152 1471 38216
rect 1535 38152 1551 38216
rect 1615 38152 1631 38216
rect 1695 38152 1711 38216
rect 1775 38152 1791 38216
rect 1855 38152 1871 38216
rect 1935 38152 1951 38216
rect 2015 38152 2031 38216
rect 2095 38152 2111 38216
rect 2175 38152 2191 38216
rect 2255 38152 2271 38216
rect 2335 38152 2351 38216
rect 2415 38152 2431 38216
rect 2495 38152 2511 38216
rect 2575 38152 12416 38216
rect 12480 38152 12498 38216
rect 12562 38152 12580 38216
rect 12644 38152 12662 38216
rect 12726 38152 12744 38216
rect 12808 38152 12826 38216
rect 12890 38152 12908 38216
rect 12972 38152 12990 38216
rect 13054 38152 13072 38216
rect 13136 38152 13154 38216
rect 13218 38152 13236 38216
rect 13300 38152 13318 38216
rect 13382 38152 13400 38216
rect 13464 38152 13482 38216
rect 13546 38152 13564 38216
rect 13628 38152 13646 38216
rect 13710 38152 13728 38216
rect 13792 38152 13810 38216
rect 13874 38152 13892 38216
rect 13956 38152 13974 38216
rect 14038 38152 14056 38216
rect 14120 38152 14138 38216
rect 14202 38152 14220 38216
rect 14284 38152 14302 38216
rect 14366 38152 14384 38216
rect 14448 38152 14466 38216
rect 14530 38152 14548 38216
rect 14612 38152 14630 38216
rect 14694 38152 14712 38216
rect 14776 38152 14794 38216
rect 14858 38152 14876 38216
rect 14940 38152 15000 38216
rect 0 38135 15000 38152
rect 0 38071 111 38135
rect 175 38071 191 38135
rect 255 38071 271 38135
rect 335 38071 351 38135
rect 415 38071 431 38135
rect 495 38071 511 38135
rect 575 38071 591 38135
rect 655 38071 671 38135
rect 735 38071 751 38135
rect 815 38071 831 38135
rect 895 38071 911 38135
rect 975 38071 991 38135
rect 1055 38071 1071 38135
rect 1135 38071 1151 38135
rect 1215 38071 1231 38135
rect 1295 38071 1311 38135
rect 1375 38071 1391 38135
rect 1455 38071 1471 38135
rect 1535 38071 1551 38135
rect 1615 38071 1631 38135
rect 1695 38071 1711 38135
rect 1775 38071 1791 38135
rect 1855 38071 1871 38135
rect 1935 38071 1951 38135
rect 2015 38071 2031 38135
rect 2095 38071 2111 38135
rect 2175 38071 2191 38135
rect 2255 38071 2271 38135
rect 2335 38071 2351 38135
rect 2415 38071 2431 38135
rect 2495 38071 2511 38135
rect 2575 38071 12416 38135
rect 12480 38071 12498 38135
rect 12562 38071 12580 38135
rect 12644 38071 12662 38135
rect 12726 38071 12744 38135
rect 12808 38071 12826 38135
rect 12890 38071 12908 38135
rect 12972 38071 12990 38135
rect 13054 38071 13072 38135
rect 13136 38071 13154 38135
rect 13218 38071 13236 38135
rect 13300 38071 13318 38135
rect 13382 38071 13400 38135
rect 13464 38071 13482 38135
rect 13546 38071 13564 38135
rect 13628 38071 13646 38135
rect 13710 38071 13728 38135
rect 13792 38071 13810 38135
rect 13874 38071 13892 38135
rect 13956 38071 13974 38135
rect 14038 38071 14056 38135
rect 14120 38071 14138 38135
rect 14202 38071 14220 38135
rect 14284 38071 14302 38135
rect 14366 38071 14384 38135
rect 14448 38071 14466 38135
rect 14530 38071 14548 38135
rect 14612 38071 14630 38135
rect 14694 38071 14712 38135
rect 14776 38071 14794 38135
rect 14858 38071 14876 38135
rect 14940 38071 15000 38135
rect 0 38054 15000 38071
rect 0 37990 111 38054
rect 175 37990 191 38054
rect 255 37990 271 38054
rect 335 37990 351 38054
rect 415 37990 431 38054
rect 495 37990 511 38054
rect 575 37990 591 38054
rect 655 37990 671 38054
rect 735 37990 751 38054
rect 815 37990 831 38054
rect 895 37990 911 38054
rect 975 37990 991 38054
rect 1055 37990 1071 38054
rect 1135 37990 1151 38054
rect 1215 37990 1231 38054
rect 1295 37990 1311 38054
rect 1375 37990 1391 38054
rect 1455 37990 1471 38054
rect 1535 37990 1551 38054
rect 1615 37990 1631 38054
rect 1695 37990 1711 38054
rect 1775 37990 1791 38054
rect 1855 37990 1871 38054
rect 1935 37990 1951 38054
rect 2015 37990 2031 38054
rect 2095 37990 2111 38054
rect 2175 37990 2191 38054
rect 2255 37990 2271 38054
rect 2335 37990 2351 38054
rect 2415 37990 2431 38054
rect 2495 37990 2511 38054
rect 2575 37990 12416 38054
rect 12480 37990 12498 38054
rect 12562 37990 12580 38054
rect 12644 37990 12662 38054
rect 12726 37990 12744 38054
rect 12808 37990 12826 38054
rect 12890 37990 12908 38054
rect 12972 37990 12990 38054
rect 13054 37990 13072 38054
rect 13136 37990 13154 38054
rect 13218 37990 13236 38054
rect 13300 37990 13318 38054
rect 13382 37990 13400 38054
rect 13464 37990 13482 38054
rect 13546 37990 13564 38054
rect 13628 37990 13646 38054
rect 13710 37990 13728 38054
rect 13792 37990 13810 38054
rect 13874 37990 13892 38054
rect 13956 37990 13974 38054
rect 14038 37990 14056 38054
rect 14120 37990 14138 38054
rect 14202 37990 14220 38054
rect 14284 37990 14302 38054
rect 14366 37990 14384 38054
rect 14448 37990 14466 38054
rect 14530 37990 14548 38054
rect 14612 37990 14630 38054
rect 14694 37990 14712 38054
rect 14776 37990 14794 38054
rect 14858 37990 14876 38054
rect 14940 37990 15000 38054
rect 0 37973 15000 37990
rect 0 37909 111 37973
rect 175 37909 191 37973
rect 255 37909 271 37973
rect 335 37909 351 37973
rect 415 37909 431 37973
rect 495 37909 511 37973
rect 575 37909 591 37973
rect 655 37909 671 37973
rect 735 37909 751 37973
rect 815 37909 831 37973
rect 895 37909 911 37973
rect 975 37909 991 37973
rect 1055 37909 1071 37973
rect 1135 37909 1151 37973
rect 1215 37909 1231 37973
rect 1295 37909 1311 37973
rect 1375 37909 1391 37973
rect 1455 37909 1471 37973
rect 1535 37909 1551 37973
rect 1615 37909 1631 37973
rect 1695 37909 1711 37973
rect 1775 37909 1791 37973
rect 1855 37909 1871 37973
rect 1935 37909 1951 37973
rect 2015 37909 2031 37973
rect 2095 37909 2111 37973
rect 2175 37909 2191 37973
rect 2255 37909 2271 37973
rect 2335 37909 2351 37973
rect 2415 37909 2431 37973
rect 2495 37909 2511 37973
rect 2575 37909 12416 37973
rect 12480 37909 12498 37973
rect 12562 37909 12580 37973
rect 12644 37909 12662 37973
rect 12726 37909 12744 37973
rect 12808 37909 12826 37973
rect 12890 37909 12908 37973
rect 12972 37909 12990 37973
rect 13054 37909 13072 37973
rect 13136 37909 13154 37973
rect 13218 37909 13236 37973
rect 13300 37909 13318 37973
rect 13382 37909 13400 37973
rect 13464 37909 13482 37973
rect 13546 37909 13564 37973
rect 13628 37909 13646 37973
rect 13710 37909 13728 37973
rect 13792 37909 13810 37973
rect 13874 37909 13892 37973
rect 13956 37909 13974 37973
rect 14038 37909 14056 37973
rect 14120 37909 14138 37973
rect 14202 37909 14220 37973
rect 14284 37909 14302 37973
rect 14366 37909 14384 37973
rect 14448 37909 14466 37973
rect 14530 37909 14548 37973
rect 14612 37909 14630 37973
rect 14694 37909 14712 37973
rect 14776 37909 14794 37973
rect 14858 37909 14876 37973
rect 14940 37909 15000 37973
rect 0 37892 15000 37909
rect 0 37828 111 37892
rect 175 37828 191 37892
rect 255 37828 271 37892
rect 335 37828 351 37892
rect 415 37828 431 37892
rect 495 37828 511 37892
rect 575 37828 591 37892
rect 655 37828 671 37892
rect 735 37828 751 37892
rect 815 37828 831 37892
rect 895 37828 911 37892
rect 975 37828 991 37892
rect 1055 37828 1071 37892
rect 1135 37828 1151 37892
rect 1215 37828 1231 37892
rect 1295 37828 1311 37892
rect 1375 37828 1391 37892
rect 1455 37828 1471 37892
rect 1535 37828 1551 37892
rect 1615 37828 1631 37892
rect 1695 37828 1711 37892
rect 1775 37828 1791 37892
rect 1855 37828 1871 37892
rect 1935 37828 1951 37892
rect 2015 37828 2031 37892
rect 2095 37828 2111 37892
rect 2175 37828 2191 37892
rect 2255 37828 2271 37892
rect 2335 37828 2351 37892
rect 2415 37828 2431 37892
rect 2495 37828 2511 37892
rect 2575 37828 12416 37892
rect 12480 37828 12498 37892
rect 12562 37828 12580 37892
rect 12644 37828 12662 37892
rect 12726 37828 12744 37892
rect 12808 37828 12826 37892
rect 12890 37828 12908 37892
rect 12972 37828 12990 37892
rect 13054 37828 13072 37892
rect 13136 37828 13154 37892
rect 13218 37828 13236 37892
rect 13300 37828 13318 37892
rect 13382 37828 13400 37892
rect 13464 37828 13482 37892
rect 13546 37828 13564 37892
rect 13628 37828 13646 37892
rect 13710 37828 13728 37892
rect 13792 37828 13810 37892
rect 13874 37828 13892 37892
rect 13956 37828 13974 37892
rect 14038 37828 14056 37892
rect 14120 37828 14138 37892
rect 14202 37828 14220 37892
rect 14284 37828 14302 37892
rect 14366 37828 14384 37892
rect 14448 37828 14466 37892
rect 14530 37828 14548 37892
rect 14612 37828 14630 37892
rect 14694 37828 14712 37892
rect 14776 37828 14794 37892
rect 14858 37828 14876 37892
rect 14940 37828 15000 37892
rect 0 37811 15000 37828
rect 0 37747 111 37811
rect 175 37747 191 37811
rect 255 37747 271 37811
rect 335 37747 351 37811
rect 415 37747 431 37811
rect 495 37747 511 37811
rect 575 37747 591 37811
rect 655 37747 671 37811
rect 735 37747 751 37811
rect 815 37747 831 37811
rect 895 37747 911 37811
rect 975 37747 991 37811
rect 1055 37747 1071 37811
rect 1135 37747 1151 37811
rect 1215 37747 1231 37811
rect 1295 37747 1311 37811
rect 1375 37747 1391 37811
rect 1455 37747 1471 37811
rect 1535 37747 1551 37811
rect 1615 37747 1631 37811
rect 1695 37747 1711 37811
rect 1775 37747 1791 37811
rect 1855 37747 1871 37811
rect 1935 37747 1951 37811
rect 2015 37747 2031 37811
rect 2095 37747 2111 37811
rect 2175 37747 2191 37811
rect 2255 37747 2271 37811
rect 2335 37747 2351 37811
rect 2415 37747 2431 37811
rect 2495 37747 2511 37811
rect 2575 37747 12416 37811
rect 12480 37747 12498 37811
rect 12562 37747 12580 37811
rect 12644 37747 12662 37811
rect 12726 37747 12744 37811
rect 12808 37747 12826 37811
rect 12890 37747 12908 37811
rect 12972 37747 12990 37811
rect 13054 37747 13072 37811
rect 13136 37747 13154 37811
rect 13218 37747 13236 37811
rect 13300 37747 13318 37811
rect 13382 37747 13400 37811
rect 13464 37747 13482 37811
rect 13546 37747 13564 37811
rect 13628 37747 13646 37811
rect 13710 37747 13728 37811
rect 13792 37747 13810 37811
rect 13874 37747 13892 37811
rect 13956 37747 13974 37811
rect 14038 37747 14056 37811
rect 14120 37747 14138 37811
rect 14202 37747 14220 37811
rect 14284 37747 14302 37811
rect 14366 37747 14384 37811
rect 14448 37747 14466 37811
rect 14530 37747 14548 37811
rect 14612 37747 14630 37811
rect 14694 37747 14712 37811
rect 14776 37747 14794 37811
rect 14858 37747 14876 37811
rect 14940 37747 15000 37811
rect 0 37730 15000 37747
rect 0 37666 111 37730
rect 175 37666 191 37730
rect 255 37666 271 37730
rect 335 37666 351 37730
rect 415 37666 431 37730
rect 495 37666 511 37730
rect 575 37666 591 37730
rect 655 37666 671 37730
rect 735 37666 751 37730
rect 815 37666 831 37730
rect 895 37666 911 37730
rect 975 37666 991 37730
rect 1055 37666 1071 37730
rect 1135 37666 1151 37730
rect 1215 37666 1231 37730
rect 1295 37666 1311 37730
rect 1375 37666 1391 37730
rect 1455 37666 1471 37730
rect 1535 37666 1551 37730
rect 1615 37666 1631 37730
rect 1695 37666 1711 37730
rect 1775 37666 1791 37730
rect 1855 37666 1871 37730
rect 1935 37666 1951 37730
rect 2015 37666 2031 37730
rect 2095 37666 2111 37730
rect 2175 37666 2191 37730
rect 2255 37666 2271 37730
rect 2335 37666 2351 37730
rect 2415 37666 2431 37730
rect 2495 37666 2511 37730
rect 2575 37666 12416 37730
rect 12480 37666 12498 37730
rect 12562 37666 12580 37730
rect 12644 37666 12662 37730
rect 12726 37666 12744 37730
rect 12808 37666 12826 37730
rect 12890 37666 12908 37730
rect 12972 37666 12990 37730
rect 13054 37666 13072 37730
rect 13136 37666 13154 37730
rect 13218 37666 13236 37730
rect 13300 37666 13318 37730
rect 13382 37666 13400 37730
rect 13464 37666 13482 37730
rect 13546 37666 13564 37730
rect 13628 37666 13646 37730
rect 13710 37666 13728 37730
rect 13792 37666 13810 37730
rect 13874 37666 13892 37730
rect 13956 37666 13974 37730
rect 14038 37666 14056 37730
rect 14120 37666 14138 37730
rect 14202 37666 14220 37730
rect 14284 37666 14302 37730
rect 14366 37666 14384 37730
rect 14448 37666 14466 37730
rect 14530 37666 14548 37730
rect 14612 37666 14630 37730
rect 14694 37666 14712 37730
rect 14776 37666 14794 37730
rect 14858 37666 14876 37730
rect 14940 37666 15000 37730
rect 0 37649 15000 37666
rect 0 37585 111 37649
rect 175 37585 191 37649
rect 255 37585 271 37649
rect 335 37585 351 37649
rect 415 37585 431 37649
rect 495 37585 511 37649
rect 575 37585 591 37649
rect 655 37585 671 37649
rect 735 37585 751 37649
rect 815 37585 831 37649
rect 895 37585 911 37649
rect 975 37585 991 37649
rect 1055 37585 1071 37649
rect 1135 37585 1151 37649
rect 1215 37585 1231 37649
rect 1295 37585 1311 37649
rect 1375 37585 1391 37649
rect 1455 37585 1471 37649
rect 1535 37585 1551 37649
rect 1615 37585 1631 37649
rect 1695 37585 1711 37649
rect 1775 37585 1791 37649
rect 1855 37585 1871 37649
rect 1935 37585 1951 37649
rect 2015 37585 2031 37649
rect 2095 37585 2111 37649
rect 2175 37585 2191 37649
rect 2255 37585 2271 37649
rect 2335 37585 2351 37649
rect 2415 37585 2431 37649
rect 2495 37585 2511 37649
rect 2575 37585 12416 37649
rect 12480 37585 12498 37649
rect 12562 37585 12580 37649
rect 12644 37585 12662 37649
rect 12726 37585 12744 37649
rect 12808 37585 12826 37649
rect 12890 37585 12908 37649
rect 12972 37585 12990 37649
rect 13054 37585 13072 37649
rect 13136 37585 13154 37649
rect 13218 37585 13236 37649
rect 13300 37585 13318 37649
rect 13382 37585 13400 37649
rect 13464 37585 13482 37649
rect 13546 37585 13564 37649
rect 13628 37585 13646 37649
rect 13710 37585 13728 37649
rect 13792 37585 13810 37649
rect 13874 37585 13892 37649
rect 13956 37585 13974 37649
rect 14038 37585 14056 37649
rect 14120 37585 14138 37649
rect 14202 37585 14220 37649
rect 14284 37585 14302 37649
rect 14366 37585 14384 37649
rect 14448 37585 14466 37649
rect 14530 37585 14548 37649
rect 14612 37585 14630 37649
rect 14694 37585 14712 37649
rect 14776 37585 14794 37649
rect 14858 37585 14876 37649
rect 14940 37585 15000 37649
rect 0 37568 15000 37585
rect 0 37504 111 37568
rect 175 37504 191 37568
rect 255 37504 271 37568
rect 335 37504 351 37568
rect 415 37504 431 37568
rect 495 37504 511 37568
rect 575 37504 591 37568
rect 655 37504 671 37568
rect 735 37504 751 37568
rect 815 37504 831 37568
rect 895 37504 911 37568
rect 975 37504 991 37568
rect 1055 37504 1071 37568
rect 1135 37504 1151 37568
rect 1215 37504 1231 37568
rect 1295 37504 1311 37568
rect 1375 37504 1391 37568
rect 1455 37504 1471 37568
rect 1535 37504 1551 37568
rect 1615 37504 1631 37568
rect 1695 37504 1711 37568
rect 1775 37504 1791 37568
rect 1855 37504 1871 37568
rect 1935 37504 1951 37568
rect 2015 37504 2031 37568
rect 2095 37504 2111 37568
rect 2175 37504 2191 37568
rect 2255 37504 2271 37568
rect 2335 37504 2351 37568
rect 2415 37504 2431 37568
rect 2495 37504 2511 37568
rect 2575 37504 12416 37568
rect 12480 37504 12498 37568
rect 12562 37504 12580 37568
rect 12644 37504 12662 37568
rect 12726 37504 12744 37568
rect 12808 37504 12826 37568
rect 12890 37504 12908 37568
rect 12972 37504 12990 37568
rect 13054 37504 13072 37568
rect 13136 37504 13154 37568
rect 13218 37504 13236 37568
rect 13300 37504 13318 37568
rect 13382 37504 13400 37568
rect 13464 37504 13482 37568
rect 13546 37504 13564 37568
rect 13628 37504 13646 37568
rect 13710 37504 13728 37568
rect 13792 37504 13810 37568
rect 13874 37504 13892 37568
rect 13956 37504 13974 37568
rect 14038 37504 14056 37568
rect 14120 37504 14138 37568
rect 14202 37504 14220 37568
rect 14284 37504 14302 37568
rect 14366 37504 14384 37568
rect 14448 37504 14466 37568
rect 14530 37504 14548 37568
rect 14612 37504 14630 37568
rect 14694 37504 14712 37568
rect 14776 37504 14794 37568
rect 14858 37504 14876 37568
rect 14940 37504 15000 37568
rect 0 37487 15000 37504
rect 0 37423 111 37487
rect 175 37423 191 37487
rect 255 37423 271 37487
rect 335 37423 351 37487
rect 415 37423 431 37487
rect 495 37423 511 37487
rect 575 37423 591 37487
rect 655 37423 671 37487
rect 735 37423 751 37487
rect 815 37423 831 37487
rect 895 37423 911 37487
rect 975 37423 991 37487
rect 1055 37423 1071 37487
rect 1135 37423 1151 37487
rect 1215 37423 1231 37487
rect 1295 37423 1311 37487
rect 1375 37423 1391 37487
rect 1455 37423 1471 37487
rect 1535 37423 1551 37487
rect 1615 37423 1631 37487
rect 1695 37423 1711 37487
rect 1775 37423 1791 37487
rect 1855 37423 1871 37487
rect 1935 37423 1951 37487
rect 2015 37423 2031 37487
rect 2095 37423 2111 37487
rect 2175 37423 2191 37487
rect 2255 37423 2271 37487
rect 2335 37423 2351 37487
rect 2415 37423 2431 37487
rect 2495 37423 2511 37487
rect 2575 37423 12416 37487
rect 12480 37423 12498 37487
rect 12562 37423 12580 37487
rect 12644 37423 12662 37487
rect 12726 37423 12744 37487
rect 12808 37423 12826 37487
rect 12890 37423 12908 37487
rect 12972 37423 12990 37487
rect 13054 37423 13072 37487
rect 13136 37423 13154 37487
rect 13218 37423 13236 37487
rect 13300 37423 13318 37487
rect 13382 37423 13400 37487
rect 13464 37423 13482 37487
rect 13546 37423 13564 37487
rect 13628 37423 13646 37487
rect 13710 37423 13728 37487
rect 13792 37423 13810 37487
rect 13874 37423 13892 37487
rect 13956 37423 13974 37487
rect 14038 37423 14056 37487
rect 14120 37423 14138 37487
rect 14202 37423 14220 37487
rect 14284 37423 14302 37487
rect 14366 37423 14384 37487
rect 14448 37423 14466 37487
rect 14530 37423 14548 37487
rect 14612 37423 14630 37487
rect 14694 37423 14712 37487
rect 14776 37423 14794 37487
rect 14858 37423 14876 37487
rect 14940 37423 15000 37487
rect 0 37406 15000 37423
rect 0 37342 111 37406
rect 175 37342 191 37406
rect 255 37342 271 37406
rect 335 37342 351 37406
rect 415 37342 431 37406
rect 495 37342 511 37406
rect 575 37342 591 37406
rect 655 37342 671 37406
rect 735 37342 751 37406
rect 815 37342 831 37406
rect 895 37342 911 37406
rect 975 37342 991 37406
rect 1055 37342 1071 37406
rect 1135 37342 1151 37406
rect 1215 37342 1231 37406
rect 1295 37342 1311 37406
rect 1375 37342 1391 37406
rect 1455 37342 1471 37406
rect 1535 37342 1551 37406
rect 1615 37342 1631 37406
rect 1695 37342 1711 37406
rect 1775 37342 1791 37406
rect 1855 37342 1871 37406
rect 1935 37342 1951 37406
rect 2015 37342 2031 37406
rect 2095 37342 2111 37406
rect 2175 37342 2191 37406
rect 2255 37342 2271 37406
rect 2335 37342 2351 37406
rect 2415 37342 2431 37406
rect 2495 37342 2511 37406
rect 2575 37342 12416 37406
rect 12480 37342 12498 37406
rect 12562 37342 12580 37406
rect 12644 37342 12662 37406
rect 12726 37342 12744 37406
rect 12808 37342 12826 37406
rect 12890 37342 12908 37406
rect 12972 37342 12990 37406
rect 13054 37342 13072 37406
rect 13136 37342 13154 37406
rect 13218 37342 13236 37406
rect 13300 37342 13318 37406
rect 13382 37342 13400 37406
rect 13464 37342 13482 37406
rect 13546 37342 13564 37406
rect 13628 37342 13646 37406
rect 13710 37342 13728 37406
rect 13792 37342 13810 37406
rect 13874 37342 13892 37406
rect 13956 37342 13974 37406
rect 14038 37342 14056 37406
rect 14120 37342 14138 37406
rect 14202 37342 14220 37406
rect 14284 37342 14302 37406
rect 14366 37342 14384 37406
rect 14448 37342 14466 37406
rect 14530 37342 14548 37406
rect 14612 37342 14630 37406
rect 14694 37342 14712 37406
rect 14776 37342 14794 37406
rect 14858 37342 14876 37406
rect 14940 37342 15000 37406
rect 0 37325 15000 37342
rect 0 37261 111 37325
rect 175 37261 191 37325
rect 255 37261 271 37325
rect 335 37261 351 37325
rect 415 37261 431 37325
rect 495 37261 511 37325
rect 575 37261 591 37325
rect 655 37261 671 37325
rect 735 37261 751 37325
rect 815 37261 831 37325
rect 895 37261 911 37325
rect 975 37261 991 37325
rect 1055 37261 1071 37325
rect 1135 37261 1151 37325
rect 1215 37261 1231 37325
rect 1295 37261 1311 37325
rect 1375 37261 1391 37325
rect 1455 37261 1471 37325
rect 1535 37261 1551 37325
rect 1615 37261 1631 37325
rect 1695 37261 1711 37325
rect 1775 37261 1791 37325
rect 1855 37261 1871 37325
rect 1935 37261 1951 37325
rect 2015 37261 2031 37325
rect 2095 37261 2111 37325
rect 2175 37261 2191 37325
rect 2255 37261 2271 37325
rect 2335 37261 2351 37325
rect 2415 37261 2431 37325
rect 2495 37261 2511 37325
rect 2575 37261 12416 37325
rect 12480 37261 12498 37325
rect 12562 37261 12580 37325
rect 12644 37261 12662 37325
rect 12726 37261 12744 37325
rect 12808 37261 12826 37325
rect 12890 37261 12908 37325
rect 12972 37261 12990 37325
rect 13054 37261 13072 37325
rect 13136 37261 13154 37325
rect 13218 37261 13236 37325
rect 13300 37261 13318 37325
rect 13382 37261 13400 37325
rect 13464 37261 13482 37325
rect 13546 37261 13564 37325
rect 13628 37261 13646 37325
rect 13710 37261 13728 37325
rect 13792 37261 13810 37325
rect 13874 37261 13892 37325
rect 13956 37261 13974 37325
rect 14038 37261 14056 37325
rect 14120 37261 14138 37325
rect 14202 37261 14220 37325
rect 14284 37261 14302 37325
rect 14366 37261 14384 37325
rect 14448 37261 14466 37325
rect 14530 37261 14548 37325
rect 14612 37261 14630 37325
rect 14694 37261 14712 37325
rect 14776 37261 14794 37325
rect 14858 37261 14876 37325
rect 14940 37261 15000 37325
rect 0 37244 15000 37261
rect 0 37180 111 37244
rect 175 37180 191 37244
rect 255 37180 271 37244
rect 335 37180 351 37244
rect 415 37180 431 37244
rect 495 37180 511 37244
rect 575 37180 591 37244
rect 655 37180 671 37244
rect 735 37180 751 37244
rect 815 37180 831 37244
rect 895 37180 911 37244
rect 975 37180 991 37244
rect 1055 37180 1071 37244
rect 1135 37180 1151 37244
rect 1215 37180 1231 37244
rect 1295 37180 1311 37244
rect 1375 37180 1391 37244
rect 1455 37180 1471 37244
rect 1535 37180 1551 37244
rect 1615 37180 1631 37244
rect 1695 37180 1711 37244
rect 1775 37180 1791 37244
rect 1855 37180 1871 37244
rect 1935 37180 1951 37244
rect 2015 37180 2031 37244
rect 2095 37180 2111 37244
rect 2175 37180 2191 37244
rect 2255 37180 2271 37244
rect 2335 37180 2351 37244
rect 2415 37180 2431 37244
rect 2495 37180 2511 37244
rect 2575 37180 12416 37244
rect 12480 37180 12498 37244
rect 12562 37180 12580 37244
rect 12644 37180 12662 37244
rect 12726 37180 12744 37244
rect 12808 37180 12826 37244
rect 12890 37180 12908 37244
rect 12972 37180 12990 37244
rect 13054 37180 13072 37244
rect 13136 37180 13154 37244
rect 13218 37180 13236 37244
rect 13300 37180 13318 37244
rect 13382 37180 13400 37244
rect 13464 37180 13482 37244
rect 13546 37180 13564 37244
rect 13628 37180 13646 37244
rect 13710 37180 13728 37244
rect 13792 37180 13810 37244
rect 13874 37180 13892 37244
rect 13956 37180 13974 37244
rect 14038 37180 14056 37244
rect 14120 37180 14138 37244
rect 14202 37180 14220 37244
rect 14284 37180 14302 37244
rect 14366 37180 14384 37244
rect 14448 37180 14466 37244
rect 14530 37180 14548 37244
rect 14612 37180 14630 37244
rect 14694 37180 14712 37244
rect 14776 37180 14794 37244
rect 14858 37180 14876 37244
rect 14940 37180 15000 37244
rect 0 37163 15000 37180
rect 0 37099 111 37163
rect 175 37099 191 37163
rect 255 37099 271 37163
rect 335 37099 351 37163
rect 415 37099 431 37163
rect 495 37099 511 37163
rect 575 37099 591 37163
rect 655 37099 671 37163
rect 735 37099 751 37163
rect 815 37099 831 37163
rect 895 37099 911 37163
rect 975 37099 991 37163
rect 1055 37099 1071 37163
rect 1135 37099 1151 37163
rect 1215 37099 1231 37163
rect 1295 37099 1311 37163
rect 1375 37099 1391 37163
rect 1455 37099 1471 37163
rect 1535 37099 1551 37163
rect 1615 37099 1631 37163
rect 1695 37099 1711 37163
rect 1775 37099 1791 37163
rect 1855 37099 1871 37163
rect 1935 37099 1951 37163
rect 2015 37099 2031 37163
rect 2095 37099 2111 37163
rect 2175 37099 2191 37163
rect 2255 37099 2271 37163
rect 2335 37099 2351 37163
rect 2415 37099 2431 37163
rect 2495 37099 2511 37163
rect 2575 37099 12416 37163
rect 12480 37099 12498 37163
rect 12562 37099 12580 37163
rect 12644 37099 12662 37163
rect 12726 37099 12744 37163
rect 12808 37099 12826 37163
rect 12890 37099 12908 37163
rect 12972 37099 12990 37163
rect 13054 37099 13072 37163
rect 13136 37099 13154 37163
rect 13218 37099 13236 37163
rect 13300 37099 13318 37163
rect 13382 37099 13400 37163
rect 13464 37099 13482 37163
rect 13546 37099 13564 37163
rect 13628 37099 13646 37163
rect 13710 37099 13728 37163
rect 13792 37099 13810 37163
rect 13874 37099 13892 37163
rect 13956 37099 13974 37163
rect 14038 37099 14056 37163
rect 14120 37099 14138 37163
rect 14202 37099 14220 37163
rect 14284 37099 14302 37163
rect 14366 37099 14384 37163
rect 14448 37099 14466 37163
rect 14530 37099 14548 37163
rect 14612 37099 14630 37163
rect 14694 37099 14712 37163
rect 14776 37099 14794 37163
rect 14858 37099 14876 37163
rect 14940 37099 15000 37163
rect 0 37082 15000 37099
rect 0 37018 111 37082
rect 175 37018 191 37082
rect 255 37018 271 37082
rect 335 37018 351 37082
rect 415 37018 431 37082
rect 495 37018 511 37082
rect 575 37018 591 37082
rect 655 37018 671 37082
rect 735 37018 751 37082
rect 815 37018 831 37082
rect 895 37018 911 37082
rect 975 37018 991 37082
rect 1055 37018 1071 37082
rect 1135 37018 1151 37082
rect 1215 37018 1231 37082
rect 1295 37018 1311 37082
rect 1375 37018 1391 37082
rect 1455 37018 1471 37082
rect 1535 37018 1551 37082
rect 1615 37018 1631 37082
rect 1695 37018 1711 37082
rect 1775 37018 1791 37082
rect 1855 37018 1871 37082
rect 1935 37018 1951 37082
rect 2015 37018 2031 37082
rect 2095 37018 2111 37082
rect 2175 37018 2191 37082
rect 2255 37018 2271 37082
rect 2335 37018 2351 37082
rect 2415 37018 2431 37082
rect 2495 37018 2511 37082
rect 2575 37018 12416 37082
rect 12480 37018 12498 37082
rect 12562 37018 12580 37082
rect 12644 37018 12662 37082
rect 12726 37018 12744 37082
rect 12808 37018 12826 37082
rect 12890 37018 12908 37082
rect 12972 37018 12990 37082
rect 13054 37018 13072 37082
rect 13136 37018 13154 37082
rect 13218 37018 13236 37082
rect 13300 37018 13318 37082
rect 13382 37018 13400 37082
rect 13464 37018 13482 37082
rect 13546 37018 13564 37082
rect 13628 37018 13646 37082
rect 13710 37018 13728 37082
rect 13792 37018 13810 37082
rect 13874 37018 13892 37082
rect 13956 37018 13974 37082
rect 14038 37018 14056 37082
rect 14120 37018 14138 37082
rect 14202 37018 14220 37082
rect 14284 37018 14302 37082
rect 14366 37018 14384 37082
rect 14448 37018 14466 37082
rect 14530 37018 14548 37082
rect 14612 37018 14630 37082
rect 14694 37018 14712 37082
rect 14776 37018 14794 37082
rect 14858 37018 14876 37082
rect 14940 37018 15000 37082
rect 0 37001 15000 37018
rect 0 36937 111 37001
rect 175 36937 191 37001
rect 255 36937 271 37001
rect 335 36937 351 37001
rect 415 36937 431 37001
rect 495 36937 511 37001
rect 575 36937 591 37001
rect 655 36937 671 37001
rect 735 36937 751 37001
rect 815 36937 831 37001
rect 895 36937 911 37001
rect 975 36937 991 37001
rect 1055 36937 1071 37001
rect 1135 36937 1151 37001
rect 1215 36937 1231 37001
rect 1295 36937 1311 37001
rect 1375 36937 1391 37001
rect 1455 36937 1471 37001
rect 1535 36937 1551 37001
rect 1615 36937 1631 37001
rect 1695 36937 1711 37001
rect 1775 36937 1791 37001
rect 1855 36937 1871 37001
rect 1935 36937 1951 37001
rect 2015 36937 2031 37001
rect 2095 36937 2111 37001
rect 2175 36937 2191 37001
rect 2255 36937 2271 37001
rect 2335 36937 2351 37001
rect 2415 36937 2431 37001
rect 2495 36937 2511 37001
rect 2575 36937 12416 37001
rect 12480 36937 12498 37001
rect 12562 36937 12580 37001
rect 12644 36937 12662 37001
rect 12726 36937 12744 37001
rect 12808 36937 12826 37001
rect 12890 36937 12908 37001
rect 12972 36937 12990 37001
rect 13054 36937 13072 37001
rect 13136 36937 13154 37001
rect 13218 36937 13236 37001
rect 13300 36937 13318 37001
rect 13382 36937 13400 37001
rect 13464 36937 13482 37001
rect 13546 36937 13564 37001
rect 13628 36937 13646 37001
rect 13710 36937 13728 37001
rect 13792 36937 13810 37001
rect 13874 36937 13892 37001
rect 13956 36937 13974 37001
rect 14038 36937 14056 37001
rect 14120 36937 14138 37001
rect 14202 36937 14220 37001
rect 14284 36937 14302 37001
rect 14366 36937 14384 37001
rect 14448 36937 14466 37001
rect 14530 36937 14548 37001
rect 14612 36937 14630 37001
rect 14694 36937 14712 37001
rect 14776 36937 14794 37001
rect 14858 36937 14876 37001
rect 14940 36937 15000 37001
rect 0 36920 15000 36937
rect 0 36856 111 36920
rect 175 36856 191 36920
rect 255 36856 271 36920
rect 335 36856 351 36920
rect 415 36856 431 36920
rect 495 36856 511 36920
rect 575 36856 591 36920
rect 655 36856 671 36920
rect 735 36856 751 36920
rect 815 36856 831 36920
rect 895 36856 911 36920
rect 975 36856 991 36920
rect 1055 36856 1071 36920
rect 1135 36856 1151 36920
rect 1215 36856 1231 36920
rect 1295 36856 1311 36920
rect 1375 36856 1391 36920
rect 1455 36856 1471 36920
rect 1535 36856 1551 36920
rect 1615 36856 1631 36920
rect 1695 36856 1711 36920
rect 1775 36856 1791 36920
rect 1855 36856 1871 36920
rect 1935 36856 1951 36920
rect 2015 36856 2031 36920
rect 2095 36856 2111 36920
rect 2175 36856 2191 36920
rect 2255 36856 2271 36920
rect 2335 36856 2351 36920
rect 2415 36856 2431 36920
rect 2495 36856 2511 36920
rect 2575 36856 12416 36920
rect 12480 36856 12498 36920
rect 12562 36856 12580 36920
rect 12644 36856 12662 36920
rect 12726 36856 12744 36920
rect 12808 36856 12826 36920
rect 12890 36856 12908 36920
rect 12972 36856 12990 36920
rect 13054 36856 13072 36920
rect 13136 36856 13154 36920
rect 13218 36856 13236 36920
rect 13300 36856 13318 36920
rect 13382 36856 13400 36920
rect 13464 36856 13482 36920
rect 13546 36856 13564 36920
rect 13628 36856 13646 36920
rect 13710 36856 13728 36920
rect 13792 36856 13810 36920
rect 13874 36856 13892 36920
rect 13956 36856 13974 36920
rect 14038 36856 14056 36920
rect 14120 36856 14138 36920
rect 14202 36856 14220 36920
rect 14284 36856 14302 36920
rect 14366 36856 14384 36920
rect 14448 36856 14466 36920
rect 14530 36856 14548 36920
rect 14612 36856 14630 36920
rect 14694 36856 14712 36920
rect 14776 36856 14794 36920
rect 14858 36856 14876 36920
rect 14940 36856 15000 36920
rect 0 36839 15000 36856
rect 0 36775 111 36839
rect 175 36775 191 36839
rect 255 36775 271 36839
rect 335 36775 351 36839
rect 415 36775 431 36839
rect 495 36775 511 36839
rect 575 36775 591 36839
rect 655 36775 671 36839
rect 735 36775 751 36839
rect 815 36775 831 36839
rect 895 36775 911 36839
rect 975 36775 991 36839
rect 1055 36775 1071 36839
rect 1135 36775 1151 36839
rect 1215 36775 1231 36839
rect 1295 36775 1311 36839
rect 1375 36775 1391 36839
rect 1455 36775 1471 36839
rect 1535 36775 1551 36839
rect 1615 36775 1631 36839
rect 1695 36775 1711 36839
rect 1775 36775 1791 36839
rect 1855 36775 1871 36839
rect 1935 36775 1951 36839
rect 2015 36775 2031 36839
rect 2095 36775 2111 36839
rect 2175 36775 2191 36839
rect 2255 36775 2271 36839
rect 2335 36775 2351 36839
rect 2415 36775 2431 36839
rect 2495 36775 2511 36839
rect 2575 36775 12416 36839
rect 12480 36775 12498 36839
rect 12562 36775 12580 36839
rect 12644 36775 12662 36839
rect 12726 36775 12744 36839
rect 12808 36775 12826 36839
rect 12890 36775 12908 36839
rect 12972 36775 12990 36839
rect 13054 36775 13072 36839
rect 13136 36775 13154 36839
rect 13218 36775 13236 36839
rect 13300 36775 13318 36839
rect 13382 36775 13400 36839
rect 13464 36775 13482 36839
rect 13546 36775 13564 36839
rect 13628 36775 13646 36839
rect 13710 36775 13728 36839
rect 13792 36775 13810 36839
rect 13874 36775 13892 36839
rect 13956 36775 13974 36839
rect 14038 36775 14056 36839
rect 14120 36775 14138 36839
rect 14202 36775 14220 36839
rect 14284 36775 14302 36839
rect 14366 36775 14384 36839
rect 14448 36775 14466 36839
rect 14530 36775 14548 36839
rect 14612 36775 14630 36839
rect 14694 36775 14712 36839
rect 14776 36775 14794 36839
rect 14858 36775 14876 36839
rect 14940 36775 15000 36839
rect 0 36758 15000 36775
rect 0 36694 111 36758
rect 175 36694 191 36758
rect 255 36694 271 36758
rect 335 36694 351 36758
rect 415 36694 431 36758
rect 495 36694 511 36758
rect 575 36694 591 36758
rect 655 36694 671 36758
rect 735 36694 751 36758
rect 815 36694 831 36758
rect 895 36694 911 36758
rect 975 36694 991 36758
rect 1055 36694 1071 36758
rect 1135 36694 1151 36758
rect 1215 36694 1231 36758
rect 1295 36694 1311 36758
rect 1375 36694 1391 36758
rect 1455 36694 1471 36758
rect 1535 36694 1551 36758
rect 1615 36694 1631 36758
rect 1695 36694 1711 36758
rect 1775 36694 1791 36758
rect 1855 36694 1871 36758
rect 1935 36694 1951 36758
rect 2015 36694 2031 36758
rect 2095 36694 2111 36758
rect 2175 36694 2191 36758
rect 2255 36694 2271 36758
rect 2335 36694 2351 36758
rect 2415 36694 2431 36758
rect 2495 36694 2511 36758
rect 2575 36694 12416 36758
rect 12480 36694 12498 36758
rect 12562 36694 12580 36758
rect 12644 36694 12662 36758
rect 12726 36694 12744 36758
rect 12808 36694 12826 36758
rect 12890 36694 12908 36758
rect 12972 36694 12990 36758
rect 13054 36694 13072 36758
rect 13136 36694 13154 36758
rect 13218 36694 13236 36758
rect 13300 36694 13318 36758
rect 13382 36694 13400 36758
rect 13464 36694 13482 36758
rect 13546 36694 13564 36758
rect 13628 36694 13646 36758
rect 13710 36694 13728 36758
rect 13792 36694 13810 36758
rect 13874 36694 13892 36758
rect 13956 36694 13974 36758
rect 14038 36694 14056 36758
rect 14120 36694 14138 36758
rect 14202 36694 14220 36758
rect 14284 36694 14302 36758
rect 14366 36694 14384 36758
rect 14448 36694 14466 36758
rect 14530 36694 14548 36758
rect 14612 36694 14630 36758
rect 14694 36694 14712 36758
rect 14776 36694 14794 36758
rect 14858 36694 14876 36758
rect 14940 36694 15000 36758
rect 0 36677 15000 36694
rect 0 36613 111 36677
rect 175 36613 191 36677
rect 255 36613 271 36677
rect 335 36613 351 36677
rect 415 36613 431 36677
rect 495 36613 511 36677
rect 575 36613 591 36677
rect 655 36613 671 36677
rect 735 36613 751 36677
rect 815 36613 831 36677
rect 895 36613 911 36677
rect 975 36613 991 36677
rect 1055 36613 1071 36677
rect 1135 36613 1151 36677
rect 1215 36613 1231 36677
rect 1295 36613 1311 36677
rect 1375 36613 1391 36677
rect 1455 36613 1471 36677
rect 1535 36613 1551 36677
rect 1615 36613 1631 36677
rect 1695 36613 1711 36677
rect 1775 36613 1791 36677
rect 1855 36613 1871 36677
rect 1935 36613 1951 36677
rect 2015 36613 2031 36677
rect 2095 36613 2111 36677
rect 2175 36613 2191 36677
rect 2255 36613 2271 36677
rect 2335 36613 2351 36677
rect 2415 36613 2431 36677
rect 2495 36613 2511 36677
rect 2575 36613 12416 36677
rect 12480 36613 12498 36677
rect 12562 36613 12580 36677
rect 12644 36613 12662 36677
rect 12726 36613 12744 36677
rect 12808 36613 12826 36677
rect 12890 36613 12908 36677
rect 12972 36613 12990 36677
rect 13054 36613 13072 36677
rect 13136 36613 13154 36677
rect 13218 36613 13236 36677
rect 13300 36613 13318 36677
rect 13382 36613 13400 36677
rect 13464 36613 13482 36677
rect 13546 36613 13564 36677
rect 13628 36613 13646 36677
rect 13710 36613 13728 36677
rect 13792 36613 13810 36677
rect 13874 36613 13892 36677
rect 13956 36613 13974 36677
rect 14038 36613 14056 36677
rect 14120 36613 14138 36677
rect 14202 36613 14220 36677
rect 14284 36613 14302 36677
rect 14366 36613 14384 36677
rect 14448 36613 14466 36677
rect 14530 36613 14548 36677
rect 14612 36613 14630 36677
rect 14694 36613 14712 36677
rect 14776 36613 14794 36677
rect 14858 36613 14876 36677
rect 14940 36613 15000 36677
rect 0 36596 15000 36613
rect 0 36532 111 36596
rect 175 36532 191 36596
rect 255 36532 271 36596
rect 335 36532 351 36596
rect 415 36532 431 36596
rect 495 36532 511 36596
rect 575 36532 591 36596
rect 655 36532 671 36596
rect 735 36532 751 36596
rect 815 36532 831 36596
rect 895 36532 911 36596
rect 975 36532 991 36596
rect 1055 36532 1071 36596
rect 1135 36532 1151 36596
rect 1215 36532 1231 36596
rect 1295 36532 1311 36596
rect 1375 36532 1391 36596
rect 1455 36532 1471 36596
rect 1535 36532 1551 36596
rect 1615 36532 1631 36596
rect 1695 36532 1711 36596
rect 1775 36532 1791 36596
rect 1855 36532 1871 36596
rect 1935 36532 1951 36596
rect 2015 36532 2031 36596
rect 2095 36532 2111 36596
rect 2175 36532 2191 36596
rect 2255 36532 2271 36596
rect 2335 36532 2351 36596
rect 2415 36532 2431 36596
rect 2495 36532 2511 36596
rect 2575 36532 12416 36596
rect 12480 36532 12498 36596
rect 12562 36532 12580 36596
rect 12644 36532 12662 36596
rect 12726 36532 12744 36596
rect 12808 36532 12826 36596
rect 12890 36532 12908 36596
rect 12972 36532 12990 36596
rect 13054 36532 13072 36596
rect 13136 36532 13154 36596
rect 13218 36532 13236 36596
rect 13300 36532 13318 36596
rect 13382 36532 13400 36596
rect 13464 36532 13482 36596
rect 13546 36532 13564 36596
rect 13628 36532 13646 36596
rect 13710 36532 13728 36596
rect 13792 36532 13810 36596
rect 13874 36532 13892 36596
rect 13956 36532 13974 36596
rect 14038 36532 14056 36596
rect 14120 36532 14138 36596
rect 14202 36532 14220 36596
rect 14284 36532 14302 36596
rect 14366 36532 14384 36596
rect 14448 36532 14466 36596
rect 14530 36532 14548 36596
rect 14612 36532 14630 36596
rect 14694 36532 14712 36596
rect 14776 36532 14794 36596
rect 14858 36532 14876 36596
rect 14940 36532 15000 36596
rect 0 36515 15000 36532
rect 0 36451 111 36515
rect 175 36451 191 36515
rect 255 36451 271 36515
rect 335 36451 351 36515
rect 415 36451 431 36515
rect 495 36451 511 36515
rect 575 36451 591 36515
rect 655 36451 671 36515
rect 735 36451 751 36515
rect 815 36451 831 36515
rect 895 36451 911 36515
rect 975 36451 991 36515
rect 1055 36451 1071 36515
rect 1135 36451 1151 36515
rect 1215 36451 1231 36515
rect 1295 36451 1311 36515
rect 1375 36451 1391 36515
rect 1455 36451 1471 36515
rect 1535 36451 1551 36515
rect 1615 36451 1631 36515
rect 1695 36451 1711 36515
rect 1775 36451 1791 36515
rect 1855 36451 1871 36515
rect 1935 36451 1951 36515
rect 2015 36451 2031 36515
rect 2095 36451 2111 36515
rect 2175 36451 2191 36515
rect 2255 36451 2271 36515
rect 2335 36451 2351 36515
rect 2415 36451 2431 36515
rect 2495 36451 2511 36515
rect 2575 36451 12416 36515
rect 12480 36451 12498 36515
rect 12562 36451 12580 36515
rect 12644 36451 12662 36515
rect 12726 36451 12744 36515
rect 12808 36451 12826 36515
rect 12890 36451 12908 36515
rect 12972 36451 12990 36515
rect 13054 36451 13072 36515
rect 13136 36451 13154 36515
rect 13218 36451 13236 36515
rect 13300 36451 13318 36515
rect 13382 36451 13400 36515
rect 13464 36451 13482 36515
rect 13546 36451 13564 36515
rect 13628 36451 13646 36515
rect 13710 36451 13728 36515
rect 13792 36451 13810 36515
rect 13874 36451 13892 36515
rect 13956 36451 13974 36515
rect 14038 36451 14056 36515
rect 14120 36451 14138 36515
rect 14202 36451 14220 36515
rect 14284 36451 14302 36515
rect 14366 36451 14384 36515
rect 14448 36451 14466 36515
rect 14530 36451 14548 36515
rect 14612 36451 14630 36515
rect 14694 36451 14712 36515
rect 14776 36451 14794 36515
rect 14858 36451 14876 36515
rect 14940 36451 15000 36515
rect 0 36434 15000 36451
rect 0 36370 111 36434
rect 175 36370 191 36434
rect 255 36370 271 36434
rect 335 36370 351 36434
rect 415 36370 431 36434
rect 495 36370 511 36434
rect 575 36370 591 36434
rect 655 36370 671 36434
rect 735 36370 751 36434
rect 815 36370 831 36434
rect 895 36370 911 36434
rect 975 36370 991 36434
rect 1055 36370 1071 36434
rect 1135 36370 1151 36434
rect 1215 36370 1231 36434
rect 1295 36370 1311 36434
rect 1375 36370 1391 36434
rect 1455 36370 1471 36434
rect 1535 36370 1551 36434
rect 1615 36370 1631 36434
rect 1695 36370 1711 36434
rect 1775 36370 1791 36434
rect 1855 36370 1871 36434
rect 1935 36370 1951 36434
rect 2015 36370 2031 36434
rect 2095 36370 2111 36434
rect 2175 36370 2191 36434
rect 2255 36370 2271 36434
rect 2335 36370 2351 36434
rect 2415 36370 2431 36434
rect 2495 36370 2511 36434
rect 2575 36370 12416 36434
rect 12480 36370 12498 36434
rect 12562 36370 12580 36434
rect 12644 36370 12662 36434
rect 12726 36370 12744 36434
rect 12808 36370 12826 36434
rect 12890 36370 12908 36434
rect 12972 36370 12990 36434
rect 13054 36370 13072 36434
rect 13136 36370 13154 36434
rect 13218 36370 13236 36434
rect 13300 36370 13318 36434
rect 13382 36370 13400 36434
rect 13464 36370 13482 36434
rect 13546 36370 13564 36434
rect 13628 36370 13646 36434
rect 13710 36370 13728 36434
rect 13792 36370 13810 36434
rect 13874 36370 13892 36434
rect 13956 36370 13974 36434
rect 14038 36370 14056 36434
rect 14120 36370 14138 36434
rect 14202 36370 14220 36434
rect 14284 36370 14302 36434
rect 14366 36370 14384 36434
rect 14448 36370 14466 36434
rect 14530 36370 14548 36434
rect 14612 36370 14630 36434
rect 14694 36370 14712 36434
rect 14776 36370 14794 36434
rect 14858 36370 14876 36434
rect 14940 36370 15000 36434
rect 0 36353 15000 36370
rect 0 36289 111 36353
rect 175 36289 191 36353
rect 255 36289 271 36353
rect 335 36289 351 36353
rect 415 36289 431 36353
rect 495 36289 511 36353
rect 575 36289 591 36353
rect 655 36289 671 36353
rect 735 36289 751 36353
rect 815 36289 831 36353
rect 895 36289 911 36353
rect 975 36289 991 36353
rect 1055 36289 1071 36353
rect 1135 36289 1151 36353
rect 1215 36289 1231 36353
rect 1295 36289 1311 36353
rect 1375 36289 1391 36353
rect 1455 36289 1471 36353
rect 1535 36289 1551 36353
rect 1615 36289 1631 36353
rect 1695 36289 1711 36353
rect 1775 36289 1791 36353
rect 1855 36289 1871 36353
rect 1935 36289 1951 36353
rect 2015 36289 2031 36353
rect 2095 36289 2111 36353
rect 2175 36289 2191 36353
rect 2255 36289 2271 36353
rect 2335 36289 2351 36353
rect 2415 36289 2431 36353
rect 2495 36289 2511 36353
rect 2575 36289 12416 36353
rect 12480 36289 12498 36353
rect 12562 36289 12580 36353
rect 12644 36289 12662 36353
rect 12726 36289 12744 36353
rect 12808 36289 12826 36353
rect 12890 36289 12908 36353
rect 12972 36289 12990 36353
rect 13054 36289 13072 36353
rect 13136 36289 13154 36353
rect 13218 36289 13236 36353
rect 13300 36289 13318 36353
rect 13382 36289 13400 36353
rect 13464 36289 13482 36353
rect 13546 36289 13564 36353
rect 13628 36289 13646 36353
rect 13710 36289 13728 36353
rect 13792 36289 13810 36353
rect 13874 36289 13892 36353
rect 13956 36289 13974 36353
rect 14038 36289 14056 36353
rect 14120 36289 14138 36353
rect 14202 36289 14220 36353
rect 14284 36289 14302 36353
rect 14366 36289 14384 36353
rect 14448 36289 14466 36353
rect 14530 36289 14548 36353
rect 14612 36289 14630 36353
rect 14694 36289 14712 36353
rect 14776 36289 14794 36353
rect 14858 36289 14876 36353
rect 14940 36289 15000 36353
rect 0 36272 15000 36289
rect 0 34768 111 36272
rect 2575 36208 12416 36272
rect 12480 36208 12498 36272
rect 12562 36208 12580 36272
rect 12644 36208 12662 36272
rect 12726 36208 12744 36272
rect 12808 36208 12826 36272
rect 12890 36208 12908 36272
rect 12972 36208 12990 36272
rect 13054 36208 13072 36272
rect 13136 36208 13154 36272
rect 13218 36208 13236 36272
rect 13300 36208 13318 36272
rect 13382 36208 13400 36272
rect 13464 36208 13482 36272
rect 13546 36208 13564 36272
rect 13628 36208 13646 36272
rect 13710 36208 13728 36272
rect 13792 36208 13810 36272
rect 13874 36208 13892 36272
rect 13956 36208 13974 36272
rect 14038 36208 14056 36272
rect 14120 36208 14138 36272
rect 14202 36208 14220 36272
rect 14284 36208 14302 36272
rect 14366 36208 14384 36272
rect 14448 36208 14466 36272
rect 14530 36208 14548 36272
rect 14612 36208 14630 36272
rect 14694 36208 14712 36272
rect 14776 36208 14794 36272
rect 14858 36208 14876 36272
rect 14940 36208 15000 36272
rect 2575 36192 15000 36208
rect 2575 36128 12416 36192
rect 12480 36128 12498 36192
rect 12562 36128 12580 36192
rect 12644 36128 12662 36192
rect 12726 36128 12744 36192
rect 12808 36128 12826 36192
rect 12890 36128 12908 36192
rect 12972 36128 12990 36192
rect 13054 36128 13072 36192
rect 13136 36128 13154 36192
rect 13218 36128 13236 36192
rect 13300 36128 13318 36192
rect 13382 36128 13400 36192
rect 13464 36128 13482 36192
rect 13546 36128 13564 36192
rect 13628 36128 13646 36192
rect 13710 36128 13728 36192
rect 13792 36128 13810 36192
rect 13874 36128 13892 36192
rect 13956 36128 13974 36192
rect 14038 36128 14056 36192
rect 14120 36128 14138 36192
rect 14202 36128 14220 36192
rect 14284 36128 14302 36192
rect 14366 36128 14384 36192
rect 14448 36128 14466 36192
rect 14530 36128 14548 36192
rect 14612 36128 14630 36192
rect 14694 36128 14712 36192
rect 14776 36128 14794 36192
rect 14858 36128 14876 36192
rect 14940 36128 15000 36192
rect 2575 36112 15000 36128
rect 2575 36048 12416 36112
rect 12480 36048 12498 36112
rect 12562 36048 12580 36112
rect 12644 36048 12662 36112
rect 12726 36048 12744 36112
rect 12808 36048 12826 36112
rect 12890 36048 12908 36112
rect 12972 36048 12990 36112
rect 13054 36048 13072 36112
rect 13136 36048 13154 36112
rect 13218 36048 13236 36112
rect 13300 36048 13318 36112
rect 13382 36048 13400 36112
rect 13464 36048 13482 36112
rect 13546 36048 13564 36112
rect 13628 36048 13646 36112
rect 13710 36048 13728 36112
rect 13792 36048 13810 36112
rect 13874 36048 13892 36112
rect 13956 36048 13974 36112
rect 14038 36048 14056 36112
rect 14120 36048 14138 36112
rect 14202 36048 14220 36112
rect 14284 36048 14302 36112
rect 14366 36048 14384 36112
rect 14448 36048 14466 36112
rect 14530 36048 14548 36112
rect 14612 36048 14630 36112
rect 14694 36048 14712 36112
rect 14776 36048 14794 36112
rect 14858 36048 14876 36112
rect 14940 36048 15000 36112
rect 2575 36032 15000 36048
rect 2575 35968 12416 36032
rect 12480 35968 12498 36032
rect 12562 35968 12580 36032
rect 12644 35968 12662 36032
rect 12726 35968 12744 36032
rect 12808 35968 12826 36032
rect 12890 35968 12908 36032
rect 12972 35968 12990 36032
rect 13054 35968 13072 36032
rect 13136 35968 13154 36032
rect 13218 35968 13236 36032
rect 13300 35968 13318 36032
rect 13382 35968 13400 36032
rect 13464 35968 13482 36032
rect 13546 35968 13564 36032
rect 13628 35968 13646 36032
rect 13710 35968 13728 36032
rect 13792 35968 13810 36032
rect 13874 35968 13892 36032
rect 13956 35968 13974 36032
rect 14038 35968 14056 36032
rect 14120 35968 14138 36032
rect 14202 35968 14220 36032
rect 14284 35968 14302 36032
rect 14366 35968 14384 36032
rect 14448 35968 14466 36032
rect 14530 35968 14548 36032
rect 14612 35968 14630 36032
rect 14694 35968 14712 36032
rect 14776 35968 14794 36032
rect 14858 35968 14876 36032
rect 14940 35968 15000 36032
rect 2575 35952 15000 35968
rect 2575 35888 12416 35952
rect 12480 35888 12498 35952
rect 12562 35888 12580 35952
rect 12644 35888 12662 35952
rect 12726 35888 12744 35952
rect 12808 35888 12826 35952
rect 12890 35888 12908 35952
rect 12972 35888 12990 35952
rect 13054 35888 13072 35952
rect 13136 35888 13154 35952
rect 13218 35888 13236 35952
rect 13300 35888 13318 35952
rect 13382 35888 13400 35952
rect 13464 35888 13482 35952
rect 13546 35888 13564 35952
rect 13628 35888 13646 35952
rect 13710 35888 13728 35952
rect 13792 35888 13810 35952
rect 13874 35888 13892 35952
rect 13956 35888 13974 35952
rect 14038 35888 14056 35952
rect 14120 35888 14138 35952
rect 14202 35888 14220 35952
rect 14284 35888 14302 35952
rect 14366 35888 14384 35952
rect 14448 35888 14466 35952
rect 14530 35888 14548 35952
rect 14612 35888 14630 35952
rect 14694 35888 14712 35952
rect 14776 35888 14794 35952
rect 14858 35888 14876 35952
rect 14940 35888 15000 35952
rect 2575 35872 15000 35888
rect 2575 35808 12416 35872
rect 12480 35808 12498 35872
rect 12562 35808 12580 35872
rect 12644 35808 12662 35872
rect 12726 35808 12744 35872
rect 12808 35808 12826 35872
rect 12890 35808 12908 35872
rect 12972 35808 12990 35872
rect 13054 35808 13072 35872
rect 13136 35808 13154 35872
rect 13218 35808 13236 35872
rect 13300 35808 13318 35872
rect 13382 35808 13400 35872
rect 13464 35808 13482 35872
rect 13546 35808 13564 35872
rect 13628 35808 13646 35872
rect 13710 35808 13728 35872
rect 13792 35808 13810 35872
rect 13874 35808 13892 35872
rect 13956 35808 13974 35872
rect 14038 35808 14056 35872
rect 14120 35808 14138 35872
rect 14202 35808 14220 35872
rect 14284 35808 14302 35872
rect 14366 35808 14384 35872
rect 14448 35808 14466 35872
rect 14530 35808 14548 35872
rect 14612 35808 14630 35872
rect 14694 35808 14712 35872
rect 14776 35808 14794 35872
rect 14858 35808 14876 35872
rect 14940 35808 15000 35872
rect 2575 35792 15000 35808
rect 2575 35728 12416 35792
rect 12480 35728 12498 35792
rect 12562 35728 12580 35792
rect 12644 35728 12662 35792
rect 12726 35728 12744 35792
rect 12808 35728 12826 35792
rect 12890 35728 12908 35792
rect 12972 35728 12990 35792
rect 13054 35728 13072 35792
rect 13136 35728 13154 35792
rect 13218 35728 13236 35792
rect 13300 35728 13318 35792
rect 13382 35728 13400 35792
rect 13464 35728 13482 35792
rect 13546 35728 13564 35792
rect 13628 35728 13646 35792
rect 13710 35728 13728 35792
rect 13792 35728 13810 35792
rect 13874 35728 13892 35792
rect 13956 35728 13974 35792
rect 14038 35728 14056 35792
rect 14120 35728 14138 35792
rect 14202 35728 14220 35792
rect 14284 35728 14302 35792
rect 14366 35728 14384 35792
rect 14448 35728 14466 35792
rect 14530 35728 14548 35792
rect 14612 35728 14630 35792
rect 14694 35728 14712 35792
rect 14776 35728 14794 35792
rect 14858 35728 14876 35792
rect 14940 35728 15000 35792
rect 2575 35712 15000 35728
rect 2575 35648 12416 35712
rect 12480 35648 12498 35712
rect 12562 35648 12580 35712
rect 12644 35648 12662 35712
rect 12726 35648 12744 35712
rect 12808 35648 12826 35712
rect 12890 35648 12908 35712
rect 12972 35648 12990 35712
rect 13054 35648 13072 35712
rect 13136 35648 13154 35712
rect 13218 35648 13236 35712
rect 13300 35648 13318 35712
rect 13382 35648 13400 35712
rect 13464 35648 13482 35712
rect 13546 35648 13564 35712
rect 13628 35648 13646 35712
rect 13710 35648 13728 35712
rect 13792 35648 13810 35712
rect 13874 35648 13892 35712
rect 13956 35648 13974 35712
rect 14038 35648 14056 35712
rect 14120 35648 14138 35712
rect 14202 35648 14220 35712
rect 14284 35648 14302 35712
rect 14366 35648 14384 35712
rect 14448 35648 14466 35712
rect 14530 35648 14548 35712
rect 14612 35648 14630 35712
rect 14694 35648 14712 35712
rect 14776 35648 14794 35712
rect 14858 35648 14876 35712
rect 14940 35648 15000 35712
rect 2575 35632 15000 35648
rect 2575 35568 12416 35632
rect 12480 35568 12498 35632
rect 12562 35568 12580 35632
rect 12644 35568 12662 35632
rect 12726 35568 12744 35632
rect 12808 35568 12826 35632
rect 12890 35568 12908 35632
rect 12972 35568 12990 35632
rect 13054 35568 13072 35632
rect 13136 35568 13154 35632
rect 13218 35568 13236 35632
rect 13300 35568 13318 35632
rect 13382 35568 13400 35632
rect 13464 35568 13482 35632
rect 13546 35568 13564 35632
rect 13628 35568 13646 35632
rect 13710 35568 13728 35632
rect 13792 35568 13810 35632
rect 13874 35568 13892 35632
rect 13956 35568 13974 35632
rect 14038 35568 14056 35632
rect 14120 35568 14138 35632
rect 14202 35568 14220 35632
rect 14284 35568 14302 35632
rect 14366 35568 14384 35632
rect 14448 35568 14466 35632
rect 14530 35568 14548 35632
rect 14612 35568 14630 35632
rect 14694 35568 14712 35632
rect 14776 35568 14794 35632
rect 14858 35568 14876 35632
rect 14940 35568 15000 35632
rect 2575 35552 15000 35568
rect 2575 35488 12416 35552
rect 12480 35488 12498 35552
rect 12562 35488 12580 35552
rect 12644 35488 12662 35552
rect 12726 35488 12744 35552
rect 12808 35488 12826 35552
rect 12890 35488 12908 35552
rect 12972 35488 12990 35552
rect 13054 35488 13072 35552
rect 13136 35488 13154 35552
rect 13218 35488 13236 35552
rect 13300 35488 13318 35552
rect 13382 35488 13400 35552
rect 13464 35488 13482 35552
rect 13546 35488 13564 35552
rect 13628 35488 13646 35552
rect 13710 35488 13728 35552
rect 13792 35488 13810 35552
rect 13874 35488 13892 35552
rect 13956 35488 13974 35552
rect 14038 35488 14056 35552
rect 14120 35488 14138 35552
rect 14202 35488 14220 35552
rect 14284 35488 14302 35552
rect 14366 35488 14384 35552
rect 14448 35488 14466 35552
rect 14530 35488 14548 35552
rect 14612 35488 14630 35552
rect 14694 35488 14712 35552
rect 14776 35488 14794 35552
rect 14858 35488 14876 35552
rect 14940 35488 15000 35552
rect 2575 35472 15000 35488
rect 2575 35408 12416 35472
rect 12480 35408 12498 35472
rect 12562 35408 12580 35472
rect 12644 35408 12662 35472
rect 12726 35408 12744 35472
rect 12808 35408 12826 35472
rect 12890 35408 12908 35472
rect 12972 35408 12990 35472
rect 13054 35408 13072 35472
rect 13136 35408 13154 35472
rect 13218 35408 13236 35472
rect 13300 35408 13318 35472
rect 13382 35408 13400 35472
rect 13464 35408 13482 35472
rect 13546 35408 13564 35472
rect 13628 35408 13646 35472
rect 13710 35408 13728 35472
rect 13792 35408 13810 35472
rect 13874 35408 13892 35472
rect 13956 35408 13974 35472
rect 14038 35408 14056 35472
rect 14120 35408 14138 35472
rect 14202 35408 14220 35472
rect 14284 35408 14302 35472
rect 14366 35408 14384 35472
rect 14448 35408 14466 35472
rect 14530 35408 14548 35472
rect 14612 35408 14630 35472
rect 14694 35408 14712 35472
rect 14776 35408 14794 35472
rect 14858 35408 14876 35472
rect 14940 35408 15000 35472
rect 2575 35392 15000 35408
rect 2575 35328 12416 35392
rect 12480 35328 12498 35392
rect 12562 35328 12580 35392
rect 12644 35328 12662 35392
rect 12726 35328 12744 35392
rect 12808 35328 12826 35392
rect 12890 35328 12908 35392
rect 12972 35328 12990 35392
rect 13054 35328 13072 35392
rect 13136 35328 13154 35392
rect 13218 35328 13236 35392
rect 13300 35328 13318 35392
rect 13382 35328 13400 35392
rect 13464 35328 13482 35392
rect 13546 35328 13564 35392
rect 13628 35328 13646 35392
rect 13710 35328 13728 35392
rect 13792 35328 13810 35392
rect 13874 35328 13892 35392
rect 13956 35328 13974 35392
rect 14038 35328 14056 35392
rect 14120 35328 14138 35392
rect 14202 35328 14220 35392
rect 14284 35328 14302 35392
rect 14366 35328 14384 35392
rect 14448 35328 14466 35392
rect 14530 35328 14548 35392
rect 14612 35328 14630 35392
rect 14694 35328 14712 35392
rect 14776 35328 14794 35392
rect 14858 35328 14876 35392
rect 14940 35328 15000 35392
rect 2575 35312 15000 35328
rect 2575 35248 12416 35312
rect 12480 35248 12498 35312
rect 12562 35248 12580 35312
rect 12644 35248 12662 35312
rect 12726 35248 12744 35312
rect 12808 35248 12826 35312
rect 12890 35248 12908 35312
rect 12972 35248 12990 35312
rect 13054 35248 13072 35312
rect 13136 35248 13154 35312
rect 13218 35248 13236 35312
rect 13300 35248 13318 35312
rect 13382 35248 13400 35312
rect 13464 35248 13482 35312
rect 13546 35248 13564 35312
rect 13628 35248 13646 35312
rect 13710 35248 13728 35312
rect 13792 35248 13810 35312
rect 13874 35248 13892 35312
rect 13956 35248 13974 35312
rect 14038 35248 14056 35312
rect 14120 35248 14138 35312
rect 14202 35248 14220 35312
rect 14284 35248 14302 35312
rect 14366 35248 14384 35312
rect 14448 35248 14466 35312
rect 14530 35248 14548 35312
rect 14612 35248 14630 35312
rect 14694 35248 14712 35312
rect 14776 35248 14794 35312
rect 14858 35248 14876 35312
rect 14940 35248 15000 35312
rect 2575 35232 15000 35248
rect 2575 35168 12416 35232
rect 12480 35168 12498 35232
rect 12562 35168 12580 35232
rect 12644 35168 12662 35232
rect 12726 35168 12744 35232
rect 12808 35168 12826 35232
rect 12890 35168 12908 35232
rect 12972 35168 12990 35232
rect 13054 35168 13072 35232
rect 13136 35168 13154 35232
rect 13218 35168 13236 35232
rect 13300 35168 13318 35232
rect 13382 35168 13400 35232
rect 13464 35168 13482 35232
rect 13546 35168 13564 35232
rect 13628 35168 13646 35232
rect 13710 35168 13728 35232
rect 13792 35168 13810 35232
rect 13874 35168 13892 35232
rect 13956 35168 13974 35232
rect 14038 35168 14056 35232
rect 14120 35168 14138 35232
rect 14202 35168 14220 35232
rect 14284 35168 14302 35232
rect 14366 35168 14384 35232
rect 14448 35168 14466 35232
rect 14530 35168 14548 35232
rect 14612 35168 14630 35232
rect 14694 35168 14712 35232
rect 14776 35168 14794 35232
rect 14858 35168 14876 35232
rect 14940 35168 15000 35232
rect 2575 35152 15000 35168
rect 2575 35088 12416 35152
rect 12480 35088 12498 35152
rect 12562 35088 12580 35152
rect 12644 35088 12662 35152
rect 12726 35088 12744 35152
rect 12808 35088 12826 35152
rect 12890 35088 12908 35152
rect 12972 35088 12990 35152
rect 13054 35088 13072 35152
rect 13136 35088 13154 35152
rect 13218 35088 13236 35152
rect 13300 35088 13318 35152
rect 13382 35088 13400 35152
rect 13464 35088 13482 35152
rect 13546 35088 13564 35152
rect 13628 35088 13646 35152
rect 13710 35088 13728 35152
rect 13792 35088 13810 35152
rect 13874 35088 13892 35152
rect 13956 35088 13974 35152
rect 14038 35088 14056 35152
rect 14120 35088 14138 35152
rect 14202 35088 14220 35152
rect 14284 35088 14302 35152
rect 14366 35088 14384 35152
rect 14448 35088 14466 35152
rect 14530 35088 14548 35152
rect 14612 35088 14630 35152
rect 14694 35088 14712 35152
rect 14776 35088 14794 35152
rect 14858 35088 14876 35152
rect 14940 35088 15000 35152
rect 2575 35072 15000 35088
rect 2575 35008 12416 35072
rect 12480 35008 12498 35072
rect 12562 35008 12580 35072
rect 12644 35008 12662 35072
rect 12726 35008 12744 35072
rect 12808 35008 12826 35072
rect 12890 35008 12908 35072
rect 12972 35008 12990 35072
rect 13054 35008 13072 35072
rect 13136 35008 13154 35072
rect 13218 35008 13236 35072
rect 13300 35008 13318 35072
rect 13382 35008 13400 35072
rect 13464 35008 13482 35072
rect 13546 35008 13564 35072
rect 13628 35008 13646 35072
rect 13710 35008 13728 35072
rect 13792 35008 13810 35072
rect 13874 35008 13892 35072
rect 13956 35008 13974 35072
rect 14038 35008 14056 35072
rect 14120 35008 14138 35072
rect 14202 35008 14220 35072
rect 14284 35008 14302 35072
rect 14366 35008 14384 35072
rect 14448 35008 14466 35072
rect 14530 35008 14548 35072
rect 14612 35008 14630 35072
rect 14694 35008 14712 35072
rect 14776 35008 14794 35072
rect 14858 35008 14876 35072
rect 14940 35008 15000 35072
rect 2575 34992 15000 35008
rect 2575 34928 12416 34992
rect 12480 34928 12498 34992
rect 12562 34928 12580 34992
rect 12644 34928 12662 34992
rect 12726 34928 12744 34992
rect 12808 34928 12826 34992
rect 12890 34928 12908 34992
rect 12972 34928 12990 34992
rect 13054 34928 13072 34992
rect 13136 34928 13154 34992
rect 13218 34928 13236 34992
rect 13300 34928 13318 34992
rect 13382 34928 13400 34992
rect 13464 34928 13482 34992
rect 13546 34928 13564 34992
rect 13628 34928 13646 34992
rect 13710 34928 13728 34992
rect 13792 34928 13810 34992
rect 13874 34928 13892 34992
rect 13956 34928 13974 34992
rect 14038 34928 14056 34992
rect 14120 34928 14138 34992
rect 14202 34928 14220 34992
rect 14284 34928 14302 34992
rect 14366 34928 14384 34992
rect 14448 34928 14466 34992
rect 14530 34928 14548 34992
rect 14612 34928 14630 34992
rect 14694 34928 14712 34992
rect 14776 34928 14794 34992
rect 14858 34928 14876 34992
rect 14940 34928 15000 34992
rect 2575 34912 15000 34928
rect 2575 34848 12416 34912
rect 12480 34848 12498 34912
rect 12562 34848 12580 34912
rect 12644 34848 12662 34912
rect 12726 34848 12744 34912
rect 12808 34848 12826 34912
rect 12890 34848 12908 34912
rect 12972 34848 12990 34912
rect 13054 34848 13072 34912
rect 13136 34848 13154 34912
rect 13218 34848 13236 34912
rect 13300 34848 13318 34912
rect 13382 34848 13400 34912
rect 13464 34848 13482 34912
rect 13546 34848 13564 34912
rect 13628 34848 13646 34912
rect 13710 34848 13728 34912
rect 13792 34848 13810 34912
rect 13874 34848 13892 34912
rect 13956 34848 13974 34912
rect 14038 34848 14056 34912
rect 14120 34848 14138 34912
rect 14202 34848 14220 34912
rect 14284 34848 14302 34912
rect 14366 34848 14384 34912
rect 14448 34848 14466 34912
rect 14530 34848 14548 34912
rect 14612 34848 14630 34912
rect 14694 34848 14712 34912
rect 14776 34848 14794 34912
rect 14858 34848 14876 34912
rect 14940 34848 15000 34912
rect 2575 34832 15000 34848
rect 2575 34768 12416 34832
rect 12480 34768 12498 34832
rect 12562 34768 12580 34832
rect 12644 34768 12662 34832
rect 12726 34768 12744 34832
rect 12808 34768 12826 34832
rect 12890 34768 12908 34832
rect 12972 34768 12990 34832
rect 13054 34768 13072 34832
rect 13136 34768 13154 34832
rect 13218 34768 13236 34832
rect 13300 34768 13318 34832
rect 13382 34768 13400 34832
rect 13464 34768 13482 34832
rect 13546 34768 13564 34832
rect 13628 34768 13646 34832
rect 13710 34768 13728 34832
rect 13792 34768 13810 34832
rect 13874 34768 13892 34832
rect 13956 34768 13974 34832
rect 14038 34768 14056 34832
rect 14120 34768 14138 34832
rect 14202 34768 14220 34832
rect 14284 34768 14302 34832
rect 14366 34768 14384 34832
rect 14448 34768 14466 34832
rect 14530 34768 14548 34832
rect 14612 34768 14630 34832
rect 14694 34768 14712 34832
rect 14776 34768 14794 34832
rect 14858 34768 14876 34832
rect 14940 34768 15000 34832
rect 0 12134 15000 34768
rect 0 12070 106 12134
rect 170 12070 188 12134
rect 252 12070 270 12134
rect 334 12070 352 12134
rect 416 12070 434 12134
rect 498 12070 516 12134
rect 580 12070 598 12134
rect 662 12070 679 12134
rect 743 12070 760 12134
rect 824 12070 841 12134
rect 905 12070 922 12134
rect 986 12070 1003 12134
rect 1067 12070 1084 12134
rect 1148 12070 1165 12134
rect 1229 12070 1246 12134
rect 1310 12070 1327 12134
rect 1391 12070 1408 12134
rect 1472 12070 1489 12134
rect 1553 12070 1570 12134
rect 1634 12070 1651 12134
rect 1715 12070 1732 12134
rect 1796 12070 1813 12134
rect 1877 12070 1894 12134
rect 1958 12070 1975 12134
rect 2039 12070 2056 12134
rect 2120 12070 2137 12134
rect 2201 12070 2218 12134
rect 2282 12070 2299 12134
rect 2363 12070 2380 12134
rect 2444 12070 2461 12134
rect 2525 12070 2542 12134
rect 2606 12070 2623 12134
rect 2687 12070 2704 12134
rect 2768 12070 2785 12134
rect 2849 12070 2866 12134
rect 2930 12070 2947 12134
rect 3011 12070 3028 12134
rect 3092 12070 3109 12134
rect 3173 12070 3190 12134
rect 3254 12070 3271 12134
rect 3335 12070 3352 12134
rect 3416 12070 3433 12134
rect 3497 12070 3514 12134
rect 3578 12070 3595 12134
rect 3659 12070 3676 12134
rect 3740 12070 3757 12134
rect 3821 12070 3838 12134
rect 3902 12070 3919 12134
rect 3983 12070 4000 12134
rect 4064 12070 4081 12134
rect 4145 12070 4162 12134
rect 4226 12070 4243 12134
rect 4307 12070 4324 12134
rect 4388 12070 4405 12134
rect 4469 12070 4486 12134
rect 4550 12070 4567 12134
rect 4631 12070 4648 12134
rect 4712 12070 4729 12134
rect 4793 12070 4810 12134
rect 4874 12070 10157 12134
rect 10221 12070 10239 12134
rect 10303 12070 10321 12134
rect 10385 12070 10403 12134
rect 10467 12070 10485 12134
rect 10549 12070 10567 12134
rect 10631 12070 10649 12134
rect 10713 12070 10731 12134
rect 10795 12070 10813 12134
rect 10877 12070 10895 12134
rect 10959 12070 10977 12134
rect 11041 12070 11059 12134
rect 11123 12070 11141 12134
rect 11205 12070 11223 12134
rect 11287 12070 11305 12134
rect 11369 12070 11386 12134
rect 11450 12070 11467 12134
rect 11531 12070 11548 12134
rect 11612 12070 11629 12134
rect 11693 12070 11710 12134
rect 11774 12070 11791 12134
rect 11855 12070 11872 12134
rect 11936 12070 11953 12134
rect 12017 12070 12034 12134
rect 12098 12070 12115 12134
rect 12179 12070 12196 12134
rect 12260 12070 12277 12134
rect 12341 12070 12358 12134
rect 12422 12070 12439 12134
rect 12503 12070 12520 12134
rect 12584 12070 12601 12134
rect 12665 12070 12682 12134
rect 12746 12070 12763 12134
rect 12827 12070 12844 12134
rect 12908 12070 12925 12134
rect 12989 12070 13006 12134
rect 13070 12070 13087 12134
rect 13151 12070 13168 12134
rect 13232 12070 13249 12134
rect 13313 12070 13330 12134
rect 13394 12070 13411 12134
rect 13475 12070 13492 12134
rect 13556 12070 13573 12134
rect 13637 12070 13654 12134
rect 13718 12070 13735 12134
rect 13799 12070 13816 12134
rect 13880 12070 13897 12134
rect 13961 12070 13978 12134
rect 14042 12070 14059 12134
rect 14123 12070 14140 12134
rect 14204 12070 14221 12134
rect 14285 12070 14302 12134
rect 14366 12070 14383 12134
rect 14447 12070 14464 12134
rect 14528 12070 14545 12134
rect 14609 12070 14626 12134
rect 14690 12070 14707 12134
rect 14771 12070 14788 12134
rect 14852 12070 15000 12134
rect 0 12052 15000 12070
rect 0 11988 106 12052
rect 170 11988 188 12052
rect 252 11988 270 12052
rect 334 11988 352 12052
rect 416 11988 434 12052
rect 498 11988 516 12052
rect 580 11988 598 12052
rect 662 11988 679 12052
rect 743 11988 760 12052
rect 824 11988 841 12052
rect 905 11988 922 12052
rect 986 11988 1003 12052
rect 1067 11988 1084 12052
rect 1148 11988 1165 12052
rect 1229 11988 1246 12052
rect 1310 11988 1327 12052
rect 1391 11988 1408 12052
rect 1472 11988 1489 12052
rect 1553 11988 1570 12052
rect 1634 11988 1651 12052
rect 1715 11988 1732 12052
rect 1796 11988 1813 12052
rect 1877 11988 1894 12052
rect 1958 11988 1975 12052
rect 2039 11988 2056 12052
rect 2120 11988 2137 12052
rect 2201 11988 2218 12052
rect 2282 11988 2299 12052
rect 2363 11988 2380 12052
rect 2444 11988 2461 12052
rect 2525 11988 2542 12052
rect 2606 11988 2623 12052
rect 2687 11988 2704 12052
rect 2768 11988 2785 12052
rect 2849 11988 2866 12052
rect 2930 11988 2947 12052
rect 3011 11988 3028 12052
rect 3092 11988 3109 12052
rect 3173 11988 3190 12052
rect 3254 11988 3271 12052
rect 3335 11988 3352 12052
rect 3416 11988 3433 12052
rect 3497 11988 3514 12052
rect 3578 11988 3595 12052
rect 3659 11988 3676 12052
rect 3740 11988 3757 12052
rect 3821 11988 3838 12052
rect 3902 11988 3919 12052
rect 3983 11988 4000 12052
rect 4064 11988 4081 12052
rect 4145 11988 4162 12052
rect 4226 11988 4243 12052
rect 4307 11988 4324 12052
rect 4388 11988 4405 12052
rect 4469 11988 4486 12052
rect 4550 11988 4567 12052
rect 4631 11988 4648 12052
rect 4712 11988 4729 12052
rect 4793 11988 4810 12052
rect 4874 11988 10157 12052
rect 10221 11988 10239 12052
rect 10303 11988 10321 12052
rect 10385 11988 10403 12052
rect 10467 11988 10485 12052
rect 10549 11988 10567 12052
rect 10631 11988 10649 12052
rect 10713 11988 10731 12052
rect 10795 11988 10813 12052
rect 10877 11988 10895 12052
rect 10959 11988 10977 12052
rect 11041 11988 11059 12052
rect 11123 11988 11141 12052
rect 11205 11988 11223 12052
rect 11287 11988 11305 12052
rect 11369 11988 11386 12052
rect 11450 11988 11467 12052
rect 11531 11988 11548 12052
rect 11612 11988 11629 12052
rect 11693 11988 11710 12052
rect 11774 11988 11791 12052
rect 11855 11988 11872 12052
rect 11936 11988 11953 12052
rect 12017 11988 12034 12052
rect 12098 11988 12115 12052
rect 12179 11988 12196 12052
rect 12260 11988 12277 12052
rect 12341 11988 12358 12052
rect 12422 11988 12439 12052
rect 12503 11988 12520 12052
rect 12584 11988 12601 12052
rect 12665 11988 12682 12052
rect 12746 11988 12763 12052
rect 12827 11988 12844 12052
rect 12908 11988 12925 12052
rect 12989 11988 13006 12052
rect 13070 11988 13087 12052
rect 13151 11988 13168 12052
rect 13232 11988 13249 12052
rect 13313 11988 13330 12052
rect 13394 11988 13411 12052
rect 13475 11988 13492 12052
rect 13556 11988 13573 12052
rect 13637 11988 13654 12052
rect 13718 11988 13735 12052
rect 13799 11988 13816 12052
rect 13880 11988 13897 12052
rect 13961 11988 13978 12052
rect 14042 11988 14059 12052
rect 14123 11988 14140 12052
rect 14204 11988 14221 12052
rect 14285 11988 14302 12052
rect 14366 11988 14383 12052
rect 14447 11988 14464 12052
rect 14528 11988 14545 12052
rect 14609 11988 14626 12052
rect 14690 11988 14707 12052
rect 14771 11988 14788 12052
rect 14852 11988 15000 12052
rect 0 11970 15000 11988
rect 0 11906 106 11970
rect 170 11906 188 11970
rect 252 11906 270 11970
rect 334 11906 352 11970
rect 416 11906 434 11970
rect 498 11906 516 11970
rect 580 11906 598 11970
rect 662 11906 679 11970
rect 743 11906 760 11970
rect 824 11906 841 11970
rect 905 11906 922 11970
rect 986 11906 1003 11970
rect 1067 11906 1084 11970
rect 1148 11906 1165 11970
rect 1229 11906 1246 11970
rect 1310 11906 1327 11970
rect 1391 11906 1408 11970
rect 1472 11906 1489 11970
rect 1553 11906 1570 11970
rect 1634 11906 1651 11970
rect 1715 11906 1732 11970
rect 1796 11906 1813 11970
rect 1877 11906 1894 11970
rect 1958 11906 1975 11970
rect 2039 11906 2056 11970
rect 2120 11906 2137 11970
rect 2201 11906 2218 11970
rect 2282 11906 2299 11970
rect 2363 11906 2380 11970
rect 2444 11906 2461 11970
rect 2525 11906 2542 11970
rect 2606 11906 2623 11970
rect 2687 11906 2704 11970
rect 2768 11906 2785 11970
rect 2849 11906 2866 11970
rect 2930 11906 2947 11970
rect 3011 11906 3028 11970
rect 3092 11906 3109 11970
rect 3173 11906 3190 11970
rect 3254 11906 3271 11970
rect 3335 11906 3352 11970
rect 3416 11906 3433 11970
rect 3497 11906 3514 11970
rect 3578 11906 3595 11970
rect 3659 11906 3676 11970
rect 3740 11906 3757 11970
rect 3821 11906 3838 11970
rect 3902 11906 3919 11970
rect 3983 11906 4000 11970
rect 4064 11906 4081 11970
rect 4145 11906 4162 11970
rect 4226 11906 4243 11970
rect 4307 11906 4324 11970
rect 4388 11906 4405 11970
rect 4469 11906 4486 11970
rect 4550 11906 4567 11970
rect 4631 11906 4648 11970
rect 4712 11906 4729 11970
rect 4793 11906 4810 11970
rect 4874 11906 10157 11970
rect 10221 11906 10239 11970
rect 10303 11906 10321 11970
rect 10385 11906 10403 11970
rect 10467 11906 10485 11970
rect 10549 11906 10567 11970
rect 10631 11906 10649 11970
rect 10713 11906 10731 11970
rect 10795 11906 10813 11970
rect 10877 11906 10895 11970
rect 10959 11906 10977 11970
rect 11041 11906 11059 11970
rect 11123 11906 11141 11970
rect 11205 11906 11223 11970
rect 11287 11906 11305 11970
rect 11369 11906 11386 11970
rect 11450 11906 11467 11970
rect 11531 11906 11548 11970
rect 11612 11906 11629 11970
rect 11693 11906 11710 11970
rect 11774 11906 11791 11970
rect 11855 11906 11872 11970
rect 11936 11906 11953 11970
rect 12017 11906 12034 11970
rect 12098 11906 12115 11970
rect 12179 11906 12196 11970
rect 12260 11906 12277 11970
rect 12341 11906 12358 11970
rect 12422 11906 12439 11970
rect 12503 11906 12520 11970
rect 12584 11906 12601 11970
rect 12665 11906 12682 11970
rect 12746 11906 12763 11970
rect 12827 11906 12844 11970
rect 12908 11906 12925 11970
rect 12989 11906 13006 11970
rect 13070 11906 13087 11970
rect 13151 11906 13168 11970
rect 13232 11906 13249 11970
rect 13313 11906 13330 11970
rect 13394 11906 13411 11970
rect 13475 11906 13492 11970
rect 13556 11906 13573 11970
rect 13637 11906 13654 11970
rect 13718 11906 13735 11970
rect 13799 11906 13816 11970
rect 13880 11906 13897 11970
rect 13961 11906 13978 11970
rect 14042 11906 14059 11970
rect 14123 11906 14140 11970
rect 14204 11906 14221 11970
rect 14285 11906 14302 11970
rect 14366 11906 14383 11970
rect 14447 11906 14464 11970
rect 14528 11906 14545 11970
rect 14609 11906 14626 11970
rect 14690 11906 14707 11970
rect 14771 11906 14788 11970
rect 14852 11906 15000 11970
rect 0 11888 15000 11906
rect 0 11824 106 11888
rect 170 11824 188 11888
rect 252 11824 270 11888
rect 334 11824 352 11888
rect 416 11824 434 11888
rect 498 11824 516 11888
rect 580 11824 598 11888
rect 662 11824 679 11888
rect 743 11824 760 11888
rect 824 11824 841 11888
rect 905 11824 922 11888
rect 986 11824 1003 11888
rect 1067 11824 1084 11888
rect 1148 11824 1165 11888
rect 1229 11824 1246 11888
rect 1310 11824 1327 11888
rect 1391 11824 1408 11888
rect 1472 11824 1489 11888
rect 1553 11824 1570 11888
rect 1634 11824 1651 11888
rect 1715 11824 1732 11888
rect 1796 11824 1813 11888
rect 1877 11824 1894 11888
rect 1958 11824 1975 11888
rect 2039 11824 2056 11888
rect 2120 11824 2137 11888
rect 2201 11824 2218 11888
rect 2282 11824 2299 11888
rect 2363 11824 2380 11888
rect 2444 11824 2461 11888
rect 2525 11824 2542 11888
rect 2606 11824 2623 11888
rect 2687 11824 2704 11888
rect 2768 11824 2785 11888
rect 2849 11824 2866 11888
rect 2930 11824 2947 11888
rect 3011 11824 3028 11888
rect 3092 11824 3109 11888
rect 3173 11824 3190 11888
rect 3254 11824 3271 11888
rect 3335 11824 3352 11888
rect 3416 11824 3433 11888
rect 3497 11824 3514 11888
rect 3578 11824 3595 11888
rect 3659 11824 3676 11888
rect 3740 11824 3757 11888
rect 3821 11824 3838 11888
rect 3902 11824 3919 11888
rect 3983 11824 4000 11888
rect 4064 11824 4081 11888
rect 4145 11824 4162 11888
rect 4226 11824 4243 11888
rect 4307 11824 4324 11888
rect 4388 11824 4405 11888
rect 4469 11824 4486 11888
rect 4550 11824 4567 11888
rect 4631 11824 4648 11888
rect 4712 11824 4729 11888
rect 4793 11824 4810 11888
rect 4874 11824 10157 11888
rect 10221 11824 10239 11888
rect 10303 11824 10321 11888
rect 10385 11824 10403 11888
rect 10467 11824 10485 11888
rect 10549 11824 10567 11888
rect 10631 11824 10649 11888
rect 10713 11824 10731 11888
rect 10795 11824 10813 11888
rect 10877 11824 10895 11888
rect 10959 11824 10977 11888
rect 11041 11824 11059 11888
rect 11123 11824 11141 11888
rect 11205 11824 11223 11888
rect 11287 11824 11305 11888
rect 11369 11824 11386 11888
rect 11450 11824 11467 11888
rect 11531 11824 11548 11888
rect 11612 11824 11629 11888
rect 11693 11824 11710 11888
rect 11774 11824 11791 11888
rect 11855 11824 11872 11888
rect 11936 11824 11953 11888
rect 12017 11824 12034 11888
rect 12098 11824 12115 11888
rect 12179 11824 12196 11888
rect 12260 11824 12277 11888
rect 12341 11824 12358 11888
rect 12422 11824 12439 11888
rect 12503 11824 12520 11888
rect 12584 11824 12601 11888
rect 12665 11824 12682 11888
rect 12746 11824 12763 11888
rect 12827 11824 12844 11888
rect 12908 11824 12925 11888
rect 12989 11824 13006 11888
rect 13070 11824 13087 11888
rect 13151 11824 13168 11888
rect 13232 11824 13249 11888
rect 13313 11824 13330 11888
rect 13394 11824 13411 11888
rect 13475 11824 13492 11888
rect 13556 11824 13573 11888
rect 13637 11824 13654 11888
rect 13718 11824 13735 11888
rect 13799 11824 13816 11888
rect 13880 11824 13897 11888
rect 13961 11824 13978 11888
rect 14042 11824 14059 11888
rect 14123 11824 14140 11888
rect 14204 11824 14221 11888
rect 14285 11824 14302 11888
rect 14366 11824 14383 11888
rect 14447 11824 14464 11888
rect 14528 11824 14545 11888
rect 14609 11824 14626 11888
rect 14690 11824 14707 11888
rect 14771 11824 14788 11888
rect 14852 11824 15000 11888
rect 0 11806 15000 11824
rect 0 11742 106 11806
rect 170 11742 188 11806
rect 252 11742 270 11806
rect 334 11742 352 11806
rect 416 11742 434 11806
rect 498 11742 516 11806
rect 580 11742 598 11806
rect 662 11742 679 11806
rect 743 11742 760 11806
rect 824 11742 841 11806
rect 905 11742 922 11806
rect 986 11742 1003 11806
rect 1067 11742 1084 11806
rect 1148 11742 1165 11806
rect 1229 11742 1246 11806
rect 1310 11742 1327 11806
rect 1391 11742 1408 11806
rect 1472 11742 1489 11806
rect 1553 11742 1570 11806
rect 1634 11742 1651 11806
rect 1715 11742 1732 11806
rect 1796 11742 1813 11806
rect 1877 11742 1894 11806
rect 1958 11742 1975 11806
rect 2039 11742 2056 11806
rect 2120 11742 2137 11806
rect 2201 11742 2218 11806
rect 2282 11742 2299 11806
rect 2363 11742 2380 11806
rect 2444 11742 2461 11806
rect 2525 11742 2542 11806
rect 2606 11742 2623 11806
rect 2687 11742 2704 11806
rect 2768 11742 2785 11806
rect 2849 11742 2866 11806
rect 2930 11742 2947 11806
rect 3011 11742 3028 11806
rect 3092 11742 3109 11806
rect 3173 11742 3190 11806
rect 3254 11742 3271 11806
rect 3335 11742 3352 11806
rect 3416 11742 3433 11806
rect 3497 11742 3514 11806
rect 3578 11742 3595 11806
rect 3659 11742 3676 11806
rect 3740 11742 3757 11806
rect 3821 11742 3838 11806
rect 3902 11742 3919 11806
rect 3983 11742 4000 11806
rect 4064 11742 4081 11806
rect 4145 11742 4162 11806
rect 4226 11742 4243 11806
rect 4307 11742 4324 11806
rect 4388 11742 4405 11806
rect 4469 11742 4486 11806
rect 4550 11742 4567 11806
rect 4631 11742 4648 11806
rect 4712 11742 4729 11806
rect 4793 11742 4810 11806
rect 4874 11742 10157 11806
rect 10221 11742 10239 11806
rect 10303 11742 10321 11806
rect 10385 11742 10403 11806
rect 10467 11742 10485 11806
rect 10549 11742 10567 11806
rect 10631 11742 10649 11806
rect 10713 11742 10731 11806
rect 10795 11742 10813 11806
rect 10877 11742 10895 11806
rect 10959 11742 10977 11806
rect 11041 11742 11059 11806
rect 11123 11742 11141 11806
rect 11205 11742 11223 11806
rect 11287 11742 11305 11806
rect 11369 11742 11386 11806
rect 11450 11742 11467 11806
rect 11531 11742 11548 11806
rect 11612 11742 11629 11806
rect 11693 11742 11710 11806
rect 11774 11742 11791 11806
rect 11855 11742 11872 11806
rect 11936 11742 11953 11806
rect 12017 11742 12034 11806
rect 12098 11742 12115 11806
rect 12179 11742 12196 11806
rect 12260 11742 12277 11806
rect 12341 11742 12358 11806
rect 12422 11742 12439 11806
rect 12503 11742 12520 11806
rect 12584 11742 12601 11806
rect 12665 11742 12682 11806
rect 12746 11742 12763 11806
rect 12827 11742 12844 11806
rect 12908 11742 12925 11806
rect 12989 11742 13006 11806
rect 13070 11742 13087 11806
rect 13151 11742 13168 11806
rect 13232 11742 13249 11806
rect 13313 11742 13330 11806
rect 13394 11742 13411 11806
rect 13475 11742 13492 11806
rect 13556 11742 13573 11806
rect 13637 11742 13654 11806
rect 13718 11742 13735 11806
rect 13799 11742 13816 11806
rect 13880 11742 13897 11806
rect 13961 11742 13978 11806
rect 14042 11742 14059 11806
rect 14123 11742 14140 11806
rect 14204 11742 14221 11806
rect 14285 11742 14302 11806
rect 14366 11742 14383 11806
rect 14447 11742 14464 11806
rect 14528 11742 14545 11806
rect 14609 11742 14626 11806
rect 14690 11742 14707 11806
rect 14771 11742 14788 11806
rect 14852 11742 15000 11806
rect 0 11724 15000 11742
rect 0 11660 106 11724
rect 170 11660 188 11724
rect 252 11660 270 11724
rect 334 11660 352 11724
rect 416 11660 434 11724
rect 498 11660 516 11724
rect 580 11660 598 11724
rect 662 11660 679 11724
rect 743 11660 760 11724
rect 824 11660 841 11724
rect 905 11660 922 11724
rect 986 11660 1003 11724
rect 1067 11660 1084 11724
rect 1148 11660 1165 11724
rect 1229 11660 1246 11724
rect 1310 11660 1327 11724
rect 1391 11660 1408 11724
rect 1472 11660 1489 11724
rect 1553 11660 1570 11724
rect 1634 11660 1651 11724
rect 1715 11660 1732 11724
rect 1796 11660 1813 11724
rect 1877 11660 1894 11724
rect 1958 11660 1975 11724
rect 2039 11660 2056 11724
rect 2120 11660 2137 11724
rect 2201 11660 2218 11724
rect 2282 11660 2299 11724
rect 2363 11660 2380 11724
rect 2444 11660 2461 11724
rect 2525 11660 2542 11724
rect 2606 11660 2623 11724
rect 2687 11660 2704 11724
rect 2768 11660 2785 11724
rect 2849 11660 2866 11724
rect 2930 11660 2947 11724
rect 3011 11660 3028 11724
rect 3092 11660 3109 11724
rect 3173 11660 3190 11724
rect 3254 11660 3271 11724
rect 3335 11660 3352 11724
rect 3416 11660 3433 11724
rect 3497 11660 3514 11724
rect 3578 11660 3595 11724
rect 3659 11660 3676 11724
rect 3740 11660 3757 11724
rect 3821 11660 3838 11724
rect 3902 11660 3919 11724
rect 3983 11660 4000 11724
rect 4064 11660 4081 11724
rect 4145 11660 4162 11724
rect 4226 11660 4243 11724
rect 4307 11660 4324 11724
rect 4388 11660 4405 11724
rect 4469 11660 4486 11724
rect 4550 11660 4567 11724
rect 4631 11660 4648 11724
rect 4712 11660 4729 11724
rect 4793 11660 4810 11724
rect 4874 11660 10157 11724
rect 10221 11660 10239 11724
rect 10303 11660 10321 11724
rect 10385 11660 10403 11724
rect 10467 11660 10485 11724
rect 10549 11660 10567 11724
rect 10631 11660 10649 11724
rect 10713 11660 10731 11724
rect 10795 11660 10813 11724
rect 10877 11660 10895 11724
rect 10959 11660 10977 11724
rect 11041 11660 11059 11724
rect 11123 11660 11141 11724
rect 11205 11660 11223 11724
rect 11287 11660 11305 11724
rect 11369 11660 11386 11724
rect 11450 11660 11467 11724
rect 11531 11660 11548 11724
rect 11612 11660 11629 11724
rect 11693 11660 11710 11724
rect 11774 11660 11791 11724
rect 11855 11660 11872 11724
rect 11936 11660 11953 11724
rect 12017 11660 12034 11724
rect 12098 11660 12115 11724
rect 12179 11660 12196 11724
rect 12260 11660 12277 11724
rect 12341 11660 12358 11724
rect 12422 11660 12439 11724
rect 12503 11660 12520 11724
rect 12584 11660 12601 11724
rect 12665 11660 12682 11724
rect 12746 11660 12763 11724
rect 12827 11660 12844 11724
rect 12908 11660 12925 11724
rect 12989 11660 13006 11724
rect 13070 11660 13087 11724
rect 13151 11660 13168 11724
rect 13232 11660 13249 11724
rect 13313 11660 13330 11724
rect 13394 11660 13411 11724
rect 13475 11660 13492 11724
rect 13556 11660 13573 11724
rect 13637 11660 13654 11724
rect 13718 11660 13735 11724
rect 13799 11660 13816 11724
rect 13880 11660 13897 11724
rect 13961 11660 13978 11724
rect 14042 11660 14059 11724
rect 14123 11660 14140 11724
rect 14204 11660 14221 11724
rect 14285 11660 14302 11724
rect 14366 11660 14383 11724
rect 14447 11660 14464 11724
rect 14528 11660 14545 11724
rect 14609 11660 14626 11724
rect 14690 11660 14707 11724
rect 14771 11660 14788 11724
rect 14852 11660 15000 11724
rect 0 11642 15000 11660
rect 0 11578 106 11642
rect 170 11578 188 11642
rect 252 11578 270 11642
rect 334 11578 352 11642
rect 416 11578 434 11642
rect 498 11578 516 11642
rect 580 11578 598 11642
rect 662 11578 679 11642
rect 743 11578 760 11642
rect 824 11578 841 11642
rect 905 11578 922 11642
rect 986 11578 1003 11642
rect 1067 11578 1084 11642
rect 1148 11578 1165 11642
rect 1229 11578 1246 11642
rect 1310 11578 1327 11642
rect 1391 11578 1408 11642
rect 1472 11578 1489 11642
rect 1553 11578 1570 11642
rect 1634 11578 1651 11642
rect 1715 11578 1732 11642
rect 1796 11578 1813 11642
rect 1877 11578 1894 11642
rect 1958 11578 1975 11642
rect 2039 11578 2056 11642
rect 2120 11578 2137 11642
rect 2201 11578 2218 11642
rect 2282 11578 2299 11642
rect 2363 11578 2380 11642
rect 2444 11578 2461 11642
rect 2525 11578 2542 11642
rect 2606 11578 2623 11642
rect 2687 11578 2704 11642
rect 2768 11578 2785 11642
rect 2849 11578 2866 11642
rect 2930 11578 2947 11642
rect 3011 11578 3028 11642
rect 3092 11578 3109 11642
rect 3173 11578 3190 11642
rect 3254 11578 3271 11642
rect 3335 11578 3352 11642
rect 3416 11578 3433 11642
rect 3497 11578 3514 11642
rect 3578 11578 3595 11642
rect 3659 11578 3676 11642
rect 3740 11578 3757 11642
rect 3821 11578 3838 11642
rect 3902 11578 3919 11642
rect 3983 11578 4000 11642
rect 4064 11578 4081 11642
rect 4145 11578 4162 11642
rect 4226 11578 4243 11642
rect 4307 11578 4324 11642
rect 4388 11578 4405 11642
rect 4469 11578 4486 11642
rect 4550 11578 4567 11642
rect 4631 11578 4648 11642
rect 4712 11578 4729 11642
rect 4793 11578 4810 11642
rect 4874 11578 10157 11642
rect 10221 11578 10239 11642
rect 10303 11578 10321 11642
rect 10385 11578 10403 11642
rect 10467 11578 10485 11642
rect 10549 11578 10567 11642
rect 10631 11578 10649 11642
rect 10713 11578 10731 11642
rect 10795 11578 10813 11642
rect 10877 11578 10895 11642
rect 10959 11578 10977 11642
rect 11041 11578 11059 11642
rect 11123 11578 11141 11642
rect 11205 11578 11223 11642
rect 11287 11578 11305 11642
rect 11369 11578 11386 11642
rect 11450 11578 11467 11642
rect 11531 11578 11548 11642
rect 11612 11578 11629 11642
rect 11693 11578 11710 11642
rect 11774 11578 11791 11642
rect 11855 11578 11872 11642
rect 11936 11578 11953 11642
rect 12017 11578 12034 11642
rect 12098 11578 12115 11642
rect 12179 11578 12196 11642
rect 12260 11578 12277 11642
rect 12341 11578 12358 11642
rect 12422 11578 12439 11642
rect 12503 11578 12520 11642
rect 12584 11578 12601 11642
rect 12665 11578 12682 11642
rect 12746 11578 12763 11642
rect 12827 11578 12844 11642
rect 12908 11578 12925 11642
rect 12989 11578 13006 11642
rect 13070 11578 13087 11642
rect 13151 11578 13168 11642
rect 13232 11578 13249 11642
rect 13313 11578 13330 11642
rect 13394 11578 13411 11642
rect 13475 11578 13492 11642
rect 13556 11578 13573 11642
rect 13637 11578 13654 11642
rect 13718 11578 13735 11642
rect 13799 11578 13816 11642
rect 13880 11578 13897 11642
rect 13961 11578 13978 11642
rect 14042 11578 14059 11642
rect 14123 11578 14140 11642
rect 14204 11578 14221 11642
rect 14285 11578 14302 11642
rect 14366 11578 14383 11642
rect 14447 11578 14464 11642
rect 14528 11578 14545 11642
rect 14609 11578 14626 11642
rect 14690 11578 14707 11642
rect 14771 11578 14788 11642
rect 14852 11578 15000 11642
rect 0 11560 15000 11578
rect 0 11496 106 11560
rect 170 11496 188 11560
rect 252 11496 270 11560
rect 334 11496 352 11560
rect 416 11496 434 11560
rect 498 11496 516 11560
rect 580 11496 598 11560
rect 662 11496 679 11560
rect 743 11496 760 11560
rect 824 11496 841 11560
rect 905 11496 922 11560
rect 986 11496 1003 11560
rect 1067 11496 1084 11560
rect 1148 11496 1165 11560
rect 1229 11496 1246 11560
rect 1310 11496 1327 11560
rect 1391 11496 1408 11560
rect 1472 11496 1489 11560
rect 1553 11496 1570 11560
rect 1634 11496 1651 11560
rect 1715 11496 1732 11560
rect 1796 11496 1813 11560
rect 1877 11496 1894 11560
rect 1958 11496 1975 11560
rect 2039 11496 2056 11560
rect 2120 11496 2137 11560
rect 2201 11496 2218 11560
rect 2282 11496 2299 11560
rect 2363 11496 2380 11560
rect 2444 11496 2461 11560
rect 2525 11496 2542 11560
rect 2606 11496 2623 11560
rect 2687 11496 2704 11560
rect 2768 11496 2785 11560
rect 2849 11496 2866 11560
rect 2930 11496 2947 11560
rect 3011 11496 3028 11560
rect 3092 11496 3109 11560
rect 3173 11496 3190 11560
rect 3254 11496 3271 11560
rect 3335 11496 3352 11560
rect 3416 11496 3433 11560
rect 3497 11496 3514 11560
rect 3578 11496 3595 11560
rect 3659 11496 3676 11560
rect 3740 11496 3757 11560
rect 3821 11496 3838 11560
rect 3902 11496 3919 11560
rect 3983 11496 4000 11560
rect 4064 11496 4081 11560
rect 4145 11496 4162 11560
rect 4226 11496 4243 11560
rect 4307 11496 4324 11560
rect 4388 11496 4405 11560
rect 4469 11496 4486 11560
rect 4550 11496 4567 11560
rect 4631 11496 4648 11560
rect 4712 11496 4729 11560
rect 4793 11496 4810 11560
rect 4874 11496 10157 11560
rect 10221 11496 10239 11560
rect 10303 11496 10321 11560
rect 10385 11496 10403 11560
rect 10467 11496 10485 11560
rect 10549 11496 10567 11560
rect 10631 11496 10649 11560
rect 10713 11496 10731 11560
rect 10795 11496 10813 11560
rect 10877 11496 10895 11560
rect 10959 11496 10977 11560
rect 11041 11496 11059 11560
rect 11123 11496 11141 11560
rect 11205 11496 11223 11560
rect 11287 11496 11305 11560
rect 11369 11496 11386 11560
rect 11450 11496 11467 11560
rect 11531 11496 11548 11560
rect 11612 11496 11629 11560
rect 11693 11496 11710 11560
rect 11774 11496 11791 11560
rect 11855 11496 11872 11560
rect 11936 11496 11953 11560
rect 12017 11496 12034 11560
rect 12098 11496 12115 11560
rect 12179 11496 12196 11560
rect 12260 11496 12277 11560
rect 12341 11496 12358 11560
rect 12422 11496 12439 11560
rect 12503 11496 12520 11560
rect 12584 11496 12601 11560
rect 12665 11496 12682 11560
rect 12746 11496 12763 11560
rect 12827 11496 12844 11560
rect 12908 11496 12925 11560
rect 12989 11496 13006 11560
rect 13070 11496 13087 11560
rect 13151 11496 13168 11560
rect 13232 11496 13249 11560
rect 13313 11496 13330 11560
rect 13394 11496 13411 11560
rect 13475 11496 13492 11560
rect 13556 11496 13573 11560
rect 13637 11496 13654 11560
rect 13718 11496 13735 11560
rect 13799 11496 13816 11560
rect 13880 11496 13897 11560
rect 13961 11496 13978 11560
rect 14042 11496 14059 11560
rect 14123 11496 14140 11560
rect 14204 11496 14221 11560
rect 14285 11496 14302 11560
rect 14366 11496 14383 11560
rect 14447 11496 14464 11560
rect 14528 11496 14545 11560
rect 14609 11496 14626 11560
rect 14690 11496 14707 11560
rect 14771 11496 14788 11560
rect 14852 11496 15000 11560
rect 0 11478 15000 11496
rect 0 11414 106 11478
rect 170 11414 188 11478
rect 252 11414 270 11478
rect 334 11414 352 11478
rect 416 11414 434 11478
rect 498 11414 516 11478
rect 580 11414 598 11478
rect 662 11414 679 11478
rect 743 11414 760 11478
rect 824 11414 841 11478
rect 905 11414 922 11478
rect 986 11414 1003 11478
rect 1067 11414 1084 11478
rect 1148 11414 1165 11478
rect 1229 11414 1246 11478
rect 1310 11414 1327 11478
rect 1391 11414 1408 11478
rect 1472 11414 1489 11478
rect 1553 11414 1570 11478
rect 1634 11414 1651 11478
rect 1715 11414 1732 11478
rect 1796 11414 1813 11478
rect 1877 11414 1894 11478
rect 1958 11414 1975 11478
rect 2039 11414 2056 11478
rect 2120 11414 2137 11478
rect 2201 11414 2218 11478
rect 2282 11414 2299 11478
rect 2363 11414 2380 11478
rect 2444 11414 2461 11478
rect 2525 11414 2542 11478
rect 2606 11414 2623 11478
rect 2687 11414 2704 11478
rect 2768 11414 2785 11478
rect 2849 11414 2866 11478
rect 2930 11414 2947 11478
rect 3011 11414 3028 11478
rect 3092 11414 3109 11478
rect 3173 11414 3190 11478
rect 3254 11414 3271 11478
rect 3335 11414 3352 11478
rect 3416 11414 3433 11478
rect 3497 11414 3514 11478
rect 3578 11414 3595 11478
rect 3659 11414 3676 11478
rect 3740 11414 3757 11478
rect 3821 11414 3838 11478
rect 3902 11414 3919 11478
rect 3983 11414 4000 11478
rect 4064 11414 4081 11478
rect 4145 11414 4162 11478
rect 4226 11414 4243 11478
rect 4307 11414 4324 11478
rect 4388 11414 4405 11478
rect 4469 11414 4486 11478
rect 4550 11414 4567 11478
rect 4631 11414 4648 11478
rect 4712 11414 4729 11478
rect 4793 11414 4810 11478
rect 4874 11414 10157 11478
rect 10221 11414 10239 11478
rect 10303 11414 10321 11478
rect 10385 11414 10403 11478
rect 10467 11414 10485 11478
rect 10549 11414 10567 11478
rect 10631 11414 10649 11478
rect 10713 11414 10731 11478
rect 10795 11414 10813 11478
rect 10877 11414 10895 11478
rect 10959 11414 10977 11478
rect 11041 11414 11059 11478
rect 11123 11414 11141 11478
rect 11205 11414 11223 11478
rect 11287 11414 11305 11478
rect 11369 11414 11386 11478
rect 11450 11414 11467 11478
rect 11531 11414 11548 11478
rect 11612 11414 11629 11478
rect 11693 11414 11710 11478
rect 11774 11414 11791 11478
rect 11855 11414 11872 11478
rect 11936 11414 11953 11478
rect 12017 11414 12034 11478
rect 12098 11414 12115 11478
rect 12179 11414 12196 11478
rect 12260 11414 12277 11478
rect 12341 11414 12358 11478
rect 12422 11414 12439 11478
rect 12503 11414 12520 11478
rect 12584 11414 12601 11478
rect 12665 11414 12682 11478
rect 12746 11414 12763 11478
rect 12827 11414 12844 11478
rect 12908 11414 12925 11478
rect 12989 11414 13006 11478
rect 13070 11414 13087 11478
rect 13151 11414 13168 11478
rect 13232 11414 13249 11478
rect 13313 11414 13330 11478
rect 13394 11414 13411 11478
rect 13475 11414 13492 11478
rect 13556 11414 13573 11478
rect 13637 11414 13654 11478
rect 13718 11414 13735 11478
rect 13799 11414 13816 11478
rect 13880 11414 13897 11478
rect 13961 11414 13978 11478
rect 14042 11414 14059 11478
rect 14123 11414 14140 11478
rect 14204 11414 14221 11478
rect 14285 11414 14302 11478
rect 14366 11414 14383 11478
rect 14447 11414 14464 11478
rect 14528 11414 14545 11478
rect 14609 11414 14626 11478
rect 14690 11414 14707 11478
rect 14771 11414 14788 11478
rect 14852 11414 15000 11478
rect 0 11396 15000 11414
rect 0 11332 106 11396
rect 170 11332 188 11396
rect 252 11332 270 11396
rect 334 11332 352 11396
rect 416 11332 434 11396
rect 498 11332 516 11396
rect 580 11332 598 11396
rect 662 11332 679 11396
rect 743 11332 760 11396
rect 824 11332 841 11396
rect 905 11332 922 11396
rect 986 11332 1003 11396
rect 1067 11332 1084 11396
rect 1148 11332 1165 11396
rect 1229 11332 1246 11396
rect 1310 11332 1327 11396
rect 1391 11332 1408 11396
rect 1472 11332 1489 11396
rect 1553 11332 1570 11396
rect 1634 11332 1651 11396
rect 1715 11332 1732 11396
rect 1796 11332 1813 11396
rect 1877 11332 1894 11396
rect 1958 11332 1975 11396
rect 2039 11332 2056 11396
rect 2120 11332 2137 11396
rect 2201 11332 2218 11396
rect 2282 11332 2299 11396
rect 2363 11332 2380 11396
rect 2444 11332 2461 11396
rect 2525 11332 2542 11396
rect 2606 11332 2623 11396
rect 2687 11332 2704 11396
rect 2768 11332 2785 11396
rect 2849 11332 2866 11396
rect 2930 11332 2947 11396
rect 3011 11332 3028 11396
rect 3092 11332 3109 11396
rect 3173 11332 3190 11396
rect 3254 11332 3271 11396
rect 3335 11332 3352 11396
rect 3416 11332 3433 11396
rect 3497 11332 3514 11396
rect 3578 11332 3595 11396
rect 3659 11332 3676 11396
rect 3740 11332 3757 11396
rect 3821 11332 3838 11396
rect 3902 11332 3919 11396
rect 3983 11332 4000 11396
rect 4064 11332 4081 11396
rect 4145 11332 4162 11396
rect 4226 11332 4243 11396
rect 4307 11332 4324 11396
rect 4388 11332 4405 11396
rect 4469 11332 4486 11396
rect 4550 11332 4567 11396
rect 4631 11332 4648 11396
rect 4712 11332 4729 11396
rect 4793 11332 4810 11396
rect 4874 11332 10157 11396
rect 10221 11332 10239 11396
rect 10303 11332 10321 11396
rect 10385 11332 10403 11396
rect 10467 11332 10485 11396
rect 10549 11332 10567 11396
rect 10631 11332 10649 11396
rect 10713 11332 10731 11396
rect 10795 11332 10813 11396
rect 10877 11332 10895 11396
rect 10959 11332 10977 11396
rect 11041 11332 11059 11396
rect 11123 11332 11141 11396
rect 11205 11332 11223 11396
rect 11287 11332 11305 11396
rect 11369 11332 11386 11396
rect 11450 11332 11467 11396
rect 11531 11332 11548 11396
rect 11612 11332 11629 11396
rect 11693 11332 11710 11396
rect 11774 11332 11791 11396
rect 11855 11332 11872 11396
rect 11936 11332 11953 11396
rect 12017 11332 12034 11396
rect 12098 11332 12115 11396
rect 12179 11332 12196 11396
rect 12260 11332 12277 11396
rect 12341 11332 12358 11396
rect 12422 11332 12439 11396
rect 12503 11332 12520 11396
rect 12584 11332 12601 11396
rect 12665 11332 12682 11396
rect 12746 11332 12763 11396
rect 12827 11332 12844 11396
rect 12908 11332 12925 11396
rect 12989 11332 13006 11396
rect 13070 11332 13087 11396
rect 13151 11332 13168 11396
rect 13232 11332 13249 11396
rect 13313 11332 13330 11396
rect 13394 11332 13411 11396
rect 13475 11332 13492 11396
rect 13556 11332 13573 11396
rect 13637 11332 13654 11396
rect 13718 11332 13735 11396
rect 13799 11332 13816 11396
rect 13880 11332 13897 11396
rect 13961 11332 13978 11396
rect 14042 11332 14059 11396
rect 14123 11332 14140 11396
rect 14204 11332 14221 11396
rect 14285 11332 14302 11396
rect 14366 11332 14383 11396
rect 14447 11332 14464 11396
rect 14528 11332 14545 11396
rect 14609 11332 14626 11396
rect 14690 11332 14707 11396
rect 14771 11332 14788 11396
rect 14852 11332 15000 11396
rect 0 11314 15000 11332
rect 0 11250 106 11314
rect 170 11250 188 11314
rect 252 11250 270 11314
rect 334 11250 352 11314
rect 416 11250 434 11314
rect 498 11250 516 11314
rect 580 11250 598 11314
rect 662 11250 679 11314
rect 743 11250 760 11314
rect 824 11250 841 11314
rect 905 11250 922 11314
rect 986 11250 1003 11314
rect 1067 11250 1084 11314
rect 1148 11250 1165 11314
rect 1229 11250 1246 11314
rect 1310 11250 1327 11314
rect 1391 11250 1408 11314
rect 1472 11250 1489 11314
rect 1553 11250 1570 11314
rect 1634 11250 1651 11314
rect 1715 11250 1732 11314
rect 1796 11250 1813 11314
rect 1877 11250 1894 11314
rect 1958 11250 1975 11314
rect 2039 11250 2056 11314
rect 2120 11250 2137 11314
rect 2201 11250 2218 11314
rect 2282 11250 2299 11314
rect 2363 11250 2380 11314
rect 2444 11250 2461 11314
rect 2525 11250 2542 11314
rect 2606 11250 2623 11314
rect 2687 11250 2704 11314
rect 2768 11250 2785 11314
rect 2849 11250 2866 11314
rect 2930 11250 2947 11314
rect 3011 11250 3028 11314
rect 3092 11250 3109 11314
rect 3173 11250 3190 11314
rect 3254 11250 3271 11314
rect 3335 11250 3352 11314
rect 3416 11250 3433 11314
rect 3497 11250 3514 11314
rect 3578 11250 3595 11314
rect 3659 11250 3676 11314
rect 3740 11250 3757 11314
rect 3821 11250 3838 11314
rect 3902 11250 3919 11314
rect 3983 11250 4000 11314
rect 4064 11250 4081 11314
rect 4145 11250 4162 11314
rect 4226 11250 4243 11314
rect 4307 11250 4324 11314
rect 4388 11250 4405 11314
rect 4469 11250 4486 11314
rect 4550 11250 4567 11314
rect 4631 11250 4648 11314
rect 4712 11250 4729 11314
rect 4793 11250 4810 11314
rect 4874 11250 10157 11314
rect 10221 11250 10239 11314
rect 10303 11250 10321 11314
rect 10385 11250 10403 11314
rect 10467 11250 10485 11314
rect 10549 11250 10567 11314
rect 10631 11250 10649 11314
rect 10713 11250 10731 11314
rect 10795 11250 10813 11314
rect 10877 11250 10895 11314
rect 10959 11250 10977 11314
rect 11041 11250 11059 11314
rect 11123 11250 11141 11314
rect 11205 11250 11223 11314
rect 11287 11250 11305 11314
rect 11369 11250 11386 11314
rect 11450 11250 11467 11314
rect 11531 11250 11548 11314
rect 11612 11250 11629 11314
rect 11693 11250 11710 11314
rect 11774 11250 11791 11314
rect 11855 11250 11872 11314
rect 11936 11250 11953 11314
rect 12017 11250 12034 11314
rect 12098 11250 12115 11314
rect 12179 11250 12196 11314
rect 12260 11250 12277 11314
rect 12341 11250 12358 11314
rect 12422 11250 12439 11314
rect 12503 11250 12520 11314
rect 12584 11250 12601 11314
rect 12665 11250 12682 11314
rect 12746 11250 12763 11314
rect 12827 11250 12844 11314
rect 12908 11250 12925 11314
rect 12989 11250 13006 11314
rect 13070 11250 13087 11314
rect 13151 11250 13168 11314
rect 13232 11250 13249 11314
rect 13313 11250 13330 11314
rect 13394 11250 13411 11314
rect 13475 11250 13492 11314
rect 13556 11250 13573 11314
rect 13637 11250 13654 11314
rect 13718 11250 13735 11314
rect 13799 11250 13816 11314
rect 13880 11250 13897 11314
rect 13961 11250 13978 11314
rect 14042 11250 14059 11314
rect 14123 11250 14140 11314
rect 14204 11250 14221 11314
rect 14285 11250 14302 11314
rect 14366 11250 14383 11314
rect 14447 11250 14464 11314
rect 14528 11250 14545 11314
rect 14609 11250 14626 11314
rect 14690 11250 14707 11314
rect 14771 11250 14788 11314
rect 14852 11250 15000 11314
rect 0 10901 15000 11250
rect 0 9949 15000 10145
rect 0 5694 15000 9193
rect 0 5630 106 5694
rect 170 5630 188 5694
rect 252 5630 270 5694
rect 334 5630 352 5694
rect 416 5630 434 5694
rect 498 5630 516 5694
rect 580 5630 598 5694
rect 662 5630 679 5694
rect 743 5630 760 5694
rect 824 5630 841 5694
rect 905 5630 922 5694
rect 986 5630 1003 5694
rect 1067 5630 1084 5694
rect 1148 5630 1165 5694
rect 1229 5630 1246 5694
rect 1310 5630 1327 5694
rect 1391 5630 1408 5694
rect 1472 5630 1489 5694
rect 1553 5630 1570 5694
rect 1634 5630 1651 5694
rect 1715 5630 1732 5694
rect 1796 5630 1813 5694
rect 1877 5630 1894 5694
rect 1958 5630 1975 5694
rect 2039 5630 2056 5694
rect 2120 5630 2137 5694
rect 2201 5630 2218 5694
rect 2282 5630 2299 5694
rect 2363 5630 2380 5694
rect 2444 5630 2461 5694
rect 2525 5630 2542 5694
rect 2606 5630 2623 5694
rect 2687 5630 2704 5694
rect 2768 5630 2785 5694
rect 2849 5630 2866 5694
rect 2930 5630 2947 5694
rect 3011 5630 3028 5694
rect 3092 5630 3109 5694
rect 3173 5630 3190 5694
rect 3254 5630 3271 5694
rect 3335 5630 3352 5694
rect 3416 5630 3433 5694
rect 3497 5630 3514 5694
rect 3578 5630 3595 5694
rect 3659 5630 3676 5694
rect 3740 5630 3757 5694
rect 3821 5630 3838 5694
rect 3902 5630 3919 5694
rect 3983 5630 4000 5694
rect 4064 5630 4081 5694
rect 4145 5630 4162 5694
rect 4226 5630 4243 5694
rect 4307 5630 4324 5694
rect 4388 5630 4405 5694
rect 4469 5630 4486 5694
rect 4550 5630 4567 5694
rect 4631 5630 4648 5694
rect 4712 5630 4729 5694
rect 4793 5630 4810 5694
rect 4874 5630 10157 5694
rect 10221 5630 10239 5694
rect 10303 5630 10321 5694
rect 10385 5630 10403 5694
rect 10467 5630 10485 5694
rect 10549 5630 10567 5694
rect 10631 5630 10649 5694
rect 10713 5630 10731 5694
rect 10795 5630 10813 5694
rect 10877 5630 10895 5694
rect 10959 5630 10977 5694
rect 11041 5630 11059 5694
rect 11123 5630 11141 5694
rect 11205 5630 11223 5694
rect 11287 5630 11305 5694
rect 11369 5630 11386 5694
rect 11450 5630 11467 5694
rect 11531 5630 11548 5694
rect 11612 5630 11629 5694
rect 11693 5630 11710 5694
rect 11774 5630 11791 5694
rect 11855 5630 11872 5694
rect 11936 5630 11953 5694
rect 12017 5630 12034 5694
rect 12098 5630 12115 5694
rect 12179 5630 12196 5694
rect 12260 5630 12277 5694
rect 12341 5630 12358 5694
rect 12422 5630 12439 5694
rect 12503 5630 12520 5694
rect 12584 5630 12601 5694
rect 12665 5630 12682 5694
rect 12746 5630 12763 5694
rect 12827 5630 12844 5694
rect 12908 5630 12925 5694
rect 12989 5630 13006 5694
rect 13070 5630 13087 5694
rect 13151 5630 13168 5694
rect 13232 5630 13249 5694
rect 13313 5630 13330 5694
rect 13394 5630 13411 5694
rect 13475 5630 13492 5694
rect 13556 5630 13573 5694
rect 13637 5630 13654 5694
rect 13718 5630 13735 5694
rect 13799 5630 13816 5694
rect 13880 5630 13897 5694
rect 13961 5630 13978 5694
rect 14042 5630 14059 5694
rect 14123 5630 14140 5694
rect 14204 5630 14221 5694
rect 14285 5630 14302 5694
rect 14366 5630 14383 5694
rect 14447 5630 14464 5694
rect 14528 5630 14545 5694
rect 14609 5630 14626 5694
rect 14690 5630 14707 5694
rect 14771 5630 14788 5694
rect 14852 5630 15000 5694
rect 0 5608 15000 5630
rect 0 5544 106 5608
rect 170 5544 188 5608
rect 252 5544 270 5608
rect 334 5544 352 5608
rect 416 5544 434 5608
rect 498 5544 516 5608
rect 580 5544 598 5608
rect 662 5544 679 5608
rect 743 5544 760 5608
rect 824 5544 841 5608
rect 905 5544 922 5608
rect 986 5544 1003 5608
rect 1067 5544 1084 5608
rect 1148 5544 1165 5608
rect 1229 5544 1246 5608
rect 1310 5544 1327 5608
rect 1391 5544 1408 5608
rect 1472 5544 1489 5608
rect 1553 5544 1570 5608
rect 1634 5544 1651 5608
rect 1715 5544 1732 5608
rect 1796 5544 1813 5608
rect 1877 5544 1894 5608
rect 1958 5544 1975 5608
rect 2039 5544 2056 5608
rect 2120 5544 2137 5608
rect 2201 5544 2218 5608
rect 2282 5544 2299 5608
rect 2363 5544 2380 5608
rect 2444 5544 2461 5608
rect 2525 5544 2542 5608
rect 2606 5544 2623 5608
rect 2687 5544 2704 5608
rect 2768 5544 2785 5608
rect 2849 5544 2866 5608
rect 2930 5544 2947 5608
rect 3011 5544 3028 5608
rect 3092 5544 3109 5608
rect 3173 5544 3190 5608
rect 3254 5544 3271 5608
rect 3335 5544 3352 5608
rect 3416 5544 3433 5608
rect 3497 5544 3514 5608
rect 3578 5544 3595 5608
rect 3659 5544 3676 5608
rect 3740 5544 3757 5608
rect 3821 5544 3838 5608
rect 3902 5544 3919 5608
rect 3983 5544 4000 5608
rect 4064 5544 4081 5608
rect 4145 5544 4162 5608
rect 4226 5544 4243 5608
rect 4307 5544 4324 5608
rect 4388 5544 4405 5608
rect 4469 5544 4486 5608
rect 4550 5544 4567 5608
rect 4631 5544 4648 5608
rect 4712 5544 4729 5608
rect 4793 5544 4810 5608
rect 4874 5544 10157 5608
rect 10221 5544 10239 5608
rect 10303 5544 10321 5608
rect 10385 5544 10403 5608
rect 10467 5544 10485 5608
rect 10549 5544 10567 5608
rect 10631 5544 10649 5608
rect 10713 5544 10731 5608
rect 10795 5544 10813 5608
rect 10877 5544 10895 5608
rect 10959 5544 10977 5608
rect 11041 5544 11059 5608
rect 11123 5544 11141 5608
rect 11205 5544 11223 5608
rect 11287 5544 11305 5608
rect 11369 5544 11386 5608
rect 11450 5544 11467 5608
rect 11531 5544 11548 5608
rect 11612 5544 11629 5608
rect 11693 5544 11710 5608
rect 11774 5544 11791 5608
rect 11855 5544 11872 5608
rect 11936 5544 11953 5608
rect 12017 5544 12034 5608
rect 12098 5544 12115 5608
rect 12179 5544 12196 5608
rect 12260 5544 12277 5608
rect 12341 5544 12358 5608
rect 12422 5544 12439 5608
rect 12503 5544 12520 5608
rect 12584 5544 12601 5608
rect 12665 5544 12682 5608
rect 12746 5544 12763 5608
rect 12827 5544 12844 5608
rect 12908 5544 12925 5608
rect 12989 5544 13006 5608
rect 13070 5544 13087 5608
rect 13151 5544 13168 5608
rect 13232 5544 13249 5608
rect 13313 5544 13330 5608
rect 13394 5544 13411 5608
rect 13475 5544 13492 5608
rect 13556 5544 13573 5608
rect 13637 5544 13654 5608
rect 13718 5544 13735 5608
rect 13799 5544 13816 5608
rect 13880 5544 13897 5608
rect 13961 5544 13978 5608
rect 14042 5544 14059 5608
rect 14123 5544 14140 5608
rect 14204 5544 14221 5608
rect 14285 5544 14302 5608
rect 14366 5544 14383 5608
rect 14447 5544 14464 5608
rect 14528 5544 14545 5608
rect 14609 5544 14626 5608
rect 14690 5544 14707 5608
rect 14771 5544 14788 5608
rect 14852 5544 15000 5608
rect 0 5522 15000 5544
rect 0 5458 106 5522
rect 170 5458 188 5522
rect 252 5458 270 5522
rect 334 5458 352 5522
rect 416 5458 434 5522
rect 498 5458 516 5522
rect 580 5458 598 5522
rect 662 5458 679 5522
rect 743 5458 760 5522
rect 824 5458 841 5522
rect 905 5458 922 5522
rect 986 5458 1003 5522
rect 1067 5458 1084 5522
rect 1148 5458 1165 5522
rect 1229 5458 1246 5522
rect 1310 5458 1327 5522
rect 1391 5458 1408 5522
rect 1472 5458 1489 5522
rect 1553 5458 1570 5522
rect 1634 5458 1651 5522
rect 1715 5458 1732 5522
rect 1796 5458 1813 5522
rect 1877 5458 1894 5522
rect 1958 5458 1975 5522
rect 2039 5458 2056 5522
rect 2120 5458 2137 5522
rect 2201 5458 2218 5522
rect 2282 5458 2299 5522
rect 2363 5458 2380 5522
rect 2444 5458 2461 5522
rect 2525 5458 2542 5522
rect 2606 5458 2623 5522
rect 2687 5458 2704 5522
rect 2768 5458 2785 5522
rect 2849 5458 2866 5522
rect 2930 5458 2947 5522
rect 3011 5458 3028 5522
rect 3092 5458 3109 5522
rect 3173 5458 3190 5522
rect 3254 5458 3271 5522
rect 3335 5458 3352 5522
rect 3416 5458 3433 5522
rect 3497 5458 3514 5522
rect 3578 5458 3595 5522
rect 3659 5458 3676 5522
rect 3740 5458 3757 5522
rect 3821 5458 3838 5522
rect 3902 5458 3919 5522
rect 3983 5458 4000 5522
rect 4064 5458 4081 5522
rect 4145 5458 4162 5522
rect 4226 5458 4243 5522
rect 4307 5458 4324 5522
rect 4388 5458 4405 5522
rect 4469 5458 4486 5522
rect 4550 5458 4567 5522
rect 4631 5458 4648 5522
rect 4712 5458 4729 5522
rect 4793 5458 4810 5522
rect 4874 5458 10157 5522
rect 10221 5458 10239 5522
rect 10303 5458 10321 5522
rect 10385 5458 10403 5522
rect 10467 5458 10485 5522
rect 10549 5458 10567 5522
rect 10631 5458 10649 5522
rect 10713 5458 10731 5522
rect 10795 5458 10813 5522
rect 10877 5458 10895 5522
rect 10959 5458 10977 5522
rect 11041 5458 11059 5522
rect 11123 5458 11141 5522
rect 11205 5458 11223 5522
rect 11287 5458 11305 5522
rect 11369 5458 11386 5522
rect 11450 5458 11467 5522
rect 11531 5458 11548 5522
rect 11612 5458 11629 5522
rect 11693 5458 11710 5522
rect 11774 5458 11791 5522
rect 11855 5458 11872 5522
rect 11936 5458 11953 5522
rect 12017 5458 12034 5522
rect 12098 5458 12115 5522
rect 12179 5458 12196 5522
rect 12260 5458 12277 5522
rect 12341 5458 12358 5522
rect 12422 5458 12439 5522
rect 12503 5458 12520 5522
rect 12584 5458 12601 5522
rect 12665 5458 12682 5522
rect 12746 5458 12763 5522
rect 12827 5458 12844 5522
rect 12908 5458 12925 5522
rect 12989 5458 13006 5522
rect 13070 5458 13087 5522
rect 13151 5458 13168 5522
rect 13232 5458 13249 5522
rect 13313 5458 13330 5522
rect 13394 5458 13411 5522
rect 13475 5458 13492 5522
rect 13556 5458 13573 5522
rect 13637 5458 13654 5522
rect 13718 5458 13735 5522
rect 13799 5458 13816 5522
rect 13880 5458 13897 5522
rect 13961 5458 13978 5522
rect 14042 5458 14059 5522
rect 14123 5458 14140 5522
rect 14204 5458 14221 5522
rect 14285 5458 14302 5522
rect 14366 5458 14383 5522
rect 14447 5458 14464 5522
rect 14528 5458 14545 5522
rect 14609 5458 14626 5522
rect 14690 5458 14707 5522
rect 14771 5458 14788 5522
rect 14852 5458 15000 5522
rect 0 5436 15000 5458
rect 0 5372 106 5436
rect 170 5372 188 5436
rect 252 5372 270 5436
rect 334 5372 352 5436
rect 416 5372 434 5436
rect 498 5372 516 5436
rect 580 5372 598 5436
rect 662 5372 679 5436
rect 743 5372 760 5436
rect 824 5372 841 5436
rect 905 5372 922 5436
rect 986 5372 1003 5436
rect 1067 5372 1084 5436
rect 1148 5372 1165 5436
rect 1229 5372 1246 5436
rect 1310 5372 1327 5436
rect 1391 5372 1408 5436
rect 1472 5372 1489 5436
rect 1553 5372 1570 5436
rect 1634 5372 1651 5436
rect 1715 5372 1732 5436
rect 1796 5372 1813 5436
rect 1877 5372 1894 5436
rect 1958 5372 1975 5436
rect 2039 5372 2056 5436
rect 2120 5372 2137 5436
rect 2201 5372 2218 5436
rect 2282 5372 2299 5436
rect 2363 5372 2380 5436
rect 2444 5372 2461 5436
rect 2525 5372 2542 5436
rect 2606 5372 2623 5436
rect 2687 5372 2704 5436
rect 2768 5372 2785 5436
rect 2849 5372 2866 5436
rect 2930 5372 2947 5436
rect 3011 5372 3028 5436
rect 3092 5372 3109 5436
rect 3173 5372 3190 5436
rect 3254 5372 3271 5436
rect 3335 5372 3352 5436
rect 3416 5372 3433 5436
rect 3497 5372 3514 5436
rect 3578 5372 3595 5436
rect 3659 5372 3676 5436
rect 3740 5372 3757 5436
rect 3821 5372 3838 5436
rect 3902 5372 3919 5436
rect 3983 5372 4000 5436
rect 4064 5372 4081 5436
rect 4145 5372 4162 5436
rect 4226 5372 4243 5436
rect 4307 5372 4324 5436
rect 4388 5372 4405 5436
rect 4469 5372 4486 5436
rect 4550 5372 4567 5436
rect 4631 5372 4648 5436
rect 4712 5372 4729 5436
rect 4793 5372 4810 5436
rect 4874 5372 10157 5436
rect 10221 5372 10239 5436
rect 10303 5372 10321 5436
rect 10385 5372 10403 5436
rect 10467 5372 10485 5436
rect 10549 5372 10567 5436
rect 10631 5372 10649 5436
rect 10713 5372 10731 5436
rect 10795 5372 10813 5436
rect 10877 5372 10895 5436
rect 10959 5372 10977 5436
rect 11041 5372 11059 5436
rect 11123 5372 11141 5436
rect 11205 5372 11223 5436
rect 11287 5372 11305 5436
rect 11369 5372 11386 5436
rect 11450 5372 11467 5436
rect 11531 5372 11548 5436
rect 11612 5372 11629 5436
rect 11693 5372 11710 5436
rect 11774 5372 11791 5436
rect 11855 5372 11872 5436
rect 11936 5372 11953 5436
rect 12017 5372 12034 5436
rect 12098 5372 12115 5436
rect 12179 5372 12196 5436
rect 12260 5372 12277 5436
rect 12341 5372 12358 5436
rect 12422 5372 12439 5436
rect 12503 5372 12520 5436
rect 12584 5372 12601 5436
rect 12665 5372 12682 5436
rect 12746 5372 12763 5436
rect 12827 5372 12844 5436
rect 12908 5372 12925 5436
rect 12989 5372 13006 5436
rect 13070 5372 13087 5436
rect 13151 5372 13168 5436
rect 13232 5372 13249 5436
rect 13313 5372 13330 5436
rect 13394 5372 13411 5436
rect 13475 5372 13492 5436
rect 13556 5372 13573 5436
rect 13637 5372 13654 5436
rect 13718 5372 13735 5436
rect 13799 5372 13816 5436
rect 13880 5372 13897 5436
rect 13961 5372 13978 5436
rect 14042 5372 14059 5436
rect 14123 5372 14140 5436
rect 14204 5372 14221 5436
rect 14285 5372 14302 5436
rect 14366 5372 14383 5436
rect 14447 5372 14464 5436
rect 14528 5372 14545 5436
rect 14609 5372 14626 5436
rect 14690 5372 14707 5436
rect 14771 5372 14788 5436
rect 14852 5372 15000 5436
rect 0 5350 15000 5372
rect 0 5286 106 5350
rect 170 5286 188 5350
rect 252 5286 270 5350
rect 334 5286 352 5350
rect 416 5286 434 5350
rect 498 5286 516 5350
rect 580 5286 598 5350
rect 662 5286 679 5350
rect 743 5286 760 5350
rect 824 5286 841 5350
rect 905 5286 922 5350
rect 986 5286 1003 5350
rect 1067 5286 1084 5350
rect 1148 5286 1165 5350
rect 1229 5286 1246 5350
rect 1310 5286 1327 5350
rect 1391 5286 1408 5350
rect 1472 5286 1489 5350
rect 1553 5286 1570 5350
rect 1634 5286 1651 5350
rect 1715 5286 1732 5350
rect 1796 5286 1813 5350
rect 1877 5286 1894 5350
rect 1958 5286 1975 5350
rect 2039 5286 2056 5350
rect 2120 5286 2137 5350
rect 2201 5286 2218 5350
rect 2282 5286 2299 5350
rect 2363 5286 2380 5350
rect 2444 5286 2461 5350
rect 2525 5286 2542 5350
rect 2606 5286 2623 5350
rect 2687 5286 2704 5350
rect 2768 5286 2785 5350
rect 2849 5286 2866 5350
rect 2930 5286 2947 5350
rect 3011 5286 3028 5350
rect 3092 5286 3109 5350
rect 3173 5286 3190 5350
rect 3254 5286 3271 5350
rect 3335 5286 3352 5350
rect 3416 5286 3433 5350
rect 3497 5286 3514 5350
rect 3578 5286 3595 5350
rect 3659 5286 3676 5350
rect 3740 5286 3757 5350
rect 3821 5286 3838 5350
rect 3902 5286 3919 5350
rect 3983 5286 4000 5350
rect 4064 5286 4081 5350
rect 4145 5286 4162 5350
rect 4226 5286 4243 5350
rect 4307 5286 4324 5350
rect 4388 5286 4405 5350
rect 4469 5286 4486 5350
rect 4550 5286 4567 5350
rect 4631 5286 4648 5350
rect 4712 5286 4729 5350
rect 4793 5286 4810 5350
rect 4874 5286 10157 5350
rect 10221 5286 10239 5350
rect 10303 5286 10321 5350
rect 10385 5286 10403 5350
rect 10467 5286 10485 5350
rect 10549 5286 10567 5350
rect 10631 5286 10649 5350
rect 10713 5286 10731 5350
rect 10795 5286 10813 5350
rect 10877 5286 10895 5350
rect 10959 5286 10977 5350
rect 11041 5286 11059 5350
rect 11123 5286 11141 5350
rect 11205 5286 11223 5350
rect 11287 5286 11305 5350
rect 11369 5286 11386 5350
rect 11450 5286 11467 5350
rect 11531 5286 11548 5350
rect 11612 5286 11629 5350
rect 11693 5286 11710 5350
rect 11774 5286 11791 5350
rect 11855 5286 11872 5350
rect 11936 5286 11953 5350
rect 12017 5286 12034 5350
rect 12098 5286 12115 5350
rect 12179 5286 12196 5350
rect 12260 5286 12277 5350
rect 12341 5286 12358 5350
rect 12422 5286 12439 5350
rect 12503 5286 12520 5350
rect 12584 5286 12601 5350
rect 12665 5286 12682 5350
rect 12746 5286 12763 5350
rect 12827 5286 12844 5350
rect 12908 5286 12925 5350
rect 12989 5286 13006 5350
rect 13070 5286 13087 5350
rect 13151 5286 13168 5350
rect 13232 5286 13249 5350
rect 13313 5286 13330 5350
rect 13394 5286 13411 5350
rect 13475 5286 13492 5350
rect 13556 5286 13573 5350
rect 13637 5286 13654 5350
rect 13718 5286 13735 5350
rect 13799 5286 13816 5350
rect 13880 5286 13897 5350
rect 13961 5286 13978 5350
rect 14042 5286 14059 5350
rect 14123 5286 14140 5350
rect 14204 5286 14221 5350
rect 14285 5286 14302 5350
rect 14366 5286 14383 5350
rect 14447 5286 14464 5350
rect 14528 5286 14545 5350
rect 14609 5286 14626 5350
rect 14690 5286 14707 5350
rect 14771 5286 14788 5350
rect 14852 5286 15000 5350
rect 0 5264 15000 5286
rect 0 5200 106 5264
rect 170 5200 188 5264
rect 252 5200 270 5264
rect 334 5200 352 5264
rect 416 5200 434 5264
rect 498 5200 516 5264
rect 580 5200 598 5264
rect 662 5200 679 5264
rect 743 5200 760 5264
rect 824 5200 841 5264
rect 905 5200 922 5264
rect 986 5200 1003 5264
rect 1067 5200 1084 5264
rect 1148 5200 1165 5264
rect 1229 5200 1246 5264
rect 1310 5200 1327 5264
rect 1391 5200 1408 5264
rect 1472 5200 1489 5264
rect 1553 5200 1570 5264
rect 1634 5200 1651 5264
rect 1715 5200 1732 5264
rect 1796 5200 1813 5264
rect 1877 5200 1894 5264
rect 1958 5200 1975 5264
rect 2039 5200 2056 5264
rect 2120 5200 2137 5264
rect 2201 5200 2218 5264
rect 2282 5200 2299 5264
rect 2363 5200 2380 5264
rect 2444 5200 2461 5264
rect 2525 5200 2542 5264
rect 2606 5200 2623 5264
rect 2687 5200 2704 5264
rect 2768 5200 2785 5264
rect 2849 5200 2866 5264
rect 2930 5200 2947 5264
rect 3011 5200 3028 5264
rect 3092 5200 3109 5264
rect 3173 5200 3190 5264
rect 3254 5200 3271 5264
rect 3335 5200 3352 5264
rect 3416 5200 3433 5264
rect 3497 5200 3514 5264
rect 3578 5200 3595 5264
rect 3659 5200 3676 5264
rect 3740 5200 3757 5264
rect 3821 5200 3838 5264
rect 3902 5200 3919 5264
rect 3983 5200 4000 5264
rect 4064 5200 4081 5264
rect 4145 5200 4162 5264
rect 4226 5200 4243 5264
rect 4307 5200 4324 5264
rect 4388 5200 4405 5264
rect 4469 5200 4486 5264
rect 4550 5200 4567 5264
rect 4631 5200 4648 5264
rect 4712 5200 4729 5264
rect 4793 5200 4810 5264
rect 4874 5200 10157 5264
rect 10221 5200 10239 5264
rect 10303 5200 10321 5264
rect 10385 5200 10403 5264
rect 10467 5200 10485 5264
rect 10549 5200 10567 5264
rect 10631 5200 10649 5264
rect 10713 5200 10731 5264
rect 10795 5200 10813 5264
rect 10877 5200 10895 5264
rect 10959 5200 10977 5264
rect 11041 5200 11059 5264
rect 11123 5200 11141 5264
rect 11205 5200 11223 5264
rect 11287 5200 11305 5264
rect 11369 5200 11386 5264
rect 11450 5200 11467 5264
rect 11531 5200 11548 5264
rect 11612 5200 11629 5264
rect 11693 5200 11710 5264
rect 11774 5200 11791 5264
rect 11855 5200 11872 5264
rect 11936 5200 11953 5264
rect 12017 5200 12034 5264
rect 12098 5200 12115 5264
rect 12179 5200 12196 5264
rect 12260 5200 12277 5264
rect 12341 5200 12358 5264
rect 12422 5200 12439 5264
rect 12503 5200 12520 5264
rect 12584 5200 12601 5264
rect 12665 5200 12682 5264
rect 12746 5200 12763 5264
rect 12827 5200 12844 5264
rect 12908 5200 12925 5264
rect 12989 5200 13006 5264
rect 13070 5200 13087 5264
rect 13151 5200 13168 5264
rect 13232 5200 13249 5264
rect 13313 5200 13330 5264
rect 13394 5200 13411 5264
rect 13475 5200 13492 5264
rect 13556 5200 13573 5264
rect 13637 5200 13654 5264
rect 13718 5200 13735 5264
rect 13799 5200 13816 5264
rect 13880 5200 13897 5264
rect 13961 5200 13978 5264
rect 14042 5200 14059 5264
rect 14123 5200 14140 5264
rect 14204 5200 14221 5264
rect 14285 5200 14302 5264
rect 14366 5200 14383 5264
rect 14447 5200 14464 5264
rect 14528 5200 14545 5264
rect 14609 5200 14626 5264
rect 14690 5200 14707 5264
rect 14771 5200 14788 5264
rect 14852 5200 15000 5264
rect 0 5178 15000 5200
rect 0 5114 106 5178
rect 170 5114 188 5178
rect 252 5114 270 5178
rect 334 5114 352 5178
rect 416 5114 434 5178
rect 498 5114 516 5178
rect 580 5114 598 5178
rect 662 5114 679 5178
rect 743 5114 760 5178
rect 824 5114 841 5178
rect 905 5114 922 5178
rect 986 5114 1003 5178
rect 1067 5114 1084 5178
rect 1148 5114 1165 5178
rect 1229 5114 1246 5178
rect 1310 5114 1327 5178
rect 1391 5114 1408 5178
rect 1472 5114 1489 5178
rect 1553 5114 1570 5178
rect 1634 5114 1651 5178
rect 1715 5114 1732 5178
rect 1796 5114 1813 5178
rect 1877 5114 1894 5178
rect 1958 5114 1975 5178
rect 2039 5114 2056 5178
rect 2120 5114 2137 5178
rect 2201 5114 2218 5178
rect 2282 5114 2299 5178
rect 2363 5114 2380 5178
rect 2444 5114 2461 5178
rect 2525 5114 2542 5178
rect 2606 5114 2623 5178
rect 2687 5114 2704 5178
rect 2768 5114 2785 5178
rect 2849 5114 2866 5178
rect 2930 5114 2947 5178
rect 3011 5114 3028 5178
rect 3092 5114 3109 5178
rect 3173 5114 3190 5178
rect 3254 5114 3271 5178
rect 3335 5114 3352 5178
rect 3416 5114 3433 5178
rect 3497 5114 3514 5178
rect 3578 5114 3595 5178
rect 3659 5114 3676 5178
rect 3740 5114 3757 5178
rect 3821 5114 3838 5178
rect 3902 5114 3919 5178
rect 3983 5114 4000 5178
rect 4064 5114 4081 5178
rect 4145 5114 4162 5178
rect 4226 5114 4243 5178
rect 4307 5114 4324 5178
rect 4388 5114 4405 5178
rect 4469 5114 4486 5178
rect 4550 5114 4567 5178
rect 4631 5114 4648 5178
rect 4712 5114 4729 5178
rect 4793 5114 4810 5178
rect 4874 5114 10157 5178
rect 10221 5114 10239 5178
rect 10303 5114 10321 5178
rect 10385 5114 10403 5178
rect 10467 5114 10485 5178
rect 10549 5114 10567 5178
rect 10631 5114 10649 5178
rect 10713 5114 10731 5178
rect 10795 5114 10813 5178
rect 10877 5114 10895 5178
rect 10959 5114 10977 5178
rect 11041 5114 11059 5178
rect 11123 5114 11141 5178
rect 11205 5114 11223 5178
rect 11287 5114 11305 5178
rect 11369 5114 11386 5178
rect 11450 5114 11467 5178
rect 11531 5114 11548 5178
rect 11612 5114 11629 5178
rect 11693 5114 11710 5178
rect 11774 5114 11791 5178
rect 11855 5114 11872 5178
rect 11936 5114 11953 5178
rect 12017 5114 12034 5178
rect 12098 5114 12115 5178
rect 12179 5114 12196 5178
rect 12260 5114 12277 5178
rect 12341 5114 12358 5178
rect 12422 5114 12439 5178
rect 12503 5114 12520 5178
rect 12584 5114 12601 5178
rect 12665 5114 12682 5178
rect 12746 5114 12763 5178
rect 12827 5114 12844 5178
rect 12908 5114 12925 5178
rect 12989 5114 13006 5178
rect 13070 5114 13087 5178
rect 13151 5114 13168 5178
rect 13232 5114 13249 5178
rect 13313 5114 13330 5178
rect 13394 5114 13411 5178
rect 13475 5114 13492 5178
rect 13556 5114 13573 5178
rect 13637 5114 13654 5178
rect 13718 5114 13735 5178
rect 13799 5114 13816 5178
rect 13880 5114 13897 5178
rect 13961 5114 13978 5178
rect 14042 5114 14059 5178
rect 14123 5114 14140 5178
rect 14204 5114 14221 5178
rect 14285 5114 14302 5178
rect 14366 5114 14383 5178
rect 14447 5114 14464 5178
rect 14528 5114 14545 5178
rect 14609 5114 14626 5178
rect 14690 5114 14707 5178
rect 14771 5114 14788 5178
rect 14852 5114 15000 5178
rect 0 5092 15000 5114
rect 0 5028 106 5092
rect 170 5028 188 5092
rect 252 5028 270 5092
rect 334 5028 352 5092
rect 416 5028 434 5092
rect 498 5028 516 5092
rect 580 5028 598 5092
rect 662 5028 679 5092
rect 743 5028 760 5092
rect 824 5028 841 5092
rect 905 5028 922 5092
rect 986 5028 1003 5092
rect 1067 5028 1084 5092
rect 1148 5028 1165 5092
rect 1229 5028 1246 5092
rect 1310 5028 1327 5092
rect 1391 5028 1408 5092
rect 1472 5028 1489 5092
rect 1553 5028 1570 5092
rect 1634 5028 1651 5092
rect 1715 5028 1732 5092
rect 1796 5028 1813 5092
rect 1877 5028 1894 5092
rect 1958 5028 1975 5092
rect 2039 5028 2056 5092
rect 2120 5028 2137 5092
rect 2201 5028 2218 5092
rect 2282 5028 2299 5092
rect 2363 5028 2380 5092
rect 2444 5028 2461 5092
rect 2525 5028 2542 5092
rect 2606 5028 2623 5092
rect 2687 5028 2704 5092
rect 2768 5028 2785 5092
rect 2849 5028 2866 5092
rect 2930 5028 2947 5092
rect 3011 5028 3028 5092
rect 3092 5028 3109 5092
rect 3173 5028 3190 5092
rect 3254 5028 3271 5092
rect 3335 5028 3352 5092
rect 3416 5028 3433 5092
rect 3497 5028 3514 5092
rect 3578 5028 3595 5092
rect 3659 5028 3676 5092
rect 3740 5028 3757 5092
rect 3821 5028 3838 5092
rect 3902 5028 3919 5092
rect 3983 5028 4000 5092
rect 4064 5028 4081 5092
rect 4145 5028 4162 5092
rect 4226 5028 4243 5092
rect 4307 5028 4324 5092
rect 4388 5028 4405 5092
rect 4469 5028 4486 5092
rect 4550 5028 4567 5092
rect 4631 5028 4648 5092
rect 4712 5028 4729 5092
rect 4793 5028 4810 5092
rect 4874 5028 10157 5092
rect 10221 5028 10239 5092
rect 10303 5028 10321 5092
rect 10385 5028 10403 5092
rect 10467 5028 10485 5092
rect 10549 5028 10567 5092
rect 10631 5028 10649 5092
rect 10713 5028 10731 5092
rect 10795 5028 10813 5092
rect 10877 5028 10895 5092
rect 10959 5028 10977 5092
rect 11041 5028 11059 5092
rect 11123 5028 11141 5092
rect 11205 5028 11223 5092
rect 11287 5028 11305 5092
rect 11369 5028 11386 5092
rect 11450 5028 11467 5092
rect 11531 5028 11548 5092
rect 11612 5028 11629 5092
rect 11693 5028 11710 5092
rect 11774 5028 11791 5092
rect 11855 5028 11872 5092
rect 11936 5028 11953 5092
rect 12017 5028 12034 5092
rect 12098 5028 12115 5092
rect 12179 5028 12196 5092
rect 12260 5028 12277 5092
rect 12341 5028 12358 5092
rect 12422 5028 12439 5092
rect 12503 5028 12520 5092
rect 12584 5028 12601 5092
rect 12665 5028 12682 5092
rect 12746 5028 12763 5092
rect 12827 5028 12844 5092
rect 12908 5028 12925 5092
rect 12989 5028 13006 5092
rect 13070 5028 13087 5092
rect 13151 5028 13168 5092
rect 13232 5028 13249 5092
rect 13313 5028 13330 5092
rect 13394 5028 13411 5092
rect 13475 5028 13492 5092
rect 13556 5028 13573 5092
rect 13637 5028 13654 5092
rect 13718 5028 13735 5092
rect 13799 5028 13816 5092
rect 13880 5028 13897 5092
rect 13961 5028 13978 5092
rect 14042 5028 14059 5092
rect 14123 5028 14140 5092
rect 14204 5028 14221 5092
rect 14285 5028 14302 5092
rect 14366 5028 14383 5092
rect 14447 5028 14464 5092
rect 14528 5028 14545 5092
rect 14609 5028 14626 5092
rect 14690 5028 14707 5092
rect 14771 5028 14788 5092
rect 14852 5028 15000 5092
rect 0 5006 15000 5028
rect 0 4942 106 5006
rect 170 4942 188 5006
rect 252 4942 270 5006
rect 334 4942 352 5006
rect 416 4942 434 5006
rect 498 4942 516 5006
rect 580 4942 598 5006
rect 662 4942 679 5006
rect 743 4942 760 5006
rect 824 4942 841 5006
rect 905 4942 922 5006
rect 986 4942 1003 5006
rect 1067 4942 1084 5006
rect 1148 4942 1165 5006
rect 1229 4942 1246 5006
rect 1310 4942 1327 5006
rect 1391 4942 1408 5006
rect 1472 4942 1489 5006
rect 1553 4942 1570 5006
rect 1634 4942 1651 5006
rect 1715 4942 1732 5006
rect 1796 4942 1813 5006
rect 1877 4942 1894 5006
rect 1958 4942 1975 5006
rect 2039 4942 2056 5006
rect 2120 4942 2137 5006
rect 2201 4942 2218 5006
rect 2282 4942 2299 5006
rect 2363 4942 2380 5006
rect 2444 4942 2461 5006
rect 2525 4942 2542 5006
rect 2606 4942 2623 5006
rect 2687 4942 2704 5006
rect 2768 4942 2785 5006
rect 2849 4942 2866 5006
rect 2930 4942 2947 5006
rect 3011 4942 3028 5006
rect 3092 4942 3109 5006
rect 3173 4942 3190 5006
rect 3254 4942 3271 5006
rect 3335 4942 3352 5006
rect 3416 4942 3433 5006
rect 3497 4942 3514 5006
rect 3578 4942 3595 5006
rect 3659 4942 3676 5006
rect 3740 4942 3757 5006
rect 3821 4942 3838 5006
rect 3902 4942 3919 5006
rect 3983 4942 4000 5006
rect 4064 4942 4081 5006
rect 4145 4942 4162 5006
rect 4226 4942 4243 5006
rect 4307 4942 4324 5006
rect 4388 4942 4405 5006
rect 4469 4942 4486 5006
rect 4550 4942 4567 5006
rect 4631 4942 4648 5006
rect 4712 4942 4729 5006
rect 4793 4942 4810 5006
rect 4874 4942 10157 5006
rect 10221 4942 10239 5006
rect 10303 4942 10321 5006
rect 10385 4942 10403 5006
rect 10467 4942 10485 5006
rect 10549 4942 10567 5006
rect 10631 4942 10649 5006
rect 10713 4942 10731 5006
rect 10795 4942 10813 5006
rect 10877 4942 10895 5006
rect 10959 4942 10977 5006
rect 11041 4942 11059 5006
rect 11123 4942 11141 5006
rect 11205 4942 11223 5006
rect 11287 4942 11305 5006
rect 11369 4942 11386 5006
rect 11450 4942 11467 5006
rect 11531 4942 11548 5006
rect 11612 4942 11629 5006
rect 11693 4942 11710 5006
rect 11774 4942 11791 5006
rect 11855 4942 11872 5006
rect 11936 4942 11953 5006
rect 12017 4942 12034 5006
rect 12098 4942 12115 5006
rect 12179 4942 12196 5006
rect 12260 4942 12277 5006
rect 12341 4942 12358 5006
rect 12422 4942 12439 5006
rect 12503 4942 12520 5006
rect 12584 4942 12601 5006
rect 12665 4942 12682 5006
rect 12746 4942 12763 5006
rect 12827 4942 12844 5006
rect 12908 4942 12925 5006
rect 12989 4942 13006 5006
rect 13070 4942 13087 5006
rect 13151 4942 13168 5006
rect 13232 4942 13249 5006
rect 13313 4942 13330 5006
rect 13394 4942 13411 5006
rect 13475 4942 13492 5006
rect 13556 4942 13573 5006
rect 13637 4942 13654 5006
rect 13718 4942 13735 5006
rect 13799 4942 13816 5006
rect 13880 4942 13897 5006
rect 13961 4942 13978 5006
rect 14042 4942 14059 5006
rect 14123 4942 14140 5006
rect 14204 4942 14221 5006
rect 14285 4942 14302 5006
rect 14366 4942 14383 5006
rect 14447 4942 14464 5006
rect 14528 4942 14545 5006
rect 14609 4942 14626 5006
rect 14690 4942 14707 5006
rect 14771 4942 14788 5006
rect 14852 4942 15000 5006
rect 0 4920 15000 4942
rect 0 4856 106 4920
rect 170 4856 188 4920
rect 252 4856 270 4920
rect 334 4856 352 4920
rect 416 4856 434 4920
rect 498 4856 516 4920
rect 580 4856 598 4920
rect 662 4856 679 4920
rect 743 4856 760 4920
rect 824 4856 841 4920
rect 905 4856 922 4920
rect 986 4856 1003 4920
rect 1067 4856 1084 4920
rect 1148 4856 1165 4920
rect 1229 4856 1246 4920
rect 1310 4856 1327 4920
rect 1391 4856 1408 4920
rect 1472 4856 1489 4920
rect 1553 4856 1570 4920
rect 1634 4856 1651 4920
rect 1715 4856 1732 4920
rect 1796 4856 1813 4920
rect 1877 4856 1894 4920
rect 1958 4856 1975 4920
rect 2039 4856 2056 4920
rect 2120 4856 2137 4920
rect 2201 4856 2218 4920
rect 2282 4856 2299 4920
rect 2363 4856 2380 4920
rect 2444 4856 2461 4920
rect 2525 4856 2542 4920
rect 2606 4856 2623 4920
rect 2687 4856 2704 4920
rect 2768 4856 2785 4920
rect 2849 4856 2866 4920
rect 2930 4856 2947 4920
rect 3011 4856 3028 4920
rect 3092 4856 3109 4920
rect 3173 4856 3190 4920
rect 3254 4856 3271 4920
rect 3335 4856 3352 4920
rect 3416 4856 3433 4920
rect 3497 4856 3514 4920
rect 3578 4856 3595 4920
rect 3659 4856 3676 4920
rect 3740 4856 3757 4920
rect 3821 4856 3838 4920
rect 3902 4856 3919 4920
rect 3983 4856 4000 4920
rect 4064 4856 4081 4920
rect 4145 4856 4162 4920
rect 4226 4856 4243 4920
rect 4307 4856 4324 4920
rect 4388 4856 4405 4920
rect 4469 4856 4486 4920
rect 4550 4856 4567 4920
rect 4631 4856 4648 4920
rect 4712 4856 4729 4920
rect 4793 4856 4810 4920
rect 4874 4856 10157 4920
rect 10221 4856 10239 4920
rect 10303 4856 10321 4920
rect 10385 4856 10403 4920
rect 10467 4856 10485 4920
rect 10549 4856 10567 4920
rect 10631 4856 10649 4920
rect 10713 4856 10731 4920
rect 10795 4856 10813 4920
rect 10877 4856 10895 4920
rect 10959 4856 10977 4920
rect 11041 4856 11059 4920
rect 11123 4856 11141 4920
rect 11205 4856 11223 4920
rect 11287 4856 11305 4920
rect 11369 4856 11386 4920
rect 11450 4856 11467 4920
rect 11531 4856 11548 4920
rect 11612 4856 11629 4920
rect 11693 4856 11710 4920
rect 11774 4856 11791 4920
rect 11855 4856 11872 4920
rect 11936 4856 11953 4920
rect 12017 4856 12034 4920
rect 12098 4856 12115 4920
rect 12179 4856 12196 4920
rect 12260 4856 12277 4920
rect 12341 4856 12358 4920
rect 12422 4856 12439 4920
rect 12503 4856 12520 4920
rect 12584 4856 12601 4920
rect 12665 4856 12682 4920
rect 12746 4856 12763 4920
rect 12827 4856 12844 4920
rect 12908 4856 12925 4920
rect 12989 4856 13006 4920
rect 13070 4856 13087 4920
rect 13151 4856 13168 4920
rect 13232 4856 13249 4920
rect 13313 4856 13330 4920
rect 13394 4856 13411 4920
rect 13475 4856 13492 4920
rect 13556 4856 13573 4920
rect 13637 4856 13654 4920
rect 13718 4856 13735 4920
rect 13799 4856 13816 4920
rect 13880 4856 13897 4920
rect 13961 4856 13978 4920
rect 14042 4856 14059 4920
rect 14123 4856 14140 4920
rect 14204 4856 14221 4920
rect 14285 4856 14302 4920
rect 14366 4856 14383 4920
rect 14447 4856 14464 4920
rect 14528 4856 14545 4920
rect 14609 4856 14626 4920
rect 14690 4856 14707 4920
rect 14771 4856 14788 4920
rect 14852 4856 15000 4920
rect 0 4834 15000 4856
rect 0 4770 106 4834
rect 170 4770 188 4834
rect 252 4770 270 4834
rect 334 4770 352 4834
rect 416 4770 434 4834
rect 498 4770 516 4834
rect 580 4770 598 4834
rect 662 4770 679 4834
rect 743 4770 760 4834
rect 824 4770 841 4834
rect 905 4770 922 4834
rect 986 4770 1003 4834
rect 1067 4770 1084 4834
rect 1148 4770 1165 4834
rect 1229 4770 1246 4834
rect 1310 4770 1327 4834
rect 1391 4770 1408 4834
rect 1472 4770 1489 4834
rect 1553 4770 1570 4834
rect 1634 4770 1651 4834
rect 1715 4770 1732 4834
rect 1796 4770 1813 4834
rect 1877 4770 1894 4834
rect 1958 4770 1975 4834
rect 2039 4770 2056 4834
rect 2120 4770 2137 4834
rect 2201 4770 2218 4834
rect 2282 4770 2299 4834
rect 2363 4770 2380 4834
rect 2444 4770 2461 4834
rect 2525 4770 2542 4834
rect 2606 4770 2623 4834
rect 2687 4770 2704 4834
rect 2768 4770 2785 4834
rect 2849 4770 2866 4834
rect 2930 4770 2947 4834
rect 3011 4770 3028 4834
rect 3092 4770 3109 4834
rect 3173 4770 3190 4834
rect 3254 4770 3271 4834
rect 3335 4770 3352 4834
rect 3416 4770 3433 4834
rect 3497 4770 3514 4834
rect 3578 4770 3595 4834
rect 3659 4770 3676 4834
rect 3740 4770 3757 4834
rect 3821 4770 3838 4834
rect 3902 4770 3919 4834
rect 3983 4770 4000 4834
rect 4064 4770 4081 4834
rect 4145 4770 4162 4834
rect 4226 4770 4243 4834
rect 4307 4770 4324 4834
rect 4388 4770 4405 4834
rect 4469 4770 4486 4834
rect 4550 4770 4567 4834
rect 4631 4770 4648 4834
rect 4712 4770 4729 4834
rect 4793 4770 4810 4834
rect 4874 4770 10157 4834
rect 10221 4770 10239 4834
rect 10303 4770 10321 4834
rect 10385 4770 10403 4834
rect 10467 4770 10485 4834
rect 10549 4770 10567 4834
rect 10631 4770 10649 4834
rect 10713 4770 10731 4834
rect 10795 4770 10813 4834
rect 10877 4770 10895 4834
rect 10959 4770 10977 4834
rect 11041 4770 11059 4834
rect 11123 4770 11141 4834
rect 11205 4770 11223 4834
rect 11287 4770 11305 4834
rect 11369 4770 11386 4834
rect 11450 4770 11467 4834
rect 11531 4770 11548 4834
rect 11612 4770 11629 4834
rect 11693 4770 11710 4834
rect 11774 4770 11791 4834
rect 11855 4770 11872 4834
rect 11936 4770 11953 4834
rect 12017 4770 12034 4834
rect 12098 4770 12115 4834
rect 12179 4770 12196 4834
rect 12260 4770 12277 4834
rect 12341 4770 12358 4834
rect 12422 4770 12439 4834
rect 12503 4770 12520 4834
rect 12584 4770 12601 4834
rect 12665 4770 12682 4834
rect 12746 4770 12763 4834
rect 12827 4770 12844 4834
rect 12908 4770 12925 4834
rect 12989 4770 13006 4834
rect 13070 4770 13087 4834
rect 13151 4770 13168 4834
rect 13232 4770 13249 4834
rect 13313 4770 13330 4834
rect 13394 4770 13411 4834
rect 13475 4770 13492 4834
rect 13556 4770 13573 4834
rect 13637 4770 13654 4834
rect 13718 4770 13735 4834
rect 13799 4770 13816 4834
rect 13880 4770 13897 4834
rect 13961 4770 13978 4834
rect 14042 4770 14059 4834
rect 14123 4770 14140 4834
rect 14204 4770 14221 4834
rect 14285 4770 14302 4834
rect 14366 4770 14383 4834
rect 14447 4770 14464 4834
rect 14528 4770 14545 4834
rect 14609 4770 14626 4834
rect 14690 4770 14707 4834
rect 14771 4770 14788 4834
rect 14852 4770 15000 4834
rect 0 7 15000 4770
<< metal5 >>
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 5997 15000 6647
rect 14807 2607 15000 3257
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 0 18917 15000 39600
rect 0 12117 14426 18917
rect 0 11267 15000 12117
rect 0 7617 14426 11267
rect 0 6967 15000 7617
rect 0 5677 14426 6967
rect 0 3577 15000 5677
rect 0 2607 14487 3577
rect 0 27 14426 2607
<< labels >>
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 3 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 4770 170 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 4770 170 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 4856 170 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 4856 170 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 4942 170 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 4942 170 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 5028 170 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 5028 170 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 5114 170 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 5114 170 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 5200 170 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 5200 170 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 5286 170 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 5286 170 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 5372 170 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 5372 170 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 5458 170 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 5458 170 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 5544 170 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 5544 170 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 5630 170 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 106 5630 170 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 34768 2575 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 34768 2575 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36289 175 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36289 175 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36370 175 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36370 175 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36451 175 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36451 175 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36532 175 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36532 175 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36613 175 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36613 175 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36694 175 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36694 175 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36775 175 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36775 175 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36856 175 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36856 175 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 36937 175 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 36937 175 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37018 175 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37018 175 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37099 175 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37099 175 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37180 175 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37180 175 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37261 175 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37261 175 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37342 175 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37342 175 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37423 175 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37423 175 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37504 175 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37504 175 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37585 175 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37585 175 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37666 175 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37666 175 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37747 175 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37747 175 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37828 175 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37828 175 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37909 175 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37909 175 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 37990 175 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 37990 175 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38071 175 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38071 175 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38152 175 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38152 175 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38233 175 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38233 175 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38314 175 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38314 175 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38395 175 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38395 175 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38476 175 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38476 175 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38557 175 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38557 175 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38638 175 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38638 175 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38719 175 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38719 175 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38800 175 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38800 175 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38881 175 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38881 175 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 38962 175 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 38962 175 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 39043 175 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 39043 175 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 39124 175 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 39124 175 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 39205 175 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 39205 175 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 39286 175 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 39286 175 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 39367 175 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 39367 175 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 39448 175 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 39448 175 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 111 39529 175 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 111 39529 175 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 34780 163 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 34860 163 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 34940 163 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35020 163 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35100 163 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35180 163 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35260 163 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35340 163 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35420 163 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35500 163 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35580 163 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35660 163 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35740 163 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35820 163 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35900 163 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 35980 163 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 36060 163 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 36140 163 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 123 36220 163 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 4770 252 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 4770 252 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 4856 252 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 4856 252 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 4942 252 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 4942 252 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 5028 252 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 5028 252 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 5114 252 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 5114 252 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 5200 252 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 5200 252 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 5286 252 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 5286 252 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 5372 252 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 5372 252 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 5458 252 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 5458 252 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 5544 252 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 5544 252 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 188 5630 252 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 188 5630 252 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36289 255 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36289 255 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36370 255 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36370 255 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36451 255 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36451 255 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36532 255 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36532 255 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36613 255 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36613 255 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36694 255 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36694 255 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36775 255 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36775 255 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36856 255 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36856 255 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 36937 255 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 36937 255 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37018 255 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37018 255 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37099 255 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37099 255 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37180 255 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37180 255 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37261 255 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37261 255 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37342 255 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37342 255 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37423 255 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37423 255 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37504 255 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37504 255 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37585 255 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37585 255 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37666 255 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37666 255 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37747 255 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37747 255 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37828 255 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37828 255 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37909 255 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37909 255 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 37990 255 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 37990 255 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38071 255 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38071 255 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38152 255 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38152 255 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38233 255 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38233 255 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38314 255 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38314 255 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38395 255 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38395 255 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38476 255 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38476 255 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38557 255 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38557 255 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38638 255 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38638 255 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38719 255 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38719 255 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38800 255 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38800 255 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38881 255 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38881 255 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 38962 255 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 38962 255 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 39043 255 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 39043 255 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 39124 255 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 39124 255 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 39205 255 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 39205 255 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 39286 255 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 39286 255 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 39367 255 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 39367 255 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 39448 255 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 39448 255 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 191 39529 255 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 191 39529 255 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 34780 243 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 34860 243 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 34940 243 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35020 243 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35100 243 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35180 243 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35260 243 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35340 243 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35420 243 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35500 243 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35580 243 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35660 243 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35740 243 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35820 243 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35900 243 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 35980 243 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 36060 243 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 36140 243 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 203 36220 243 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 4770 334 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 4770 334 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 4856 334 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 4856 334 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 4942 334 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 4942 334 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 5028 334 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 5028 334 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 5114 334 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 5114 334 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 5200 334 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 5200 334 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 5286 334 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 5286 334 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 5372 334 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 5372 334 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 5458 334 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 5458 334 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 5544 334 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 5544 334 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 270 5630 334 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 270 5630 334 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36289 335 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36289 335 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36370 335 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36370 335 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36451 335 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36451 335 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36532 335 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36532 335 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36613 335 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36613 335 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36694 335 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36694 335 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36775 335 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36775 335 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36856 335 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36856 335 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 36937 335 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 36937 335 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37018 335 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37018 335 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37099 335 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37099 335 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37180 335 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37180 335 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37261 335 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37261 335 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37342 335 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37342 335 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37423 335 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37423 335 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37504 335 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37504 335 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37585 335 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37585 335 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37666 335 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37666 335 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37747 335 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37747 335 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37828 335 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37828 335 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37909 335 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37909 335 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 37990 335 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 37990 335 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38071 335 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38071 335 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38152 335 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38152 335 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38233 335 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38233 335 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38314 335 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38314 335 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38395 335 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38395 335 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38476 335 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38476 335 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38557 335 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38557 335 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38638 335 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38638 335 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38719 335 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38719 335 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38800 335 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38800 335 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38881 335 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38881 335 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 38962 335 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 38962 335 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 39043 335 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 39043 335 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 39124 335 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 39124 335 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 39205 335 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 39205 335 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 39286 335 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 39286 335 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 39367 335 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 39367 335 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 39448 335 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 39448 335 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 271 39529 335 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 271 39529 335 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 34780 323 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 34860 323 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 34940 323 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35020 323 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35100 323 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35180 323 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35260 323 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35340 323 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35420 323 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35500 323 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35580 323 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35660 323 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35740 323 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35820 323 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35900 323 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 35980 323 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 36060 323 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 36140 323 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 283 36220 323 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36289 415 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36289 415 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36370 415 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36370 415 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36451 415 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36451 415 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36532 415 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36532 415 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36613 415 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36613 415 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36694 415 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36694 415 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36775 415 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36775 415 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36856 415 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36856 415 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 36937 415 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 36937 415 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37018 415 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37018 415 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37099 415 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37099 415 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37180 415 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37180 415 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37261 415 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37261 415 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37342 415 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37342 415 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37423 415 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37423 415 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37504 415 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37504 415 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37585 415 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37585 415 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37666 415 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37666 415 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37747 415 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37747 415 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37828 415 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37828 415 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37909 415 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37909 415 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 37990 415 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 37990 415 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38071 415 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38071 415 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38152 415 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38152 415 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38233 415 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38233 415 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38314 415 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38314 415 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38395 415 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38395 415 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38476 415 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38476 415 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38557 415 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38557 415 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38638 415 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38638 415 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38719 415 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38719 415 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38800 415 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38800 415 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38881 415 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38881 415 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 38962 415 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 38962 415 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 39043 415 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 39043 415 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 39124 415 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 39124 415 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 39205 415 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 39205 415 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 39286 415 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 39286 415 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 39367 415 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 39367 415 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 39448 415 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 39448 415 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 351 39529 415 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 351 39529 415 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 4770 416 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 4770 416 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 4856 416 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 4856 416 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 4942 416 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 4942 416 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 5028 416 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 5028 416 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 5114 416 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 5114 416 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 5200 416 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 5200 416 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 5286 416 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 5286 416 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 5372 416 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 5372 416 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 5458 416 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 5458 416 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 5544 416 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 5544 416 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 352 5630 416 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 352 5630 416 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 34780 403 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 34860 403 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 34940 403 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35020 403 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35100 403 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35180 403 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35260 403 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35340 403 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35420 403 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35500 403 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35580 403 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35660 403 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35740 403 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35820 403 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35900 403 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 35980 403 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 36060 403 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 36140 403 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 363 36220 403 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36289 2095 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36289 2095 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36370 2095 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36370 2095 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36451 2095 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36451 2095 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36532 2095 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36532 2095 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36613 2095 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36613 2095 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36694 2095 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36694 2095 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36775 2095 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36775 2095 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36856 2095 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36856 2095 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 36937 2095 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 36937 2095 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37018 2095 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37018 2095 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37099 2095 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37099 2095 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37180 2095 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37180 2095 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37261 2095 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37261 2095 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37342 2095 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37342 2095 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37423 2095 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37423 2095 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37504 2095 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37504 2095 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37585 2095 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37585 2095 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37666 2095 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37666 2095 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37747 2095 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37747 2095 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37828 2095 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37828 2095 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37909 2095 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37909 2095 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 37990 2095 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 37990 2095 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38071 2095 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38071 2095 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38152 2095 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38152 2095 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38233 2095 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38233 2095 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38314 2095 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38314 2095 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38395 2095 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38395 2095 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38476 2095 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38476 2095 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38557 2095 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38557 2095 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38638 2095 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38638 2095 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38719 2095 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38719 2095 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38800 2095 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38800 2095 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38881 2095 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38881 2095 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 38962 2095 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 38962 2095 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 39043 2095 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 39043 2095 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 39124 2095 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 39124 2095 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 39205 2095 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 39205 2095 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 39286 2095 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 39286 2095 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 39367 2095 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 39367 2095 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 39448 2095 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 39448 2095 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2031 39529 2095 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2031 39529 2095 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 34780 2083 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 34860 2083 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 34940 2083 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35020 2083 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35100 2083 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35180 2083 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35260 2083 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35340 2083 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35420 2083 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35500 2083 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35580 2083 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35660 2083 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35740 2083 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35820 2083 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35900 2083 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 35980 2083 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 36060 2083 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 36140 2083 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2043 36220 2083 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 4770 2120 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 4770 2120 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 4856 2120 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 4856 2120 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 4942 2120 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 4942 2120 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 5028 2120 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 5028 2120 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 5114 2120 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 5114 2120 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 5200 2120 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 5200 2120 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 5286 2120 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 5286 2120 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 5372 2120 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 5372 2120 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 5458 2120 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 5458 2120 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 5544 2120 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 5544 2120 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2056 5630 2120 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2056 5630 2120 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36289 2175 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36289 2175 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36370 2175 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36370 2175 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36451 2175 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36451 2175 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36532 2175 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36532 2175 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36613 2175 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36613 2175 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36694 2175 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36694 2175 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36775 2175 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36775 2175 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36856 2175 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36856 2175 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 36937 2175 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 36937 2175 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37018 2175 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37018 2175 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37099 2175 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37099 2175 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37180 2175 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37180 2175 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37261 2175 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37261 2175 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37342 2175 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37342 2175 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37423 2175 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37423 2175 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37504 2175 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37504 2175 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37585 2175 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37585 2175 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37666 2175 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37666 2175 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37747 2175 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37747 2175 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37828 2175 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37828 2175 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37909 2175 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37909 2175 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 37990 2175 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 37990 2175 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38071 2175 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38071 2175 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38152 2175 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38152 2175 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38233 2175 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38233 2175 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38314 2175 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38314 2175 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38395 2175 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38395 2175 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38476 2175 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38476 2175 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38557 2175 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38557 2175 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38638 2175 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38638 2175 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38719 2175 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38719 2175 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38800 2175 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38800 2175 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38881 2175 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38881 2175 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 38962 2175 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 38962 2175 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 39043 2175 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 39043 2175 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 39124 2175 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 39124 2175 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 39205 2175 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 39205 2175 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 39286 2175 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 39286 2175 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 39367 2175 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 39367 2175 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 39448 2175 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 39448 2175 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2111 39529 2175 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2111 39529 2175 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 34780 2163 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 34860 2163 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 34940 2163 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35020 2163 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35100 2163 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35180 2163 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35260 2163 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35340 2163 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35420 2163 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35500 2163 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35580 2163 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35660 2163 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35740 2163 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35820 2163 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35900 2163 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 35980 2163 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 36060 2163 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 36140 2163 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2123 36220 2163 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 4770 2201 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 4770 2201 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 4856 2201 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 4856 2201 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 4942 2201 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 4942 2201 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 5028 2201 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 5028 2201 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 5114 2201 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 5114 2201 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 5200 2201 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 5200 2201 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 5286 2201 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 5286 2201 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 5372 2201 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 5372 2201 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 5458 2201 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 5458 2201 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 5544 2201 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 5544 2201 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2137 5630 2201 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2137 5630 2201 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36289 2255 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36289 2255 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36370 2255 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36370 2255 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36451 2255 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36451 2255 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36532 2255 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36532 2255 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36613 2255 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36613 2255 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36694 2255 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36694 2255 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36775 2255 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36775 2255 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36856 2255 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36856 2255 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 36937 2255 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 36937 2255 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37018 2255 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37018 2255 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37099 2255 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37099 2255 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37180 2255 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37180 2255 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37261 2255 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37261 2255 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37342 2255 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37342 2255 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37423 2255 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37423 2255 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37504 2255 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37504 2255 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37585 2255 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37585 2255 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37666 2255 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37666 2255 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37747 2255 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37747 2255 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37828 2255 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37828 2255 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37909 2255 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37909 2255 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 37990 2255 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 37990 2255 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38071 2255 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38071 2255 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38152 2255 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38152 2255 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38233 2255 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38233 2255 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38314 2255 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38314 2255 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38395 2255 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38395 2255 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38476 2255 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38476 2255 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38557 2255 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38557 2255 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38638 2255 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38638 2255 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38719 2255 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38719 2255 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38800 2255 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38800 2255 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38881 2255 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38881 2255 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 38962 2255 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 38962 2255 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 39043 2255 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 39043 2255 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 39124 2255 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 39124 2255 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 39205 2255 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 39205 2255 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 39286 2255 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 39286 2255 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 39367 2255 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 39367 2255 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 39448 2255 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 39448 2255 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2191 39529 2255 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2191 39529 2255 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 34780 2243 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 34860 2243 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 34940 2243 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35020 2243 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35100 2243 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35180 2243 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35260 2243 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35340 2243 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35420 2243 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35500 2243 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35580 2243 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35660 2243 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35740 2243 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35820 2243 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35900 2243 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 35980 2243 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 36060 2243 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 36140 2243 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2203 36220 2243 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 4770 2282 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 4770 2282 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 4856 2282 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 4856 2282 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 4942 2282 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 4942 2282 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 5028 2282 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 5028 2282 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 5114 2282 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 5114 2282 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 5200 2282 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 5200 2282 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 5286 2282 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 5286 2282 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 5372 2282 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 5372 2282 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 5458 2282 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 5458 2282 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 5544 2282 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 5544 2282 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2218 5630 2282 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2218 5630 2282 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36289 2335 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36289 2335 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36370 2335 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36370 2335 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36451 2335 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36451 2335 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36532 2335 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36532 2335 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36613 2335 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36613 2335 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36694 2335 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36694 2335 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36775 2335 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36775 2335 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36856 2335 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36856 2335 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 36937 2335 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 36937 2335 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37018 2335 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37018 2335 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37099 2335 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37099 2335 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37180 2335 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37180 2335 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37261 2335 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37261 2335 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37342 2335 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37342 2335 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37423 2335 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37423 2335 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37504 2335 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37504 2335 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37585 2335 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37585 2335 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37666 2335 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37666 2335 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37747 2335 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37747 2335 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37828 2335 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37828 2335 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37909 2335 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37909 2335 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 37990 2335 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 37990 2335 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38071 2335 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38071 2335 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38152 2335 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38152 2335 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38233 2335 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38233 2335 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38314 2335 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38314 2335 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38395 2335 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38395 2335 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38476 2335 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38476 2335 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38557 2335 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38557 2335 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38638 2335 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38638 2335 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38719 2335 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38719 2335 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38800 2335 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38800 2335 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38881 2335 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38881 2335 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 38962 2335 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 38962 2335 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 39043 2335 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 39043 2335 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 39124 2335 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 39124 2335 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 39205 2335 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 39205 2335 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 39286 2335 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 39286 2335 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 39367 2335 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 39367 2335 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 39448 2335 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 39448 2335 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2271 39529 2335 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2271 39529 2335 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 34780 2323 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 34860 2323 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 34940 2323 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35020 2323 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35100 2323 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35180 2323 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35260 2323 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35340 2323 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35420 2323 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35500 2323 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35580 2323 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35660 2323 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35740 2323 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35820 2323 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35900 2323 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 35980 2323 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 36060 2323 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 36140 2323 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2283 36220 2323 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 4770 2363 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 4770 2363 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 4856 2363 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 4856 2363 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 4942 2363 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 4942 2363 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 5028 2363 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 5028 2363 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 5114 2363 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 5114 2363 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 5200 2363 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 5200 2363 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 5286 2363 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 5286 2363 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 5372 2363 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 5372 2363 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 5458 2363 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 5458 2363 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 5544 2363 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 5544 2363 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2299 5630 2363 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2299 5630 2363 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36289 2415 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36289 2415 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36370 2415 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36370 2415 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36451 2415 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36451 2415 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36532 2415 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36532 2415 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36613 2415 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36613 2415 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36694 2415 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36694 2415 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36775 2415 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36775 2415 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36856 2415 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36856 2415 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 36937 2415 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 36937 2415 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37018 2415 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37018 2415 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37099 2415 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37099 2415 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37180 2415 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37180 2415 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37261 2415 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37261 2415 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37342 2415 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37342 2415 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37423 2415 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37423 2415 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37504 2415 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37504 2415 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37585 2415 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37585 2415 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37666 2415 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37666 2415 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37747 2415 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37747 2415 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37828 2415 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37828 2415 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37909 2415 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37909 2415 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 37990 2415 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 37990 2415 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38071 2415 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38071 2415 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38152 2415 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38152 2415 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38233 2415 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38233 2415 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38314 2415 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38314 2415 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38395 2415 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38395 2415 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38476 2415 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38476 2415 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38557 2415 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38557 2415 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38638 2415 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38638 2415 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38719 2415 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38719 2415 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38800 2415 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38800 2415 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38881 2415 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38881 2415 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 38962 2415 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 38962 2415 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 39043 2415 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 39043 2415 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 39124 2415 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 39124 2415 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 39205 2415 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 39205 2415 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 39286 2415 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 39286 2415 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 39367 2415 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 39367 2415 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 39448 2415 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 39448 2415 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2351 39529 2415 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2351 39529 2415 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 34780 2403 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 34860 2403 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 34940 2403 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35020 2403 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35100 2403 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35180 2403 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35260 2403 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35340 2403 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35420 2403 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35500 2403 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35580 2403 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35660 2403 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35740 2403 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35820 2403 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35900 2403 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 35980 2403 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 36060 2403 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 36140 2403 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2363 36220 2403 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 4770 2444 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 4770 2444 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 4856 2444 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 4856 2444 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 4942 2444 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 4942 2444 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 5028 2444 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 5028 2444 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 5114 2444 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 5114 2444 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 5200 2444 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 5200 2444 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 5286 2444 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 5286 2444 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 5372 2444 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 5372 2444 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 5458 2444 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 5458 2444 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 5544 2444 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 5544 2444 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2380 5630 2444 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2380 5630 2444 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36289 2495 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36289 2495 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36370 2495 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36370 2495 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36451 2495 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36451 2495 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36532 2495 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36532 2495 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36613 2495 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36613 2495 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36694 2495 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36694 2495 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36775 2495 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36775 2495 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36856 2495 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36856 2495 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 36937 2495 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 36937 2495 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37018 2495 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37018 2495 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37099 2495 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37099 2495 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37180 2495 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37180 2495 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37261 2495 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37261 2495 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37342 2495 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37342 2495 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37423 2495 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37423 2495 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37504 2495 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37504 2495 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37585 2495 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37585 2495 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37666 2495 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37666 2495 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37747 2495 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37747 2495 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37828 2495 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37828 2495 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37909 2495 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37909 2495 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 37990 2495 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 37990 2495 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38071 2495 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38071 2495 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38152 2495 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38152 2495 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38233 2495 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38233 2495 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38314 2495 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38314 2495 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38395 2495 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38395 2495 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38476 2495 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38476 2495 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38557 2495 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38557 2495 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38638 2495 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38638 2495 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38719 2495 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38719 2495 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38800 2495 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38800 2495 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38881 2495 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38881 2495 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 38962 2495 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 38962 2495 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 39043 2495 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 39043 2495 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 39124 2495 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 39124 2495 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 39205 2495 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 39205 2495 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 39286 2495 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 39286 2495 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 39367 2495 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 39367 2495 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 39448 2495 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 39448 2495 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2431 39529 2495 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2431 39529 2495 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 34780 2483 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 34860 2483 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 34940 2483 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35020 2483 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35100 2483 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35180 2483 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35260 2483 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35340 2483 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35420 2483 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35500 2483 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35580 2483 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35660 2483 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35740 2483 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35820 2483 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35900 2483 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 35980 2483 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 36060 2483 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 36140 2483 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2443 36220 2483 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 4770 2525 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 4770 2525 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 4856 2525 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 4856 2525 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 4942 2525 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 4942 2525 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 5028 2525 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 5028 2525 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 5114 2525 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 5114 2525 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 5200 2525 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 5200 2525 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 5286 2525 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 5286 2525 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 5372 2525 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 5372 2525 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 5458 2525 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 5458 2525 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 5544 2525 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 5544 2525 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2461 5630 2525 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2461 5630 2525 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36289 2575 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36289 2575 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36370 2575 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36370 2575 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36451 2575 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36451 2575 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36532 2575 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36532 2575 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36613 2575 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36613 2575 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36694 2575 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36694 2575 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36775 2575 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36775 2575 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36856 2575 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36856 2575 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 36937 2575 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 36937 2575 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37018 2575 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37018 2575 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37099 2575 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37099 2575 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37180 2575 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37180 2575 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37261 2575 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37261 2575 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37342 2575 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37342 2575 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37423 2575 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37423 2575 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37504 2575 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37504 2575 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37585 2575 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37585 2575 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37666 2575 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37666 2575 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37747 2575 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37747 2575 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37828 2575 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37828 2575 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37909 2575 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37909 2575 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 37990 2575 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 37990 2575 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38071 2575 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38071 2575 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38152 2575 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38152 2575 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38233 2575 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38233 2575 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38314 2575 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38314 2575 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38395 2575 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38395 2575 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38476 2575 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38476 2575 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38557 2575 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38557 2575 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38638 2575 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38638 2575 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38719 2575 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38719 2575 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38800 2575 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38800 2575 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38881 2575 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38881 2575 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 38962 2575 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 38962 2575 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 39043 2575 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 39043 2575 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 39124 2575 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 39124 2575 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 39205 2575 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 39205 2575 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 39286 2575 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 39286 2575 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 39367 2575 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 39367 2575 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 39448 2575 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 39448 2575 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2511 39529 2575 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2511 39529 2575 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 34780 2563 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 34860 2563 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 34940 2563 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35020 2563 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35100 2563 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35180 2563 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35260 2563 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35340 2563 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35420 2563 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35500 2563 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35580 2563 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35660 2563 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35740 2563 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35820 2563 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35900 2563 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 35980 2563 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 36060 2563 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2523 36140 2563 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 4770 2606 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 4770 2606 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 4856 2606 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 4856 2606 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 4942 2606 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 4942 2606 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 5028 2606 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 5028 2606 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 5114 2606 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 5114 2606 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 5200 2606 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 5200 2606 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 5286 2606 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 5286 2606 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 5372 2606 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 5372 2606 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 5458 2606 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 5458 2606 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 5544 2606 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 5544 2606 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2542 5630 2606 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2542 5630 2606 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 4770 2687 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 4770 2687 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 4856 2687 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 4856 2687 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 4942 2687 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 4942 2687 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 5028 2687 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 5028 2687 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 5114 2687 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 5114 2687 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 5200 2687 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 5200 2687 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 5286 2687 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 5286 2687 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 5372 2687 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 5372 2687 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 5458 2687 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 5458 2687 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 5544 2687 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 5544 2687 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2623 5630 2687 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2623 5630 2687 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 4770 2768 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 4770 2768 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 4856 2768 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 4856 2768 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 4942 2768 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 4942 2768 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 5028 2768 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 5028 2768 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 5114 2768 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 5114 2768 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 5200 2768 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 5200 2768 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 5286 2768 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 5286 2768 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 5372 2768 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 5372 2768 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 5458 2768 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 5458 2768 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 5544 2768 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 5544 2768 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2704 5630 2768 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2704 5630 2768 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 4770 2849 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 4770 2849 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 4856 2849 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 4856 2849 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 4942 2849 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 4942 2849 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 5028 2849 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 5028 2849 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 5114 2849 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 5114 2849 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 5200 2849 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 5200 2849 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 5286 2849 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 5286 2849 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 5372 2849 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 5372 2849 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 5458 2849 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 5458 2849 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 5544 2849 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 5544 2849 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2785 5630 2849 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2785 5630 2849 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 4770 2930 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 4770 2930 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 4856 2930 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 4856 2930 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 4942 2930 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 4942 2930 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 5028 2930 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 5028 2930 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 5114 2930 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 5114 2930 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 5200 2930 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 5200 2930 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 5286 2930 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 5286 2930 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 5372 2930 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 5372 2930 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 5458 2930 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 5458 2930 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 5544 2930 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 5544 2930 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2866 5630 2930 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2866 5630 2930 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 4770 3011 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 4770 3011 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 4856 3011 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 4856 3011 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 4942 3011 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 4942 3011 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 5028 3011 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 5028 3011 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 5114 3011 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 5114 3011 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 5200 3011 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 5200 3011 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 5286 3011 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 5286 3011 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 5372 3011 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 5372 3011 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 5458 3011 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 5458 3011 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 5544 3011 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 5544 3011 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 2947 5630 3011 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 2947 5630 3011 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 4770 3092 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 4770 3092 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 4856 3092 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 4856 3092 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 4942 3092 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 4942 3092 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 5028 3092 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 5028 3092 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 5114 3092 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 5114 3092 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 5200 3092 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 5200 3092 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 5286 3092 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 5286 3092 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 5372 3092 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 5372 3092 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 5458 3092 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 5458 3092 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 5544 3092 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 5544 3092 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3028 5630 3092 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3028 5630 3092 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 4770 3173 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 4770 3173 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 4856 3173 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 4856 3173 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 4942 3173 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 4942 3173 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 5028 3173 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 5028 3173 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 5114 3173 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 5114 3173 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 5200 3173 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 5200 3173 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 5286 3173 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 5286 3173 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 5372 3173 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 5372 3173 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 5458 3173 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 5458 3173 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 5544 3173 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 5544 3173 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3109 5630 3173 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3109 5630 3173 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 4770 3254 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 4770 3254 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 4856 3254 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 4856 3254 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 4942 3254 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 4942 3254 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 5028 3254 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 5028 3254 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 5114 3254 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 5114 3254 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 5200 3254 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 5200 3254 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 5286 3254 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 5286 3254 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 5372 3254 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 5372 3254 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 5458 3254 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 5458 3254 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 5544 3254 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 5544 3254 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3190 5630 3254 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3190 5630 3254 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 4770 3335 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 4770 3335 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 4856 3335 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 4856 3335 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 4942 3335 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 4942 3335 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 5028 3335 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 5028 3335 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 5114 3335 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 5114 3335 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 5200 3335 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 5200 3335 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 5286 3335 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 5286 3335 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 5372 3335 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 5372 3335 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 5458 3335 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 5458 3335 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 5544 3335 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 5544 3335 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3271 5630 3335 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3271 5630 3335 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 4770 3416 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 4770 3416 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 4856 3416 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 4856 3416 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 4942 3416 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 4942 3416 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 5028 3416 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 5028 3416 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 5114 3416 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 5114 3416 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 5200 3416 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 5200 3416 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 5286 3416 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 5286 3416 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 5372 3416 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 5372 3416 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 5458 3416 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 5458 3416 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 5544 3416 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 5544 3416 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3352 5630 3416 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3352 5630 3416 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 4770 3497 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 4770 3497 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 4856 3497 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 4856 3497 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 4942 3497 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 4942 3497 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 5028 3497 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 5028 3497 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 5114 3497 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 5114 3497 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 5200 3497 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 5200 3497 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 5286 3497 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 5286 3497 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 5372 3497 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 5372 3497 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 5458 3497 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 5458 3497 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 5544 3497 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 5544 3497 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3433 5630 3497 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3433 5630 3497 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 4770 3578 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 4770 3578 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 4856 3578 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 4856 3578 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 4942 3578 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 4942 3578 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 5028 3578 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 5028 3578 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 5114 3578 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 5114 3578 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 5200 3578 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 5200 3578 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 5286 3578 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 5286 3578 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 5372 3578 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 5372 3578 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 5458 3578 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 5458 3578 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 5544 3578 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 5544 3578 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3514 5630 3578 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3514 5630 3578 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 4770 3659 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 4770 3659 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 4856 3659 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 4856 3659 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 4942 3659 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 4942 3659 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 5028 3659 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 5028 3659 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 5114 3659 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 5114 3659 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 5200 3659 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 5200 3659 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 5286 3659 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 5286 3659 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 5372 3659 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 5372 3659 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 5458 3659 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 5458 3659 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 5544 3659 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 5544 3659 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3595 5630 3659 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3595 5630 3659 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 4770 3740 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 4770 3740 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 4856 3740 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 4856 3740 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 4942 3740 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 4942 3740 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 5028 3740 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 5028 3740 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 5114 3740 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 5114 3740 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 5200 3740 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 5200 3740 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 5286 3740 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 5286 3740 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 5372 3740 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 5372 3740 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 5458 3740 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 5458 3740 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 5544 3740 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 5544 3740 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3676 5630 3740 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3676 5630 3740 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 4770 3821 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 4770 3821 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 4856 3821 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 4856 3821 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 4942 3821 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 4942 3821 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 5028 3821 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 5028 3821 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 5114 3821 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 5114 3821 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 5200 3821 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 5200 3821 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 5286 3821 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 5286 3821 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 5372 3821 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 5372 3821 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 5458 3821 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 5458 3821 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 5544 3821 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 5544 3821 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3757 5630 3821 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3757 5630 3821 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 4770 3902 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 4770 3902 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 4856 3902 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 4856 3902 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 4942 3902 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 4942 3902 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 5028 3902 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 5028 3902 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 5114 3902 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 5114 3902 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 5200 3902 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 5200 3902 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 5286 3902 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 5286 3902 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 5372 3902 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 5372 3902 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 5458 3902 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 5458 3902 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 5544 3902 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 5544 3902 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3838 5630 3902 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3838 5630 3902 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 4770 3983 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 4770 3983 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 4856 3983 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 4856 3983 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 4942 3983 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 4942 3983 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 5028 3983 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 5028 3983 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 5114 3983 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 5114 3983 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 5200 3983 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 5200 3983 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 5286 3983 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 5286 3983 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 5372 3983 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 5372 3983 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 5458 3983 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 5458 3983 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 5544 3983 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 5544 3983 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 3919 5630 3983 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 3919 5630 3983 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36289 495 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36289 495 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36370 495 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36370 495 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36451 495 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36451 495 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36532 495 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36532 495 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36613 495 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36613 495 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36694 495 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36694 495 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36775 495 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36775 495 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36856 495 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36856 495 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 36937 495 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 36937 495 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37018 495 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37018 495 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37099 495 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37099 495 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37180 495 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37180 495 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37261 495 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37261 495 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37342 495 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37342 495 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37423 495 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37423 495 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37504 495 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37504 495 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37585 495 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37585 495 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37666 495 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37666 495 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37747 495 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37747 495 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37828 495 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37828 495 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37909 495 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37909 495 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 37990 495 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 37990 495 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38071 495 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38071 495 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38152 495 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38152 495 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38233 495 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38233 495 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38314 495 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38314 495 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38395 495 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38395 495 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38476 495 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38476 495 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38557 495 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38557 495 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38638 495 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38638 495 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38719 495 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38719 495 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38800 495 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38800 495 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38881 495 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38881 495 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 38962 495 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 38962 495 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 39043 495 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 39043 495 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 39124 495 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 39124 495 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 39205 495 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 39205 495 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 39286 495 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 39286 495 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 39367 495 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 39367 495 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 39448 495 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 39448 495 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 431 39529 495 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 431 39529 495 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 4770 498 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 4770 498 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 4856 498 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 4856 498 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 4942 498 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 4942 498 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 5028 498 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 5028 498 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 5114 498 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 5114 498 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 5200 498 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 5200 498 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 5286 498 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 5286 498 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 5372 498 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 5372 498 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 5458 498 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 5458 498 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 5544 498 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 5544 498 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 434 5630 498 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 434 5630 498 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 34780 483 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 34860 483 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 34940 483 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35020 483 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35100 483 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35180 483 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35260 483 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35340 483 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35420 483 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35500 483 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35580 483 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35660 483 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35740 483 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35820 483 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35900 483 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 35980 483 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 36060 483 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 36140 483 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 443 36220 483 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36289 575 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36289 575 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36370 575 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36370 575 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36451 575 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36451 575 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36532 575 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36532 575 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36613 575 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36613 575 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36694 575 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36694 575 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36775 575 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36775 575 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36856 575 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36856 575 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 36937 575 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 36937 575 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37018 575 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37018 575 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37099 575 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37099 575 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37180 575 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37180 575 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37261 575 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37261 575 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37342 575 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37342 575 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37423 575 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37423 575 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37504 575 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37504 575 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37585 575 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37585 575 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37666 575 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37666 575 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37747 575 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37747 575 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37828 575 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37828 575 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37909 575 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37909 575 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 37990 575 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 37990 575 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38071 575 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38071 575 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38152 575 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38152 575 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38233 575 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38233 575 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38314 575 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38314 575 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38395 575 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38395 575 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38476 575 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38476 575 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38557 575 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38557 575 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38638 575 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38638 575 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38719 575 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38719 575 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38800 575 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38800 575 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38881 575 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38881 575 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 38962 575 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 38962 575 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 39043 575 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 39043 575 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 39124 575 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 39124 575 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 39205 575 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 39205 575 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 39286 575 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 39286 575 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 39367 575 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 39367 575 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 39448 575 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 39448 575 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 511 39529 575 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 511 39529 575 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 4770 580 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 4770 580 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 4856 580 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 4856 580 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 4942 580 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 4942 580 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 5028 580 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 5028 580 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 5114 580 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 5114 580 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 5200 580 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 5200 580 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 5286 580 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 5286 580 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 5372 580 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 5372 580 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 5458 580 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 5458 580 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 5544 580 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 5544 580 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 516 5630 580 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 516 5630 580 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 34780 563 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 34860 563 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 34940 563 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35020 563 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35100 563 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35180 563 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35260 563 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35340 563 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35420 563 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35500 563 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35580 563 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35660 563 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35740 563 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35820 563 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35900 563 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 35980 563 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 36060 563 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 36140 563 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 523 36220 563 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36289 655 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36289 655 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36370 655 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36370 655 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36451 655 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36451 655 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36532 655 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36532 655 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36613 655 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36613 655 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36694 655 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36694 655 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36775 655 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36775 655 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36856 655 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36856 655 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 36937 655 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 36937 655 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37018 655 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37018 655 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37099 655 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37099 655 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37180 655 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37180 655 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37261 655 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37261 655 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37342 655 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37342 655 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37423 655 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37423 655 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37504 655 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37504 655 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37585 655 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37585 655 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37666 655 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37666 655 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37747 655 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37747 655 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37828 655 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37828 655 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37909 655 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37909 655 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 37990 655 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 37990 655 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38071 655 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38071 655 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38152 655 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38152 655 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38233 655 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38233 655 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38314 655 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38314 655 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38395 655 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38395 655 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38476 655 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38476 655 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38557 655 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38557 655 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38638 655 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38638 655 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38719 655 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38719 655 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38800 655 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38800 655 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38881 655 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38881 655 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 38962 655 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 38962 655 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 39043 655 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 39043 655 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 39124 655 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 39124 655 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 39205 655 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 39205 655 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 39286 655 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 39286 655 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 39367 655 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 39367 655 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 39448 655 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 39448 655 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 591 39529 655 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 591 39529 655 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 4770 662 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 4770 662 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 4856 662 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 4856 662 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 4942 662 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 4942 662 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 5028 662 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 5028 662 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 5114 662 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 5114 662 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 5200 662 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 5200 662 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 5286 662 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 5286 662 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 5372 662 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 5372 662 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 5458 662 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 5458 662 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 5544 662 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 5544 662 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 598 5630 662 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 598 5630 662 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 4770 4064 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 4770 4064 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 4856 4064 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 4856 4064 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 4942 4064 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 4942 4064 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 5028 4064 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 5028 4064 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 5114 4064 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 5114 4064 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 5200 4064 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 5200 4064 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 5286 4064 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 5286 4064 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 5372 4064 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 5372 4064 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 5458 4064 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 5458 4064 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 5544 4064 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 5544 4064 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4000 5630 4064 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4000 5630 4064 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 4770 4145 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 4770 4145 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 4856 4145 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 4856 4145 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 4942 4145 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 4942 4145 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 5028 4145 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 5028 4145 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 5114 4145 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 5114 4145 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 5200 4145 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 5200 4145 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 5286 4145 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 5286 4145 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 5372 4145 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 5372 4145 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 5458 4145 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 5458 4145 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 5544 4145 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 5544 4145 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4081 5630 4145 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4081 5630 4145 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 4770 4226 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 4770 4226 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 4856 4226 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 4856 4226 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 4942 4226 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 4942 4226 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 5028 4226 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 5028 4226 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 5114 4226 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 5114 4226 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 5200 4226 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 5200 4226 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 5286 4226 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 5286 4226 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 5372 4226 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 5372 4226 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 5458 4226 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 5458 4226 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 5544 4226 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 5544 4226 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4162 5630 4226 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4162 5630 4226 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 4770 4307 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 4770 4307 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 4856 4307 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 4856 4307 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 4942 4307 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 4942 4307 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 5028 4307 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 5028 4307 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 5114 4307 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 5114 4307 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 5200 4307 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 5200 4307 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 5286 4307 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 5286 4307 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 5372 4307 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 5372 4307 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 5458 4307 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 5458 4307 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 5544 4307 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 5544 4307 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4243 5630 4307 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4243 5630 4307 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 4770 4388 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 4770 4388 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 4856 4388 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 4856 4388 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 4942 4388 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 4942 4388 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 5028 4388 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 5028 4388 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 5114 4388 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 5114 4388 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 5200 4388 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 5200 4388 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 5286 4388 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 5286 4388 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 5372 4388 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 5372 4388 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 5458 4388 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 5458 4388 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 5544 4388 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 5544 4388 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4324 5630 4388 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4324 5630 4388 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 4770 4469 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 4770 4469 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 4856 4469 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 4856 4469 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 4942 4469 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 4942 4469 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 5028 4469 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 5028 4469 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 5114 4469 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 5114 4469 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 5200 4469 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 5200 4469 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 5286 4469 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 5286 4469 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 5372 4469 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 5372 4469 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 5458 4469 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 5458 4469 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 5544 4469 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 5544 4469 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4405 5630 4469 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4405 5630 4469 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 4770 4550 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 4770 4550 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 4856 4550 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 4856 4550 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 4942 4550 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 4942 4550 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 5028 4550 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 5028 4550 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 5114 4550 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 5114 4550 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 5200 4550 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 5200 4550 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 5286 4550 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 5286 4550 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 5372 4550 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 5372 4550 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 5458 4550 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 5458 4550 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 5544 4550 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 5544 4550 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4486 5630 4550 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4486 5630 4550 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 4770 4631 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 4770 4631 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 4856 4631 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 4856 4631 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 4942 4631 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 4942 4631 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 5028 4631 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 5028 4631 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 5114 4631 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 5114 4631 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 5200 4631 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 5200 4631 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 5286 4631 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 5286 4631 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 5372 4631 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 5372 4631 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 5458 4631 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 5458 4631 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 5544 4631 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 5544 4631 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4567 5630 4631 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4567 5630 4631 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 4770 4712 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 4770 4712 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 4856 4712 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 4856 4712 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 4942 4712 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 4942 4712 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 5028 4712 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 5028 4712 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 5114 4712 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 5114 4712 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 5200 4712 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 5200 4712 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 5286 4712 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 5286 4712 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 5372 4712 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 5372 4712 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 5458 4712 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 5458 4712 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 5544 4712 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 5544 4712 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4648 5630 4712 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4648 5630 4712 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 4770 4793 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 4770 4793 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 4856 4793 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 4856 4793 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 4942 4793 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 4942 4793 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 5028 4793 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 5028 4793 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 5114 4793 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 5114 4793 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 5200 4793 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 5200 4793 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 5286 4793 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 5286 4793 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 5372 4793 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 5372 4793 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 5458 4793 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 5458 4793 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 5544 4793 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 5544 4793 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4729 5630 4793 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4729 5630 4793 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 4770 4874 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 4770 4874 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 4856 4874 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 4856 4874 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 4942 4874 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 4942 4874 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 5028 4874 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 5028 4874 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 5114 4874 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 5114 4874 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 5200 4874 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 5200 4874 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 5286 4874 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 5286 4874 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 5372 4874 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 5372 4874 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 5458 4874 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 5458 4874 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 5544 4874 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 5544 4874 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 4810 5630 4874 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 4810 5630 4874 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 34780 643 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 34860 643 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 34940 643 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35020 643 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35100 643 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35180 643 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35260 643 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35340 643 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35420 643 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35500 643 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35580 643 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35660 643 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35740 643 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35820 643 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35900 643 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 35980 643 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 36060 643 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 36140 643 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 603 36220 643 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36289 735 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36289 735 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36370 735 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36370 735 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36451 735 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36451 735 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36532 735 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36532 735 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36613 735 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36613 735 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36694 735 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36694 735 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36775 735 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36775 735 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36856 735 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36856 735 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 36937 735 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 36937 735 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37018 735 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37018 735 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37099 735 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37099 735 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37180 735 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37180 735 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37261 735 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37261 735 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37342 735 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37342 735 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37423 735 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37423 735 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37504 735 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37504 735 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37585 735 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37585 735 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37666 735 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37666 735 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37747 735 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37747 735 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37828 735 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37828 735 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37909 735 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37909 735 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 37990 735 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 37990 735 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38071 735 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38071 735 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38152 735 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38152 735 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38233 735 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38233 735 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38314 735 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38314 735 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38395 735 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38395 735 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38476 735 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38476 735 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38557 735 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38557 735 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38638 735 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38638 735 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38719 735 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38719 735 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38800 735 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38800 735 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38881 735 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38881 735 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 38962 735 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 38962 735 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 39043 735 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 39043 735 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 39124 735 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 39124 735 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 39205 735 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 39205 735 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 39286 735 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 39286 735 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 39367 735 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 39367 735 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 39448 735 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 39448 735 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 671 39529 735 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 671 39529 735 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 4770 743 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 4770 743 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 4856 743 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 4856 743 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 4942 743 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 4942 743 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 5028 743 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 5028 743 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 5114 743 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 5114 743 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 5200 743 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 5200 743 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 5286 743 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 5286 743 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 5372 743 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 5372 743 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 5458 743 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 5458 743 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 5544 743 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 5544 743 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 679 5630 743 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 679 5630 743 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 34780 723 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 34860 723 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 34940 723 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35020 723 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35100 723 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35180 723 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35260 723 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35340 723 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35420 723 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35500 723 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35580 723 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35660 723 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35740 723 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35820 723 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35900 723 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 35980 723 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 36060 723 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 36140 723 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 683 36220 723 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36289 815 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36289 815 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36370 815 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36370 815 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36451 815 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36451 815 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36532 815 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36532 815 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36613 815 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36613 815 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36694 815 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36694 815 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36775 815 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36775 815 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36856 815 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36856 815 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 36937 815 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 36937 815 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37018 815 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37018 815 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37099 815 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37099 815 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37180 815 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37180 815 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37261 815 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37261 815 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37342 815 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37342 815 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37423 815 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37423 815 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37504 815 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37504 815 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37585 815 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37585 815 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37666 815 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37666 815 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37747 815 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37747 815 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37828 815 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37828 815 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37909 815 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37909 815 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 37990 815 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 37990 815 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38071 815 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38071 815 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38152 815 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38152 815 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38233 815 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38233 815 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38314 815 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38314 815 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38395 815 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38395 815 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38476 815 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38476 815 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38557 815 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38557 815 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38638 815 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38638 815 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38719 815 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38719 815 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38800 815 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38800 815 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38881 815 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38881 815 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 38962 815 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 38962 815 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 39043 815 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 39043 815 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 39124 815 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 39124 815 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 39205 815 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 39205 815 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 39286 815 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 39286 815 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 39367 815 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 39367 815 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 39448 815 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 39448 815 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 751 39529 815 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 751 39529 815 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 4770 824 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 4770 824 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 4856 824 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 4856 824 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 4942 824 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 4942 824 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 5028 824 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 5028 824 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 5114 824 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 5114 824 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 5200 824 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 5200 824 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 5286 824 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 5286 824 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 5372 824 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 5372 824 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 5458 824 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 5458 824 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 5544 824 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 5544 824 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 760 5630 824 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 760 5630 824 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 34780 803 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 34860 803 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 34940 803 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35020 803 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35100 803 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35180 803 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35260 803 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35340 803 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35420 803 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35500 803 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35580 803 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35660 803 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35740 803 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35820 803 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35900 803 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 35980 803 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 36060 803 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 36140 803 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 763 36220 803 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36289 895 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36289 895 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36370 895 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36370 895 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36451 895 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36451 895 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36532 895 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36532 895 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36613 895 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36613 895 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36694 895 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36694 895 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36775 895 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36775 895 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36856 895 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36856 895 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 36937 895 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 36937 895 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37018 895 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37018 895 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37099 895 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37099 895 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37180 895 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37180 895 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37261 895 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37261 895 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37342 895 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37342 895 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37423 895 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37423 895 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37504 895 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37504 895 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37585 895 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37585 895 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37666 895 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37666 895 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37747 895 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37747 895 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37828 895 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37828 895 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37909 895 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37909 895 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 37990 895 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 37990 895 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38071 895 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38071 895 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38152 895 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38152 895 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38233 895 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38233 895 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38314 895 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38314 895 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38395 895 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38395 895 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38476 895 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38476 895 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38557 895 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38557 895 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38638 895 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38638 895 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38719 895 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38719 895 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38800 895 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38800 895 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38881 895 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38881 895 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 38962 895 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 38962 895 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 39043 895 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 39043 895 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 39124 895 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 39124 895 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 39205 895 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 39205 895 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 39286 895 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 39286 895 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 39367 895 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 39367 895 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 39448 895 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 39448 895 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 831 39529 895 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 831 39529 895 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 4770 905 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 4770 905 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 4856 905 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 4856 905 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 4942 905 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 4942 905 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 5028 905 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 5028 905 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 5114 905 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 5114 905 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 5200 905 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 5200 905 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 5286 905 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 5286 905 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 5372 905 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 5372 905 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 5458 905 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 5458 905 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 5544 905 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 5544 905 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 841 5630 905 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 841 5630 905 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 34780 883 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 34860 883 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 34940 883 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35020 883 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35100 883 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35180 883 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35260 883 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35340 883 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35420 883 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35500 883 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35580 883 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35660 883 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35740 883 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35820 883 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35900 883 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 35980 883 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 36060 883 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 36140 883 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 843 36220 883 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36289 975 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36289 975 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36370 975 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36370 975 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36451 975 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36451 975 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36532 975 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36532 975 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36613 975 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36613 975 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36694 975 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36694 975 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36775 975 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36775 975 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36856 975 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36856 975 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 36937 975 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 36937 975 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37018 975 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37018 975 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37099 975 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37099 975 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37180 975 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37180 975 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37261 975 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37261 975 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37342 975 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37342 975 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37423 975 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37423 975 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37504 975 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37504 975 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37585 975 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37585 975 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37666 975 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37666 975 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37747 975 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37747 975 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37828 975 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37828 975 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37909 975 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37909 975 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 37990 975 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 37990 975 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38071 975 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38071 975 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38152 975 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38152 975 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38233 975 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38233 975 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38314 975 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38314 975 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38395 975 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38395 975 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38476 975 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38476 975 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38557 975 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38557 975 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38638 975 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38638 975 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38719 975 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38719 975 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38800 975 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38800 975 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38881 975 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38881 975 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 38962 975 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 38962 975 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 39043 975 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 39043 975 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 39124 975 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 39124 975 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 39205 975 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 39205 975 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 39286 975 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 39286 975 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 39367 975 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 39367 975 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 39448 975 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 39448 975 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 911 39529 975 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 911 39529 975 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 4770 986 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 4770 986 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 4856 986 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 4856 986 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 4942 986 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 4942 986 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 5028 986 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 5028 986 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 5114 986 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 5114 986 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 5200 986 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 5200 986 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 5286 986 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 5286 986 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 5372 986 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 5372 986 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 5458 986 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 5458 986 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 5544 986 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 5544 986 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 922 5630 986 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 922 5630 986 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 34780 963 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 34860 963 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 34940 963 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35020 963 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35100 963 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35180 963 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35260 963 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35340 963 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35420 963 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35500 963 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35580 963 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35660 963 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35740 963 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35820 963 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35900 963 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 35980 963 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 36060 963 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 36140 963 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 923 36220 963 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36289 1055 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36289 1055 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36370 1055 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36370 1055 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36451 1055 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36451 1055 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36532 1055 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36532 1055 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36613 1055 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36613 1055 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36694 1055 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36694 1055 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36775 1055 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36775 1055 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36856 1055 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36856 1055 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 36937 1055 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 36937 1055 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37018 1055 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37018 1055 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37099 1055 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37099 1055 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37180 1055 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37180 1055 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37261 1055 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37261 1055 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37342 1055 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37342 1055 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37423 1055 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37423 1055 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37504 1055 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37504 1055 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37585 1055 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37585 1055 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37666 1055 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37666 1055 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37747 1055 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37747 1055 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37828 1055 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37828 1055 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37909 1055 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37909 1055 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 37990 1055 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 37990 1055 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38071 1055 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38071 1055 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38152 1055 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38152 1055 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38233 1055 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38233 1055 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38314 1055 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38314 1055 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38395 1055 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38395 1055 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38476 1055 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38476 1055 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38557 1055 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38557 1055 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38638 1055 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38638 1055 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38719 1055 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38719 1055 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38800 1055 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38800 1055 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38881 1055 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38881 1055 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 38962 1055 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 38962 1055 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 39043 1055 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 39043 1055 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 39124 1055 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 39124 1055 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 39205 1055 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 39205 1055 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 39286 1055 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 39286 1055 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 39367 1055 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 39367 1055 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 39448 1055 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 39448 1055 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 991 39529 1055 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 991 39529 1055 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 34780 1043 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 34860 1043 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 34940 1043 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35020 1043 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35100 1043 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35180 1043 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35260 1043 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35340 1043 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35420 1043 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35500 1043 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35580 1043 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35660 1043 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35740 1043 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35820 1043 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35900 1043 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 35980 1043 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 36060 1043 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 36140 1043 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 36220 1043 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 4770 1067 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 4770 1067 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 4856 1067 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 4856 1067 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 4942 1067 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 4942 1067 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 5028 1067 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 5028 1067 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 5114 1067 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 5114 1067 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 5200 1067 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 5200 1067 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 5286 1067 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 5286 1067 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 5372 1067 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 5372 1067 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 5458 1067 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 5458 1067 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 5544 1067 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 5544 1067 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1003 5630 1067 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1003 5630 1067 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36289 1135 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36289 1135 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36370 1135 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36370 1135 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36451 1135 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36451 1135 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36532 1135 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36532 1135 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36613 1135 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36613 1135 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36694 1135 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36694 1135 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36775 1135 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36775 1135 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36856 1135 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36856 1135 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 36937 1135 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 36937 1135 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37018 1135 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37018 1135 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37099 1135 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37099 1135 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37180 1135 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37180 1135 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37261 1135 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37261 1135 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37342 1135 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37342 1135 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37423 1135 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37423 1135 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37504 1135 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37504 1135 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37585 1135 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37585 1135 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37666 1135 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37666 1135 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37747 1135 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37747 1135 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37828 1135 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37828 1135 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37909 1135 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37909 1135 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 37990 1135 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 37990 1135 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38071 1135 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38071 1135 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38152 1135 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38152 1135 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38233 1135 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38233 1135 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38314 1135 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38314 1135 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38395 1135 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38395 1135 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38476 1135 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38476 1135 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38557 1135 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38557 1135 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38638 1135 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38638 1135 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38719 1135 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38719 1135 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38800 1135 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38800 1135 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38881 1135 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38881 1135 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 38962 1135 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 38962 1135 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 39043 1135 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 39043 1135 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 39124 1135 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 39124 1135 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 39205 1135 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 39205 1135 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 39286 1135 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 39286 1135 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 39367 1135 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 39367 1135 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 39448 1135 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 39448 1135 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1071 39529 1135 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1071 39529 1135 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 34780 1123 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 34860 1123 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 34940 1123 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35020 1123 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35100 1123 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35180 1123 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35260 1123 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35340 1123 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35420 1123 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35500 1123 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35580 1123 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35660 1123 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35740 1123 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35820 1123 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35900 1123 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 35980 1123 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 36060 1123 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 36140 1123 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1083 36220 1123 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 4770 1148 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 4770 1148 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 4856 1148 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 4856 1148 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 4942 1148 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 4942 1148 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 5028 1148 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 5028 1148 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 5114 1148 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 5114 1148 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 5200 1148 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 5200 1148 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 5286 1148 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 5286 1148 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 5372 1148 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 5372 1148 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 5458 1148 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 5458 1148 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 5544 1148 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 5544 1148 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1084 5630 1148 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1084 5630 1148 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36289 1215 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36289 1215 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36370 1215 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36370 1215 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36451 1215 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36451 1215 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36532 1215 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36532 1215 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36613 1215 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36613 1215 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36694 1215 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36694 1215 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36775 1215 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36775 1215 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36856 1215 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36856 1215 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 36937 1215 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 36937 1215 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37018 1215 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37018 1215 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37099 1215 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37099 1215 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37180 1215 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37180 1215 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37261 1215 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37261 1215 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37342 1215 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37342 1215 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37423 1215 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37423 1215 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37504 1215 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37504 1215 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37585 1215 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37585 1215 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37666 1215 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37666 1215 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37747 1215 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37747 1215 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37828 1215 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37828 1215 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37909 1215 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37909 1215 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 37990 1215 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 37990 1215 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38071 1215 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38071 1215 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38152 1215 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38152 1215 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38233 1215 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38233 1215 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38314 1215 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38314 1215 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38395 1215 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38395 1215 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38476 1215 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38476 1215 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38557 1215 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38557 1215 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38638 1215 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38638 1215 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38719 1215 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38719 1215 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38800 1215 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38800 1215 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38881 1215 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38881 1215 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 38962 1215 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 38962 1215 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 39043 1215 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 39043 1215 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 39124 1215 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 39124 1215 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 39205 1215 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 39205 1215 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 39286 1215 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 39286 1215 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 39367 1215 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 39367 1215 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 39448 1215 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 39448 1215 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1151 39529 1215 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1151 39529 1215 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 34780 1203 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 34860 1203 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 34940 1203 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35020 1203 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35100 1203 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35180 1203 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35260 1203 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35340 1203 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35420 1203 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35500 1203 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35580 1203 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35660 1203 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35740 1203 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35820 1203 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35900 1203 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 35980 1203 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 36060 1203 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 36140 1203 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1163 36220 1203 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 4770 1229 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 4770 1229 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 4856 1229 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 4856 1229 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 4942 1229 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 4942 1229 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 5028 1229 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 5028 1229 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 5114 1229 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 5114 1229 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 5200 1229 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 5200 1229 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 5286 1229 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 5286 1229 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 5372 1229 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 5372 1229 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 5458 1229 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 5458 1229 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 5544 1229 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 5544 1229 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1165 5630 1229 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1165 5630 1229 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 4770 10221 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 4770 10221 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 4856 10221 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 4856 10221 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 4942 10221 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 4942 10221 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 5028 10221 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 5028 10221 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 5114 10221 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 5114 10221 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 5200 10221 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 5200 10221 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 5286 10221 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 5286 10221 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 5372 10221 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 5372 10221 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 5458 10221 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 5458 10221 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 5544 10221 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 5544 10221 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10157 5630 10221 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10157 5630 10221 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 4770 10303 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 4770 10303 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 4856 10303 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 4856 10303 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 4942 10303 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 4942 10303 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 5028 10303 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 5028 10303 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 5114 10303 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 5114 10303 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 5200 10303 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 5200 10303 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 5286 10303 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 5286 10303 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 5372 10303 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 5372 10303 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 5458 10303 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 5458 10303 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 5544 10303 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 5544 10303 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10239 5630 10303 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10239 5630 10303 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 4770 10385 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 4770 10385 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 4856 10385 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 4856 10385 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 4942 10385 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 4942 10385 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 5028 10385 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 5028 10385 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 5114 10385 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 5114 10385 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 5200 10385 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 5200 10385 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 5286 10385 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 5286 10385 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 5372 10385 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 5372 10385 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 5458 10385 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 5458 10385 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 5544 10385 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 5544 10385 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10321 5630 10385 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10321 5630 10385 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 4770 10467 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 4770 10467 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 4856 10467 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 4856 10467 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 4942 10467 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 4942 10467 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 5028 10467 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 5028 10467 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 5114 10467 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 5114 10467 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 5200 10467 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 5200 10467 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 5286 10467 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 5286 10467 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 5372 10467 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 5372 10467 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 5458 10467 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 5458 10467 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 5544 10467 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 5544 10467 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10403 5630 10467 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10403 5630 10467 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 4770 10549 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 4770 10549 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 4856 10549 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 4856 10549 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 4942 10549 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 4942 10549 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 5028 10549 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 5028 10549 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 5114 10549 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 5114 10549 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 5200 10549 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 5200 10549 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 5286 10549 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 5286 10549 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 5372 10549 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 5372 10549 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 5458 10549 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 5458 10549 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 5544 10549 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 5544 10549 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10485 5630 10549 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10485 5630 10549 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 4770 10631 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 4770 10631 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 4856 10631 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 4856 10631 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 4942 10631 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 4942 10631 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 5028 10631 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 5028 10631 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 5114 10631 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 5114 10631 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 5200 10631 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 5200 10631 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 5286 10631 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 5286 10631 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 5372 10631 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 5372 10631 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 5458 10631 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 5458 10631 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 5544 10631 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 5544 10631 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10567 5630 10631 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10567 5630 10631 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 4770 10713 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 4770 10713 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 4856 10713 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 4856 10713 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 4942 10713 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 4942 10713 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 5028 10713 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 5028 10713 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 5114 10713 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 5114 10713 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 5200 10713 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 5200 10713 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 5286 10713 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 5286 10713 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 5372 10713 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 5372 10713 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 5458 10713 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 5458 10713 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 5544 10713 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 5544 10713 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10649 5630 10713 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10649 5630 10713 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 4770 10795 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 4770 10795 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 4856 10795 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 4856 10795 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 4942 10795 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 4942 10795 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 5028 10795 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 5028 10795 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 5114 10795 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 5114 10795 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 5200 10795 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 5200 10795 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 5286 10795 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 5286 10795 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 5372 10795 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 5372 10795 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 5458 10795 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 5458 10795 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 5544 10795 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 5544 10795 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10731 5630 10795 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10731 5630 10795 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 4770 10877 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 4770 10877 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 4856 10877 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 4856 10877 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 4942 10877 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 4942 10877 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 5028 10877 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 5028 10877 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 5114 10877 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 5114 10877 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 5200 10877 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 5200 10877 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 5286 10877 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 5286 10877 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 5372 10877 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 5372 10877 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 5458 10877 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 5458 10877 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 5544 10877 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 5544 10877 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10813 5630 10877 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10813 5630 10877 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 4770 10959 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 4770 10959 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 4856 10959 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 4856 10959 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 4942 10959 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 4942 10959 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 5028 10959 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 5028 10959 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 5114 10959 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 5114 10959 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 5200 10959 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 5200 10959 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 5286 10959 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 5286 10959 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 5372 10959 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 5372 10959 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 5458 10959 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 5458 10959 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 5544 10959 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 5544 10959 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10895 5630 10959 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10895 5630 10959 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 4770 11041 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 4770 11041 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 4856 11041 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 4856 11041 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 4942 11041 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 4942 11041 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 5028 11041 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 5028 11041 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 5114 11041 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 5114 11041 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 5200 11041 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 5200 11041 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 5286 11041 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 5286 11041 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 5372 11041 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 5372 11041 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 5458 11041 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 5458 11041 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 5544 11041 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 5544 11041 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 10977 5630 11041 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 10977 5630 11041 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 4770 11123 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 4770 11123 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 4856 11123 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 4856 11123 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 4942 11123 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 4942 11123 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 5028 11123 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 5028 11123 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 5114 11123 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 5114 11123 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 5200 11123 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 5200 11123 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 5286 11123 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 5286 11123 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 5372 11123 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 5372 11123 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 5458 11123 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 5458 11123 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 5544 11123 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 5544 11123 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11059 5630 11123 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11059 5630 11123 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 4770 11205 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 4770 11205 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 4856 11205 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 4856 11205 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 4942 11205 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 4942 11205 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 5028 11205 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 5028 11205 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 5114 11205 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 5114 11205 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 5200 11205 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 5200 11205 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 5286 11205 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 5286 11205 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 5372 11205 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 5372 11205 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 5458 11205 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 5458 11205 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 5544 11205 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 5544 11205 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11141 5630 11205 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11141 5630 11205 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 4770 11287 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 4770 11287 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 4856 11287 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 4856 11287 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 4942 11287 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 4942 11287 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 5028 11287 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 5028 11287 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 5114 11287 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 5114 11287 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 5200 11287 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 5200 11287 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 5286 11287 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 5286 11287 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 5372 11287 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 5372 11287 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 5458 11287 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 5458 11287 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 5544 11287 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 5544 11287 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11223 5630 11287 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11223 5630 11287 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 4770 11369 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 4770 11369 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 4856 11369 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 4856 11369 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 4942 11369 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 4942 11369 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 5028 11369 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 5028 11369 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 5114 11369 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 5114 11369 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 5200 11369 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 5200 11369 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 5286 11369 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 5286 11369 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 5372 11369 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 5372 11369 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 5458 11369 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 5458 11369 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 5544 11369 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 5544 11369 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11305 5630 11369 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11305 5630 11369 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 4770 11450 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 4770 11450 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 4856 11450 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 4856 11450 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 4942 11450 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 4942 11450 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 5028 11450 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 5028 11450 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 5114 11450 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 5114 11450 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 5200 11450 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 5200 11450 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 5286 11450 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 5286 11450 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 5372 11450 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 5372 11450 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 5458 11450 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 5458 11450 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 5544 11450 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 5544 11450 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11386 5630 11450 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11386 5630 11450 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 4770 11531 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 4770 11531 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 4856 11531 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 4856 11531 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 4942 11531 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 4942 11531 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 5028 11531 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 5028 11531 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 5114 11531 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 5114 11531 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 5200 11531 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 5200 11531 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 5286 11531 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 5286 11531 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 5372 11531 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 5372 11531 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 5458 11531 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 5458 11531 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 5544 11531 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 5544 11531 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11467 5630 11531 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11467 5630 11531 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 4770 11612 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 4770 11612 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 4856 11612 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 4856 11612 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 4942 11612 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 4942 11612 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 5028 11612 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 5028 11612 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 5114 11612 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 5114 11612 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 5200 11612 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 5200 11612 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 5286 11612 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 5286 11612 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 5372 11612 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 5372 11612 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 5458 11612 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 5458 11612 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 5544 11612 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 5544 11612 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11548 5630 11612 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11548 5630 11612 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 4770 11693 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 4770 11693 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 4856 11693 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 4856 11693 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 4942 11693 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 4942 11693 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 5028 11693 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 5028 11693 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 5114 11693 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 5114 11693 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 5200 11693 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 5200 11693 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 5286 11693 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 5286 11693 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 5372 11693 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 5372 11693 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 5458 11693 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 5458 11693 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 5544 11693 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 5544 11693 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11629 5630 11693 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11629 5630 11693 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 4770 11774 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 4770 11774 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 4856 11774 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 4856 11774 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 4942 11774 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 4942 11774 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 5028 11774 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 5028 11774 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 5114 11774 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 5114 11774 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 5200 11774 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 5200 11774 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 5286 11774 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 5286 11774 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 5372 11774 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 5372 11774 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 5458 11774 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 5458 11774 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 5544 11774 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 5544 11774 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11710 5630 11774 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11710 5630 11774 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 4770 11855 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 4770 11855 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 4856 11855 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 4856 11855 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 4942 11855 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 4942 11855 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 5028 11855 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 5028 11855 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 5114 11855 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 5114 11855 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 5200 11855 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 5200 11855 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 5286 11855 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 5286 11855 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 5372 11855 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 5372 11855 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 5458 11855 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 5458 11855 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 5544 11855 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 5544 11855 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11791 5630 11855 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11791 5630 11855 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 4770 11936 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 4770 11936 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 4856 11936 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 4856 11936 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 4942 11936 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 4942 11936 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 5028 11936 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 5028 11936 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 5114 11936 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 5114 11936 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 5200 11936 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 5200 11936 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 5286 11936 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 5286 11936 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 5372 11936 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 5372 11936 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 5458 11936 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 5458 11936 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 5544 11936 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 5544 11936 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11872 5630 11936 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11872 5630 11936 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 4770 12017 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 4770 12017 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 4856 12017 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 4856 12017 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 4942 12017 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 4942 12017 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 5028 12017 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 5028 12017 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 5114 12017 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 5114 12017 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 5200 12017 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 5200 12017 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 5286 12017 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 5286 12017 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 5372 12017 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 5372 12017 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 5458 12017 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 5458 12017 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 5544 12017 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 5544 12017 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 11953 5630 12017 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 11953 5630 12017 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36289 1295 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36289 1295 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36370 1295 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36370 1295 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36451 1295 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36451 1295 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36532 1295 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36532 1295 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36613 1295 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36613 1295 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36694 1295 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36694 1295 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36775 1295 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36775 1295 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36856 1295 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36856 1295 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 36937 1295 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 36937 1295 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37018 1295 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37018 1295 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37099 1295 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37099 1295 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37180 1295 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37180 1295 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37261 1295 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37261 1295 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37342 1295 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37342 1295 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37423 1295 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37423 1295 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37504 1295 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37504 1295 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37585 1295 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37585 1295 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37666 1295 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37666 1295 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37747 1295 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37747 1295 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37828 1295 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37828 1295 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37909 1295 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37909 1295 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 37990 1295 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 37990 1295 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38071 1295 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38071 1295 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38152 1295 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38152 1295 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38233 1295 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38233 1295 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38314 1295 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38314 1295 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38395 1295 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38395 1295 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38476 1295 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38476 1295 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38557 1295 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38557 1295 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38638 1295 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38638 1295 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38719 1295 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38719 1295 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38800 1295 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38800 1295 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38881 1295 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38881 1295 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 38962 1295 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 38962 1295 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 39043 1295 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 39043 1295 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 39124 1295 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 39124 1295 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 39205 1295 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 39205 1295 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 39286 1295 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 39286 1295 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 39367 1295 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 39367 1295 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 39448 1295 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 39448 1295 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1231 39529 1295 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1231 39529 1295 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 34780 1283 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 34860 1283 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 34940 1283 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35020 1283 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35100 1283 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35180 1283 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35260 1283 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35340 1283 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35420 1283 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35500 1283 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35580 1283 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35660 1283 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35740 1283 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35820 1283 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35900 1283 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 35980 1283 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 36060 1283 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 36140 1283 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1243 36220 1283 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 4770 1310 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 4770 1310 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 4856 1310 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 4856 1310 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 4942 1310 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 4942 1310 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 5028 1310 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 5028 1310 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 5114 1310 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 5114 1310 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 5200 1310 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 5200 1310 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 5286 1310 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 5286 1310 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 5372 1310 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 5372 1310 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 5458 1310 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 5458 1310 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 5544 1310 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 5544 1310 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1246 5630 1310 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1246 5630 1310 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36289 1375 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36289 1375 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36370 1375 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36370 1375 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36451 1375 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36451 1375 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36532 1375 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36532 1375 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36613 1375 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36613 1375 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36694 1375 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36694 1375 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36775 1375 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36775 1375 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36856 1375 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36856 1375 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 36937 1375 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 36937 1375 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37018 1375 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37018 1375 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37099 1375 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37099 1375 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37180 1375 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37180 1375 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37261 1375 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37261 1375 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37342 1375 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37342 1375 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37423 1375 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37423 1375 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37504 1375 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37504 1375 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37585 1375 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37585 1375 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37666 1375 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37666 1375 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37747 1375 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37747 1375 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37828 1375 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37828 1375 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37909 1375 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37909 1375 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 37990 1375 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 37990 1375 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38071 1375 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38071 1375 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38152 1375 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38152 1375 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38233 1375 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38233 1375 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38314 1375 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38314 1375 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38395 1375 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38395 1375 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38476 1375 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38476 1375 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38557 1375 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38557 1375 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38638 1375 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38638 1375 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38719 1375 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38719 1375 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38800 1375 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38800 1375 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38881 1375 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38881 1375 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 38962 1375 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 38962 1375 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 39043 1375 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 39043 1375 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 39124 1375 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 39124 1375 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 39205 1375 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 39205 1375 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 39286 1375 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 39286 1375 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 39367 1375 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 39367 1375 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 39448 1375 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 39448 1375 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1311 39529 1375 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1311 39529 1375 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 34780 1363 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 34860 1363 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 34940 1363 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35020 1363 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35100 1363 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35180 1363 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35260 1363 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35340 1363 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35420 1363 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35500 1363 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35580 1363 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35660 1363 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35740 1363 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35820 1363 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35900 1363 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 35980 1363 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 36060 1363 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 36140 1363 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1323 36220 1363 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 4770 1391 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 4770 1391 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 4856 1391 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 4856 1391 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 4942 1391 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 4942 1391 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 5028 1391 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 5028 1391 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 5114 1391 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 5114 1391 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 5200 1391 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 5200 1391 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 5286 1391 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 5286 1391 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 5372 1391 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 5372 1391 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 5458 1391 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 5458 1391 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 5544 1391 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 5544 1391 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1327 5630 1391 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1327 5630 1391 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36289 1455 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36289 1455 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36370 1455 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36370 1455 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36451 1455 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36451 1455 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36532 1455 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36532 1455 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36613 1455 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36613 1455 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36694 1455 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36694 1455 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36775 1455 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36775 1455 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36856 1455 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36856 1455 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 36937 1455 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 36937 1455 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37018 1455 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37018 1455 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37099 1455 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37099 1455 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37180 1455 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37180 1455 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37261 1455 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37261 1455 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37342 1455 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37342 1455 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37423 1455 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37423 1455 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37504 1455 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37504 1455 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37585 1455 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37585 1455 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37666 1455 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37666 1455 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37747 1455 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37747 1455 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37828 1455 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37828 1455 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37909 1455 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37909 1455 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 37990 1455 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 37990 1455 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38071 1455 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38071 1455 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38152 1455 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38152 1455 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38233 1455 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38233 1455 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38314 1455 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38314 1455 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38395 1455 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38395 1455 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38476 1455 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38476 1455 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38557 1455 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38557 1455 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38638 1455 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38638 1455 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38719 1455 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38719 1455 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38800 1455 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38800 1455 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38881 1455 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38881 1455 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 38962 1455 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 38962 1455 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 39043 1455 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 39043 1455 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 39124 1455 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 39124 1455 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 39205 1455 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 39205 1455 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 39286 1455 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 39286 1455 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 39367 1455 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 39367 1455 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 39448 1455 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 39448 1455 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1391 39529 1455 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1391 39529 1455 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 4770 12098 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 4770 12098 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 4856 12098 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 4856 12098 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 4942 12098 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 4942 12098 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 5028 12098 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 5028 12098 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 5114 12098 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 5114 12098 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 5200 12098 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 5200 12098 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 5286 12098 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 5286 12098 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 5372 12098 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 5372 12098 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 5458 12098 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 5458 12098 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 5544 12098 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 5544 12098 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12034 5630 12098 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12034 5630 12098 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 4770 12179 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 4770 12179 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 4856 12179 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 4856 12179 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 4942 12179 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 4942 12179 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 5028 12179 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 5028 12179 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 5114 12179 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 5114 12179 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 5200 12179 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 5200 12179 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 5286 12179 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 5286 12179 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 5372 12179 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 5372 12179 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 5458 12179 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 5458 12179 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 5544 12179 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 5544 12179 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12115 5630 12179 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12115 5630 12179 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 4770 12260 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 4770 12260 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 4856 12260 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 4856 12260 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 4942 12260 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 4942 12260 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 5028 12260 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 5028 12260 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 5114 12260 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 5114 12260 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 5200 12260 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 5200 12260 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 5286 12260 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 5286 12260 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 5372 12260 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 5372 12260 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 5458 12260 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 5458 12260 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 5544 12260 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 5544 12260 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12196 5630 12260 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12196 5630 12260 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 4770 12341 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 4770 12341 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 4856 12341 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 4856 12341 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 4942 12341 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 4942 12341 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 5028 12341 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 5028 12341 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 5114 12341 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 5114 12341 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 5200 12341 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 5200 12341 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 5286 12341 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 5286 12341 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 5372 12341 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 5372 12341 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 5458 12341 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 5458 12341 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 5544 12341 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 5544 12341 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12277 5630 12341 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12277 5630 12341 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 4770 12422 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 4770 12422 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 4856 12422 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 4856 12422 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 4942 12422 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 4942 12422 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 5028 12422 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 5028 12422 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 5114 12422 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 5114 12422 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 5200 12422 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 5200 12422 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 5286 12422 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 5286 12422 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 5372 12422 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 5372 12422 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 5458 12422 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 5458 12422 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 5544 12422 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 5544 12422 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12358 5630 12422 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12358 5630 12422 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 34768 12480 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 34768 12480 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 34848 12480 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 34848 12480 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 34928 12480 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 34928 12480 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35008 12480 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35008 12480 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35088 12480 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35088 12480 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35168 12480 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35168 12480 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35248 12480 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35248 12480 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35328 12480 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35328 12480 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35408 12480 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35408 12480 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35488 12480 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35488 12480 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35568 12480 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35568 12480 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35648 12480 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35648 12480 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35728 12480 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35728 12480 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35808 12480 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35808 12480 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35888 12480 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35888 12480 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 35968 12480 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 35968 12480 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36048 12480 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36048 12480 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36128 12480 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36128 12480 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36208 12480 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36208 12480 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36289 12480 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36289 12480 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36370 12480 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36370 12480 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36451 12480 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36451 12480 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36532 12480 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36532 12480 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36613 12480 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36613 12480 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36694 12480 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36694 12480 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36775 12480 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36775 12480 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36856 12480 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36856 12480 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 36937 12480 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 36937 12480 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37018 12480 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37018 12480 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37099 12480 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37099 12480 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37180 12480 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37180 12480 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37261 12480 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37261 12480 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37342 12480 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37342 12480 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37423 12480 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37423 12480 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37504 12480 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37504 12480 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37585 12480 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37585 12480 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37666 12480 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37666 12480 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37747 12480 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37747 12480 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37828 12480 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37828 12480 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37909 12480 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37909 12480 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 37990 12480 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 37990 12480 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38071 12480 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38071 12480 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38152 12480 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38152 12480 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38233 12480 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38233 12480 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38314 12480 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38314 12480 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38395 12480 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38395 12480 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38476 12480 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38476 12480 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38557 12480 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38557 12480 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38638 12480 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38638 12480 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38719 12480 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38719 12480 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38800 12480 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38800 12480 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38881 12480 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38881 12480 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 38962 12480 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 38962 12480 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 39043 12480 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 39043 12480 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 39124 12480 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 39124 12480 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 39205 12480 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 39205 12480 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 39286 12480 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 39286 12480 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 39367 12480 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 39367 12480 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 39448 12480 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 39448 12480 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12416 39529 12480 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12416 39529 12480 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 4770 12503 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 4770 12503 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 4856 12503 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 4856 12503 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 4942 12503 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 4942 12503 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 5028 12503 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 5028 12503 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 5114 12503 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 5114 12503 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 5200 12503 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 5200 12503 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 5286 12503 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 5286 12503 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 5372 12503 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 5372 12503 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 5458 12503 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 5458 12503 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 5544 12503 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 5544 12503 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12439 5630 12503 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12439 5630 12503 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 34768 12562 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 34768 12562 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 34848 12562 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 34848 12562 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 34928 12562 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 34928 12562 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35008 12562 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35008 12562 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35088 12562 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35088 12562 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35168 12562 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35168 12562 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35248 12562 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35248 12562 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35328 12562 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35328 12562 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35408 12562 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35408 12562 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35488 12562 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35488 12562 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35568 12562 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35568 12562 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35648 12562 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35648 12562 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35728 12562 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35728 12562 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35808 12562 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35808 12562 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35888 12562 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35888 12562 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 35968 12562 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 35968 12562 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36048 12562 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36048 12562 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36128 12562 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36128 12562 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36208 12562 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36208 12562 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36289 12562 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36289 12562 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36370 12562 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36370 12562 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36451 12562 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36451 12562 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36532 12562 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36532 12562 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36613 12562 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36613 12562 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36694 12562 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36694 12562 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36775 12562 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36775 12562 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36856 12562 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36856 12562 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 36937 12562 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 36937 12562 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37018 12562 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37018 12562 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37099 12562 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37099 12562 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37180 12562 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37180 12562 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37261 12562 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37261 12562 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37342 12562 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37342 12562 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37423 12562 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37423 12562 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37504 12562 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37504 12562 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37585 12562 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37585 12562 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37666 12562 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37666 12562 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37747 12562 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37747 12562 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37828 12562 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37828 12562 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37909 12562 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37909 12562 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 37990 12562 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 37990 12562 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38071 12562 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38071 12562 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38152 12562 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38152 12562 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38233 12562 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38233 12562 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38314 12562 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38314 12562 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38395 12562 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38395 12562 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38476 12562 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38476 12562 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38557 12562 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38557 12562 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38638 12562 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38638 12562 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38719 12562 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38719 12562 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38800 12562 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38800 12562 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38881 12562 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38881 12562 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 38962 12562 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 38962 12562 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 39043 12562 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 39043 12562 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 39124 12562 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 39124 12562 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 39205 12562 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 39205 12562 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 39286 12562 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 39286 12562 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 39367 12562 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 39367 12562 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 39448 12562 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 39448 12562 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12498 39529 12562 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12498 39529 12562 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 4770 12584 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 4770 12584 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 4856 12584 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 4856 12584 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 4942 12584 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 4942 12584 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 5028 12584 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 5028 12584 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 5114 12584 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 5114 12584 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 5200 12584 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 5200 12584 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 5286 12584 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 5286 12584 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 5372 12584 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 5372 12584 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 5458 12584 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 5458 12584 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 5544 12584 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 5544 12584 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12520 5630 12584 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12520 5630 12584 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 34768 12644 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 34768 12644 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 34848 12644 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 34848 12644 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 34928 12644 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 34928 12644 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35008 12644 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35008 12644 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35088 12644 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35088 12644 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35168 12644 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35168 12644 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35248 12644 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35248 12644 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35328 12644 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35328 12644 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35408 12644 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35408 12644 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35488 12644 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35488 12644 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35568 12644 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35568 12644 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35648 12644 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35648 12644 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35728 12644 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35728 12644 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35808 12644 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35808 12644 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35888 12644 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35888 12644 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 35968 12644 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 35968 12644 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36048 12644 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36048 12644 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36128 12644 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36128 12644 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36208 12644 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36208 12644 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36289 12644 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36289 12644 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36370 12644 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36370 12644 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36451 12644 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36451 12644 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36532 12644 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36532 12644 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36613 12644 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36613 12644 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36694 12644 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36694 12644 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36775 12644 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36775 12644 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36856 12644 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36856 12644 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 36937 12644 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 36937 12644 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37018 12644 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37018 12644 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37099 12644 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37099 12644 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37180 12644 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37180 12644 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37261 12644 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37261 12644 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37342 12644 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37342 12644 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37423 12644 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37423 12644 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37504 12644 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37504 12644 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37585 12644 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37585 12644 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37666 12644 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37666 12644 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37747 12644 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37747 12644 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37828 12644 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37828 12644 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37909 12644 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37909 12644 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 37990 12644 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 37990 12644 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38071 12644 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38071 12644 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38152 12644 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38152 12644 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38233 12644 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38233 12644 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38314 12644 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38314 12644 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38395 12644 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38395 12644 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38476 12644 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38476 12644 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38557 12644 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38557 12644 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38638 12644 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38638 12644 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38719 12644 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38719 12644 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38800 12644 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38800 12644 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38881 12644 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38881 12644 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 38962 12644 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 38962 12644 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 39043 12644 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 39043 12644 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 39124 12644 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 39124 12644 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 39205 12644 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 39205 12644 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 39286 12644 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 39286 12644 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 39367 12644 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 39367 12644 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 39448 12644 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 39448 12644 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12580 39529 12644 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12580 39529 12644 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 4770 12665 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 4770 12665 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 4856 12665 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 4856 12665 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 4942 12665 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 4942 12665 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 5028 12665 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 5028 12665 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 5114 12665 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 5114 12665 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 5200 12665 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 5200 12665 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 5286 12665 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 5286 12665 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 5372 12665 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 5372 12665 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 5458 12665 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 5458 12665 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 5544 12665 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 5544 12665 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12601 5630 12665 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12601 5630 12665 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 34768 12726 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 34768 12726 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 34848 12726 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 34848 12726 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 34928 12726 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 34928 12726 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35008 12726 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35008 12726 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35088 12726 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35088 12726 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35168 12726 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35168 12726 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35248 12726 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35248 12726 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35328 12726 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35328 12726 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35408 12726 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35408 12726 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35488 12726 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35488 12726 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35568 12726 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35568 12726 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35648 12726 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35648 12726 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35728 12726 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35728 12726 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35808 12726 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35808 12726 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35888 12726 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35888 12726 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 35968 12726 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 35968 12726 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36048 12726 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36048 12726 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36128 12726 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36128 12726 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36208 12726 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36208 12726 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36289 12726 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36289 12726 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36370 12726 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36370 12726 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36451 12726 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36451 12726 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36532 12726 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36532 12726 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36613 12726 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36613 12726 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36694 12726 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36694 12726 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36775 12726 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36775 12726 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36856 12726 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36856 12726 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 36937 12726 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 36937 12726 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37018 12726 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37018 12726 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37099 12726 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37099 12726 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37180 12726 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37180 12726 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37261 12726 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37261 12726 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37342 12726 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37342 12726 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37423 12726 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37423 12726 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37504 12726 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37504 12726 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37585 12726 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37585 12726 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37666 12726 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37666 12726 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37747 12726 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37747 12726 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37828 12726 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37828 12726 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37909 12726 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37909 12726 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 37990 12726 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 37990 12726 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38071 12726 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38071 12726 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38152 12726 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38152 12726 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38233 12726 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38233 12726 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38314 12726 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38314 12726 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38395 12726 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38395 12726 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38476 12726 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38476 12726 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38557 12726 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38557 12726 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38638 12726 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38638 12726 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38719 12726 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38719 12726 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38800 12726 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38800 12726 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38881 12726 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38881 12726 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 38962 12726 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 38962 12726 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 39043 12726 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 39043 12726 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 39124 12726 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 39124 12726 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 39205 12726 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 39205 12726 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 39286 12726 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 39286 12726 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 39367 12726 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 39367 12726 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 39448 12726 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 39448 12726 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12662 39529 12726 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12662 39529 12726 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 4770 12746 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 4770 12746 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 4856 12746 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 4856 12746 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 4942 12746 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 4942 12746 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 5028 12746 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 5028 12746 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 5114 12746 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 5114 12746 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 5200 12746 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 5200 12746 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 5286 12746 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 5286 12746 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 5372 12746 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 5372 12746 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 5458 12746 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 5458 12746 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 5544 12746 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 5544 12746 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12682 5630 12746 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12682 5630 12746 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 34768 12808 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 34768 12808 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 34848 12808 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 34848 12808 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 34928 12808 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 34928 12808 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35008 12808 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35008 12808 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35088 12808 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35088 12808 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35168 12808 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35168 12808 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35248 12808 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35248 12808 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35328 12808 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35328 12808 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35408 12808 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35408 12808 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35488 12808 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35488 12808 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35568 12808 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35568 12808 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35648 12808 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35648 12808 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35728 12808 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35728 12808 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35808 12808 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35808 12808 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35888 12808 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35888 12808 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 35968 12808 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 35968 12808 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36048 12808 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36048 12808 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36128 12808 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36128 12808 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36208 12808 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36208 12808 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36289 12808 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36289 12808 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36370 12808 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36370 12808 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36451 12808 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36451 12808 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36532 12808 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36532 12808 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36613 12808 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36613 12808 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36694 12808 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36694 12808 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36775 12808 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36775 12808 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36856 12808 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36856 12808 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 36937 12808 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 36937 12808 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37018 12808 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37018 12808 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37099 12808 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37099 12808 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37180 12808 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37180 12808 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37261 12808 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37261 12808 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37342 12808 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37342 12808 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37423 12808 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37423 12808 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37504 12808 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37504 12808 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37585 12808 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37585 12808 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37666 12808 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37666 12808 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37747 12808 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37747 12808 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37828 12808 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37828 12808 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37909 12808 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37909 12808 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 37990 12808 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 37990 12808 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38071 12808 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38071 12808 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38152 12808 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38152 12808 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38233 12808 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38233 12808 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38314 12808 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38314 12808 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38395 12808 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38395 12808 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38476 12808 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38476 12808 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38557 12808 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38557 12808 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38638 12808 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38638 12808 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38719 12808 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38719 12808 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38800 12808 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38800 12808 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38881 12808 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38881 12808 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 38962 12808 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 38962 12808 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 39043 12808 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 39043 12808 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 39124 12808 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 39124 12808 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 39205 12808 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 39205 12808 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 39286 12808 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 39286 12808 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 39367 12808 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 39367 12808 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 39448 12808 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 39448 12808 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12744 39529 12808 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12744 39529 12808 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 4770 12827 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 4770 12827 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 4856 12827 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 4856 12827 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 4942 12827 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 4942 12827 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 5028 12827 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 5028 12827 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 5114 12827 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 5114 12827 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 5200 12827 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 5200 12827 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 5286 12827 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 5286 12827 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 5372 12827 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 5372 12827 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 5458 12827 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 5458 12827 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 5544 12827 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 5544 12827 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12763 5630 12827 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12763 5630 12827 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 34768 12890 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 34768 12890 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 34848 12890 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 34848 12890 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 34928 12890 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 34928 12890 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35008 12890 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35008 12890 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35088 12890 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35088 12890 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35168 12890 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35168 12890 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35248 12890 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35248 12890 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35328 12890 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35328 12890 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35408 12890 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35408 12890 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35488 12890 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35488 12890 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35568 12890 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35568 12890 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35648 12890 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35648 12890 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35728 12890 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35728 12890 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35808 12890 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35808 12890 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35888 12890 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35888 12890 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 35968 12890 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 35968 12890 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36048 12890 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36048 12890 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36128 12890 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36128 12890 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36208 12890 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36208 12890 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36289 12890 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36289 12890 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36370 12890 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36370 12890 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36451 12890 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36451 12890 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36532 12890 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36532 12890 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36613 12890 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36613 12890 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36694 12890 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36694 12890 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36775 12890 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36775 12890 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36856 12890 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36856 12890 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 36937 12890 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 36937 12890 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37018 12890 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37018 12890 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37099 12890 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37099 12890 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37180 12890 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37180 12890 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37261 12890 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37261 12890 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37342 12890 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37342 12890 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37423 12890 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37423 12890 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37504 12890 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37504 12890 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37585 12890 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37585 12890 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37666 12890 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37666 12890 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37747 12890 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37747 12890 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37828 12890 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37828 12890 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37909 12890 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37909 12890 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 37990 12890 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 37990 12890 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38071 12890 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38071 12890 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38152 12890 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38152 12890 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38233 12890 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38233 12890 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38314 12890 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38314 12890 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38395 12890 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38395 12890 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38476 12890 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38476 12890 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38557 12890 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38557 12890 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38638 12890 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38638 12890 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38719 12890 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38719 12890 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38800 12890 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38800 12890 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38881 12890 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38881 12890 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 38962 12890 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 38962 12890 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 39043 12890 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 39043 12890 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 39124 12890 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 39124 12890 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 39205 12890 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 39205 12890 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 39286 12890 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 39286 12890 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 39367 12890 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 39367 12890 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 39448 12890 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 39448 12890 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12826 39529 12890 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12826 39529 12890 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 4770 12908 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 4770 12908 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 4856 12908 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 4856 12908 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 4942 12908 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 4942 12908 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 5028 12908 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 5028 12908 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 5114 12908 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 5114 12908 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 5200 12908 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 5200 12908 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 5286 12908 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 5286 12908 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 5372 12908 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 5372 12908 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 5458 12908 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 5458 12908 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 5544 12908 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 5544 12908 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12844 5630 12908 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12844 5630 12908 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 34768 12972 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 34768 12972 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 34848 12972 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 34848 12972 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 34928 12972 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 34928 12972 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35008 12972 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35008 12972 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35088 12972 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35088 12972 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35168 12972 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35168 12972 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35248 12972 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35248 12972 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35328 12972 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35328 12972 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35408 12972 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35408 12972 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35488 12972 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35488 12972 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35568 12972 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35568 12972 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35648 12972 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35648 12972 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35728 12972 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35728 12972 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35808 12972 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35808 12972 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35888 12972 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35888 12972 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 35968 12972 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 35968 12972 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36048 12972 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36048 12972 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36128 12972 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36128 12972 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36208 12972 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36208 12972 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36289 12972 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36289 12972 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36370 12972 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36370 12972 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36451 12972 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36451 12972 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36532 12972 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36532 12972 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36613 12972 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36613 12972 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36694 12972 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36694 12972 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36775 12972 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36775 12972 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36856 12972 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36856 12972 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 36937 12972 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 36937 12972 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37018 12972 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37018 12972 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37099 12972 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37099 12972 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37180 12972 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37180 12972 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37261 12972 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37261 12972 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37342 12972 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37342 12972 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37423 12972 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37423 12972 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37504 12972 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37504 12972 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37585 12972 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37585 12972 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37666 12972 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37666 12972 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37747 12972 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37747 12972 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37828 12972 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37828 12972 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37909 12972 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37909 12972 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 37990 12972 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 37990 12972 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38071 12972 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38071 12972 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38152 12972 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38152 12972 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38233 12972 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38233 12972 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38314 12972 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38314 12972 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38395 12972 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38395 12972 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38476 12972 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38476 12972 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38557 12972 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38557 12972 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38638 12972 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38638 12972 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38719 12972 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38719 12972 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38800 12972 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38800 12972 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38881 12972 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38881 12972 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 38962 12972 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 38962 12972 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 39043 12972 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 39043 12972 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 39124 12972 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 39124 12972 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 39205 12972 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 39205 12972 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 39286 12972 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 39286 12972 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 39367 12972 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 39367 12972 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 39448 12972 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 39448 12972 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12908 39529 12972 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12908 39529 12972 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 4770 12989 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 4770 12989 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 4856 12989 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 4856 12989 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 4942 12989 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 4942 12989 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 5028 12989 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 5028 12989 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 5114 12989 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 5114 12989 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 5200 12989 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 5200 12989 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 5286 12989 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 5286 12989 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 5372 12989 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 5372 12989 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 5458 12989 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 5458 12989 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 5544 12989 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 5544 12989 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12925 5630 12989 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12925 5630 12989 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 34768 13054 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 34768 13054 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 34848 13054 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 34848 13054 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 34928 13054 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 34928 13054 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35008 13054 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35008 13054 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35088 13054 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35088 13054 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35168 13054 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35168 13054 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35248 13054 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35248 13054 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35328 13054 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35328 13054 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35408 13054 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35408 13054 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35488 13054 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35488 13054 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35568 13054 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35568 13054 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35648 13054 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35648 13054 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35728 13054 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35728 13054 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35808 13054 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35808 13054 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35888 13054 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35888 13054 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 35968 13054 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 35968 13054 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36048 13054 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36048 13054 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36128 13054 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36128 13054 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36208 13054 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36208 13054 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36289 13054 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36289 13054 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36370 13054 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36370 13054 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36451 13054 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36451 13054 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36532 13054 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36532 13054 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36613 13054 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36613 13054 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36694 13054 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36694 13054 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36775 13054 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36775 13054 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36856 13054 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36856 13054 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 36937 13054 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 36937 13054 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37018 13054 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37018 13054 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37099 13054 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37099 13054 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37180 13054 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37180 13054 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37261 13054 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37261 13054 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37342 13054 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37342 13054 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37423 13054 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37423 13054 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37504 13054 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37504 13054 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37585 13054 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37585 13054 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37666 13054 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37666 13054 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37747 13054 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37747 13054 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37828 13054 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37828 13054 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37909 13054 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37909 13054 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 37990 13054 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 37990 13054 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38071 13054 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38071 13054 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38152 13054 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38152 13054 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38233 13054 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38233 13054 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38314 13054 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38314 13054 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38395 13054 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38395 13054 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38476 13054 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38476 13054 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38557 13054 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38557 13054 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38638 13054 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38638 13054 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38719 13054 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38719 13054 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38800 13054 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38800 13054 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38881 13054 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38881 13054 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 38962 13054 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 38962 13054 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 39043 13054 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 39043 13054 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 39124 13054 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 39124 13054 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 39205 13054 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 39205 13054 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 39286 13054 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 39286 13054 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 39367 13054 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 39367 13054 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 39448 13054 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 39448 13054 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 12990 39529 13054 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 12990 39529 13054 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 4770 13070 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 4770 13070 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 4856 13070 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 4856 13070 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 4942 13070 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 4942 13070 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 5028 13070 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 5028 13070 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 5114 13070 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 5114 13070 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 5200 13070 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 5200 13070 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 5286 13070 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 5286 13070 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 5372 13070 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 5372 13070 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 5458 13070 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 5458 13070 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 5544 13070 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 5544 13070 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13006 5630 13070 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13006 5630 13070 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 34768 13136 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 34768 13136 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 34848 13136 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 34848 13136 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 34928 13136 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 34928 13136 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35008 13136 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35008 13136 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35088 13136 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35088 13136 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35168 13136 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35168 13136 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35248 13136 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35248 13136 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35328 13136 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35328 13136 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35408 13136 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35408 13136 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35488 13136 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35488 13136 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35568 13136 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35568 13136 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35648 13136 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35648 13136 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35728 13136 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35728 13136 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35808 13136 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35808 13136 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35888 13136 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35888 13136 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 35968 13136 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 35968 13136 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36048 13136 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36048 13136 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36128 13136 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36128 13136 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36208 13136 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36208 13136 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36289 13136 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36289 13136 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36370 13136 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36370 13136 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36451 13136 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36451 13136 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36532 13136 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36532 13136 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36613 13136 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36613 13136 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36694 13136 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36694 13136 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36775 13136 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36775 13136 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36856 13136 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36856 13136 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 36937 13136 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 36937 13136 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37018 13136 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37018 13136 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37099 13136 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37099 13136 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37180 13136 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37180 13136 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37261 13136 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37261 13136 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37342 13136 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37342 13136 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37423 13136 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37423 13136 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37504 13136 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37504 13136 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37585 13136 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37585 13136 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37666 13136 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37666 13136 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37747 13136 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37747 13136 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37828 13136 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37828 13136 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37909 13136 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37909 13136 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 37990 13136 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 37990 13136 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38071 13136 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38071 13136 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38152 13136 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38152 13136 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38233 13136 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38233 13136 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38314 13136 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38314 13136 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38395 13136 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38395 13136 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38476 13136 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38476 13136 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38557 13136 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38557 13136 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38638 13136 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38638 13136 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38719 13136 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38719 13136 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38800 13136 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38800 13136 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38881 13136 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38881 13136 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 38962 13136 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 38962 13136 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 39043 13136 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 39043 13136 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 39124 13136 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 39124 13136 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 39205 13136 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 39205 13136 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 39286 13136 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 39286 13136 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 39367 13136 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 39367 13136 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 39448 13136 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 39448 13136 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13072 39529 13136 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13072 39529 13136 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 4770 13151 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 4770 13151 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 4856 13151 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 4856 13151 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 4942 13151 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 4942 13151 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 5028 13151 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 5028 13151 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 5114 13151 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 5114 13151 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 5200 13151 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 5200 13151 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 5286 13151 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 5286 13151 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 5372 13151 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 5372 13151 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 5458 13151 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 5458 13151 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 5544 13151 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 5544 13151 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13087 5630 13151 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13087 5630 13151 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 34768 13218 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 34768 13218 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 34848 13218 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 34848 13218 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 34928 13218 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 34928 13218 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35008 13218 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35008 13218 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35088 13218 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35088 13218 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35168 13218 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35168 13218 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35248 13218 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35248 13218 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35328 13218 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35328 13218 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35408 13218 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35408 13218 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35488 13218 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35488 13218 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35568 13218 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35568 13218 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35648 13218 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35648 13218 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35728 13218 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35728 13218 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35808 13218 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35808 13218 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35888 13218 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35888 13218 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 35968 13218 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 35968 13218 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36048 13218 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36048 13218 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36128 13218 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36128 13218 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36208 13218 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36208 13218 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36289 13218 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36289 13218 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36370 13218 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36370 13218 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36451 13218 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36451 13218 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36532 13218 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36532 13218 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36613 13218 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36613 13218 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36694 13218 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36694 13218 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36775 13218 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36775 13218 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36856 13218 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36856 13218 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 36937 13218 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 36937 13218 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37018 13218 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37018 13218 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37099 13218 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37099 13218 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37180 13218 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37180 13218 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37261 13218 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37261 13218 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37342 13218 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37342 13218 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37423 13218 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37423 13218 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37504 13218 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37504 13218 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37585 13218 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37585 13218 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37666 13218 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37666 13218 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37747 13218 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37747 13218 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37828 13218 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37828 13218 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37909 13218 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37909 13218 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 37990 13218 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 37990 13218 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38071 13218 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38071 13218 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38152 13218 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38152 13218 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38233 13218 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38233 13218 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38314 13218 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38314 13218 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38395 13218 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38395 13218 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38476 13218 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38476 13218 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38557 13218 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38557 13218 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38638 13218 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38638 13218 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38719 13218 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38719 13218 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38800 13218 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38800 13218 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38881 13218 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38881 13218 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 38962 13218 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 38962 13218 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 39043 13218 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 39043 13218 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 39124 13218 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 39124 13218 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 39205 13218 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 39205 13218 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 39286 13218 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 39286 13218 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 39367 13218 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 39367 13218 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 39448 13218 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 39448 13218 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13154 39529 13218 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13154 39529 13218 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 4770 13232 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 4770 13232 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 4856 13232 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 4856 13232 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 4942 13232 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 4942 13232 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 5028 13232 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 5028 13232 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 5114 13232 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 5114 13232 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 5200 13232 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 5200 13232 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 5286 13232 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 5286 13232 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 5372 13232 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 5372 13232 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 5458 13232 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 5458 13232 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 5544 13232 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 5544 13232 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13168 5630 13232 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13168 5630 13232 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 34768 13300 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 34768 13300 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 34848 13300 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 34848 13300 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 34928 13300 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 34928 13300 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35008 13300 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35008 13300 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35088 13300 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35088 13300 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35168 13300 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35168 13300 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35248 13300 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35248 13300 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35328 13300 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35328 13300 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35408 13300 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35408 13300 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35488 13300 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35488 13300 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35568 13300 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35568 13300 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35648 13300 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35648 13300 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35728 13300 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35728 13300 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35808 13300 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35808 13300 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35888 13300 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35888 13300 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 35968 13300 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 35968 13300 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36048 13300 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36048 13300 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36128 13300 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36128 13300 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36208 13300 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36208 13300 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36289 13300 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36289 13300 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36370 13300 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36370 13300 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36451 13300 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36451 13300 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36532 13300 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36532 13300 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36613 13300 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36613 13300 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36694 13300 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36694 13300 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36775 13300 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36775 13300 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36856 13300 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36856 13300 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 36937 13300 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 36937 13300 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37018 13300 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37018 13300 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37099 13300 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37099 13300 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37180 13300 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37180 13300 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37261 13300 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37261 13300 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37342 13300 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37342 13300 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37423 13300 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37423 13300 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37504 13300 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37504 13300 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37585 13300 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37585 13300 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37666 13300 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37666 13300 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37747 13300 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37747 13300 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37828 13300 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37828 13300 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37909 13300 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37909 13300 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 37990 13300 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 37990 13300 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38071 13300 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38071 13300 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38152 13300 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38152 13300 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38233 13300 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38233 13300 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38314 13300 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38314 13300 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38395 13300 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38395 13300 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38476 13300 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38476 13300 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38557 13300 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38557 13300 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38638 13300 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38638 13300 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38719 13300 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38719 13300 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38800 13300 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38800 13300 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38881 13300 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38881 13300 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 38962 13300 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 38962 13300 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 39043 13300 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 39043 13300 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 39124 13300 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 39124 13300 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 39205 13300 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 39205 13300 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 39286 13300 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 39286 13300 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 39367 13300 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 39367 13300 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 39448 13300 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 39448 13300 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13236 39529 13300 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13236 39529 13300 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 4770 13313 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 4770 13313 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 4856 13313 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 4856 13313 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 4942 13313 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 4942 13313 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 5028 13313 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 5028 13313 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 5114 13313 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 5114 13313 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 5200 13313 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 5200 13313 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 5286 13313 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 5286 13313 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 5372 13313 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 5372 13313 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 5458 13313 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 5458 13313 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 5544 13313 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 5544 13313 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13249 5630 13313 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13249 5630 13313 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 34768 13382 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 34768 13382 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 34848 13382 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 34848 13382 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 34928 13382 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 34928 13382 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35008 13382 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35008 13382 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35088 13382 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35088 13382 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35168 13382 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35168 13382 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35248 13382 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35248 13382 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35328 13382 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35328 13382 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35408 13382 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35408 13382 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35488 13382 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35488 13382 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35568 13382 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35568 13382 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35648 13382 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35648 13382 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35728 13382 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35728 13382 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35808 13382 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35808 13382 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35888 13382 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35888 13382 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 35968 13382 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 35968 13382 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36048 13382 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36048 13382 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36128 13382 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36128 13382 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36208 13382 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36208 13382 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36289 13382 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36289 13382 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36370 13382 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36370 13382 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36451 13382 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36451 13382 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36532 13382 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36532 13382 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36613 13382 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36613 13382 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36694 13382 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36694 13382 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36775 13382 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36775 13382 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36856 13382 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36856 13382 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 36937 13382 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 36937 13382 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37018 13382 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37018 13382 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37099 13382 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37099 13382 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37180 13382 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37180 13382 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37261 13382 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37261 13382 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37342 13382 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37342 13382 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37423 13382 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37423 13382 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37504 13382 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37504 13382 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37585 13382 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37585 13382 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37666 13382 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37666 13382 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37747 13382 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37747 13382 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37828 13382 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37828 13382 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37909 13382 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37909 13382 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 37990 13382 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 37990 13382 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38071 13382 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38071 13382 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38152 13382 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38152 13382 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38233 13382 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38233 13382 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38314 13382 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38314 13382 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38395 13382 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38395 13382 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38476 13382 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38476 13382 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38557 13382 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38557 13382 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38638 13382 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38638 13382 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38719 13382 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38719 13382 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38800 13382 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38800 13382 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38881 13382 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38881 13382 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 38962 13382 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 38962 13382 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 39043 13382 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 39043 13382 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 39124 13382 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 39124 13382 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 39205 13382 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 39205 13382 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 39286 13382 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 39286 13382 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 39367 13382 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 39367 13382 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 39448 13382 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 39448 13382 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13318 39529 13382 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13318 39529 13382 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 4770 13394 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 4770 13394 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 4856 13394 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 4856 13394 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 4942 13394 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 4942 13394 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 5028 13394 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 5028 13394 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 5114 13394 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 5114 13394 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 5200 13394 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 5200 13394 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 5286 13394 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 5286 13394 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 5372 13394 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 5372 13394 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 5458 13394 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 5458 13394 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 5544 13394 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 5544 13394 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13330 5630 13394 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13330 5630 13394 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 34768 13464 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 34768 13464 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 34848 13464 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 34848 13464 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 34928 13464 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 34928 13464 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35008 13464 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35008 13464 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35088 13464 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35088 13464 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35168 13464 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35168 13464 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35248 13464 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35248 13464 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35328 13464 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35328 13464 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35408 13464 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35408 13464 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35488 13464 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35488 13464 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35568 13464 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35568 13464 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35648 13464 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35648 13464 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35728 13464 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35728 13464 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35808 13464 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35808 13464 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35888 13464 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35888 13464 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 35968 13464 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 35968 13464 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36048 13464 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36048 13464 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36128 13464 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36128 13464 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36208 13464 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36208 13464 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36289 13464 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36289 13464 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36370 13464 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36370 13464 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36451 13464 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36451 13464 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36532 13464 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36532 13464 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36613 13464 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36613 13464 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36694 13464 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36694 13464 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36775 13464 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36775 13464 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36856 13464 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36856 13464 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 36937 13464 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 36937 13464 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37018 13464 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37018 13464 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37099 13464 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37099 13464 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37180 13464 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37180 13464 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37261 13464 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37261 13464 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37342 13464 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37342 13464 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37423 13464 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37423 13464 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37504 13464 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37504 13464 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37585 13464 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37585 13464 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37666 13464 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37666 13464 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37747 13464 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37747 13464 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37828 13464 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37828 13464 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37909 13464 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37909 13464 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 37990 13464 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 37990 13464 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38071 13464 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38071 13464 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38152 13464 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38152 13464 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38233 13464 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38233 13464 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38314 13464 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38314 13464 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38395 13464 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38395 13464 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38476 13464 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38476 13464 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38557 13464 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38557 13464 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38638 13464 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38638 13464 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38719 13464 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38719 13464 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38800 13464 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38800 13464 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38881 13464 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38881 13464 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 38962 13464 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 38962 13464 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 39043 13464 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 39043 13464 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 39124 13464 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 39124 13464 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 39205 13464 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 39205 13464 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 39286 13464 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 39286 13464 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 39367 13464 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 39367 13464 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 39448 13464 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 39448 13464 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13400 39529 13464 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13400 39529 13464 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 4770 13475 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 4770 13475 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 4856 13475 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 4856 13475 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 4942 13475 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 4942 13475 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 5028 13475 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 5028 13475 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 5114 13475 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 5114 13475 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 5200 13475 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 5200 13475 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 5286 13475 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 5286 13475 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 5372 13475 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 5372 13475 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 5458 13475 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 5458 13475 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 5544 13475 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 5544 13475 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13411 5630 13475 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13411 5630 13475 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 34768 13546 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 34768 13546 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 34848 13546 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 34848 13546 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 34928 13546 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 34928 13546 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35008 13546 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35008 13546 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35088 13546 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35088 13546 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35168 13546 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35168 13546 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35248 13546 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35248 13546 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35328 13546 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35328 13546 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35408 13546 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35408 13546 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35488 13546 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35488 13546 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35568 13546 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35568 13546 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35648 13546 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35648 13546 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35728 13546 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35728 13546 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35808 13546 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35808 13546 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35888 13546 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35888 13546 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 35968 13546 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 35968 13546 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36048 13546 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36048 13546 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36128 13546 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36128 13546 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36208 13546 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36208 13546 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36289 13546 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36289 13546 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36370 13546 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36370 13546 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36451 13546 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36451 13546 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36532 13546 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36532 13546 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36613 13546 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36613 13546 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36694 13546 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36694 13546 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36775 13546 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36775 13546 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36856 13546 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36856 13546 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 36937 13546 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 36937 13546 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37018 13546 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37018 13546 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37099 13546 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37099 13546 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37180 13546 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37180 13546 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37261 13546 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37261 13546 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37342 13546 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37342 13546 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37423 13546 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37423 13546 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37504 13546 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37504 13546 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37585 13546 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37585 13546 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37666 13546 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37666 13546 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37747 13546 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37747 13546 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37828 13546 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37828 13546 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37909 13546 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37909 13546 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 37990 13546 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 37990 13546 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38071 13546 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38071 13546 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38152 13546 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38152 13546 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38233 13546 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38233 13546 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38314 13546 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38314 13546 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38395 13546 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38395 13546 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38476 13546 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38476 13546 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38557 13546 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38557 13546 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38638 13546 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38638 13546 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38719 13546 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38719 13546 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38800 13546 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38800 13546 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38881 13546 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38881 13546 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 38962 13546 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 38962 13546 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 39043 13546 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 39043 13546 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 39124 13546 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 39124 13546 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 39205 13546 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 39205 13546 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 39286 13546 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 39286 13546 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 39367 13546 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 39367 13546 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 39448 13546 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 39448 13546 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13482 39529 13546 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13482 39529 13546 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 4770 13556 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 4770 13556 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 4856 13556 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 4856 13556 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 4942 13556 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 4942 13556 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 5028 13556 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 5028 13556 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 5114 13556 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 5114 13556 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 5200 13556 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 5200 13556 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 5286 13556 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 5286 13556 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 5372 13556 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 5372 13556 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 5458 13556 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 5458 13556 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 5544 13556 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 5544 13556 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13492 5630 13556 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13492 5630 13556 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 34768 13628 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 34768 13628 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 34848 13628 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 34848 13628 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 34928 13628 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 34928 13628 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35008 13628 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35008 13628 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35088 13628 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35088 13628 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35168 13628 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35168 13628 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35248 13628 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35248 13628 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35328 13628 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35328 13628 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35408 13628 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35408 13628 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35488 13628 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35488 13628 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35568 13628 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35568 13628 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35648 13628 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35648 13628 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35728 13628 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35728 13628 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35808 13628 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35808 13628 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35888 13628 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35888 13628 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 35968 13628 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 35968 13628 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36048 13628 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36048 13628 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36128 13628 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36128 13628 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36208 13628 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36208 13628 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36289 13628 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36289 13628 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36370 13628 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36370 13628 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36451 13628 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36451 13628 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36532 13628 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36532 13628 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36613 13628 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36613 13628 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36694 13628 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36694 13628 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36775 13628 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36775 13628 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36856 13628 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36856 13628 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 36937 13628 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 36937 13628 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37018 13628 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37018 13628 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37099 13628 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37099 13628 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37180 13628 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37180 13628 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37261 13628 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37261 13628 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37342 13628 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37342 13628 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37423 13628 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37423 13628 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37504 13628 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37504 13628 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37585 13628 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37585 13628 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37666 13628 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37666 13628 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37747 13628 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37747 13628 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37828 13628 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37828 13628 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37909 13628 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37909 13628 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 37990 13628 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 37990 13628 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38071 13628 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38071 13628 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38152 13628 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38152 13628 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38233 13628 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38233 13628 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38314 13628 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38314 13628 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38395 13628 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38395 13628 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38476 13628 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38476 13628 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38557 13628 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38557 13628 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38638 13628 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38638 13628 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38719 13628 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38719 13628 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38800 13628 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38800 13628 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38881 13628 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38881 13628 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 38962 13628 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 38962 13628 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 39043 13628 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 39043 13628 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 39124 13628 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 39124 13628 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 39205 13628 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 39205 13628 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 39286 13628 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 39286 13628 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 39367 13628 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 39367 13628 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 39448 13628 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 39448 13628 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13564 39529 13628 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13564 39529 13628 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 4770 13637 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 4770 13637 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 4856 13637 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 4856 13637 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 4942 13637 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 4942 13637 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 5028 13637 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 5028 13637 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 5114 13637 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 5114 13637 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 5200 13637 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 5200 13637 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 5286 13637 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 5286 13637 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 5372 13637 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 5372 13637 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 5458 13637 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 5458 13637 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 5544 13637 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 5544 13637 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13573 5630 13637 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13573 5630 13637 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 34768 13710 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 34768 13710 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 34848 13710 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 34848 13710 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 34928 13710 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 34928 13710 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35008 13710 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35008 13710 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35088 13710 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35088 13710 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35168 13710 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35168 13710 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35248 13710 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35248 13710 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35328 13710 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35328 13710 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35408 13710 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35408 13710 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35488 13710 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35488 13710 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35568 13710 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35568 13710 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35648 13710 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35648 13710 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35728 13710 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35728 13710 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35808 13710 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35808 13710 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35888 13710 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35888 13710 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 35968 13710 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 35968 13710 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36048 13710 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36048 13710 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36128 13710 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36128 13710 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36208 13710 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36208 13710 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36289 13710 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36289 13710 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36370 13710 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36370 13710 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36451 13710 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36451 13710 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36532 13710 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36532 13710 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36613 13710 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36613 13710 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36694 13710 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36694 13710 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36775 13710 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36775 13710 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36856 13710 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36856 13710 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 36937 13710 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 36937 13710 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37018 13710 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37018 13710 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37099 13710 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37099 13710 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37180 13710 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37180 13710 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37261 13710 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37261 13710 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37342 13710 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37342 13710 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37423 13710 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37423 13710 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37504 13710 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37504 13710 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37585 13710 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37585 13710 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37666 13710 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37666 13710 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37747 13710 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37747 13710 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37828 13710 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37828 13710 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37909 13710 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37909 13710 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 37990 13710 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 37990 13710 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38071 13710 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38071 13710 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38152 13710 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38152 13710 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38233 13710 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38233 13710 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38314 13710 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38314 13710 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38395 13710 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38395 13710 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38476 13710 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38476 13710 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38557 13710 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38557 13710 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38638 13710 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38638 13710 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38719 13710 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38719 13710 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38800 13710 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38800 13710 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38881 13710 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38881 13710 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 38962 13710 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 38962 13710 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 39043 13710 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 39043 13710 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 39124 13710 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 39124 13710 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 39205 13710 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 39205 13710 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 39286 13710 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 39286 13710 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 39367 13710 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 39367 13710 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 39448 13710 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 39448 13710 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13646 39529 13710 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13646 39529 13710 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 4770 13718 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 4770 13718 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 4856 13718 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 4856 13718 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 4942 13718 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 4942 13718 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 5028 13718 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 5028 13718 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 5114 13718 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 5114 13718 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 5200 13718 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 5200 13718 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 5286 13718 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 5286 13718 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 5372 13718 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 5372 13718 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 5458 13718 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 5458 13718 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 5544 13718 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 5544 13718 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13654 5630 13718 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13654 5630 13718 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 34768 13792 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 34768 13792 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 34848 13792 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 34848 13792 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 34928 13792 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 34928 13792 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35008 13792 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35008 13792 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35088 13792 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35088 13792 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35168 13792 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35168 13792 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35248 13792 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35248 13792 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35328 13792 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35328 13792 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35408 13792 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35408 13792 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35488 13792 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35488 13792 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35568 13792 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35568 13792 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35648 13792 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35648 13792 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35728 13792 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35728 13792 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35808 13792 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35808 13792 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35888 13792 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35888 13792 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 35968 13792 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 35968 13792 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36048 13792 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36048 13792 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36128 13792 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36128 13792 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36208 13792 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36208 13792 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36289 13792 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36289 13792 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36370 13792 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36370 13792 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36451 13792 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36451 13792 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36532 13792 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36532 13792 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36613 13792 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36613 13792 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36694 13792 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36694 13792 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36775 13792 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36775 13792 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36856 13792 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36856 13792 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 36937 13792 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 36937 13792 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37018 13792 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37018 13792 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37099 13792 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37099 13792 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37180 13792 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37180 13792 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37261 13792 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37261 13792 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37342 13792 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37342 13792 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37423 13792 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37423 13792 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37504 13792 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37504 13792 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37585 13792 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37585 13792 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37666 13792 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37666 13792 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37747 13792 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37747 13792 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37828 13792 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37828 13792 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37909 13792 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37909 13792 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 37990 13792 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 37990 13792 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38071 13792 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38071 13792 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38152 13792 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38152 13792 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38233 13792 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38233 13792 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38314 13792 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38314 13792 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38395 13792 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38395 13792 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38476 13792 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38476 13792 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38557 13792 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38557 13792 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38638 13792 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38638 13792 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38719 13792 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38719 13792 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38800 13792 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38800 13792 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38881 13792 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38881 13792 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 38962 13792 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 38962 13792 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 39043 13792 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 39043 13792 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 39124 13792 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 39124 13792 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 39205 13792 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 39205 13792 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 39286 13792 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 39286 13792 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 39367 13792 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 39367 13792 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 39448 13792 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 39448 13792 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13728 39529 13792 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13728 39529 13792 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 4770 13799 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 4770 13799 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 4856 13799 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 4856 13799 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 4942 13799 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 4942 13799 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 5028 13799 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 5028 13799 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 5114 13799 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 5114 13799 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 5200 13799 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 5200 13799 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 5286 13799 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 5286 13799 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 5372 13799 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 5372 13799 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 5458 13799 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 5458 13799 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 5544 13799 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 5544 13799 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13735 5630 13799 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13735 5630 13799 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 34768 13874 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 34768 13874 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 34848 13874 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 34848 13874 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 34928 13874 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 34928 13874 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35008 13874 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35008 13874 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35088 13874 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35088 13874 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35168 13874 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35168 13874 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35248 13874 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35248 13874 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35328 13874 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35328 13874 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35408 13874 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35408 13874 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35488 13874 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35488 13874 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35568 13874 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35568 13874 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35648 13874 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35648 13874 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35728 13874 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35728 13874 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35808 13874 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35808 13874 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35888 13874 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35888 13874 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 35968 13874 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 35968 13874 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36048 13874 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36048 13874 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36128 13874 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36128 13874 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36208 13874 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36208 13874 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36289 13874 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36289 13874 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36370 13874 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36370 13874 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36451 13874 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36451 13874 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36532 13874 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36532 13874 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36613 13874 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36613 13874 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36694 13874 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36694 13874 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36775 13874 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36775 13874 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36856 13874 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36856 13874 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 36937 13874 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 36937 13874 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37018 13874 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37018 13874 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37099 13874 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37099 13874 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37180 13874 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37180 13874 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37261 13874 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37261 13874 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37342 13874 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37342 13874 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37423 13874 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37423 13874 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37504 13874 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37504 13874 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37585 13874 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37585 13874 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37666 13874 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37666 13874 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37747 13874 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37747 13874 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37828 13874 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37828 13874 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37909 13874 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37909 13874 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 37990 13874 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 37990 13874 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38071 13874 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38071 13874 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38152 13874 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38152 13874 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38233 13874 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38233 13874 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38314 13874 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38314 13874 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38395 13874 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38395 13874 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38476 13874 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38476 13874 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38557 13874 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38557 13874 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38638 13874 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38638 13874 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38719 13874 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38719 13874 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38800 13874 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38800 13874 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38881 13874 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38881 13874 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 38962 13874 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 38962 13874 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 39043 13874 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 39043 13874 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 39124 13874 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 39124 13874 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 39205 13874 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 39205 13874 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 39286 13874 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 39286 13874 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 39367 13874 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 39367 13874 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 39448 13874 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 39448 13874 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13810 39529 13874 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13810 39529 13874 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 4770 13880 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 4770 13880 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 4856 13880 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 4856 13880 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 4942 13880 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 4942 13880 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 5028 13880 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 5028 13880 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 5114 13880 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 5114 13880 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 5200 13880 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 5200 13880 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 5286 13880 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 5286 13880 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 5372 13880 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 5372 13880 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 5458 13880 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 5458 13880 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 5544 13880 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 5544 13880 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13816 5630 13880 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13816 5630 13880 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 34768 13956 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 34768 13956 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 34848 13956 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 34848 13956 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 34928 13956 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 34928 13956 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35008 13956 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35008 13956 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35088 13956 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35088 13956 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35168 13956 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35168 13956 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35248 13956 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35248 13956 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35328 13956 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35328 13956 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35408 13956 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35408 13956 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35488 13956 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35488 13956 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35568 13956 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35568 13956 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35648 13956 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35648 13956 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35728 13956 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35728 13956 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35808 13956 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35808 13956 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35888 13956 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35888 13956 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 35968 13956 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 35968 13956 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36048 13956 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36048 13956 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36128 13956 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36128 13956 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36208 13956 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36208 13956 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36289 13956 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36289 13956 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36370 13956 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36370 13956 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36451 13956 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36451 13956 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36532 13956 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36532 13956 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36613 13956 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36613 13956 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36694 13956 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36694 13956 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36775 13956 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36775 13956 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36856 13956 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36856 13956 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 36937 13956 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 36937 13956 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37018 13956 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37018 13956 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37099 13956 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37099 13956 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37180 13956 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37180 13956 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37261 13956 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37261 13956 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37342 13956 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37342 13956 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37423 13956 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37423 13956 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37504 13956 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37504 13956 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37585 13956 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37585 13956 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37666 13956 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37666 13956 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37747 13956 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37747 13956 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37828 13956 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37828 13956 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37909 13956 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37909 13956 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 37990 13956 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 37990 13956 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38071 13956 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38071 13956 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38152 13956 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38152 13956 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38233 13956 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38233 13956 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38314 13956 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38314 13956 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38395 13956 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38395 13956 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38476 13956 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38476 13956 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38557 13956 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38557 13956 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38638 13956 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38638 13956 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38719 13956 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38719 13956 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38800 13956 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38800 13956 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38881 13956 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38881 13956 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 38962 13956 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 38962 13956 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 39043 13956 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 39043 13956 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 39124 13956 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 39124 13956 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 39205 13956 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 39205 13956 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 39286 13956 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 39286 13956 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 39367 13956 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 39367 13956 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 39448 13956 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 39448 13956 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13892 39529 13956 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13892 39529 13956 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 4770 13961 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 4770 13961 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 4856 13961 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 4856 13961 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 4942 13961 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 4942 13961 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 5028 13961 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 5028 13961 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 5114 13961 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 5114 13961 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 5200 13961 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 5200 13961 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 5286 13961 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 5286 13961 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 5372 13961 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 5372 13961 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 5458 13961 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 5458 13961 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 5544 13961 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 5544 13961 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13897 5630 13961 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13897 5630 13961 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 34768 14038 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 34768 14038 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 34848 14038 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 34848 14038 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 34928 14038 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 34928 14038 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35008 14038 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35008 14038 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35088 14038 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35088 14038 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35168 14038 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35168 14038 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35248 14038 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35248 14038 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35328 14038 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35328 14038 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35408 14038 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35408 14038 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35488 14038 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35488 14038 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35568 14038 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35568 14038 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35648 14038 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35648 14038 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35728 14038 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35728 14038 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35808 14038 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35808 14038 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35888 14038 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35888 14038 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 35968 14038 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 35968 14038 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36048 14038 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36048 14038 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36128 14038 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36128 14038 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36208 14038 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36208 14038 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36289 14038 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36289 14038 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36370 14038 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36370 14038 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36451 14038 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36451 14038 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36532 14038 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36532 14038 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36613 14038 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36613 14038 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36694 14038 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36694 14038 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36775 14038 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36775 14038 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36856 14038 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36856 14038 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 36937 14038 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 36937 14038 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37018 14038 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37018 14038 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37099 14038 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37099 14038 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37180 14038 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37180 14038 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37261 14038 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37261 14038 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37342 14038 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37342 14038 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37423 14038 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37423 14038 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37504 14038 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37504 14038 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37585 14038 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37585 14038 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37666 14038 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37666 14038 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37747 14038 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37747 14038 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37828 14038 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37828 14038 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37909 14038 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37909 14038 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 37990 14038 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 37990 14038 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38071 14038 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38071 14038 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38152 14038 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38152 14038 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38233 14038 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38233 14038 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38314 14038 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38314 14038 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38395 14038 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38395 14038 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38476 14038 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38476 14038 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38557 14038 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38557 14038 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38638 14038 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38638 14038 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38719 14038 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38719 14038 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38800 14038 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38800 14038 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38881 14038 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38881 14038 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 38962 14038 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 38962 14038 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 39043 14038 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 39043 14038 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 39124 14038 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 39124 14038 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 39205 14038 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 39205 14038 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 39286 14038 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 39286 14038 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 39367 14038 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 39367 14038 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 39448 14038 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 39448 14038 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13974 39529 14038 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13974 39529 14038 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 4770 14042 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 4770 14042 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 4856 14042 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 4856 14042 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 4942 14042 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 4942 14042 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 5028 14042 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 5028 14042 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 5114 14042 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 5114 14042 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 5200 14042 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 5200 14042 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 5286 14042 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 5286 14042 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 5372 14042 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 5372 14042 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 5458 14042 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 5458 14042 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 5544 14042 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 5544 14042 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 13978 5630 14042 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 13978 5630 14042 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 34780 1443 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 34860 1443 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 34940 1443 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35020 1443 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35100 1443 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35180 1443 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35260 1443 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35340 1443 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35420 1443 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35500 1443 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35580 1443 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35660 1443 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35740 1443 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35820 1443 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35900 1443 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 35980 1443 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 36060 1443 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 36140 1443 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1403 36220 1443 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 4770 1472 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 4770 1472 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 4856 1472 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 4856 1472 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 4942 1472 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 4942 1472 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 5028 1472 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 5028 1472 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 5114 1472 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 5114 1472 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 5200 1472 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 5200 1472 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 5286 1472 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 5286 1472 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 5372 1472 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 5372 1472 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 5458 1472 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 5458 1472 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 5544 1472 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 5544 1472 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1408 5630 1472 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1408 5630 1472 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36289 1535 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36289 1535 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36370 1535 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36370 1535 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36451 1535 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36451 1535 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36532 1535 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36532 1535 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36613 1535 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36613 1535 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36694 1535 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36694 1535 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36775 1535 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36775 1535 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36856 1535 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36856 1535 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 36937 1535 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 36937 1535 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37018 1535 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37018 1535 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37099 1535 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37099 1535 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37180 1535 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37180 1535 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37261 1535 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37261 1535 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37342 1535 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37342 1535 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37423 1535 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37423 1535 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37504 1535 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37504 1535 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37585 1535 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37585 1535 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37666 1535 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37666 1535 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37747 1535 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37747 1535 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37828 1535 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37828 1535 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37909 1535 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37909 1535 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 37990 1535 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 37990 1535 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38071 1535 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38071 1535 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38152 1535 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38152 1535 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38233 1535 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38233 1535 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38314 1535 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38314 1535 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38395 1535 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38395 1535 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38476 1535 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38476 1535 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38557 1535 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38557 1535 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38638 1535 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38638 1535 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38719 1535 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38719 1535 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38800 1535 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38800 1535 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38881 1535 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38881 1535 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 38962 1535 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 38962 1535 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 39043 1535 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 39043 1535 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 39124 1535 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 39124 1535 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 39205 1535 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 39205 1535 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 39286 1535 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 39286 1535 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 39367 1535 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 39367 1535 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 39448 1535 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 39448 1535 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1471 39529 1535 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1471 39529 1535 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 34780 1523 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 34860 1523 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 34940 1523 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35020 1523 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35100 1523 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35180 1523 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35260 1523 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35340 1523 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35420 1523 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35500 1523 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35580 1523 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35660 1523 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35740 1523 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35820 1523 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35900 1523 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 35980 1523 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 36060 1523 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 36140 1523 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1483 36220 1523 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 4770 1553 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 4770 1553 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 4856 1553 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 4856 1553 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 4942 1553 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 4942 1553 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 5028 1553 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 5028 1553 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 5114 1553 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 5114 1553 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 5200 1553 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 5200 1553 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 5286 1553 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 5286 1553 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 5372 1553 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 5372 1553 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 5458 1553 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 5458 1553 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 5544 1553 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 5544 1553 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1489 5630 1553 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1489 5630 1553 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36289 1615 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36289 1615 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36370 1615 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36370 1615 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36451 1615 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36451 1615 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36532 1615 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36532 1615 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36613 1615 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36613 1615 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36694 1615 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36694 1615 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36775 1615 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36775 1615 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36856 1615 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36856 1615 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 36937 1615 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 36937 1615 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37018 1615 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37018 1615 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37099 1615 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37099 1615 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37180 1615 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37180 1615 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37261 1615 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37261 1615 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37342 1615 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37342 1615 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37423 1615 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37423 1615 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37504 1615 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37504 1615 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37585 1615 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37585 1615 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37666 1615 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37666 1615 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37747 1615 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37747 1615 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37828 1615 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37828 1615 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37909 1615 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37909 1615 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 37990 1615 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 37990 1615 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38071 1615 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38071 1615 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38152 1615 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38152 1615 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38233 1615 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38233 1615 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38314 1615 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38314 1615 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38395 1615 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38395 1615 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38476 1615 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38476 1615 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38557 1615 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38557 1615 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38638 1615 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38638 1615 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38719 1615 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38719 1615 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38800 1615 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38800 1615 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38881 1615 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38881 1615 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 38962 1615 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 38962 1615 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 39043 1615 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 39043 1615 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 39124 1615 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 39124 1615 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 39205 1615 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 39205 1615 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 39286 1615 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 39286 1615 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 39367 1615 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 39367 1615 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 39448 1615 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 39448 1615 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1551 39529 1615 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1551 39529 1615 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 34780 1603 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 34860 1603 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 34940 1603 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35020 1603 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35100 1603 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35180 1603 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35260 1603 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35340 1603 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35420 1603 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35500 1603 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35580 1603 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35660 1603 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35740 1603 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35820 1603 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35900 1603 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 35980 1603 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 36060 1603 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 36140 1603 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1563 36220 1603 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 4770 1634 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 4770 1634 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 4856 1634 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 4856 1634 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 4942 1634 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 4942 1634 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 5028 1634 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 5028 1634 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 5114 1634 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 5114 1634 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 5200 1634 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 5200 1634 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 5286 1634 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 5286 1634 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 5372 1634 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 5372 1634 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 5458 1634 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 5458 1634 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 5544 1634 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 5544 1634 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1570 5630 1634 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1570 5630 1634 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 34768 14120 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 34768 14120 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 34848 14120 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 34848 14120 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 34928 14120 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 34928 14120 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35008 14120 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35008 14120 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35088 14120 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35088 14120 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35168 14120 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35168 14120 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35248 14120 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35248 14120 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35328 14120 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35328 14120 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35408 14120 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35408 14120 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35488 14120 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35488 14120 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35568 14120 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35568 14120 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35648 14120 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35648 14120 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35728 14120 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35728 14120 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35808 14120 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35808 14120 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35888 14120 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35888 14120 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 35968 14120 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 35968 14120 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36048 14120 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36048 14120 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36128 14120 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36128 14120 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36208 14120 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36208 14120 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36289 14120 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36289 14120 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36370 14120 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36370 14120 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36451 14120 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36451 14120 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36532 14120 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36532 14120 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36613 14120 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36613 14120 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36694 14120 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36694 14120 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36775 14120 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36775 14120 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36856 14120 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36856 14120 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 36937 14120 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 36937 14120 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37018 14120 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37018 14120 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37099 14120 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37099 14120 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37180 14120 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37180 14120 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37261 14120 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37261 14120 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37342 14120 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37342 14120 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37423 14120 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37423 14120 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37504 14120 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37504 14120 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37585 14120 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37585 14120 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37666 14120 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37666 14120 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37747 14120 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37747 14120 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37828 14120 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37828 14120 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37909 14120 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37909 14120 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 37990 14120 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 37990 14120 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38071 14120 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38071 14120 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38152 14120 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38152 14120 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38233 14120 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38233 14120 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38314 14120 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38314 14120 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38395 14120 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38395 14120 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38476 14120 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38476 14120 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38557 14120 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38557 14120 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38638 14120 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38638 14120 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38719 14120 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38719 14120 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38800 14120 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38800 14120 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38881 14120 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38881 14120 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 38962 14120 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 38962 14120 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 39043 14120 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 39043 14120 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 39124 14120 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 39124 14120 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 39205 14120 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 39205 14120 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 39286 14120 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 39286 14120 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 39367 14120 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 39367 14120 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 39448 14120 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 39448 14120 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14056 39529 14120 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14056 39529 14120 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 4770 14123 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 4770 14123 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 4856 14123 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 4856 14123 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 4942 14123 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 4942 14123 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 5028 14123 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 5028 14123 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 5114 14123 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 5114 14123 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 5200 14123 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 5200 14123 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 5286 14123 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 5286 14123 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 5372 14123 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 5372 14123 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 5458 14123 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 5458 14123 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 5544 14123 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 5544 14123 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14059 5630 14123 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14059 5630 14123 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 34768 14202 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 34768 14202 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 34848 14202 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 34848 14202 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 34928 14202 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 34928 14202 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35008 14202 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35008 14202 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35088 14202 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35088 14202 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35168 14202 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35168 14202 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35248 14202 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35248 14202 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35328 14202 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35328 14202 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35408 14202 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35408 14202 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35488 14202 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35488 14202 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35568 14202 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35568 14202 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35648 14202 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35648 14202 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35728 14202 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35728 14202 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35808 14202 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35808 14202 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35888 14202 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35888 14202 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 35968 14202 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 35968 14202 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36048 14202 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36048 14202 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36128 14202 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36128 14202 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36208 14202 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36208 14202 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36289 14202 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36289 14202 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36370 14202 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36370 14202 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36451 14202 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36451 14202 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36532 14202 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36532 14202 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36613 14202 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36613 14202 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36694 14202 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36694 14202 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36775 14202 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36775 14202 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36856 14202 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36856 14202 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 36937 14202 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 36937 14202 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37018 14202 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37018 14202 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37099 14202 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37099 14202 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37180 14202 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37180 14202 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37261 14202 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37261 14202 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37342 14202 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37342 14202 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37423 14202 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37423 14202 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37504 14202 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37504 14202 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37585 14202 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37585 14202 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37666 14202 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37666 14202 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37747 14202 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37747 14202 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37828 14202 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37828 14202 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37909 14202 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37909 14202 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 37990 14202 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 37990 14202 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38071 14202 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38071 14202 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38152 14202 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38152 14202 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38233 14202 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38233 14202 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38314 14202 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38314 14202 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38395 14202 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38395 14202 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38476 14202 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38476 14202 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38557 14202 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38557 14202 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38638 14202 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38638 14202 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38719 14202 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38719 14202 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38800 14202 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38800 14202 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38881 14202 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38881 14202 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 38962 14202 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 38962 14202 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 39043 14202 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 39043 14202 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 39124 14202 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 39124 14202 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 39205 14202 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 39205 14202 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 39286 14202 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 39286 14202 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 39367 14202 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 39367 14202 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 39448 14202 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 39448 14202 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14138 39529 14202 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14138 39529 14202 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 4770 14204 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 4770 14204 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 4856 14204 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 4856 14204 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 4942 14204 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 4942 14204 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 5028 14204 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 5028 14204 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 5114 14204 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 5114 14204 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 5200 14204 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 5200 14204 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 5286 14204 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 5286 14204 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 5372 14204 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 5372 14204 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 5458 14204 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 5458 14204 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 5544 14204 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 5544 14204 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14140 5630 14204 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14140 5630 14204 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 34768 14284 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 34768 14284 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 34848 14284 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 34848 14284 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 34928 14284 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 34928 14284 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35008 14284 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35008 14284 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35088 14284 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35088 14284 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35168 14284 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35168 14284 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35248 14284 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35248 14284 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35328 14284 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35328 14284 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35408 14284 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35408 14284 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35488 14284 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35488 14284 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35568 14284 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35568 14284 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35648 14284 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35648 14284 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35728 14284 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35728 14284 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35808 14284 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35808 14284 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35888 14284 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35888 14284 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 35968 14284 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 35968 14284 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36048 14284 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36048 14284 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36128 14284 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36128 14284 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36208 14284 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36208 14284 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36289 14284 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36289 14284 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36370 14284 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36370 14284 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36451 14284 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36451 14284 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36532 14284 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36532 14284 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36613 14284 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36613 14284 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36694 14284 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36694 14284 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36775 14284 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36775 14284 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36856 14284 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36856 14284 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 36937 14284 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 36937 14284 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37018 14284 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37018 14284 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37099 14284 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37099 14284 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37180 14284 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37180 14284 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37261 14284 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37261 14284 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37342 14284 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37342 14284 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37423 14284 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37423 14284 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37504 14284 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37504 14284 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37585 14284 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37585 14284 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37666 14284 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37666 14284 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37747 14284 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37747 14284 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37828 14284 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37828 14284 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37909 14284 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37909 14284 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 37990 14284 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 37990 14284 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38071 14284 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38071 14284 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38152 14284 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38152 14284 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38233 14284 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38233 14284 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38314 14284 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38314 14284 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38395 14284 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38395 14284 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38476 14284 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38476 14284 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38557 14284 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38557 14284 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38638 14284 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38638 14284 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38719 14284 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38719 14284 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38800 14284 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38800 14284 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38881 14284 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38881 14284 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 38962 14284 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 38962 14284 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 39043 14284 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 39043 14284 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 39124 14284 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 39124 14284 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 39205 14284 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 39205 14284 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 39286 14284 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 39286 14284 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 39367 14284 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 39367 14284 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 39448 14284 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 39448 14284 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14220 39529 14284 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14220 39529 14284 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 4770 14285 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 4770 14285 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 4856 14285 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 4856 14285 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 4942 14285 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 4942 14285 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 5028 14285 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 5028 14285 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 5114 14285 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 5114 14285 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 5200 14285 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 5200 14285 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 5286 14285 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 5286 14285 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 5372 14285 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 5372 14285 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 5458 14285 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 5458 14285 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 5544 14285 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 5544 14285 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14221 5630 14285 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14221 5630 14285 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 34768 14366 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 34768 14366 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 34848 14366 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 34848 14366 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 34928 14366 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 34928 14366 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35008 14366 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35008 14366 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35088 14366 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35088 14366 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35168 14366 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35168 14366 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35248 14366 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35248 14366 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35328 14366 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35328 14366 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35408 14366 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35408 14366 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35488 14366 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35488 14366 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35568 14366 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35568 14366 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35648 14366 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35648 14366 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35728 14366 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35728 14366 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35808 14366 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35808 14366 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35888 14366 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35888 14366 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 35968 14366 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 35968 14366 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36048 14366 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36048 14366 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36128 14366 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36128 14366 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36208 14366 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36208 14366 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36289 14366 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36289 14366 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36370 14366 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36370 14366 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36451 14366 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36451 14366 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36532 14366 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36532 14366 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36613 14366 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36613 14366 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36694 14366 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36694 14366 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36775 14366 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36775 14366 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36856 14366 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36856 14366 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 36937 14366 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 36937 14366 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37018 14366 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37018 14366 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37099 14366 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37099 14366 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37180 14366 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37180 14366 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37261 14366 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37261 14366 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37342 14366 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37342 14366 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37423 14366 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37423 14366 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37504 14366 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37504 14366 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37585 14366 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37585 14366 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37666 14366 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37666 14366 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37747 14366 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37747 14366 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37828 14366 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37828 14366 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37909 14366 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37909 14366 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 37990 14366 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 37990 14366 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38071 14366 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38071 14366 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38152 14366 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38152 14366 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38233 14366 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38233 14366 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38314 14366 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38314 14366 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38395 14366 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38395 14366 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38476 14366 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38476 14366 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38557 14366 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38557 14366 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38638 14366 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38638 14366 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38719 14366 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38719 14366 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38800 14366 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38800 14366 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38881 14366 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38881 14366 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 38962 14366 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 38962 14366 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 39043 14366 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 39043 14366 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 39124 14366 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 39124 14366 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 39205 14366 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 39205 14366 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 39286 14366 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 39286 14366 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 39367 14366 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 39367 14366 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 39448 14366 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 39448 14366 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 39529 14366 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 39529 14366 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 4770 14366 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 4770 14366 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 4856 14366 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 4856 14366 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 4942 14366 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 4942 14366 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 5028 14366 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 5028 14366 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 5114 14366 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 5114 14366 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 5200 14366 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 5200 14366 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 5286 14366 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 5286 14366 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 5372 14366 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 5372 14366 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 5458 14366 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 5458 14366 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 5544 14366 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 5544 14366 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14302 5630 14366 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14302 5630 14366 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 4770 14447 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 4770 14447 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 4856 14447 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 4856 14447 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 4942 14447 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 4942 14447 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 5028 14447 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 5028 14447 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 5114 14447 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 5114 14447 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 5200 14447 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 5200 14447 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 5286 14447 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 5286 14447 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 5372 14447 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 5372 14447 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 5458 14447 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 5458 14447 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 5544 14447 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 5544 14447 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14383 5630 14447 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14383 5630 14447 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 34768 14448 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 34768 14448 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 34848 14448 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 34848 14448 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 34928 14448 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 34928 14448 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35008 14448 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35008 14448 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35088 14448 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35088 14448 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35168 14448 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35168 14448 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35248 14448 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35248 14448 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35328 14448 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35328 14448 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35408 14448 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35408 14448 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35488 14448 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35488 14448 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35568 14448 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35568 14448 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35648 14448 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35648 14448 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35728 14448 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35728 14448 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35808 14448 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35808 14448 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35888 14448 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35888 14448 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 35968 14448 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 35968 14448 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36048 14448 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36048 14448 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36128 14448 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36128 14448 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36208 14448 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36208 14448 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36289 14448 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36289 14448 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36370 14448 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36370 14448 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36451 14448 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36451 14448 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36532 14448 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36532 14448 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36613 14448 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36613 14448 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36694 14448 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36694 14448 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36775 14448 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36775 14448 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36856 14448 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36856 14448 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 36937 14448 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 36937 14448 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37018 14448 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37018 14448 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37099 14448 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37099 14448 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37180 14448 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37180 14448 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37261 14448 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37261 14448 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37342 14448 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37342 14448 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37423 14448 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37423 14448 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37504 14448 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37504 14448 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37585 14448 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37585 14448 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37666 14448 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37666 14448 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37747 14448 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37747 14448 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37828 14448 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37828 14448 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37909 14448 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37909 14448 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 37990 14448 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 37990 14448 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38071 14448 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38071 14448 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38152 14448 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38152 14448 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38233 14448 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38233 14448 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38314 14448 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38314 14448 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38395 14448 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38395 14448 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38476 14448 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38476 14448 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38557 14448 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38557 14448 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38638 14448 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38638 14448 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38719 14448 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38719 14448 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38800 14448 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38800 14448 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38881 14448 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38881 14448 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 38962 14448 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 38962 14448 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 39043 14448 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 39043 14448 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 39124 14448 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 39124 14448 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 39205 14448 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 39205 14448 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 39286 14448 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 39286 14448 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 39367 14448 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 39367 14448 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 39448 14448 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 39448 14448 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14384 39529 14448 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14384 39529 14448 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 4770 14528 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 4770 14528 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 4856 14528 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 4856 14528 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 4942 14528 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 4942 14528 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 5028 14528 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 5028 14528 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 5114 14528 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 5114 14528 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 5200 14528 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 5200 14528 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 5286 14528 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 5286 14528 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 5372 14528 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 5372 14528 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 5458 14528 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 5458 14528 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 5544 14528 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 5544 14528 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14464 5630 14528 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14464 5630 14528 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 34768 14530 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 34768 14530 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 34848 14530 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 34848 14530 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 34928 14530 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 34928 14530 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35008 14530 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35008 14530 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35088 14530 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35088 14530 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35168 14530 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35168 14530 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35248 14530 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35248 14530 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35328 14530 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35328 14530 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35408 14530 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35408 14530 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35488 14530 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35488 14530 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35568 14530 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35568 14530 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35648 14530 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35648 14530 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35728 14530 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35728 14530 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35808 14530 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35808 14530 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35888 14530 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35888 14530 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 35968 14530 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 35968 14530 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36048 14530 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36048 14530 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36128 14530 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36128 14530 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36208 14530 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36208 14530 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36289 14530 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36289 14530 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36370 14530 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36370 14530 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36451 14530 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36451 14530 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36532 14530 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36532 14530 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36613 14530 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36613 14530 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36694 14530 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36694 14530 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36775 14530 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36775 14530 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36856 14530 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36856 14530 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 36937 14530 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 36937 14530 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37018 14530 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37018 14530 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37099 14530 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37099 14530 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37180 14530 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37180 14530 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37261 14530 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37261 14530 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37342 14530 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37342 14530 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37423 14530 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37423 14530 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37504 14530 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37504 14530 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37585 14530 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37585 14530 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37666 14530 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37666 14530 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37747 14530 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37747 14530 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37828 14530 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37828 14530 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37909 14530 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37909 14530 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 37990 14530 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 37990 14530 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38071 14530 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38071 14530 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38152 14530 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38152 14530 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38233 14530 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38233 14530 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38314 14530 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38314 14530 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38395 14530 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38395 14530 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38476 14530 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38476 14530 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38557 14530 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38557 14530 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38638 14530 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38638 14530 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38719 14530 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38719 14530 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38800 14530 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38800 14530 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38881 14530 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38881 14530 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 38962 14530 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 38962 14530 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 39043 14530 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 39043 14530 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 39124 14530 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 39124 14530 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 39205 14530 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 39205 14530 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 39286 14530 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 39286 14530 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 39367 14530 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 39367 14530 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 39448 14530 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 39448 14530 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14466 39529 14530 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14466 39529 14530 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 4770 14609 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 4770 14609 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 4856 14609 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 4856 14609 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 4942 14609 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 4942 14609 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 5028 14609 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 5028 14609 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 5114 14609 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 5114 14609 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 5200 14609 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 5200 14609 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 5286 14609 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 5286 14609 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 5372 14609 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 5372 14609 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 5458 14609 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 5458 14609 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 5544 14609 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 5544 14609 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14545 5630 14609 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14545 5630 14609 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 34768 14612 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 34768 14612 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 34848 14612 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 34848 14612 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 34928 14612 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 34928 14612 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35008 14612 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35008 14612 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35088 14612 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35088 14612 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35168 14612 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35168 14612 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35248 14612 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35248 14612 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35328 14612 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35328 14612 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35408 14612 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35408 14612 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35488 14612 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35488 14612 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35568 14612 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35568 14612 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35648 14612 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35648 14612 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35728 14612 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35728 14612 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35808 14612 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35808 14612 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35888 14612 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35888 14612 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 35968 14612 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 35968 14612 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36048 14612 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36048 14612 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36128 14612 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36128 14612 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36208 14612 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36208 14612 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36289 14612 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36289 14612 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36370 14612 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36370 14612 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36451 14612 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36451 14612 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36532 14612 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36532 14612 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36613 14612 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36613 14612 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36694 14612 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36694 14612 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36775 14612 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36775 14612 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36856 14612 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36856 14612 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 36937 14612 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 36937 14612 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37018 14612 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37018 14612 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37099 14612 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37099 14612 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37180 14612 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37180 14612 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37261 14612 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37261 14612 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37342 14612 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37342 14612 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37423 14612 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37423 14612 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37504 14612 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37504 14612 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37585 14612 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37585 14612 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37666 14612 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37666 14612 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37747 14612 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37747 14612 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37828 14612 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37828 14612 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37909 14612 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37909 14612 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 37990 14612 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 37990 14612 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38071 14612 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38071 14612 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38152 14612 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38152 14612 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38233 14612 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38233 14612 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38314 14612 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38314 14612 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38395 14612 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38395 14612 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38476 14612 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38476 14612 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38557 14612 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38557 14612 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38638 14612 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38638 14612 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38719 14612 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38719 14612 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38800 14612 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38800 14612 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38881 14612 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38881 14612 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 38962 14612 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 38962 14612 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 39043 14612 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 39043 14612 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 39124 14612 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 39124 14612 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 39205 14612 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 39205 14612 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 39286 14612 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 39286 14612 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 39367 14612 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 39367 14612 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 39448 14612 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 39448 14612 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14548 39529 14612 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14548 39529 14612 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 4770 14690 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 4770 14690 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 4856 14690 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 4856 14690 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 4942 14690 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 4942 14690 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 5028 14690 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 5028 14690 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 5114 14690 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 5114 14690 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 5200 14690 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 5200 14690 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 5286 14690 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 5286 14690 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 5372 14690 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 5372 14690 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 5458 14690 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 5458 14690 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 5544 14690 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 5544 14690 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14626 5630 14690 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14626 5630 14690 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 34768 14694 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 34768 14694 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 34848 14694 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 34848 14694 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 34928 14694 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 34928 14694 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35008 14694 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35008 14694 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35088 14694 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35088 14694 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35168 14694 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35168 14694 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35248 14694 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35248 14694 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35328 14694 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35328 14694 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35408 14694 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35408 14694 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35488 14694 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35488 14694 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35568 14694 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35568 14694 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35648 14694 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35648 14694 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35728 14694 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35728 14694 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35808 14694 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35808 14694 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35888 14694 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35888 14694 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 35968 14694 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 35968 14694 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36048 14694 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36048 14694 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36128 14694 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36128 14694 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36208 14694 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36208 14694 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36289 14694 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36289 14694 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36370 14694 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36370 14694 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36451 14694 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36451 14694 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36532 14694 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36532 14694 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36613 14694 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36613 14694 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36694 14694 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36694 14694 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36775 14694 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36775 14694 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36856 14694 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36856 14694 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 36937 14694 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 36937 14694 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37018 14694 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37018 14694 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37099 14694 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37099 14694 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37180 14694 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37180 14694 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37261 14694 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37261 14694 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37342 14694 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37342 14694 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37423 14694 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37423 14694 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37504 14694 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37504 14694 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37585 14694 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37585 14694 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37666 14694 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37666 14694 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37747 14694 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37747 14694 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37828 14694 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37828 14694 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37909 14694 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37909 14694 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 37990 14694 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 37990 14694 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38071 14694 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38071 14694 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38152 14694 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38152 14694 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38233 14694 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38233 14694 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38314 14694 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38314 14694 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38395 14694 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38395 14694 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38476 14694 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38476 14694 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38557 14694 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38557 14694 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38638 14694 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38638 14694 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38719 14694 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38719 14694 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38800 14694 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38800 14694 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38881 14694 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38881 14694 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 38962 14694 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 38962 14694 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 39043 14694 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 39043 14694 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 39124 14694 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 39124 14694 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 39205 14694 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 39205 14694 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 39286 14694 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 39286 14694 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 39367 14694 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 39367 14694 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 39448 14694 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 39448 14694 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14630 39529 14694 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14630 39529 14694 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 4770 14771 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 4770 14771 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 4856 14771 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 4856 14771 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 4942 14771 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 4942 14771 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 5028 14771 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 5028 14771 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 5114 14771 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 5114 14771 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 5200 14771 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 5200 14771 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 5286 14771 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 5286 14771 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 5372 14771 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 5372 14771 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 5458 14771 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 5458 14771 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 5544 14771 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 5544 14771 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14707 5630 14771 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14707 5630 14771 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 34768 14776 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 34768 14776 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 34848 14776 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 34848 14776 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 34928 14776 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 34928 14776 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35008 14776 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35008 14776 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35088 14776 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35088 14776 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35168 14776 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35168 14776 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35248 14776 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35248 14776 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35328 14776 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35328 14776 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35408 14776 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35408 14776 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35488 14776 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35488 14776 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35568 14776 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35568 14776 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35648 14776 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35648 14776 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35728 14776 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35728 14776 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35808 14776 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35808 14776 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35888 14776 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35888 14776 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 35968 14776 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 35968 14776 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36048 14776 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36048 14776 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36128 14776 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36128 14776 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36208 14776 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36208 14776 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36289 14776 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36289 14776 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36370 14776 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36370 14776 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36451 14776 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36451 14776 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36532 14776 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36532 14776 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36613 14776 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36613 14776 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36694 14776 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36694 14776 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36775 14776 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36775 14776 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36856 14776 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36856 14776 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 36937 14776 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 36937 14776 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37018 14776 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37018 14776 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37099 14776 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37099 14776 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37180 14776 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37180 14776 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37261 14776 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37261 14776 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37342 14776 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37342 14776 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37423 14776 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37423 14776 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37504 14776 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37504 14776 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37585 14776 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37585 14776 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37666 14776 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37666 14776 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37747 14776 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37747 14776 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37828 14776 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37828 14776 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37909 14776 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37909 14776 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 37990 14776 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 37990 14776 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38071 14776 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38071 14776 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38152 14776 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38152 14776 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38233 14776 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38233 14776 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38314 14776 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38314 14776 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38395 14776 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38395 14776 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38476 14776 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38476 14776 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38557 14776 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38557 14776 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38638 14776 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38638 14776 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38719 14776 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38719 14776 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38800 14776 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38800 14776 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38881 14776 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38881 14776 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 38962 14776 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 38962 14776 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 39043 14776 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 39043 14776 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 39124 14776 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 39124 14776 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 39205 14776 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 39205 14776 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 39286 14776 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 39286 14776 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 39367 14776 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 39367 14776 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 39448 14776 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 39448 14776 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14712 39529 14776 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14712 39529 14776 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 4770 14852 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 4770 14852 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 4856 14852 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 4856 14852 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 4942 14852 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 4942 14852 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 5028 14852 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 5028 14852 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 5114 14852 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 5114 14852 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 5200 14852 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 5200 14852 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 5286 14852 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 5286 14852 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 5372 14852 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 5372 14852 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 5458 14852 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 5458 14852 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 5544 14852 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 5544 14852 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14788 5630 14852 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14788 5630 14852 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 34768 14858 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 34768 14858 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 34848 14858 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 34848 14858 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 34928 14858 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 34928 14858 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35008 14858 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35008 14858 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35088 14858 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35088 14858 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35168 14858 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35168 14858 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35248 14858 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35248 14858 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35328 14858 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35328 14858 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35408 14858 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35408 14858 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35488 14858 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35488 14858 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35568 14858 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35568 14858 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35648 14858 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35648 14858 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35728 14858 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35728 14858 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35808 14858 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35808 14858 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35888 14858 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35888 14858 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 35968 14858 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 35968 14858 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36048 14858 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36048 14858 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36128 14858 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36128 14858 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36208 14858 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36208 14858 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36289 14858 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36289 14858 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36370 14858 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36370 14858 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36451 14858 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36451 14858 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36532 14858 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36532 14858 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36613 14858 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36613 14858 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36694 14858 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36694 14858 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36775 14858 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36775 14858 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36856 14858 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36856 14858 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 36937 14858 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 36937 14858 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37018 14858 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37018 14858 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37099 14858 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37099 14858 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37180 14858 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37180 14858 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37261 14858 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37261 14858 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37342 14858 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37342 14858 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37423 14858 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37423 14858 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37504 14858 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37504 14858 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37585 14858 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37585 14858 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37666 14858 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37666 14858 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37747 14858 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37747 14858 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37828 14858 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37828 14858 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37909 14858 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37909 14858 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 37990 14858 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 37990 14858 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38071 14858 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38071 14858 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38152 14858 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38152 14858 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38233 14858 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38233 14858 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38314 14858 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38314 14858 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38395 14858 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38395 14858 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38476 14858 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38476 14858 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38557 14858 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38557 14858 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38638 14858 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38638 14858 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38719 14858 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38719 14858 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38800 14858 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38800 14858 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38881 14858 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38881 14858 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 38962 14858 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 38962 14858 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 39043 14858 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 39043 14858 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 39124 14858 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 39124 14858 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 39205 14858 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 39205 14858 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 39286 14858 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 39286 14858 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 39367 14858 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 39367 14858 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 39448 14858 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 39448 14858 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14794 39529 14858 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14794 39529 14858 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 34768 14940 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 34768 14940 34832 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 34848 14940 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 34848 14940 34912 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 34928 14940 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 34928 14940 34992 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35008 14940 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35008 14940 35072 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35088 14940 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35088 14940 35152 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35168 14940 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35168 14940 35232 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35248 14940 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35248 14940 35312 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35328 14940 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35328 14940 35392 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35408 14940 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35408 14940 35472 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35488 14940 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35488 14940 35552 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35568 14940 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35568 14940 35632 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35648 14940 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35648 14940 35712 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35728 14940 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35728 14940 35792 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35808 14940 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35808 14940 35872 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35888 14940 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35888 14940 35952 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 35968 14940 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 35968 14940 36032 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36048 14940 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36048 14940 36112 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36128 14940 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36128 14940 36192 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36208 14940 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36208 14940 36272 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36289 14940 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36289 14940 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36370 14940 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36370 14940 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36451 14940 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36451 14940 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36532 14940 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36532 14940 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36613 14940 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36613 14940 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36694 14940 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36694 14940 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36775 14940 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36775 14940 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36856 14940 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36856 14940 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 36937 14940 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 36937 14940 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37018 14940 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37018 14940 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37099 14940 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37099 14940 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37180 14940 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37180 14940 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37261 14940 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37261 14940 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37342 14940 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37342 14940 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37423 14940 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37423 14940 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37504 14940 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37504 14940 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37585 14940 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37585 14940 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37666 14940 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37666 14940 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37747 14940 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37747 14940 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37828 14940 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37828 14940 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37909 14940 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37909 14940 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 37990 14940 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 37990 14940 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38071 14940 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38071 14940 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38152 14940 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38152 14940 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38233 14940 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38233 14940 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38314 14940 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38314 14940 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38395 14940 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38395 14940 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38476 14940 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38476 14940 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38557 14940 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38557 14940 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38638 14940 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38638 14940 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38719 14940 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38719 14940 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38800 14940 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38800 14940 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38881 14940 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38881 14940 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 38962 14940 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 38962 14940 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 39043 14940 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 39043 14940 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 39124 14940 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 39124 14940 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 39205 14940 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 39205 14940 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 39286 14940 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 39286 14940 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 39367 14940 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 39367 14940 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 39448 14940 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 39448 14940 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14876 39529 14940 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 14876 39529 14940 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36289 1695 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36289 1695 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36370 1695 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36370 1695 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36451 1695 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36451 1695 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36532 1695 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36532 1695 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36613 1695 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36613 1695 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36694 1695 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36694 1695 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36775 1695 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36775 1695 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36856 1695 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36856 1695 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 36937 1695 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 36937 1695 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37018 1695 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37018 1695 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37099 1695 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37099 1695 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37180 1695 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37180 1695 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37261 1695 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37261 1695 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37342 1695 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37342 1695 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37423 1695 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37423 1695 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37504 1695 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37504 1695 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37585 1695 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37585 1695 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37666 1695 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37666 1695 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37747 1695 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37747 1695 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37828 1695 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37828 1695 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37909 1695 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37909 1695 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 37990 1695 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 37990 1695 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38071 1695 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38071 1695 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38152 1695 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38152 1695 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38233 1695 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38233 1695 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38314 1695 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38314 1695 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38395 1695 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38395 1695 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38476 1695 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38476 1695 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38557 1695 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38557 1695 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38638 1695 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38638 1695 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38719 1695 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38719 1695 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38800 1695 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38800 1695 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38881 1695 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38881 1695 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 38962 1695 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 38962 1695 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 39043 1695 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 39043 1695 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 39124 1695 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 39124 1695 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 39205 1695 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 39205 1695 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 39286 1695 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 39286 1695 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 39367 1695 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 39367 1695 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 39448 1695 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 39448 1695 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1631 39529 1695 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1631 39529 1695 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 34780 1683 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 34860 1683 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 34940 1683 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35020 1683 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35100 1683 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35180 1683 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35260 1683 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35340 1683 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35420 1683 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35500 1683 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35580 1683 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35660 1683 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35740 1683 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35820 1683 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35900 1683 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 35980 1683 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 36060 1683 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 36140 1683 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1643 36220 1683 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 4770 1715 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 4770 1715 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 4856 1715 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 4856 1715 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 4942 1715 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 4942 1715 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 5028 1715 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 5028 1715 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 5114 1715 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 5114 1715 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 5200 1715 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 5200 1715 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 5286 1715 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 5286 1715 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 5372 1715 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 5372 1715 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 5458 1715 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 5458 1715 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 5544 1715 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 5544 1715 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1651 5630 1715 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1651 5630 1715 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36289 1775 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36289 1775 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36370 1775 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36370 1775 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36451 1775 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36451 1775 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36532 1775 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36532 1775 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36613 1775 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36613 1775 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36694 1775 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36694 1775 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36775 1775 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36775 1775 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36856 1775 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36856 1775 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 36937 1775 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 36937 1775 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37018 1775 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37018 1775 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37099 1775 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37099 1775 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37180 1775 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37180 1775 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37261 1775 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37261 1775 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37342 1775 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37342 1775 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37423 1775 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37423 1775 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37504 1775 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37504 1775 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37585 1775 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37585 1775 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37666 1775 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37666 1775 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37747 1775 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37747 1775 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37828 1775 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37828 1775 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37909 1775 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37909 1775 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 37990 1775 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 37990 1775 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38071 1775 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38071 1775 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38152 1775 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38152 1775 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38233 1775 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38233 1775 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38314 1775 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38314 1775 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38395 1775 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38395 1775 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38476 1775 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38476 1775 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38557 1775 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38557 1775 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38638 1775 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38638 1775 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38719 1775 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38719 1775 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38800 1775 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38800 1775 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38881 1775 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38881 1775 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 38962 1775 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 38962 1775 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 39043 1775 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 39043 1775 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 39124 1775 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 39124 1775 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 39205 1775 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 39205 1775 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 39286 1775 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 39286 1775 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 39367 1775 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 39367 1775 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 39448 1775 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 39448 1775 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1711 39529 1775 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1711 39529 1775 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 34780 1763 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 34860 1763 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 34940 1763 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35020 1763 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35100 1763 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35180 1763 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35260 1763 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35340 1763 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35420 1763 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35500 1763 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35580 1763 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35660 1763 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35740 1763 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35820 1763 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35900 1763 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 35980 1763 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 36060 1763 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 36140 1763 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1723 36220 1763 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 4770 1796 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 4770 1796 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 4856 1796 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 4856 1796 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 4942 1796 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 4942 1796 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 5028 1796 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 5028 1796 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 5114 1796 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 5114 1796 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 5200 1796 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 5200 1796 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 5286 1796 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 5286 1796 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 5372 1796 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 5372 1796 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 5458 1796 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 5458 1796 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 5544 1796 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 5544 1796 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1732 5630 1796 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1732 5630 1796 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36289 1855 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36289 1855 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36370 1855 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36370 1855 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36451 1855 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36451 1855 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36532 1855 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36532 1855 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36613 1855 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36613 1855 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36694 1855 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36694 1855 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36775 1855 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36775 1855 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36856 1855 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36856 1855 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 36937 1855 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 36937 1855 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37018 1855 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37018 1855 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37099 1855 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37099 1855 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37180 1855 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37180 1855 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37261 1855 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37261 1855 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37342 1855 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37342 1855 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37423 1855 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37423 1855 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37504 1855 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37504 1855 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37585 1855 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37585 1855 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37666 1855 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37666 1855 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37747 1855 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37747 1855 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37828 1855 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37828 1855 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37909 1855 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37909 1855 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 37990 1855 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 37990 1855 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38071 1855 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38071 1855 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38152 1855 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38152 1855 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38233 1855 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38233 1855 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38314 1855 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38314 1855 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38395 1855 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38395 1855 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38476 1855 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38476 1855 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38557 1855 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38557 1855 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38638 1855 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38638 1855 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38719 1855 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38719 1855 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38800 1855 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38800 1855 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38881 1855 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38881 1855 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 38962 1855 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 38962 1855 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 39043 1855 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 39043 1855 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 39124 1855 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 39124 1855 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 39205 1855 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 39205 1855 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 39286 1855 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 39286 1855 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 39367 1855 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 39367 1855 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 39448 1855 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 39448 1855 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1791 39529 1855 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1791 39529 1855 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 34780 1843 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 34860 1843 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 34940 1843 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35020 1843 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35100 1843 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35180 1843 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35260 1843 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35340 1843 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35420 1843 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35500 1843 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35580 1843 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35660 1843 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35740 1843 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35820 1843 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35900 1843 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 35980 1843 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 36060 1843 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 36140 1843 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1803 36220 1843 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 4770 1877 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 4770 1877 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 4856 1877 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 4856 1877 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 4942 1877 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 4942 1877 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 5028 1877 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 5028 1877 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 5114 1877 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 5114 1877 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 5200 1877 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 5200 1877 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 5286 1877 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 5286 1877 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 5372 1877 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 5372 1877 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 5458 1877 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 5458 1877 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 5544 1877 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 5544 1877 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1813 5630 1877 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1813 5630 1877 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36289 1935 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36289 1935 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36370 1935 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36370 1935 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36451 1935 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36451 1935 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36532 1935 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36532 1935 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36613 1935 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36613 1935 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36694 1935 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36694 1935 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36775 1935 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36775 1935 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36856 1935 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36856 1935 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 36937 1935 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 36937 1935 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37018 1935 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37018 1935 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37099 1935 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37099 1935 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37180 1935 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37180 1935 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37261 1935 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37261 1935 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37342 1935 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37342 1935 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37423 1935 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37423 1935 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37504 1935 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37504 1935 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37585 1935 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37585 1935 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37666 1935 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37666 1935 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37747 1935 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37747 1935 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37828 1935 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37828 1935 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37909 1935 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37909 1935 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 37990 1935 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 37990 1935 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38071 1935 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38071 1935 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38152 1935 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38152 1935 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38233 1935 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38233 1935 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38314 1935 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38314 1935 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38395 1935 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38395 1935 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38476 1935 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38476 1935 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38557 1935 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38557 1935 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38638 1935 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38638 1935 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38719 1935 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38719 1935 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38800 1935 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38800 1935 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38881 1935 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38881 1935 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 38962 1935 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 38962 1935 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 39043 1935 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 39043 1935 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 39124 1935 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 39124 1935 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 39205 1935 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 39205 1935 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 39286 1935 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 39286 1935 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 39367 1935 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 39367 1935 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 39448 1935 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 39448 1935 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1871 39529 1935 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1871 39529 1935 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 34780 1923 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 34860 1923 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 34940 1923 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35020 1923 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35100 1923 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35180 1923 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35260 1923 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35340 1923 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35420 1923 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35500 1923 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35580 1923 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35660 1923 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35740 1923 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35820 1923 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35900 1923 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 35980 1923 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 36060 1923 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 36140 1923 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1883 36220 1923 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 4770 1958 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 4770 1958 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 4856 1958 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 4856 1958 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 4942 1958 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 4942 1958 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 5028 1958 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 5028 1958 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 5114 1958 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 5114 1958 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 5200 1958 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 5200 1958 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 5286 1958 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 5286 1958 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 5372 1958 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 5372 1958 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 5458 1958 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 5458 1958 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 5544 1958 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 5544 1958 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1894 5630 1958 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1894 5630 1958 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36289 2015 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36289 2015 36353 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36370 2015 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36370 2015 36434 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36451 2015 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36451 2015 36515 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36532 2015 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36532 2015 36596 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36613 2015 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36613 2015 36677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36694 2015 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36694 2015 36758 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36775 2015 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36775 2015 36839 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36856 2015 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36856 2015 36920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 36937 2015 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 36937 2015 37001 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37018 2015 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37018 2015 37082 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37099 2015 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37099 2015 37163 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37180 2015 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37180 2015 37244 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37261 2015 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37261 2015 37325 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37342 2015 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37342 2015 37406 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37423 2015 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37423 2015 37487 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37504 2015 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37504 2015 37568 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37585 2015 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37585 2015 37649 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37666 2015 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37666 2015 37730 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37747 2015 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37747 2015 37811 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37828 2015 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37828 2015 37892 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37909 2015 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37909 2015 37973 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 37990 2015 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 37990 2015 38054 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38071 2015 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38071 2015 38135 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38152 2015 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38152 2015 38216 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38233 2015 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38233 2015 38297 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38314 2015 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38314 2015 38378 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38395 2015 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38395 2015 38459 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38476 2015 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38476 2015 38540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38557 2015 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38557 2015 38621 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38638 2015 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38638 2015 38702 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38719 2015 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38719 2015 38783 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38800 2015 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38800 2015 38864 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38881 2015 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38881 2015 38945 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 38962 2015 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 38962 2015 39026 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 39043 2015 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 39043 2015 39107 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 39124 2015 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 39124 2015 39188 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 39205 2015 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 39205 2015 39269 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 39286 2015 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 39286 2015 39350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 39367 2015 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 39367 2015 39431 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 39448 2015 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 39448 2015 39512 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1951 39529 2015 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1951 39529 2015 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 34780 2003 34820 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 34860 2003 34900 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 34940 2003 34980 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35020 2003 35060 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35100 2003 35140 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35180 2003 35220 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35260 2003 35300 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35340 2003 35380 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35420 2003 35460 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35500 2003 35540 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35580 2003 35620 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35660 2003 35700 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35740 2003 35780 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35820 2003 35860 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35900 2003 35940 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 35980 2003 36020 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 36060 2003 36100 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 36140 2003 36180 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1963 36220 2003 36260 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 4770 2039 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 4770 2039 4834 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 4856 2039 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 4856 2039 4920 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 4942 2039 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 4942 2039 5006 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 5028 2039 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 5028 2039 5092 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 5114 2039 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 5114 2039 5178 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 5200 2039 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 5200 2039 5264 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 5286 2039 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 5286 2039 5350 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 5372 2039 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 5372 2039 5436 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 5458 2039 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 5458 2039 5522 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 5544 2039 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 5544 2039 5608 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 1975 5630 2039 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal3 s 1975 5630 2039 5694 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 106 11250 170 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11250 170 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11332 170 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11332 170 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11414 170 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11414 170 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11496 170 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11496 170 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11578 170 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11578 170 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11660 170 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11660 170 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11742 170 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11742 170 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11824 170 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11824 170 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11906 170 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11906 170 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 11988 170 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 11988 170 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 106 12070 170 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 106 12070 170 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11250 252 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11250 252 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11332 252 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11332 252 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11414 252 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11414 252 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11496 252 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11496 252 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11578 252 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11578 252 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11660 252 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11660 252 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11742 252 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11742 252 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11824 252 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11824 252 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11906 252 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11906 252 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 11988 252 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 11988 252 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 188 12070 252 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 188 12070 252 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11250 334 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11250 334 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11332 334 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11332 334 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11414 334 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11414 334 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11496 334 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11496 334 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11578 334 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11578 334 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11660 334 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11660 334 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11742 334 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11742 334 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11824 334 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11824 334 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11906 334 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11906 334 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 11988 334 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 11988 334 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 270 12070 334 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 270 12070 334 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11250 416 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11250 416 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11332 416 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11332 416 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11414 416 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11414 416 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11496 416 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11496 416 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11578 416 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11578 416 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11660 416 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11660 416 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11742 416 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11742 416 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11824 416 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11824 416 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11906 416 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11906 416 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 11988 416 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 11988 416 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 352 12070 416 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 352 12070 416 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11250 2120 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11250 2120 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11332 2120 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11332 2120 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11414 2120 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11414 2120 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11496 2120 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11496 2120 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11578 2120 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11578 2120 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11660 2120 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11660 2120 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11742 2120 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11742 2120 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11824 2120 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11824 2120 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11906 2120 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11906 2120 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 11988 2120 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 11988 2120 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2056 12070 2120 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2056 12070 2120 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11250 2201 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11250 2201 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11332 2201 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11332 2201 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11414 2201 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11414 2201 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11496 2201 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11496 2201 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11578 2201 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11578 2201 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11660 2201 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11660 2201 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11742 2201 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11742 2201 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11824 2201 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11824 2201 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11906 2201 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11906 2201 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 11988 2201 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 11988 2201 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2137 12070 2201 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2137 12070 2201 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11250 2282 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11250 2282 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11332 2282 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11332 2282 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11414 2282 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11414 2282 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11496 2282 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11496 2282 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11578 2282 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11578 2282 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11660 2282 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11660 2282 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11742 2282 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11742 2282 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11824 2282 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11824 2282 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11906 2282 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11906 2282 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 11988 2282 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 11988 2282 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2218 12070 2282 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2218 12070 2282 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11250 2363 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11250 2363 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11332 2363 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11332 2363 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11414 2363 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11414 2363 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11496 2363 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11496 2363 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11578 2363 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11578 2363 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11660 2363 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11660 2363 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11742 2363 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11742 2363 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11824 2363 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11824 2363 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11906 2363 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11906 2363 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 11988 2363 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 11988 2363 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2299 12070 2363 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2299 12070 2363 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11250 2444 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11250 2444 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11332 2444 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11332 2444 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11414 2444 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11414 2444 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11496 2444 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11496 2444 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11578 2444 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11578 2444 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11660 2444 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11660 2444 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11742 2444 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11742 2444 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11824 2444 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11824 2444 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11906 2444 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11906 2444 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 11988 2444 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 11988 2444 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2380 12070 2444 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2380 12070 2444 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11250 2525 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11250 2525 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11332 2525 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11332 2525 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11414 2525 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11414 2525 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11496 2525 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11496 2525 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11578 2525 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11578 2525 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11660 2525 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11660 2525 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11742 2525 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11742 2525 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11824 2525 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11824 2525 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11906 2525 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11906 2525 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 11988 2525 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 11988 2525 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2461 12070 2525 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2461 12070 2525 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11250 2606 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11250 2606 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11332 2606 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11332 2606 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11414 2606 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11414 2606 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11496 2606 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11496 2606 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11578 2606 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11578 2606 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11660 2606 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11660 2606 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11742 2606 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11742 2606 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11824 2606 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11824 2606 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11906 2606 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11906 2606 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 11988 2606 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 11988 2606 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2542 12070 2606 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2542 12070 2606 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11250 2687 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11250 2687 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11332 2687 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11332 2687 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11414 2687 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11414 2687 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11496 2687 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11496 2687 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11578 2687 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11578 2687 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11660 2687 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11660 2687 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11742 2687 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11742 2687 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11824 2687 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11824 2687 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11906 2687 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11906 2687 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 11988 2687 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 11988 2687 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2623 12070 2687 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2623 12070 2687 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11250 2768 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11250 2768 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11332 2768 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11332 2768 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11414 2768 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11414 2768 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11496 2768 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11496 2768 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11578 2768 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11578 2768 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11660 2768 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11660 2768 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11742 2768 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11742 2768 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11824 2768 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11824 2768 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11906 2768 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11906 2768 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 11988 2768 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 11988 2768 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2704 12070 2768 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2704 12070 2768 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11250 2849 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11250 2849 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11332 2849 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11332 2849 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11414 2849 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11414 2849 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11496 2849 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11496 2849 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11578 2849 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11578 2849 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11660 2849 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11660 2849 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11742 2849 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11742 2849 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11824 2849 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11824 2849 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11906 2849 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11906 2849 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 11988 2849 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 11988 2849 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2785 12070 2849 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2785 12070 2849 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11250 2930 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11250 2930 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11332 2930 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11332 2930 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11414 2930 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11414 2930 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11496 2930 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11496 2930 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11578 2930 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11578 2930 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11660 2930 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11660 2930 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11742 2930 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11742 2930 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11824 2930 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11824 2930 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11906 2930 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11906 2930 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 11988 2930 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 11988 2930 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2866 12070 2930 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2866 12070 2930 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11250 3011 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11250 3011 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11332 3011 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11332 3011 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11414 3011 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11414 3011 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11496 3011 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11496 3011 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11578 3011 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11578 3011 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11660 3011 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11660 3011 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11742 3011 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11742 3011 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11824 3011 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11824 3011 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11906 3011 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11906 3011 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 11988 3011 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 11988 3011 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 2947 12070 3011 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 2947 12070 3011 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11250 3092 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11250 3092 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11332 3092 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11332 3092 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11414 3092 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11414 3092 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11496 3092 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11496 3092 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11578 3092 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11578 3092 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11660 3092 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11660 3092 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11742 3092 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11742 3092 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11824 3092 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11824 3092 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11906 3092 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11906 3092 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 11988 3092 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 11988 3092 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3028 12070 3092 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3028 12070 3092 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11250 3173 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11250 3173 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11332 3173 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11332 3173 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11414 3173 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11414 3173 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11496 3173 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11496 3173 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11578 3173 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11578 3173 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11660 3173 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11660 3173 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11742 3173 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11742 3173 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11824 3173 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11824 3173 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11906 3173 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11906 3173 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 11988 3173 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 11988 3173 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3109 12070 3173 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3109 12070 3173 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11250 3254 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11250 3254 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11332 3254 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11332 3254 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11414 3254 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11414 3254 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11496 3254 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11496 3254 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11578 3254 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11578 3254 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11660 3254 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11660 3254 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11742 3254 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11742 3254 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11824 3254 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11824 3254 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11906 3254 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11906 3254 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 11988 3254 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 11988 3254 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3190 12070 3254 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3190 12070 3254 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11250 3335 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11250 3335 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11332 3335 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11332 3335 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11414 3335 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11414 3335 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11496 3335 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11496 3335 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11578 3335 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11578 3335 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11660 3335 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11660 3335 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11742 3335 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11742 3335 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11824 3335 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11824 3335 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11906 3335 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11906 3335 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 11988 3335 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 11988 3335 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3271 12070 3335 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3271 12070 3335 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11250 3416 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11250 3416 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11332 3416 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11332 3416 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11414 3416 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11414 3416 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11496 3416 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11496 3416 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11578 3416 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11578 3416 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11660 3416 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11660 3416 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11742 3416 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11742 3416 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11824 3416 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11824 3416 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11906 3416 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11906 3416 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 11988 3416 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 11988 3416 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3352 12070 3416 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3352 12070 3416 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11250 3497 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11250 3497 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11332 3497 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11332 3497 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11414 3497 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11414 3497 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11496 3497 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11496 3497 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11578 3497 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11578 3497 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11660 3497 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11660 3497 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11742 3497 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11742 3497 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11824 3497 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11824 3497 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11906 3497 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11906 3497 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 11988 3497 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 11988 3497 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3433 12070 3497 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3433 12070 3497 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11250 3578 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11250 3578 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11332 3578 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11332 3578 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11414 3578 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11414 3578 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11496 3578 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11496 3578 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11578 3578 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11578 3578 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11660 3578 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11660 3578 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11742 3578 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11742 3578 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11824 3578 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11824 3578 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11906 3578 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11906 3578 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 11988 3578 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 11988 3578 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3514 12070 3578 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3514 12070 3578 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11250 3659 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11250 3659 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11332 3659 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11332 3659 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11414 3659 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11414 3659 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11496 3659 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11496 3659 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11578 3659 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11578 3659 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11660 3659 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11660 3659 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11742 3659 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11742 3659 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11824 3659 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11824 3659 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11906 3659 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11906 3659 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 11988 3659 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 11988 3659 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3595 12070 3659 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3595 12070 3659 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11250 3740 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11250 3740 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11332 3740 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11332 3740 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11414 3740 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11414 3740 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11496 3740 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11496 3740 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11578 3740 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11578 3740 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11660 3740 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11660 3740 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11742 3740 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11742 3740 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11824 3740 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11824 3740 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11906 3740 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11906 3740 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 11988 3740 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 11988 3740 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3676 12070 3740 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3676 12070 3740 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11250 3821 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11250 3821 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11332 3821 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11332 3821 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11414 3821 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11414 3821 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11496 3821 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11496 3821 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11578 3821 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11578 3821 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11660 3821 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11660 3821 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11742 3821 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11742 3821 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11824 3821 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11824 3821 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11906 3821 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11906 3821 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 11988 3821 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 11988 3821 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3757 12070 3821 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3757 12070 3821 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11250 3902 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11250 3902 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11332 3902 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11332 3902 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11414 3902 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11414 3902 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11496 3902 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11496 3902 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11578 3902 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11578 3902 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11660 3902 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11660 3902 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11742 3902 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11742 3902 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11824 3902 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11824 3902 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11906 3902 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11906 3902 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 11988 3902 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 11988 3902 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3838 12070 3902 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3838 12070 3902 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11250 3983 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11250 3983 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11332 3983 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11332 3983 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11414 3983 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11414 3983 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11496 3983 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11496 3983 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11578 3983 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11578 3983 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11660 3983 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11660 3983 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11742 3983 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11742 3983 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11824 3983 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11824 3983 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11906 3983 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11906 3983 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 11988 3983 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 11988 3983 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 3919 12070 3983 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 3919 12070 3983 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11250 498 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11250 498 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11332 498 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11332 498 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11414 498 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11414 498 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11496 498 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11496 498 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11578 498 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11578 498 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11660 498 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11660 498 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11742 498 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11742 498 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11824 498 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11824 498 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11906 498 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11906 498 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 11988 498 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 11988 498 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 434 12070 498 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 434 12070 498 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11250 580 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11250 580 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11332 580 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11332 580 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11414 580 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11414 580 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11496 580 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11496 580 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11578 580 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11578 580 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11660 580 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11660 580 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11742 580 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11742 580 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11824 580 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11824 580 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11906 580 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11906 580 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 11988 580 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 11988 580 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 516 12070 580 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 516 12070 580 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11250 662 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11250 662 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11332 662 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11332 662 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11414 662 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11414 662 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11496 662 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11496 662 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11578 662 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11578 662 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11660 662 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11660 662 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11742 662 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11742 662 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11824 662 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11824 662 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11906 662 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11906 662 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 11988 662 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 11988 662 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 598 12070 662 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 598 12070 662 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11250 4064 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11250 4064 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11332 4064 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11332 4064 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11414 4064 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11414 4064 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11496 4064 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11496 4064 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11578 4064 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11578 4064 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11660 4064 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11660 4064 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11742 4064 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11742 4064 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11824 4064 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11824 4064 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11906 4064 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11906 4064 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 11988 4064 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 11988 4064 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4000 12070 4064 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4000 12070 4064 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11250 4145 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11250 4145 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11332 4145 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11332 4145 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11414 4145 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11414 4145 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11496 4145 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11496 4145 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11578 4145 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11578 4145 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11660 4145 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11660 4145 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11742 4145 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11742 4145 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11824 4145 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11824 4145 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11906 4145 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11906 4145 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 11988 4145 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 11988 4145 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4081 12070 4145 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4081 12070 4145 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11250 4226 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11250 4226 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11332 4226 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11332 4226 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11414 4226 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11414 4226 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11496 4226 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11496 4226 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11578 4226 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11578 4226 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11660 4226 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11660 4226 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11742 4226 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11742 4226 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11824 4226 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11824 4226 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11906 4226 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11906 4226 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 11988 4226 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 11988 4226 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4162 12070 4226 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4162 12070 4226 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11250 4307 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11250 4307 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11332 4307 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11332 4307 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11414 4307 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11414 4307 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11496 4307 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11496 4307 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11578 4307 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11578 4307 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11660 4307 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11660 4307 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11742 4307 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11742 4307 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11824 4307 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11824 4307 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11906 4307 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11906 4307 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 11988 4307 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 11988 4307 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4243 12070 4307 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4243 12070 4307 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11250 4388 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11250 4388 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11332 4388 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11332 4388 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11414 4388 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11414 4388 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11496 4388 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11496 4388 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11578 4388 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11578 4388 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11660 4388 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11660 4388 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11742 4388 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11742 4388 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11824 4388 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11824 4388 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11906 4388 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11906 4388 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 11988 4388 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 11988 4388 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4324 12070 4388 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4324 12070 4388 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11250 4469 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11250 4469 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11332 4469 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11332 4469 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11414 4469 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11414 4469 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11496 4469 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11496 4469 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11578 4469 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11578 4469 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11660 4469 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11660 4469 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11742 4469 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11742 4469 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11824 4469 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11824 4469 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11906 4469 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11906 4469 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 11988 4469 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 11988 4469 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4405 12070 4469 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4405 12070 4469 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11250 4550 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11250 4550 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11332 4550 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11332 4550 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11414 4550 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11414 4550 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11496 4550 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11496 4550 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11578 4550 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11578 4550 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11660 4550 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11660 4550 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11742 4550 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11742 4550 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11824 4550 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11824 4550 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11906 4550 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11906 4550 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 11988 4550 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 11988 4550 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4486 12070 4550 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4486 12070 4550 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11250 4631 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11250 4631 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11332 4631 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11332 4631 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11414 4631 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11414 4631 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11496 4631 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11496 4631 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11578 4631 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11578 4631 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11660 4631 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11660 4631 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11742 4631 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11742 4631 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11824 4631 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11824 4631 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11906 4631 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11906 4631 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 11988 4631 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 11988 4631 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4567 12070 4631 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4567 12070 4631 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11250 4712 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11250 4712 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11332 4712 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11332 4712 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11414 4712 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11414 4712 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11496 4712 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11496 4712 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11578 4712 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11578 4712 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11660 4712 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11660 4712 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11742 4712 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11742 4712 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11824 4712 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11824 4712 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11906 4712 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11906 4712 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 11988 4712 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 11988 4712 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4648 12070 4712 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4648 12070 4712 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11250 4793 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11250 4793 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11332 4793 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11332 4793 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11414 4793 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11414 4793 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11496 4793 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11496 4793 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11578 4793 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11578 4793 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11660 4793 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11660 4793 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11742 4793 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11742 4793 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11824 4793 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11824 4793 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11906 4793 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11906 4793 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 11988 4793 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 11988 4793 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4729 12070 4793 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4729 12070 4793 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11250 4874 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11250 4874 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11332 4874 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11332 4874 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11414 4874 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11414 4874 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11496 4874 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11496 4874 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11578 4874 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11578 4874 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11660 4874 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11660 4874 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11742 4874 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11742 4874 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11824 4874 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11824 4874 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11906 4874 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11906 4874 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 11988 4874 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 11988 4874 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 4810 12070 4874 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 4810 12070 4874 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11250 743 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11250 743 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11332 743 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11332 743 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11414 743 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11414 743 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11496 743 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11496 743 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11578 743 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11578 743 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11660 743 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11660 743 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11742 743 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11742 743 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11824 743 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11824 743 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11906 743 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11906 743 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 11988 743 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 11988 743 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 679 12070 743 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 679 12070 743 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11250 824 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11250 824 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11332 824 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11332 824 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11414 824 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11414 824 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11496 824 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11496 824 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11578 824 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11578 824 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11660 824 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11660 824 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11742 824 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11742 824 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11824 824 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11824 824 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11906 824 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11906 824 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 11988 824 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 11988 824 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 760 12070 824 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 760 12070 824 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11250 905 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11250 905 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11332 905 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11332 905 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11414 905 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11414 905 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11496 905 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11496 905 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11578 905 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11578 905 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11660 905 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11660 905 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11742 905 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11742 905 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11824 905 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11824 905 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11906 905 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11906 905 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 11988 905 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 11988 905 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 841 12070 905 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 841 12070 905 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11250 986 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11250 986 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11332 986 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11332 986 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11414 986 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11414 986 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11496 986 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11496 986 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11578 986 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11578 986 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11660 986 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11660 986 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11742 986 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11742 986 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11824 986 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11824 986 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11906 986 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11906 986 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 11988 986 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 11988 986 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 922 12070 986 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 922 12070 986 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11250 1067 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11250 1067 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11332 1067 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11332 1067 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11414 1067 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11414 1067 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11496 1067 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11496 1067 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11578 1067 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11578 1067 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11660 1067 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11660 1067 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11742 1067 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11742 1067 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11824 1067 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11824 1067 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11906 1067 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11906 1067 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 11988 1067 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 11988 1067 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1003 12070 1067 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1003 12070 1067 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11250 1148 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11250 1148 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11332 1148 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11332 1148 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11414 1148 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11414 1148 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11496 1148 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11496 1148 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11578 1148 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11578 1148 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11660 1148 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11660 1148 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11742 1148 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11742 1148 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11824 1148 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11824 1148 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11906 1148 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11906 1148 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 11988 1148 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 11988 1148 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1084 12070 1148 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1084 12070 1148 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11250 1229 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11250 1229 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11332 1229 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11332 1229 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11414 1229 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11414 1229 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11496 1229 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11496 1229 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11578 1229 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11578 1229 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11660 1229 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11660 1229 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11742 1229 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11742 1229 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11824 1229 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11824 1229 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11906 1229 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11906 1229 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 11988 1229 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 11988 1229 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1165 12070 1229 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1165 12070 1229 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11250 10221 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11250 10221 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11332 10221 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11332 10221 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11414 10221 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11414 10221 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11496 10221 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11496 10221 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11578 10221 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11578 10221 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11660 10221 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11660 10221 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11742 10221 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11742 10221 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11824 10221 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11824 10221 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11906 10221 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11906 10221 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 11988 10221 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 11988 10221 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10157 12070 10221 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10157 12070 10221 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11250 10303 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11250 10303 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11332 10303 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11332 10303 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11414 10303 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11414 10303 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11496 10303 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11496 10303 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11578 10303 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11578 10303 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11660 10303 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11660 10303 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11742 10303 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11742 10303 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11824 10303 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11824 10303 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11906 10303 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11906 10303 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 11988 10303 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 11988 10303 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10239 12070 10303 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10239 12070 10303 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11250 10385 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11250 10385 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11332 10385 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11332 10385 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11414 10385 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11414 10385 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11496 10385 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11496 10385 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11578 10385 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11578 10385 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11660 10385 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11660 10385 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11742 10385 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11742 10385 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11824 10385 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11824 10385 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11906 10385 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11906 10385 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 11988 10385 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 11988 10385 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10321 12070 10385 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10321 12070 10385 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11250 10467 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11250 10467 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11332 10467 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11332 10467 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11414 10467 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11414 10467 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11496 10467 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11496 10467 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11578 10467 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11578 10467 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11660 10467 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11660 10467 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11742 10467 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11742 10467 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11824 10467 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11824 10467 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11906 10467 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11906 10467 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 11988 10467 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 11988 10467 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10403 12070 10467 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10403 12070 10467 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11250 10549 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11250 10549 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11332 10549 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11332 10549 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11414 10549 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11414 10549 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11496 10549 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11496 10549 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11578 10549 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11578 10549 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11660 10549 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11660 10549 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11742 10549 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11742 10549 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11824 10549 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11824 10549 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11906 10549 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11906 10549 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 11988 10549 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 11988 10549 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10485 12070 10549 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10485 12070 10549 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11250 10631 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11250 10631 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11332 10631 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11332 10631 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11414 10631 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11414 10631 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11496 10631 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11496 10631 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11578 10631 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11578 10631 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11660 10631 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11660 10631 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11742 10631 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11742 10631 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11824 10631 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11824 10631 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11906 10631 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11906 10631 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 11988 10631 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 11988 10631 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10567 12070 10631 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10567 12070 10631 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11250 10713 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11250 10713 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11332 10713 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11332 10713 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11414 10713 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11414 10713 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11496 10713 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11496 10713 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11578 10713 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11578 10713 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11660 10713 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11660 10713 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11742 10713 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11742 10713 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11824 10713 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11824 10713 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11906 10713 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11906 10713 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 11988 10713 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 11988 10713 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10649 12070 10713 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10649 12070 10713 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11250 10795 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11250 10795 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11332 10795 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11332 10795 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11414 10795 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11414 10795 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11496 10795 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11496 10795 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11578 10795 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11578 10795 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11660 10795 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11660 10795 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11742 10795 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11742 10795 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11824 10795 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11824 10795 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11906 10795 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11906 10795 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 11988 10795 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 11988 10795 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10731 12070 10795 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10731 12070 10795 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11250 10877 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11250 10877 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11332 10877 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11332 10877 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11414 10877 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11414 10877 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11496 10877 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11496 10877 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11578 10877 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11578 10877 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11660 10877 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11660 10877 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11742 10877 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11742 10877 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11824 10877 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11824 10877 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11906 10877 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11906 10877 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 11988 10877 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 11988 10877 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10813 12070 10877 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10813 12070 10877 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11250 10959 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11250 10959 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11332 10959 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11332 10959 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11414 10959 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11414 10959 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11496 10959 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11496 10959 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11578 10959 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11578 10959 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11660 10959 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11660 10959 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11742 10959 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11742 10959 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11824 10959 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11824 10959 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11906 10959 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11906 10959 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 11988 10959 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 11988 10959 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10895 12070 10959 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10895 12070 10959 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11250 11041 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11250 11041 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11332 11041 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11332 11041 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11414 11041 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11414 11041 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11496 11041 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11496 11041 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11578 11041 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11578 11041 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11660 11041 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11660 11041 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11742 11041 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11742 11041 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11824 11041 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11824 11041 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11906 11041 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11906 11041 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 11988 11041 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 11988 11041 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 10977 12070 11041 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 10977 12070 11041 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11250 11123 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11250 11123 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11332 11123 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11332 11123 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11414 11123 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11414 11123 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11496 11123 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11496 11123 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11578 11123 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11578 11123 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11660 11123 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11660 11123 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11742 11123 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11742 11123 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11824 11123 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11824 11123 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11906 11123 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11906 11123 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 11988 11123 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 11988 11123 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11059 12070 11123 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11059 12070 11123 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11250 11205 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11250 11205 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11332 11205 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11332 11205 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11414 11205 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11414 11205 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11496 11205 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11496 11205 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11578 11205 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11578 11205 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11660 11205 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11660 11205 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11742 11205 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11742 11205 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11824 11205 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11824 11205 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11906 11205 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11906 11205 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 11988 11205 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 11988 11205 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11141 12070 11205 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11141 12070 11205 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11250 11287 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11250 11287 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11332 11287 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11332 11287 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11414 11287 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11414 11287 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11496 11287 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11496 11287 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11578 11287 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11578 11287 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11660 11287 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11660 11287 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11742 11287 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11742 11287 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11824 11287 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11824 11287 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11906 11287 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11906 11287 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 11988 11287 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 11988 11287 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11223 12070 11287 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11223 12070 11287 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11250 11369 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11250 11369 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11332 11369 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11332 11369 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11414 11369 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11414 11369 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11496 11369 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11496 11369 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11578 11369 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11578 11369 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11660 11369 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11660 11369 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11742 11369 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11742 11369 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11824 11369 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11824 11369 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11906 11369 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11906 11369 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 11988 11369 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 11988 11369 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11305 12070 11369 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11305 12070 11369 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11250 11450 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11250 11450 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11332 11450 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11332 11450 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11414 11450 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11414 11450 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11496 11450 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11496 11450 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11578 11450 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11578 11450 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11660 11450 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11660 11450 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11742 11450 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11742 11450 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11824 11450 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11824 11450 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11906 11450 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11906 11450 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 11988 11450 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 11988 11450 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11386 12070 11450 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11386 12070 11450 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11250 11531 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11250 11531 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11332 11531 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11332 11531 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11414 11531 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11414 11531 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11496 11531 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11496 11531 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11578 11531 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11578 11531 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11660 11531 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11660 11531 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11742 11531 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11742 11531 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11824 11531 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11824 11531 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11906 11531 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11906 11531 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 11988 11531 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 11988 11531 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11467 12070 11531 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11467 12070 11531 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11250 11612 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11250 11612 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11332 11612 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11332 11612 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11414 11612 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11414 11612 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11496 11612 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11496 11612 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11578 11612 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11578 11612 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11660 11612 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11660 11612 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11742 11612 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11742 11612 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11824 11612 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11824 11612 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11906 11612 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11906 11612 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 11988 11612 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 11988 11612 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11548 12070 11612 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11548 12070 11612 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11250 11693 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11250 11693 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11332 11693 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11332 11693 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11414 11693 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11414 11693 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11496 11693 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11496 11693 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11578 11693 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11578 11693 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11660 11693 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11660 11693 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11742 11693 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11742 11693 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11824 11693 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11824 11693 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11906 11693 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11906 11693 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 11988 11693 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 11988 11693 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11629 12070 11693 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11629 12070 11693 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11250 11774 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11250 11774 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11332 11774 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11332 11774 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11414 11774 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11414 11774 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11496 11774 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11496 11774 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11578 11774 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11578 11774 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11660 11774 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11660 11774 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11742 11774 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11742 11774 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11824 11774 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11824 11774 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11906 11774 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11906 11774 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 11988 11774 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 11988 11774 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11710 12070 11774 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11710 12070 11774 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11250 11855 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11250 11855 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11332 11855 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11332 11855 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11414 11855 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11414 11855 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11496 11855 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11496 11855 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11578 11855 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11578 11855 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11660 11855 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11660 11855 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11742 11855 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11742 11855 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11824 11855 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11824 11855 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11906 11855 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11906 11855 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 11988 11855 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 11988 11855 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11791 12070 11855 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11791 12070 11855 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11250 11936 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11250 11936 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11332 11936 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11332 11936 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11414 11936 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11414 11936 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11496 11936 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11496 11936 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11578 11936 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11578 11936 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11660 11936 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11660 11936 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11742 11936 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11742 11936 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11824 11936 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11824 11936 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11906 11936 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11906 11936 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 11988 11936 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 11988 11936 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11872 12070 11936 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11872 12070 11936 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11250 12017 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11250 12017 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11332 12017 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11332 12017 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11414 12017 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11414 12017 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11496 12017 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11496 12017 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11578 12017 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11578 12017 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11660 12017 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11660 12017 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11742 12017 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11742 12017 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11824 12017 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11824 12017 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11906 12017 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11906 12017 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 11988 12017 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 11988 12017 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 11953 12070 12017 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 11953 12070 12017 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11250 1310 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11250 1310 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11332 1310 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11332 1310 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11414 1310 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11414 1310 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11496 1310 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11496 1310 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11578 1310 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11578 1310 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11660 1310 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11660 1310 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11742 1310 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11742 1310 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11824 1310 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11824 1310 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11906 1310 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11906 1310 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 11988 1310 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 11988 1310 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1246 12070 1310 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1246 12070 1310 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11250 1391 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11250 1391 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11332 1391 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11332 1391 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11414 1391 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11414 1391 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11496 1391 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11496 1391 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11578 1391 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11578 1391 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11660 1391 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11660 1391 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11742 1391 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11742 1391 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11824 1391 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11824 1391 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11906 1391 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11906 1391 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 11988 1391 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 11988 1391 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1327 12070 1391 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1327 12070 1391 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11250 12098 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11250 12098 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11332 12098 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11332 12098 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11414 12098 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11414 12098 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11496 12098 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11496 12098 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11578 12098 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11578 12098 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11660 12098 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11660 12098 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11742 12098 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11742 12098 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11824 12098 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11824 12098 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11906 12098 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11906 12098 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 11988 12098 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 11988 12098 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12034 12070 12098 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12034 12070 12098 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11250 12179 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11250 12179 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11332 12179 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11332 12179 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11414 12179 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11414 12179 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11496 12179 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11496 12179 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11578 12179 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11578 12179 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11660 12179 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11660 12179 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11742 12179 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11742 12179 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11824 12179 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11824 12179 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11906 12179 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11906 12179 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 11988 12179 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 11988 12179 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12115 12070 12179 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12115 12070 12179 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11250 12260 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11250 12260 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11332 12260 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11332 12260 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11414 12260 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11414 12260 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11496 12260 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11496 12260 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11578 12260 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11578 12260 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11660 12260 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11660 12260 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11742 12260 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11742 12260 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11824 12260 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11824 12260 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11906 12260 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11906 12260 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 11988 12260 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 11988 12260 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12196 12070 12260 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12196 12070 12260 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11250 12341 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11250 12341 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11332 12341 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11332 12341 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11414 12341 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11414 12341 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11496 12341 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11496 12341 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11578 12341 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11578 12341 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11660 12341 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11660 12341 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11742 12341 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11742 12341 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11824 12341 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11824 12341 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11906 12341 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11906 12341 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 11988 12341 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 11988 12341 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12277 12070 12341 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12277 12070 12341 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11250 12422 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11250 12422 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11332 12422 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11332 12422 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11414 12422 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11414 12422 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11496 12422 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11496 12422 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11578 12422 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11578 12422 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11660 12422 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11660 12422 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11742 12422 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11742 12422 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11824 12422 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11824 12422 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11906 12422 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11906 12422 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 11988 12422 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 11988 12422 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12358 12070 12422 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12358 12070 12422 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11250 12503 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11250 12503 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11332 12503 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11332 12503 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11414 12503 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11414 12503 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11496 12503 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11496 12503 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11578 12503 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11578 12503 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11660 12503 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11660 12503 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11742 12503 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11742 12503 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11824 12503 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11824 12503 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11906 12503 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11906 12503 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 11988 12503 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 11988 12503 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12439 12070 12503 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12439 12070 12503 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11250 12584 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11250 12584 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11332 12584 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11332 12584 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11414 12584 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11414 12584 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11496 12584 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11496 12584 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11578 12584 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11578 12584 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11660 12584 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11660 12584 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11742 12584 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11742 12584 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11824 12584 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11824 12584 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11906 12584 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11906 12584 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 11988 12584 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 11988 12584 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12520 12070 12584 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12520 12070 12584 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11250 12665 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11250 12665 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11332 12665 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11332 12665 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11414 12665 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11414 12665 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11496 12665 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11496 12665 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11578 12665 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11578 12665 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11660 12665 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11660 12665 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11742 12665 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11742 12665 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11824 12665 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11824 12665 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11906 12665 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11906 12665 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 11988 12665 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 11988 12665 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12601 12070 12665 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12601 12070 12665 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11250 12746 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11250 12746 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11332 12746 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11332 12746 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11414 12746 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11414 12746 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11496 12746 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11496 12746 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11578 12746 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11578 12746 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11660 12746 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11660 12746 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11742 12746 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11742 12746 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11824 12746 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11824 12746 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11906 12746 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11906 12746 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 11988 12746 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 11988 12746 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12682 12070 12746 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12682 12070 12746 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11250 12827 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11250 12827 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11332 12827 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11332 12827 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11414 12827 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11414 12827 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11496 12827 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11496 12827 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11578 12827 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11578 12827 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11660 12827 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11660 12827 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11742 12827 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11742 12827 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11824 12827 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11824 12827 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11906 12827 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11906 12827 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 11988 12827 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 11988 12827 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12763 12070 12827 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12763 12070 12827 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11250 12908 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11250 12908 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11332 12908 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11332 12908 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11414 12908 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11414 12908 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11496 12908 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11496 12908 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11578 12908 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11578 12908 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11660 12908 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11660 12908 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11742 12908 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11742 12908 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11824 12908 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11824 12908 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11906 12908 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11906 12908 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 11988 12908 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 11988 12908 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12844 12070 12908 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12844 12070 12908 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11250 12989 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11250 12989 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11332 12989 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11332 12989 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11414 12989 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11414 12989 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11496 12989 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11496 12989 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11578 12989 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11578 12989 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11660 12989 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11660 12989 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11742 12989 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11742 12989 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11824 12989 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11824 12989 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11906 12989 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11906 12989 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 11988 12989 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 11988 12989 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 12925 12070 12989 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 12925 12070 12989 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11250 13070 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11250 13070 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11332 13070 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11332 13070 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11414 13070 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11414 13070 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11496 13070 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11496 13070 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11578 13070 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11578 13070 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11660 13070 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11660 13070 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11742 13070 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11742 13070 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11824 13070 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11824 13070 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11906 13070 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11906 13070 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 11988 13070 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 11988 13070 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13006 12070 13070 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13006 12070 13070 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11250 13151 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11250 13151 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11332 13151 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11332 13151 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11414 13151 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11414 13151 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11496 13151 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11496 13151 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11578 13151 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11578 13151 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11660 13151 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11660 13151 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11742 13151 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11742 13151 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11824 13151 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11824 13151 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11906 13151 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11906 13151 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 11988 13151 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 11988 13151 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13087 12070 13151 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13087 12070 13151 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11250 13232 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11250 13232 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11332 13232 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11332 13232 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11414 13232 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11414 13232 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11496 13232 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11496 13232 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11578 13232 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11578 13232 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11660 13232 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11660 13232 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11742 13232 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11742 13232 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11824 13232 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11824 13232 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11906 13232 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11906 13232 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 11988 13232 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 11988 13232 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13168 12070 13232 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13168 12070 13232 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11250 13313 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11250 13313 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11332 13313 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11332 13313 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11414 13313 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11414 13313 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11496 13313 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11496 13313 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11578 13313 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11578 13313 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11660 13313 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11660 13313 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11742 13313 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11742 13313 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11824 13313 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11824 13313 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11906 13313 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11906 13313 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 11988 13313 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 11988 13313 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13249 12070 13313 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13249 12070 13313 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11250 13394 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11250 13394 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11332 13394 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11332 13394 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11414 13394 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11414 13394 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11496 13394 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11496 13394 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11578 13394 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11578 13394 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11660 13394 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11660 13394 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11742 13394 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11742 13394 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11824 13394 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11824 13394 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11906 13394 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11906 13394 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 11988 13394 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 11988 13394 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13330 12070 13394 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13330 12070 13394 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11250 13475 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11250 13475 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11332 13475 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11332 13475 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11414 13475 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11414 13475 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11496 13475 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11496 13475 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11578 13475 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11578 13475 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11660 13475 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11660 13475 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11742 13475 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11742 13475 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11824 13475 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11824 13475 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11906 13475 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11906 13475 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 11988 13475 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 11988 13475 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13411 12070 13475 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13411 12070 13475 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11250 13556 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11250 13556 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11332 13556 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11332 13556 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11414 13556 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11414 13556 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11496 13556 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11496 13556 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11578 13556 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11578 13556 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11660 13556 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11660 13556 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11742 13556 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11742 13556 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11824 13556 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11824 13556 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11906 13556 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11906 13556 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 11988 13556 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 11988 13556 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13492 12070 13556 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13492 12070 13556 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11250 13637 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11250 13637 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11332 13637 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11332 13637 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11414 13637 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11414 13637 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11496 13637 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11496 13637 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11578 13637 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11578 13637 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11660 13637 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11660 13637 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11742 13637 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11742 13637 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11824 13637 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11824 13637 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11906 13637 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11906 13637 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 11988 13637 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 11988 13637 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13573 12070 13637 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13573 12070 13637 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11250 13718 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11250 13718 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11332 13718 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11332 13718 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11414 13718 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11414 13718 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11496 13718 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11496 13718 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11578 13718 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11578 13718 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11660 13718 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11660 13718 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11742 13718 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11742 13718 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11824 13718 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11824 13718 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11906 13718 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11906 13718 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 11988 13718 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 11988 13718 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13654 12070 13718 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13654 12070 13718 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11250 13799 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11250 13799 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11332 13799 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11332 13799 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11414 13799 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11414 13799 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11496 13799 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11496 13799 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11578 13799 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11578 13799 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11660 13799 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11660 13799 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11742 13799 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11742 13799 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11824 13799 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11824 13799 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11906 13799 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11906 13799 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 11988 13799 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 11988 13799 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13735 12070 13799 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13735 12070 13799 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11250 13880 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11250 13880 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11332 13880 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11332 13880 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11414 13880 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11414 13880 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11496 13880 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11496 13880 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11578 13880 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11578 13880 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11660 13880 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11660 13880 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11742 13880 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11742 13880 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11824 13880 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11824 13880 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11906 13880 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11906 13880 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 11988 13880 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 11988 13880 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13816 12070 13880 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13816 12070 13880 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11250 13961 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11250 13961 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11332 13961 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11332 13961 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11414 13961 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11414 13961 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11496 13961 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11496 13961 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11578 13961 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11578 13961 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11660 13961 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11660 13961 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11742 13961 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11742 13961 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11824 13961 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11824 13961 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11906 13961 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11906 13961 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 11988 13961 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 11988 13961 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13897 12070 13961 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13897 12070 13961 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11250 14042 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11250 14042 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11332 14042 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11332 14042 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11414 14042 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11414 14042 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11496 14042 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11496 14042 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11578 14042 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11578 14042 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11660 14042 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11660 14042 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11742 14042 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11742 14042 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11824 14042 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11824 14042 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11906 14042 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11906 14042 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 11988 14042 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 11988 14042 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 13978 12070 14042 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 13978 12070 14042 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11250 1472 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11250 1472 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11332 1472 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11332 1472 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11414 1472 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11414 1472 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11496 1472 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11496 1472 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11578 1472 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11578 1472 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11660 1472 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11660 1472 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11742 1472 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11742 1472 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11824 1472 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11824 1472 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11906 1472 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11906 1472 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 11988 1472 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 11988 1472 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1408 12070 1472 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1408 12070 1472 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11250 1553 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11250 1553 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11332 1553 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11332 1553 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11414 1553 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11414 1553 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11496 1553 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11496 1553 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11578 1553 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11578 1553 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11660 1553 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11660 1553 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11742 1553 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11742 1553 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11824 1553 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11824 1553 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11906 1553 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11906 1553 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 11988 1553 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 11988 1553 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1489 12070 1553 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1489 12070 1553 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11250 1634 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11250 1634 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11332 1634 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11332 1634 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11414 1634 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11414 1634 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11496 1634 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11496 1634 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11578 1634 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11578 1634 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11660 1634 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11660 1634 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11742 1634 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11742 1634 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11824 1634 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11824 1634 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11906 1634 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11906 1634 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 11988 1634 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 11988 1634 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1570 12070 1634 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1570 12070 1634 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11250 14123 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11250 14123 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11332 14123 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11332 14123 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11414 14123 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11414 14123 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11496 14123 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11496 14123 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11578 14123 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11578 14123 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11660 14123 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11660 14123 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11742 14123 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11742 14123 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11824 14123 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11824 14123 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11906 14123 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11906 14123 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 11988 14123 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 11988 14123 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14059 12070 14123 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14059 12070 14123 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11250 14204 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11250 14204 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11332 14204 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11332 14204 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11414 14204 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11414 14204 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11496 14204 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11496 14204 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11578 14204 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11578 14204 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11660 14204 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11660 14204 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11742 14204 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11742 14204 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11824 14204 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11824 14204 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11906 14204 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11906 14204 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 11988 14204 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 11988 14204 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14140 12070 14204 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14140 12070 14204 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11250 14285 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11250 14285 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11332 14285 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11332 14285 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11414 14285 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11414 14285 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11496 14285 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11496 14285 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11578 14285 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11578 14285 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11660 14285 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11660 14285 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11742 14285 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11742 14285 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11824 14285 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11824 14285 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11906 14285 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11906 14285 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 11988 14285 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 11988 14285 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14221 12070 14285 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14221 12070 14285 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11250 14366 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11250 14366 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11332 14366 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11332 14366 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11414 14366 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11414 14366 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11496 14366 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11496 14366 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11578 14366 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11578 14366 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11660 14366 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11660 14366 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11742 14366 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11742 14366 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11824 14366 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11824 14366 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11906 14366 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11906 14366 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 11988 14366 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 11988 14366 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14302 12070 14366 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14302 12070 14366 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11250 14447 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11250 14447 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11332 14447 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11332 14447 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11414 14447 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11414 14447 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11496 14447 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11496 14447 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11578 14447 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11578 14447 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11660 14447 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11660 14447 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11742 14447 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11742 14447 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11824 14447 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11824 14447 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11906 14447 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11906 14447 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 11988 14447 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 11988 14447 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14383 12070 14447 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14383 12070 14447 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11250 14528 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11250 14528 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11332 14528 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11332 14528 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11414 14528 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11414 14528 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11496 14528 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11496 14528 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11578 14528 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11578 14528 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11660 14528 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11660 14528 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11742 14528 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11742 14528 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11824 14528 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11824 14528 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11906 14528 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11906 14528 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 11988 14528 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 11988 14528 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14464 12070 14528 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14464 12070 14528 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11250 14609 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11250 14609 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11332 14609 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11332 14609 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11414 14609 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11414 14609 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11496 14609 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11496 14609 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11578 14609 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11578 14609 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11660 14609 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11660 14609 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11742 14609 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11742 14609 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11824 14609 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11824 14609 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11906 14609 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11906 14609 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 11988 14609 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 11988 14609 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14545 12070 14609 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14545 12070 14609 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11250 14690 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11250 14690 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11332 14690 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11332 14690 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11414 14690 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11414 14690 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11496 14690 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11496 14690 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11578 14690 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11578 14690 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11660 14690 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11660 14690 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11742 14690 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11742 14690 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11824 14690 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11824 14690 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11906 14690 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11906 14690 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 11988 14690 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 11988 14690 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14626 12070 14690 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14626 12070 14690 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11250 14771 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11250 14771 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11332 14771 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11332 14771 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11414 14771 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11414 14771 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11496 14771 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11496 14771 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11578 14771 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11578 14771 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11660 14771 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11660 14771 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11742 14771 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11742 14771 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11824 14771 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11824 14771 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11906 14771 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11906 14771 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 11988 14771 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 11988 14771 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14707 12070 14771 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14707 12070 14771 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11250 14852 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11250 14852 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11332 14852 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11332 14852 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11414 14852 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11414 14852 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11496 14852 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11496 14852 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11578 14852 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11578 14852 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11660 14852 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11660 14852 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11742 14852 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11742 14852 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11824 14852 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11824 14852 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11906 14852 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11906 14852 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 11988 14852 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 11988 14852 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 14788 12070 14852 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 14788 12070 14852 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11250 1715 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11250 1715 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11332 1715 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11332 1715 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11414 1715 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11414 1715 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11496 1715 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11496 1715 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11578 1715 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11578 1715 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11660 1715 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11660 1715 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11742 1715 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11742 1715 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11824 1715 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11824 1715 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11906 1715 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11906 1715 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 11988 1715 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 11988 1715 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1651 12070 1715 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1651 12070 1715 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11250 1796 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11250 1796 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11332 1796 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11332 1796 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11414 1796 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11414 1796 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11496 1796 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11496 1796 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11578 1796 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11578 1796 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11660 1796 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11660 1796 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11742 1796 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11742 1796 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11824 1796 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11824 1796 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11906 1796 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11906 1796 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 11988 1796 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 11988 1796 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1732 12070 1796 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1732 12070 1796 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11250 1877 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11250 1877 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11332 1877 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11332 1877 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11414 1877 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11414 1877 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11496 1877 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11496 1877 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11578 1877 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11578 1877 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11660 1877 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11660 1877 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11742 1877 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11742 1877 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11824 1877 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11824 1877 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11906 1877 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11906 1877 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 11988 1877 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 11988 1877 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1813 12070 1877 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1813 12070 1877 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11250 1958 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11250 1958 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11332 1958 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11332 1958 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11414 1958 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11414 1958 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11496 1958 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11496 1958 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11578 1958 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11578 1958 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11660 1958 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11660 1958 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11742 1958 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11742 1958 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11824 1958 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11824 1958 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11906 1958 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11906 1958 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 11988 1958 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 11988 1958 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1894 12070 1958 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1894 12070 1958 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11250 2039 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11250 2039 11314 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11332 2039 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11332 2039 11396 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11414 2039 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11414 2039 11478 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11496 2039 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11496 2039 11560 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11578 2039 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11578 2039 11642 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11660 2039 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11660 2039 11724 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11742 2039 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11742 2039 11806 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11824 2039 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11824 2039 11888 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11906 2039 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11906 2039 11970 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 11988 2039 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 11988 2039 12052 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal4 s 1975 12070 2039 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal3 s 1975 12070 2039 12134 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 39600
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 13753878
string GDS_START 13341958
<< end >>
