magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 17 299 85 493
rect 17 177 52 299
rect 260 215 344 255
rect 378 215 444 255
rect 478 215 544 255
rect 17 51 85 177
rect 649 215 719 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 119 299 153 527
rect 207 367 257 527
rect 386 333 452 493
rect 512 367 578 527
rect 612 333 678 493
rect 191 299 678 333
rect 191 249 225 299
rect 86 215 225 249
rect 119 17 169 177
rect 207 147 452 181
rect 207 51 273 147
rect 307 17 352 109
rect 386 51 452 147
rect 578 173 612 299
rect 578 51 678 173
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 260 215 344 255 6 A1
port 1 nsew signal input
rlabel locali s 378 215 444 255 6 A2
port 2 nsew signal input
rlabel locali s 478 215 544 255 6 B1
port 3 nsew signal input
rlabel locali s 649 215 719 265 6 C1
port 4 nsew signal input
rlabel locali s 17 299 85 493 6 X
port 9 nsew signal output
rlabel locali s 17 177 52 299 6 X
port 9 nsew signal output
rlabel locali s 17 51 85 177 6 X
port 9 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3999992
string GDS_START 3993208
<< end >>
