magic
tech sky130A
timestamp 1624855509
<< checkpaint >>
rect -630 -630 780 2130
<< pwell >>
rect 0 0 150 1500
<< nsubdiff >>
rect 0 0 150 1500
use sky130_fd_io__gnd2gnd_strap  sky130_fd_io__gnd2gnd_strap_0
timestamp 1624855509
transform 1 0 0 0 1 0
box 0 0 150 1500
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 14498326
string GDS_START 14498142
<< end >>
