magic
tech sky130A
timestamp 1624857261
<< checkpaint >>
rect -630 -630 726 726
<< metal1 >>
rect 0 3 3 93
rect 93 3 96 93
<< via1 >>
rect 3 3 93 93
<< metal2 >>
rect 3 93 93 96
rect 3 0 93 3
<< properties >>
string FIXED_BBOX 0 0 96 96
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_8kbyte_1rw1r_32x2048_8.gds
string GDS_END 44269244
string GDS_START 44268408
<< end >>
