magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1260 -1260 16260 41260
<< metal2 >>
rect 99 0 4879 148
rect 5179 0 5579 107
rect 10078 0 14858 148
<< metal3 >>
rect 99 0 4879 391
rect 5179 0 7379 545
rect 7578 0 9778 2266
rect 10078 0 14858 18037
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 7329 27865 7594 29187
rect 0 14007 254 18997
rect 14746 14007 15000 18997
rect 0 12837 254 13687
rect 14746 12837 15000 13687
rect 0 11667 254 12517
rect 14746 11667 15000 12517
rect 0 9547 254 11347
rect 14746 9547 15000 11347
rect 0 8337 254 9227
rect 14746 8337 15000 9227
rect 0 7368 254 8017
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 14746 6397 15000 7047
rect 0 5187 254 6077
rect 14746 5187 15000 6077
rect 0 3977 254 4867
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 14746 1797 15000 2687
rect 0 427 254 1477
rect 14746 427 15000 1477
use sky130_fd_io__hvc_clampv2  sky130_fd_io__hvc_clampv2_0
timestamp 1624855509
transform 1 0 0 0 1 0
box 0 0 15000 40000
<< labels >>
flabel metal3 s 99 0 4879 391 0 FreeSans 2000 0 0 0 P_CORE
port 7 nsew default bidirectional
flabel metal3 s 7578 0 9778 318 0 FreeSans 2000 0 0 0 DRN_HVC
port 4 nsew default bidirectional
flabel metal3 s 10078 0 14858 391 0 FreeSans 2000 0 0 0 P_CORE
port 8 nsew default bidirectional
flabel metal3 s 5179 0 7379 148 2 FreeSans 2000 90 0 0 SRC_BDY_HVC
port 10 nsew default bidirectional
flabel metal2 s 10078 0 14858 148 2 FreeSans 2000 90 0 0 DRN_HVC
port 5 nsew default bidirectional
flabel metal2 s 99 0 4879 148 2 FreeSans 2000 90 0 0 SRC_BDY_HVC
port 11 nsew default bidirectional
flabel metal2 s 5179 0 5579 107 2 FreeSans 1000 90 0 0 OGC_HVC
port 6 nsew default bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 36 nsew default bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 48 nsew default bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 2 nsew default bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 0 nsew default bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 32 nsew default bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 24 nsew default bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 64 nsew default bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 52 nsew default bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 25 nsew default bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 20 nsew default bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 12 nsew default bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 16 nsew default bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 37 nsew default bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 60 nsew default bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 38 nsew default bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 39 nsew default bidirectional
flabel metal4 s 14746 7347 15000 8037 3 FreeSans 520 180 0 0 VSSA
port 40 nsew default bidirectional
flabel metal4 s 14746 8317 15000 9247 3 FreeSans 520 180 0 0 VSSD
port 49 nsew default bidirectional
flabel metal4 s 14746 9673 15000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 3 nsew default bidirectional
flabel metal4 s 14746 10625 15000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 1 nsew default bidirectional
flabel metal4 s 14746 12817 15000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 33 nsew default bidirectional
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 520 180 0 0 VDDIO
port 26 nsew default bidirectional
flabel metal4 s 14746 6377 15000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 65 nsew default bidirectional
flabel metal4 s 14746 5167 15000 6097 3 FreeSans 520 180 0 0 VSSIO
port 53 nsew default bidirectional
flabel metal4 s 14746 3957 15000 4887 3 FreeSans 520 180 0 0 VDDIO
port 27 nsew default bidirectional
flabel metal4 s 14807 2987 15000 3677 3 FreeSans 520 180 0 0 VDDA
port 21 nsew default bidirectional
flabel metal4 s 14746 1777 15000 2707 3 FreeSans 520 180 0 0 VCCD
port 13 nsew default bidirectional
flabel metal4 s 14746 407 15000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 17 nsew default bidirectional
flabel metal4 s 14746 11281 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 41 nsew default bidirectional
flabel metal4 s 14746 11647 15000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 61 nsew default bidirectional
flabel metal4 s 14746 9547 15000 9613 3 FreeSans 520 180 0 0 VSSA
port 42 nsew default bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 54 nsew default bidirectional
flabel metal4 s 127 38321 127 38321 3 FreeSans 520 0 0 0 VSSIO
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 55 nsew default bidirectional
flabel metal4 s 14873 38321 14873 38321 3 FreeSans 520 180 0 0 VSSIO
flabel metal4 s 14746 10329 15000 10565 3 FreeSans 520 180 0 0 VSSA
port 43 nsew default bidirectional
flabel metal5 s 7329 27865 7594 29187 0 FreeSans 2000 0 0 0 P_PAD
port 9 nsew default bidirectional
flabel metal5 s 14746 5187 15000 6077 3 FreeSans 520 180 0 0 VSSIO
port 56 nsew default bidirectional
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 57 nsew default bidirectional
flabel metal5 s 14746 12837 15000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 34 nsew default bidirectional
flabel metal5 s 14746 11667 15000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 62 nsew default bidirectional
flabel metal5 s 14746 6397 15000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 66 nsew default bidirectional
flabel metal5 s 14746 7368 15000 8017 3 FreeSans 520 180 0 0 VSSA
port 44 nsew default bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 58 nsew default bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 45 nsew default bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 28 nsew default bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 14 nsew default bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 18 nsew default bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 22 nsew default bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 29 nsew default bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 35 nsew default bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 46 nsew default bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 50 nsew default bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 59 nsew default bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 67 nsew default bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 63 nsew default bidirectional
flabel metal5 s 14746 9547 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 47 nsew default bidirectional
flabel metal5 s 14746 3977 15000 4867 3 FreeSans 520 180 0 0 VDDIO
port 30 nsew default bidirectional
flabel metal5 s 14746 1797 15000 2687 3 FreeSans 520 180 0 0 VCCD
port 15 nsew default bidirectional
flabel metal5 s 14746 427 15000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 19 nsew default bidirectional
flabel metal5 s 14807 3007 15000 3657 3 FreeSans 520 180 0 0 VDDA
port 23 nsew default bidirectional
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 520 180 0 0 VDDIO
port 31 nsew default bidirectional
flabel metal5 s 14746 8337 15000 9227 3 FreeSans 520 180 0 0 VSSD
port 51 nsew default bidirectional
rlabel metal4 s 14746 10625 15000 11221 1 AMUXBUS_A
port 1 nsew default bidirectional
rlabel metal4 s 14746 9673 15000 10269 1 AMUXBUS_B
port 3 nsew default bidirectional
rlabel metal3 s 7578 0 9778 2266 1 DRN_HVC
port 5 nsew default bidirectional
rlabel metal3 s 10078 0 14858 18037 1 P_CORE
port 8 nsew default bidirectional
rlabel metal3 s 5179 0 7379 545 1 SRC_BDY_HVC
port 11 nsew default bidirectional
rlabel metal4 s 14746 1777 15000 2707 1 VCCD
port 15 nsew default bidirectional
rlabel metal5 s 0 1797 254 2687 1 VCCD
port 15 nsew default bidirectional
rlabel metal5 s 14746 1797 15000 2687 1 VCCD
port 15 nsew default bidirectional
rlabel metal4 s 14746 407 15000 1497 1 VCCHIB
port 19 nsew default bidirectional
rlabel metal5 s 0 427 254 1477 1 VCCHIB
port 19 nsew default bidirectional
rlabel metal5 s 14746 427 15000 1477 1 VCCHIB
port 19 nsew default bidirectional
rlabel metal4 s 14807 2987 15000 3677 1 VDDA
port 23 nsew default bidirectional
rlabel metal5 s 0 3007 193 3657 1 VDDA
port 23 nsew default bidirectional
rlabel metal5 s 14807 3007 15000 3657 1 VDDA
port 23 nsew default bidirectional
rlabel metal4 s 0 14007 254 19000 1 VDDIO
port 31 nsew default bidirectional
rlabel metal4 s 14746 3957 15000 4887 1 VDDIO
port 31 nsew default bidirectional
rlabel metal4 s 14746 14007 15000 19000 1 VDDIO
port 31 nsew default bidirectional
rlabel metal5 s 0 3977 254 4867 1 VDDIO
port 31 nsew default bidirectional
rlabel metal5 s 0 14007 254 18997 1 VDDIO
port 31 nsew default bidirectional
rlabel metal5 s 14746 3977 15000 4867 1 VDDIO
port 31 nsew default bidirectional
rlabel metal5 s 14746 14007 15000 18997 1 VDDIO
port 31 nsew default bidirectional
rlabel metal4 s 14746 12817 15000 13707 1 VDDIO_Q
port 35 nsew default bidirectional
rlabel metal5 s 0 12837 254 13687 1 VDDIO_Q
port 35 nsew default bidirectional
rlabel metal5 s 14746 12837 15000 13687 1 VDDIO_Q
port 35 nsew default bidirectional
rlabel metal4 s 0 9547 15000 9613 1 VSSA
port 47 nsew default bidirectional
rlabel metal4 s 0 10329 254 10565 1 VSSA
port 47 nsew default bidirectional
rlabel metal4 s 0 11281 15000 11347 1 VSSA
port 47 nsew default bidirectional
rlabel metal4 s 14746 7347 15000 8037 1 VSSA
port 47 nsew default bidirectional
rlabel metal4 s 14746 9547 15000 9613 1 VSSA
port 47 nsew default bidirectional
rlabel metal4 s 14746 10329 15000 10565 1 VSSA
port 47 nsew default bidirectional
rlabel metal4 s 14746 11281 15000 11347 1 VSSA
port 47 nsew default bidirectional
rlabel metal5 s 0 7368 254 8017 1 VSSA
port 47 nsew default bidirectional
rlabel metal5 s 0 9547 254 11347 1 VSSA
port 47 nsew default bidirectional
rlabel metal5 s 14746 7368 15000 8017 1 VSSA
port 47 nsew default bidirectional
rlabel metal5 s 14746 9547 15000 11347 1 VSSA
port 47 nsew default bidirectional
rlabel metal4 s 14746 8317 15000 9247 1 VSSD
port 51 nsew default bidirectional
rlabel metal5 s 0 8337 254 9227 1 VSSD
port 51 nsew default bidirectional
rlabel metal5 s 14746 8337 15000 9227 1 VSSD
port 51 nsew default bidirectional
rlabel metal4 s 14746 35157 15000 40000 1 VSSIO
port 59 nsew default bidirectional
rlabel metal4 s 14746 5167 15000 6097 1 VSSIO
port 59 nsew default bidirectional
rlabel metal4 s 14872 38320 14874 38322 1 VSSIO
port 59 nsew default bidirectional
rlabel metal5 s 0 35157 254 40000 1 VSSIO
port 59 nsew default bidirectional
rlabel metal5 s 0 5187 254 6077 1 VSSIO
port 59 nsew default bidirectional
rlabel metal5 s 14746 35157 15000 40000 1 VSSIO
port 59 nsew default bidirectional
rlabel metal5 s 14746 5187 15000 6077 1 VSSIO
port 59 nsew default bidirectional
rlabel metal4 s 14746 11647 15000 12537 1 VSSIO_Q
port 63 nsew default bidirectional
rlabel metal5 s 0 11667 254 12517 1 VSSIO_Q
port 63 nsew default bidirectional
rlabel metal5 s 14746 11667 15000 12517 1 VSSIO_Q
port 63 nsew default bidirectional
rlabel metal4 s 14746 6377 15000 7067 1 VSWITCH
port 67 nsew default bidirectional
rlabel metal5 s 0 6397 254 7047 1 VSWITCH
port 67 nsew default bidirectional
rlabel metal5 s 14746 6397 15000 7047 1 VSWITCH
port 67 nsew default bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 15000 40000
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 5498800
string GDS_START 5489324
<< end >>
