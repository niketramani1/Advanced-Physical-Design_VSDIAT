magic
tech sky130A
magscale 1 2
timestamp 1624855602
<< nwell >>
rect -66 377 1026 897
<< pwell >>
rect 0 -17 960 17
<< locali >>
rect 244 415 294 751
rect 556 415 622 751
rect 244 381 622 415
rect 244 356 278 381
rect 25 310 278 356
rect 777 355 843 424
rect 244 275 278 310
rect 244 241 606 275
rect 244 99 294 241
rect 556 99 606 241
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 960 831
rect 18 735 208 751
rect 18 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 208 735
rect 18 435 208 701
rect 330 735 520 751
rect 330 701 336 735
rect 370 701 408 735
rect 442 701 480 735
rect 514 701 520 735
rect 330 451 520 701
rect 658 735 848 751
rect 658 701 664 735
rect 698 701 736 735
rect 770 701 808 735
rect 842 701 848 735
rect 658 460 848 701
rect 314 319 720 345
rect 884 319 934 751
rect 314 311 934 319
rect 686 285 934 311
rect 18 113 208 265
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 208 113
rect 330 113 520 205
rect 18 73 208 79
rect 330 79 336 113
rect 370 79 408 113
rect 442 79 480 113
rect 514 79 520 113
rect 642 113 832 249
rect 330 73 520 79
rect 642 79 648 113
rect 682 79 720 113
rect 754 79 792 113
rect 826 79 832 113
rect 868 99 934 285
rect 642 73 832 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 24 701 58 735
rect 96 701 130 735
rect 168 701 202 735
rect 336 701 370 735
rect 408 701 442 735
rect 480 701 514 735
rect 664 701 698 735
rect 736 701 770 735
rect 808 701 842 735
rect 24 79 58 113
rect 96 79 130 113
rect 168 79 202 113
rect 336 79 370 113
rect 408 79 442 113
rect 480 79 514 113
rect 648 79 682 113
rect 720 79 754 113
rect 792 79 826 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 831 960 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 960 831
rect 0 791 960 797
rect 0 735 960 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 336 735
rect 370 701 408 735
rect 442 701 480 735
rect 514 701 664 735
rect 698 701 736 735
rect 770 701 808 735
rect 842 701 960 735
rect 0 689 960 701
rect 0 113 960 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 336 113
rect 370 79 408 113
rect 442 79 480 113
rect 514 79 648 113
rect 682 79 720 113
rect 754 79 792 113
rect 826 79 960 113
rect 0 51 960 79
rect 0 17 960 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -23 960 -17
<< labels >>
rlabel locali s 777 355 843 424 6 A
port 1 nsew signal input
rlabel locali s 556 415 622 751 6 X
port 6 nsew signal output
rlabel locali s 556 99 606 241 6 X
port 6 nsew signal output
rlabel locali s 244 415 294 751 6 X
port 6 nsew signal output
rlabel locali s 244 381 622 415 6 X
port 6 nsew signal output
rlabel locali s 244 356 278 381 6 X
port 6 nsew signal output
rlabel locali s 244 275 278 310 6 X
port 6 nsew signal output
rlabel locali s 244 241 606 275 6 X
port 6 nsew signal output
rlabel locali s 244 99 294 241 6 X
port 6 nsew signal output
rlabel locali s 25 310 278 356 6 X
port 6 nsew signal output
rlabel metal1 s 0 51 960 125 6 VGND
port 2 nsew ground bidirectional
rlabel pwell s 0 -17 960 17 8 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 960 23 8 VNB
port 3 nsew ground bidirectional
rlabel nwell s -66 377 1026 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 791 960 837 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 960 763 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 960 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 879070
string GDS_START 867864
<< end >>
