magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 103 51 171 493
rect 301 215 367 323
rect 401 51 478 323
rect 536 215 620 323
rect 674 265 732 474
rect 660 199 732 265
rect 862 263 903 471
rect 766 201 903 263
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 27 299 69 527
rect 27 17 69 177
rect 207 439 331 527
rect 372 405 428 493
rect 465 451 531 527
rect 573 405 639 493
rect 206 357 639 405
rect 206 177 261 357
rect 206 143 361 177
rect 207 17 257 109
rect 295 51 361 143
rect 777 299 828 527
rect 573 125 843 165
rect 573 51 639 125
rect 677 17 743 91
rect 777 51 843 125
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 862 263 903 471 6 A1
port 1 nsew signal input
rlabel locali s 766 201 903 263 6 A1
port 1 nsew signal input
rlabel locali s 674 265 732 474 6 A2
port 2 nsew signal input
rlabel locali s 660 199 732 265 6 A2
port 2 nsew signal input
rlabel locali s 536 215 620 323 6 B1
port 3 nsew signal input
rlabel locali s 401 51 478 323 6 C1
port 4 nsew signal input
rlabel locali s 301 215 367 323 6 D1
port 5 nsew signal input
rlabel locali s 103 51 171 493 6 X
port 10 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3150220
string GDS_START 3142112
<< end >>
