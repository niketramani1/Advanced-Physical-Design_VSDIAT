magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1260 -1250 1794 1876
<< nwell >>
rect 0 284 534 616
<< mvnmos >>
rect 119 36 239 120
rect 295 36 415 120
<< mvpmos >>
rect 119 350 239 550
rect 295 350 415 550
<< mvndiff >>
rect 66 82 119 120
rect 66 48 74 82
rect 108 48 119 82
rect 66 36 119 48
rect 239 82 295 120
rect 239 48 250 82
rect 284 48 295 82
rect 239 36 295 48
rect 415 82 468 120
rect 415 48 426 82
rect 460 48 468 82
rect 415 36 468 48
<< mvpdiff >>
rect 66 532 119 550
rect 66 498 74 532
rect 108 498 119 532
rect 66 464 119 498
rect 66 430 74 464
rect 108 430 119 464
rect 66 396 119 430
rect 66 362 74 396
rect 108 362 119 396
rect 66 350 119 362
rect 239 532 295 550
rect 239 498 250 532
rect 284 498 295 532
rect 239 464 295 498
rect 239 430 250 464
rect 284 430 295 464
rect 239 396 295 430
rect 239 362 250 396
rect 284 362 295 396
rect 239 350 295 362
rect 415 532 468 550
rect 415 498 426 532
rect 460 498 468 532
rect 415 464 468 498
rect 415 430 426 464
rect 460 430 468 464
rect 415 396 468 430
rect 415 362 426 396
rect 460 362 468 396
rect 415 350 468 362
<< mvndiffc >>
rect 74 48 108 82
rect 250 48 284 82
rect 426 48 460 82
<< mvpdiffc >>
rect 74 498 108 532
rect 74 430 108 464
rect 74 362 108 396
rect 250 498 284 532
rect 250 430 284 464
rect 250 362 284 396
rect 426 498 460 532
rect 426 430 460 464
rect 426 362 460 396
<< poly >>
rect 119 550 239 576
rect 295 550 415 576
rect 119 324 239 350
rect 295 324 415 350
rect 119 286 415 324
rect 119 252 155 286
rect 189 252 415 286
rect 119 218 415 252
rect 119 184 155 218
rect 189 184 415 218
rect 119 146 415 184
rect 119 120 239 146
rect 295 120 415 146
rect 119 10 239 36
rect 295 10 415 36
<< polycont >>
rect 155 252 189 286
rect 155 184 189 218
<< locali >>
rect 74 486 108 498
rect 74 396 108 430
rect 74 346 108 362
rect 240 532 284 550
rect 240 498 250 532
rect 240 464 284 498
rect 240 430 250 464
rect 240 396 284 430
rect 240 362 250 396
rect 155 288 189 302
rect 155 218 189 252
rect 155 168 189 182
rect 240 288 284 362
rect 426 486 460 498
rect 426 396 460 430
rect 426 346 460 362
rect 240 254 245 288
rect 279 254 284 288
rect 240 216 284 254
rect 240 182 245 216
rect 279 182 284 216
rect 74 82 108 94
rect 240 82 284 182
rect 240 48 250 82
rect 240 32 284 48
rect 426 82 460 94
<< viali >>
rect 74 532 108 558
rect 74 524 108 532
rect 74 464 108 486
rect 74 452 108 464
rect 155 286 189 288
rect 155 254 189 286
rect 155 184 189 216
rect 155 182 189 184
rect 426 532 460 558
rect 426 524 460 532
rect 426 464 460 486
rect 426 452 460 464
rect 245 254 279 288
rect 245 182 279 216
rect 74 94 108 128
rect 74 48 108 56
rect 74 22 108 48
rect 426 94 460 128
rect 426 48 460 56
rect 426 22 460 48
<< metal1 >>
rect 68 558 466 570
rect 68 524 74 558
rect 108 524 426 558
rect 460 524 466 558
rect 68 486 466 524
rect 68 452 74 486
rect 108 452 426 486
rect 460 452 466 486
rect 68 440 466 452
rect 149 288 195 300
rect 149 254 155 288
rect 189 254 195 288
rect 149 216 195 254
rect 149 182 155 216
rect 189 182 195 216
rect 149 170 195 182
rect 239 288 285 300
rect 239 254 245 288
rect 279 254 285 288
rect 239 216 285 254
rect 239 182 245 216
rect 279 182 285 216
rect 239 170 285 182
rect 68 128 466 140
rect 68 94 74 128
rect 108 94 426 128
rect 460 94 466 128
rect 68 56 466 94
rect 68 22 74 56
rect 108 22 426 56
rect 460 22 466 56
rect 68 10 466 22
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1624855509
transform -1 0 205 0 -1 302
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808441  sky130_fd_pr__pfet_01v8__example_55959141808441_0
timestamp 1624855509
transform 1 0 119 0 1 350
box -28 0 324 97
use sky130_fd_pr__nfet_01v8__example_55959141808571  sky130_fd_pr__nfet_01v8__example_55959141808571_0
timestamp 1624855509
transform 1 0 119 0 1 36
box -28 0 324 29
<< labels >>
flabel metal1 s 164 202 189 260 3 FreeSans 520 0 0 0 A
flabel metal1 s 145 481 232 545 3 FreeSans 520 0 0 0 VDA
flabel metal1 s 146 33 242 90 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 249 209 276 267 3 FreeSans 520 0 0 0 Y
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 618090
string GDS_START 615490
<< end >>
