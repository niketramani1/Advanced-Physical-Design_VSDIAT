magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 387 425 627 473
rect 17 215 85 328
rect 187 299 266 340
rect 187 119 221 299
rect 339 215 446 323
rect 187 53 257 119
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 408 69 444
rect 110 442 182 527
rect 285 442 351 527
rect 17 391 344 408
rect 17 374 532 391
rect 17 362 153 374
rect 119 181 153 362
rect 310 357 532 374
rect 17 147 153 181
rect 17 58 69 147
rect 255 187 289 265
rect 498 265 532 357
rect 566 299 627 385
rect 498 199 558 265
rect 255 181 319 187
rect 255 165 432 181
rect 593 165 627 299
rect 255 153 627 165
rect 285 147 627 153
rect 398 131 627 147
rect 119 17 153 113
rect 304 17 338 113
rect 398 61 432 131
rect 566 121 627 131
rect 466 17 532 97
rect 566 61 617 121
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 339 215 446 323 6 A
port 1 nsew signal input
rlabel locali s 387 425 627 473 6 B
port 2 nsew signal input
rlabel locali s 17 215 85 328 6 C_N
port 3 nsew signal input
rlabel locali s 187 299 266 340 6 X
port 8 nsew signal output
rlabel locali s 187 119 221 299 6 X
port 8 nsew signal output
rlabel locali s 187 53 257 119 6 X
port 8 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3886390
string GDS_START 3880600
<< end >>
