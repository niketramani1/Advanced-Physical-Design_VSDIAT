magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 212 312 263 493
rect 17 197 88 271
rect 229 166 263 312
rect 212 51 263 166
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 35 341 69 493
rect 112 375 178 527
rect 35 307 178 341
rect 144 265 178 307
rect 144 199 195 265
rect 144 161 178 199
rect 298 297 350 527
rect 35 127 178 161
rect 35 51 69 127
rect 112 17 178 93
rect 298 17 350 185
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel locali s 17 197 88 271 6 A
port 1 nsew signal input
rlabel locali s 229 166 263 312 6 X
port 6 nsew signal output
rlabel locali s 212 312 263 493 6 X
port 6 nsew signal output
rlabel locali s 212 51 263 166 6 X
port 6 nsew signal output
rlabel metal1 s 0 -48 368 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 406 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1237440
string GDS_START 1233004
<< end >>
