magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1260 -1286 1734 1568
<< scnmos >>
rect 60 0 90 252
rect 168 0 198 252
rect 276 0 306 252
rect 384 0 414 252
<< ndiff >>
rect 0 143 60 252
rect 0 109 8 143
rect 42 109 60 143
rect 0 0 60 109
rect 90 143 168 252
rect 90 109 112 143
rect 146 109 168 143
rect 90 0 168 109
rect 198 143 276 252
rect 198 109 220 143
rect 254 109 276 143
rect 198 0 276 109
rect 306 143 384 252
rect 306 109 328 143
rect 362 109 384 143
rect 306 0 384 109
rect 414 143 474 252
rect 414 109 432 143
rect 466 109 474 143
rect 414 0 474 109
<< ndiffc >>
rect 8 109 42 143
rect 112 109 146 143
rect 220 109 254 143
rect 328 109 362 143
rect 432 109 466 143
<< poly >>
rect 60 278 414 308
rect 60 252 90 278
rect 168 252 198 278
rect 276 252 306 278
rect 384 252 414 278
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
<< locali >>
rect 112 193 362 227
rect 8 143 42 159
rect 8 93 42 109
rect 112 143 146 193
rect 112 93 146 109
rect 220 143 254 159
rect 220 93 254 109
rect 328 143 362 193
rect 328 93 362 109
rect 432 143 466 159
rect 432 93 466 109
use contact_11  contact_11_0
timestamp 1624857261
transform 1 0 424 0 1 93
box 0 0 1 1
use contact_11  contact_11_1
timestamp 1624857261
transform 1 0 320 0 1 93
box 0 0 1 1
use contact_11  contact_11_2
timestamp 1624857261
transform 1 0 212 0 1 93
box 0 0 1 1
use contact_11  contact_11_3
timestamp 1624857261
transform 1 0 104 0 1 93
box 0 0 1 1
use contact_11  contact_11_4
timestamp 1624857261
transform 1 0 0 0 1 93
box 0 0 1 1
<< labels >>
rlabel poly s 237 293 237 293 4 G
rlabel locali s 237 126 237 126 4 S
rlabel locali s 449 126 449 126 4 S
rlabel locali s 25 126 25 126 4 S
rlabel locali s 237 210 237 210 4 D
<< properties >>
string FIXED_BBOX -25 -26 499 308
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 9265636
string GDS_START 9264252
<< end >>
