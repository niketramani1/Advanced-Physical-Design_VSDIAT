magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 329 427 436 493
rect 29 199 100 323
rect 202 199 267 323
rect 373 165 436 427
rect 313 105 436 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 54 391 132 426
rect 229 425 295 527
rect 54 357 339 391
rect 134 165 168 357
rect 305 199 339 357
rect 50 17 98 165
rect 134 85 190 165
rect 236 17 279 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 202 199 267 323 6 A
port 1 nsew signal input
rlabel locali s 29 199 100 323 6 B
port 2 nsew signal input
rlabel locali s 373 165 436 427 6 X
port 7 nsew signal output
rlabel locali s 329 427 436 493 6 X
port 7 nsew signal output
rlabel locali s 313 105 436 165 6 X
port 7 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4022
string GDS_START 128
<< end >>
