magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1306 -1260 1388 1289
use sky130_fd_pr__hvdfm1sd__example_55959141808452  sky130_fd_pr__hvdfm1sd__example_55959141808452_0
timestamp 1624855509
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808122  sky130_fd_pr__hvdfl1sd__example_55959141808122_0
timestamp 1624855509
transform -1 0 -18 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 13 128 13 0 FreeSans 300 0 0 0 D
flabel comment s -46 29 -46 29 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 298462
string GDS_START 297344
<< end >>
