magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1235 -1186 1385 1335
<< labels >>
rlabel poly s 75 74 75 74 4 G
rlabel mvpsubdiff s 25 74 25 74 4 S
rlabel mvpsubdiff s 125 74 125 74 4 D
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 9197244
string GDS_START 9196596
<< end >>
