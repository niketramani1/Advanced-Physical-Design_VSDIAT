magic
tech sky130A
magscale 1 2
timestamp 1624855596
<< checkpaint >>
rect -1326 -1283 3438 2911
<< nwell >>
rect -66 377 160 1251
rect 560 403 867 865
rect 1267 493 2178 1251
rect 1960 377 2178 493
<< pwell >>
rect 0 1611 2112 1645
rect 0 -17 2112 17
<< scnmos >>
rect 656 151 686 319
rect 742 151 772 319
<< scpmoshvt >>
rect 656 439 686 607
rect 742 439 772 607
<< mvnmos >>
rect 404 1221 504 1521
rect 560 1221 660 1521
rect 716 1221 816 1521
rect 872 1221 972 1521
rect 1028 1221 1128 1521
rect 1764 1371 1864 1521
rect 1929 1371 2029 1521
rect 1097 107 1197 407
rect 1253 107 1353 407
rect 1409 107 1509 407
rect 1565 107 1665 407
rect 1721 107 1821 407
<< mvpmos >>
rect 1398 885 1598 969
rect 1764 885 1864 1185
rect 1929 885 2029 1185
rect 1406 563 1606 647
<< ndiff >>
rect 597 299 656 319
rect 597 265 611 299
rect 645 265 656 299
rect 597 197 656 265
rect 597 163 611 197
rect 645 163 656 197
rect 597 151 656 163
rect 686 299 742 319
rect 686 265 697 299
rect 731 265 742 299
rect 686 193 742 265
rect 686 159 697 193
rect 731 159 742 193
rect 686 151 742 159
rect 772 299 831 319
rect 772 265 783 299
rect 817 265 831 299
rect 772 197 831 265
rect 772 163 783 197
rect 817 163 831 197
rect 772 151 831 163
<< pdiff >>
rect 597 595 656 607
rect 597 561 611 595
rect 645 561 656 595
rect 597 483 656 561
rect 597 449 611 483
rect 645 449 656 483
rect 597 439 656 449
rect 686 595 742 607
rect 686 561 697 595
rect 731 561 742 595
rect 686 483 742 561
rect 686 449 697 483
rect 731 449 742 483
rect 686 439 742 449
rect 772 565 831 607
rect 772 531 783 565
rect 817 531 831 565
rect 772 483 831 531
rect 772 449 783 483
rect 817 449 831 483
rect 772 439 831 449
<< mvndiff >>
rect 351 1509 404 1521
rect 351 1475 359 1509
rect 393 1475 404 1509
rect 351 1429 404 1475
rect 351 1395 359 1429
rect 393 1395 404 1429
rect 351 1347 404 1395
rect 351 1313 359 1347
rect 393 1313 404 1347
rect 351 1267 404 1313
rect 351 1233 359 1267
rect 393 1233 404 1267
rect 351 1221 404 1233
rect 504 1509 560 1521
rect 504 1475 515 1509
rect 549 1475 560 1509
rect 504 1429 560 1475
rect 504 1395 515 1429
rect 549 1395 560 1429
rect 504 1347 560 1395
rect 504 1313 515 1347
rect 549 1313 560 1347
rect 504 1267 560 1313
rect 504 1233 515 1267
rect 549 1233 560 1267
rect 504 1221 560 1233
rect 660 1509 716 1521
rect 660 1475 671 1509
rect 705 1475 716 1509
rect 660 1429 716 1475
rect 660 1395 671 1429
rect 705 1395 716 1429
rect 660 1347 716 1395
rect 660 1313 671 1347
rect 705 1313 716 1347
rect 660 1267 716 1313
rect 660 1233 671 1267
rect 705 1233 716 1267
rect 660 1221 716 1233
rect 816 1509 872 1521
rect 816 1475 827 1509
rect 861 1475 872 1509
rect 816 1429 872 1475
rect 816 1395 827 1429
rect 861 1395 872 1429
rect 816 1347 872 1395
rect 816 1313 827 1347
rect 861 1313 872 1347
rect 816 1267 872 1313
rect 816 1233 827 1267
rect 861 1233 872 1267
rect 816 1221 872 1233
rect 972 1509 1028 1521
rect 972 1475 983 1509
rect 1017 1475 1028 1509
rect 972 1429 1028 1475
rect 972 1395 983 1429
rect 1017 1395 1028 1429
rect 972 1347 1028 1395
rect 972 1313 983 1347
rect 1017 1313 1028 1347
rect 972 1267 1028 1313
rect 972 1233 983 1267
rect 1017 1233 1028 1267
rect 972 1221 1028 1233
rect 1128 1509 1181 1521
rect 1128 1475 1139 1509
rect 1173 1475 1181 1509
rect 1128 1429 1181 1475
rect 1128 1395 1139 1429
rect 1173 1395 1181 1429
rect 1128 1347 1181 1395
rect 1711 1509 1764 1521
rect 1711 1475 1719 1509
rect 1753 1475 1764 1509
rect 1711 1417 1764 1475
rect 1711 1383 1719 1417
rect 1753 1383 1764 1417
rect 1711 1371 1764 1383
rect 1864 1509 1929 1521
rect 1864 1475 1884 1509
rect 1918 1475 1929 1509
rect 1864 1417 1929 1475
rect 1864 1383 1884 1417
rect 1918 1383 1929 1417
rect 1864 1371 1929 1383
rect 2029 1509 2082 1521
rect 2029 1475 2040 1509
rect 2074 1475 2082 1509
rect 2029 1417 2082 1475
rect 2029 1383 2040 1417
rect 2074 1383 2082 1417
rect 2029 1371 2082 1383
rect 1128 1313 1139 1347
rect 1173 1313 1181 1347
rect 1128 1267 1181 1313
rect 1128 1233 1139 1267
rect 1173 1233 1181 1267
rect 1128 1221 1181 1233
rect 1044 395 1097 407
rect 1044 361 1052 395
rect 1086 361 1097 395
rect 1044 315 1097 361
rect 1044 281 1052 315
rect 1086 281 1097 315
rect 1044 233 1097 281
rect 1044 199 1052 233
rect 1086 199 1097 233
rect 1044 153 1097 199
rect 1044 119 1052 153
rect 1086 119 1097 153
rect 1044 107 1097 119
rect 1197 395 1253 407
rect 1197 361 1208 395
rect 1242 361 1253 395
rect 1197 315 1253 361
rect 1197 281 1208 315
rect 1242 281 1253 315
rect 1197 233 1253 281
rect 1197 199 1208 233
rect 1242 199 1253 233
rect 1197 153 1253 199
rect 1197 119 1208 153
rect 1242 119 1253 153
rect 1197 107 1253 119
rect 1353 395 1409 407
rect 1353 361 1364 395
rect 1398 361 1409 395
rect 1353 315 1409 361
rect 1353 281 1364 315
rect 1398 281 1409 315
rect 1353 233 1409 281
rect 1353 199 1364 233
rect 1398 199 1409 233
rect 1353 153 1409 199
rect 1353 119 1364 153
rect 1398 119 1409 153
rect 1353 107 1409 119
rect 1509 395 1565 407
rect 1509 361 1520 395
rect 1554 361 1565 395
rect 1509 315 1565 361
rect 1509 281 1520 315
rect 1554 281 1565 315
rect 1509 233 1565 281
rect 1509 199 1520 233
rect 1554 199 1565 233
rect 1509 153 1565 199
rect 1509 119 1520 153
rect 1554 119 1565 153
rect 1509 107 1565 119
rect 1665 395 1721 407
rect 1665 361 1676 395
rect 1710 361 1721 395
rect 1665 315 1721 361
rect 1665 281 1676 315
rect 1710 281 1721 315
rect 1665 233 1721 281
rect 1665 199 1676 233
rect 1710 199 1721 233
rect 1665 153 1721 199
rect 1665 119 1676 153
rect 1710 119 1721 153
rect 1665 107 1721 119
rect 1821 395 1874 407
rect 1821 361 1832 395
rect 1866 361 1874 395
rect 1821 315 1874 361
rect 1821 281 1832 315
rect 1866 281 1874 315
rect 1821 233 1874 281
rect 1821 199 1832 233
rect 1866 199 1874 233
rect 1821 153 1874 199
rect 1821 119 1832 153
rect 1866 119 1874 153
rect 1821 107 1874 119
<< mvpdiff >>
rect 1711 1173 1764 1185
rect 1711 1139 1719 1173
rect 1753 1139 1764 1173
rect 1711 1093 1764 1139
rect 1711 1059 1719 1093
rect 1753 1059 1764 1093
rect 1711 1011 1764 1059
rect 1711 977 1719 1011
rect 1753 977 1764 1011
rect 1333 944 1398 969
rect 1333 910 1353 944
rect 1387 910 1398 944
rect 1333 885 1398 910
rect 1598 944 1651 969
rect 1598 910 1609 944
rect 1643 910 1651 944
rect 1598 885 1651 910
rect 1711 931 1764 977
rect 1711 897 1719 931
rect 1753 897 1764 931
rect 1711 885 1764 897
rect 1864 1173 1929 1185
rect 1864 1139 1884 1173
rect 1918 1139 1929 1173
rect 1864 1093 1929 1139
rect 1864 1059 1884 1093
rect 1918 1059 1929 1093
rect 1864 1011 1929 1059
rect 1864 977 1884 1011
rect 1918 977 1929 1011
rect 1864 931 1929 977
rect 1864 897 1884 931
rect 1918 897 1929 931
rect 1864 885 1929 897
rect 2029 1173 2082 1185
rect 2029 1139 2040 1173
rect 2074 1139 2082 1173
rect 2029 1093 2082 1139
rect 2029 1059 2040 1093
rect 2074 1059 2082 1093
rect 2029 1011 2082 1059
rect 2029 977 2040 1011
rect 2074 977 2082 1011
rect 2029 931 2082 977
rect 2029 897 2040 931
rect 2074 897 2082 931
rect 2029 885 2082 897
rect 1333 677 1391 689
rect 1333 643 1349 677
rect 1383 647 1391 677
rect 1621 677 1679 689
rect 1621 647 1629 677
rect 1383 643 1406 647
rect 1333 609 1406 643
rect 1333 575 1361 609
rect 1395 575 1406 609
rect 1333 563 1406 575
rect 1606 643 1629 647
rect 1663 643 1679 677
rect 1606 609 1679 643
rect 1606 575 1617 609
rect 1651 575 1679 609
rect 1606 563 1679 575
<< ndiffc >>
rect 611 265 645 299
rect 611 163 645 197
rect 697 265 731 299
rect 697 159 731 193
rect 783 265 817 299
rect 783 163 817 197
<< pdiffc >>
rect 611 561 645 595
rect 611 449 645 483
rect 697 561 731 595
rect 697 449 731 483
rect 783 531 817 565
rect 783 449 817 483
<< mvndiffc >>
rect 359 1475 393 1509
rect 359 1395 393 1429
rect 359 1313 393 1347
rect 359 1233 393 1267
rect 515 1475 549 1509
rect 515 1395 549 1429
rect 515 1313 549 1347
rect 515 1233 549 1267
rect 671 1475 705 1509
rect 671 1395 705 1429
rect 671 1313 705 1347
rect 671 1233 705 1267
rect 827 1475 861 1509
rect 827 1395 861 1429
rect 827 1313 861 1347
rect 827 1233 861 1267
rect 983 1475 1017 1509
rect 983 1395 1017 1429
rect 983 1313 1017 1347
rect 983 1233 1017 1267
rect 1139 1475 1173 1509
rect 1139 1395 1173 1429
rect 1719 1475 1753 1509
rect 1719 1383 1753 1417
rect 1884 1475 1918 1509
rect 1884 1383 1918 1417
rect 2040 1475 2074 1509
rect 2040 1383 2074 1417
rect 1139 1313 1173 1347
rect 1139 1233 1173 1267
rect 1052 361 1086 395
rect 1052 281 1086 315
rect 1052 199 1086 233
rect 1052 119 1086 153
rect 1208 361 1242 395
rect 1208 281 1242 315
rect 1208 199 1242 233
rect 1208 119 1242 153
rect 1364 361 1398 395
rect 1364 281 1398 315
rect 1364 199 1398 233
rect 1364 119 1398 153
rect 1520 361 1554 395
rect 1520 281 1554 315
rect 1520 199 1554 233
rect 1520 119 1554 153
rect 1676 361 1710 395
rect 1676 281 1710 315
rect 1676 199 1710 233
rect 1676 119 1710 153
rect 1832 361 1866 395
rect 1832 281 1866 315
rect 1832 199 1866 233
rect 1832 119 1866 153
<< mvpdiffc >>
rect 1719 1139 1753 1173
rect 1719 1059 1753 1093
rect 1719 977 1753 1011
rect 1353 910 1387 944
rect 1609 910 1643 944
rect 1719 897 1753 931
rect 1884 1139 1918 1173
rect 1884 1059 1918 1093
rect 1884 977 1918 1011
rect 1884 897 1918 931
rect 2040 1139 2074 1173
rect 2040 1059 2074 1093
rect 2040 977 2074 1011
rect 2040 897 2074 931
rect 1349 643 1383 677
rect 1361 575 1395 609
rect 1629 643 1663 677
rect 1617 575 1651 609
<< nsubdiff >>
rect 653 824 831 829
rect 653 790 677 824
rect 711 790 773 824
rect 807 790 831 824
rect 653 714 831 790
rect 653 680 677 714
rect 711 680 773 714
rect 807 680 831 714
rect 653 661 831 680
<< mvpsubdiff >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2112 1645
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 94 831
rect 1543 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2112 831
<< nsubdiffcont >>
rect 677 790 711 824
rect 773 790 807 824
rect 677 680 711 714
rect 773 680 807 714
<< mvpsubdiffcont >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
<< poly >>
rect 404 1521 504 1547
rect 560 1521 660 1547
rect 716 1521 816 1547
rect 872 1521 972 1547
rect 1028 1521 1128 1547
rect 1764 1521 1864 1547
rect 1929 1521 2029 1547
rect 1764 1345 1864 1371
rect 1764 1311 1848 1345
rect 1929 1311 2029 1371
rect 1532 1295 1848 1311
rect 1532 1261 1548 1295
rect 1582 1261 1848 1295
rect 1532 1245 1848 1261
rect 1890 1295 2029 1311
rect 1890 1261 1906 1295
rect 1940 1261 1974 1295
rect 2008 1261 2029 1295
rect 1890 1245 2029 1261
rect 1532 1227 1598 1245
rect 404 1199 504 1221
rect 560 1199 660 1221
rect 716 1199 816 1221
rect 872 1199 972 1221
rect 1028 1199 1128 1221
rect 404 1133 1128 1199
rect 1532 1193 1548 1227
rect 1582 1193 1598 1227
rect 1532 1159 1598 1193
rect 1764 1211 1848 1245
rect 1764 1185 1864 1211
rect 1929 1185 2029 1245
rect 573 1083 639 1133
rect 573 1049 589 1083
rect 623 1049 639 1083
rect 573 1015 639 1049
rect 573 981 589 1015
rect 623 981 639 1015
rect 1532 1125 1548 1159
rect 1582 1125 1598 1159
rect 1532 1091 1598 1125
rect 1532 1057 1548 1091
rect 1582 1057 1598 1091
rect 1532 995 1598 1057
rect 573 947 639 981
rect 1398 969 1598 995
rect 573 913 589 947
rect 623 913 639 947
rect 573 897 639 913
rect 1398 859 1598 885
rect 1764 859 1864 885
rect 1929 859 2029 885
rect 1433 729 1567 745
rect 1433 695 1449 729
rect 1483 695 1517 729
rect 1551 695 1567 729
rect 1433 673 1567 695
rect 1406 647 1606 673
rect 656 607 686 633
rect 742 607 772 633
rect 499 424 565 440
rect 1406 537 1606 563
rect 956 479 1821 495
rect 956 445 972 479
rect 1006 445 1040 479
rect 1074 445 1108 479
rect 1142 445 1821 479
rect 499 390 515 424
rect 549 407 565 424
rect 656 407 686 439
rect 742 407 772 439
rect 956 429 1821 445
rect 1097 407 1197 429
rect 1253 407 1353 429
rect 1409 407 1509 429
rect 1565 407 1665 429
rect 1721 407 1821 429
rect 549 390 686 407
rect 499 356 686 390
rect 499 322 515 356
rect 549 341 686 356
rect 728 391 862 407
rect 728 357 744 391
rect 778 357 812 391
rect 846 357 862 391
rect 728 341 862 357
rect 549 322 565 341
rect 499 306 565 322
rect 656 319 686 341
rect 742 319 772 341
rect 656 125 686 151
rect 742 125 772 151
rect 1097 81 1197 107
rect 1253 81 1353 107
rect 1409 81 1509 107
rect 1565 81 1665 107
rect 1721 81 1821 107
<< polycont >>
rect 1548 1261 1582 1295
rect 1906 1261 1940 1295
rect 1974 1261 2008 1295
rect 1548 1193 1582 1227
rect 589 1049 623 1083
rect 589 981 623 1015
rect 1548 1125 1582 1159
rect 1548 1057 1582 1091
rect 589 913 623 947
rect 1449 695 1483 729
rect 1517 695 1551 729
rect 972 445 1006 479
rect 1040 445 1074 479
rect 1108 445 1142 479
rect 515 390 549 424
rect 515 322 549 356
rect 744 357 778 391
rect 812 357 846 391
<< locali >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2112 1645
rect 317 1543 1059 1577
rect 317 1509 323 1543
rect 357 1509 395 1543
rect 429 1509 435 1543
rect 629 1509 635 1543
rect 669 1509 707 1543
rect 741 1509 747 1543
rect 941 1509 947 1543
rect 981 1509 1019 1543
rect 1053 1509 1059 1543
rect 1842 1543 1960 1549
rect 317 1475 359 1509
rect 393 1475 435 1509
rect 317 1429 435 1475
rect 317 1395 359 1429
rect 393 1395 435 1429
rect 317 1347 435 1395
rect 317 1313 359 1347
rect 393 1313 435 1347
rect 317 1267 435 1313
rect 317 1233 359 1267
rect 393 1233 435 1267
rect 317 1217 435 1233
rect 499 1475 515 1509
rect 549 1475 565 1509
rect 499 1429 565 1475
rect 499 1395 515 1429
rect 549 1395 565 1429
rect 499 1347 565 1395
rect 499 1313 515 1347
rect 549 1313 565 1347
rect 499 1267 565 1313
rect 499 1233 515 1267
rect 549 1233 565 1267
rect 629 1475 671 1509
rect 705 1475 747 1509
rect 629 1429 747 1475
rect 629 1395 671 1429
rect 705 1395 747 1429
rect 629 1347 747 1395
rect 629 1313 671 1347
rect 705 1313 747 1347
rect 629 1267 747 1313
rect 629 1233 671 1267
rect 705 1233 747 1267
rect 811 1475 827 1509
rect 861 1475 877 1509
rect 811 1429 877 1475
rect 811 1395 827 1429
rect 861 1395 877 1429
rect 811 1347 877 1395
rect 811 1313 827 1347
rect 861 1313 877 1347
rect 811 1267 877 1313
rect 811 1233 827 1267
rect 861 1233 877 1267
rect 941 1475 983 1509
rect 1017 1475 1059 1509
rect 941 1429 1059 1475
rect 941 1395 983 1429
rect 1017 1395 1059 1429
rect 941 1347 1059 1395
rect 941 1313 983 1347
rect 1017 1313 1059 1347
rect 941 1267 1059 1313
rect 941 1233 983 1267
rect 1017 1233 1059 1267
rect 1123 1509 1189 1525
rect 1123 1475 1139 1509
rect 1173 1475 1189 1509
rect 1123 1429 1189 1475
rect 1123 1395 1139 1429
rect 1173 1395 1189 1429
rect 1123 1347 1189 1395
rect 1123 1313 1139 1347
rect 1173 1313 1189 1347
rect 1123 1267 1189 1313
rect 1703 1509 1769 1525
rect 1703 1475 1719 1509
rect 1753 1475 1769 1509
rect 1703 1417 1769 1475
rect 1703 1383 1719 1417
rect 1753 1383 1769 1417
rect 1703 1311 1769 1383
rect 1842 1509 1848 1543
rect 1882 1509 1920 1543
rect 1954 1509 1960 1543
rect 1842 1475 1884 1509
rect 1918 1475 1960 1509
rect 1842 1417 1960 1475
rect 1842 1383 1884 1417
rect 1918 1383 1960 1417
rect 1842 1367 1960 1383
rect 2024 1509 2090 1525
rect 2024 1475 2040 1509
rect 2074 1475 2090 1509
rect 2024 1417 2090 1475
rect 2024 1383 2040 1417
rect 2074 1383 2090 1417
rect 2024 1345 2090 1383
rect 1123 1233 1139 1267
rect 1173 1233 1189 1267
rect 499 1199 565 1233
rect 811 1199 877 1233
rect 1123 1199 1189 1233
rect 1532 1295 1598 1311
rect 1532 1261 1548 1295
rect 1582 1261 1598 1295
rect 1532 1227 1598 1261
rect 1532 1199 1548 1227
rect 499 1193 1548 1199
rect 1582 1193 1598 1227
rect 499 1159 1598 1193
rect 499 1133 1548 1159
rect 577 1083 635 1099
rect 577 1049 589 1083
rect 623 1049 635 1083
rect 577 1015 635 1049
rect 577 981 589 1015
rect 623 981 635 1015
rect 577 947 635 981
rect 577 913 589 947
rect 623 913 635 947
rect 0 797 31 831
rect 65 797 160 831
rect 577 611 635 913
rect 669 824 823 840
rect 669 790 677 824
rect 711 790 773 824
rect 807 790 823 824
rect 669 714 823 790
rect 669 680 677 714
rect 711 680 773 714
rect 807 680 823 714
rect 669 655 823 680
rect 669 645 769 655
rect 687 644 769 645
rect 577 595 653 611
rect 577 561 611 595
rect 645 561 653 595
rect 577 553 653 561
rect 595 483 653 553
rect 595 449 611 483
rect 645 449 653 483
rect 499 424 561 440
rect 499 390 515 424
rect 549 390 561 424
rect 499 356 561 390
rect 499 322 515 356
rect 549 322 561 356
rect 499 306 561 322
rect 595 399 653 449
rect 687 610 697 644
rect 731 621 769 644
rect 803 621 823 655
rect 1237 693 1303 1133
rect 1532 1125 1548 1133
rect 1582 1125 1598 1159
rect 1532 1091 1598 1125
rect 1532 1057 1548 1091
rect 1582 1057 1598 1091
rect 1532 1041 1598 1057
rect 1703 1295 2008 1311
rect 1703 1261 1906 1295
rect 1940 1261 1974 1295
rect 1703 1245 2008 1261
rect 1703 1173 1769 1245
rect 2042 1211 2090 1345
rect 1703 1139 1719 1173
rect 1753 1139 1769 1173
rect 1703 1093 1769 1139
rect 1703 1059 1719 1093
rect 1753 1059 1769 1093
rect 1703 1011 1769 1059
rect 1703 977 1719 1011
rect 1753 977 1769 1011
rect 1337 944 1499 960
rect 1337 910 1353 944
rect 1387 910 1499 944
rect 1337 894 1499 910
rect 1433 761 1499 894
rect 1551 944 1669 960
rect 1551 933 1609 944
rect 1643 933 1669 944
rect 1551 899 1557 933
rect 1591 910 1609 933
rect 1591 899 1629 910
rect 1663 899 1669 933
rect 1551 881 1669 899
rect 1703 931 1769 977
rect 1703 897 1719 931
rect 1753 897 1769 931
rect 1703 881 1769 897
rect 1842 1173 1960 1189
rect 1842 1139 1884 1173
rect 1918 1139 1960 1173
rect 1842 1093 1960 1139
rect 1842 1059 1884 1093
rect 1918 1059 1960 1093
rect 1842 1011 1960 1059
rect 1842 977 1884 1011
rect 1918 977 1960 1011
rect 1842 933 1960 977
rect 1842 899 1848 933
rect 1882 931 1920 933
rect 1882 899 1884 931
rect 1842 897 1884 899
rect 1918 899 1920 931
rect 1954 899 1960 933
rect 1918 897 1960 899
rect 1842 881 1960 897
rect 2024 1173 2090 1211
rect 2024 1139 2040 1173
rect 2074 1139 2090 1173
rect 2024 1093 2090 1139
rect 2024 1059 2040 1093
rect 2074 1059 2090 1093
rect 2024 1011 2090 1059
rect 2024 977 2040 1011
rect 2074 977 2090 1011
rect 2024 931 2090 977
rect 2024 897 2040 931
rect 2074 897 2090 931
rect 2024 881 2090 897
rect 1551 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2112 831
rect 1433 729 1567 761
rect 1433 695 1449 729
rect 1483 695 1517 729
rect 1551 695 1567 729
rect 1237 677 1399 693
rect 1237 643 1349 677
rect 1383 643 1399 677
rect 1237 627 1399 643
rect 731 615 823 621
rect 731 610 741 615
rect 687 595 741 610
rect 687 561 697 595
rect 731 561 741 595
rect 1333 609 1399 627
rect 687 483 741 561
rect 687 449 697 483
rect 731 449 741 483
rect 687 433 741 449
rect 775 565 837 581
rect 775 531 783 565
rect 817 531 837 565
rect 1333 575 1361 609
rect 1395 575 1399 609
rect 1333 559 1399 575
rect 1433 679 1567 695
rect 1601 729 1719 741
rect 1601 695 1607 729
rect 1641 695 1679 729
rect 1713 695 1719 729
rect 775 495 837 531
rect 1433 495 1499 679
rect 1601 677 1719 695
rect 1601 643 1629 677
rect 1663 643 1719 677
rect 1601 609 1719 643
rect 1601 575 1617 609
rect 1651 575 1719 609
rect 1601 559 1719 575
rect 775 483 1158 495
rect 775 449 783 483
rect 817 479 1158 483
rect 817 449 972 479
rect 775 445 972 449
rect 1006 445 1040 479
rect 1074 445 1108 479
rect 1142 445 1158 479
rect 775 433 1158 445
rect 896 429 1158 433
rect 1192 429 1882 495
rect 595 391 862 399
rect 595 357 744 391
rect 778 357 812 391
rect 846 357 862 391
rect 595 349 862 357
rect 595 299 653 349
rect 896 315 962 429
rect 1192 395 1258 429
rect 1504 395 1570 429
rect 1816 395 1882 429
rect 595 265 611 299
rect 645 265 653 299
rect 595 197 653 265
rect 595 163 611 197
rect 645 163 653 197
rect 595 147 653 163
rect 687 299 741 315
rect 687 265 697 299
rect 731 265 741 299
rect 687 193 741 265
rect 687 159 697 193
rect 731 159 741 193
rect 687 119 741 159
rect 775 299 962 315
rect 775 265 783 299
rect 817 265 962 299
rect 775 249 962 265
rect 1010 361 1052 395
rect 1086 361 1128 395
rect 1010 315 1128 361
rect 1010 281 1052 315
rect 1086 281 1128 315
rect 775 197 837 249
rect 775 163 783 197
rect 817 163 837 197
rect 775 147 837 163
rect 1010 233 1128 281
rect 1010 199 1052 233
rect 1086 199 1128 233
rect 1010 153 1128 199
rect 687 113 697 119
rect 619 107 697 113
rect 619 73 625 107
rect 659 85 697 107
rect 731 113 741 119
rect 1010 119 1052 153
rect 1086 119 1128 153
rect 1192 361 1208 395
rect 1242 361 1258 395
rect 1192 315 1258 361
rect 1192 281 1208 315
rect 1242 281 1258 315
rect 1192 233 1258 281
rect 1192 199 1208 233
rect 1242 199 1258 233
rect 1192 153 1258 199
rect 1192 119 1208 153
rect 1242 119 1258 153
rect 1322 361 1364 395
rect 1398 361 1440 395
rect 1322 315 1440 361
rect 1322 281 1364 315
rect 1398 281 1440 315
rect 1322 233 1440 281
rect 1322 199 1364 233
rect 1398 199 1440 233
rect 1322 153 1440 199
rect 1322 119 1364 153
rect 1398 119 1440 153
rect 1504 361 1520 395
rect 1554 361 1570 395
rect 1504 315 1570 361
rect 1504 281 1520 315
rect 1554 281 1570 315
rect 1504 233 1570 281
rect 1504 199 1520 233
rect 1554 199 1570 233
rect 1504 153 1570 199
rect 1504 119 1520 153
rect 1554 119 1570 153
rect 1634 361 1676 395
rect 1710 361 1752 395
rect 1634 315 1752 361
rect 1634 281 1676 315
rect 1710 281 1752 315
rect 1634 233 1752 281
rect 1634 199 1676 233
rect 1710 199 1752 233
rect 1634 153 1752 199
rect 1634 119 1676 153
rect 1710 119 1752 153
rect 731 107 809 113
rect 731 85 769 107
rect 659 73 769 85
rect 803 73 809 107
rect 619 67 809 73
rect 1010 85 1016 119
rect 1050 85 1088 119
rect 1122 85 1128 119
rect 1322 85 1328 119
rect 1362 85 1400 119
rect 1434 85 1440 119
rect 1634 85 1640 119
rect 1674 85 1712 119
rect 1746 85 1752 119
rect 1816 361 1832 395
rect 1866 361 1882 395
rect 1816 315 1882 361
rect 1816 281 1832 315
rect 1866 281 1882 315
rect 1816 233 1882 281
rect 1816 199 1832 233
rect 1866 199 1882 233
rect 1816 153 1882 199
rect 1816 119 1832 153
rect 1866 119 1882 153
rect 1816 103 1882 119
rect 1010 51 1752 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 323 1509 357 1543
rect 395 1509 429 1543
rect 635 1509 669 1543
rect 707 1509 741 1543
rect 947 1509 981 1543
rect 1019 1509 1053 1543
rect 1848 1509 1882 1543
rect 1920 1509 1954 1543
rect 31 797 65 831
rect 697 610 731 644
rect 769 621 803 655
rect 1557 899 1591 933
rect 1629 910 1643 933
rect 1643 910 1663 933
rect 1629 899 1663 910
rect 1848 899 1882 933
rect 1920 899 1954 933
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 1607 695 1641 729
rect 1679 695 1713 729
rect 625 73 659 107
rect 697 85 731 119
rect 769 73 803 107
rect 1016 85 1050 119
rect 1088 85 1122 119
rect 1328 85 1362 119
rect 1400 85 1434 119
rect 1640 85 1674 119
rect 1712 85 1746 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 1645 2112 1651
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2112 1645
rect 0 1605 2112 1611
rect 0 1543 2112 1577
rect 0 1509 323 1543
rect 357 1509 395 1543
rect 429 1509 635 1543
rect 669 1509 707 1543
rect 741 1509 947 1543
rect 981 1509 1019 1543
rect 1053 1509 1848 1543
rect 1882 1509 1920 1543
rect 1954 1509 2112 1543
rect 0 1503 2112 1509
rect 0 933 2112 939
rect 0 899 1557 933
rect 1591 899 1629 933
rect 1663 899 1848 933
rect 1882 899 1920 933
rect 1954 899 2112 933
rect 0 865 2112 899
rect 0 831 2112 837
rect 0 797 31 831
rect 65 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2112 831
rect 0 791 2112 797
rect 0 729 2112 763
rect 0 695 1607 729
rect 1641 695 1679 729
rect 1713 695 2112 729
rect 0 689 2112 695
rect 14 655 2098 661
rect 14 644 769 655
rect 14 610 697 644
rect 731 621 769 644
rect 803 621 2098 655
rect 731 610 2098 621
rect 14 604 2098 610
rect 0 119 2112 125
rect 0 107 697 119
rect 0 73 625 107
rect 659 85 697 107
rect 731 107 1016 119
rect 731 85 769 107
rect 659 73 769 85
rect 803 85 1016 107
rect 1050 85 1088 119
rect 1122 85 1328 119
rect 1362 85 1400 119
rect 1434 85 1640 119
rect 1674 85 1712 119
rect 1746 85 2112 119
rect 803 73 2112 85
rect 0 51 2112 73
rect 0 17 2112 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -23 2112 -17
<< labels >>
rlabel comment s 0 0 0 0 4 lsbuflv2hv_1
flabel metal1 s 0 865 2112 939 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 689 2112 763 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 1503 2112 1577 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 51 2112 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 2112 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 14 604 2098 661 0 FreeSans 340 0 0 0 LVPWR
port 2 nsew power bidirectional
flabel metal1 s 0 791 2112 837 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 1605 2112 1628 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2047 1204 2081 1238 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2047 1130 2081 1164 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2047 1056 2081 1090 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2047 1278 2081 1312 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2047 1352 2081 1386 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unithvdbl
string LEFclass CORE
string FIXED_BBOX 0 0 2112 1628
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string LEFsymmetry X Y
string GDS_END 326888
string GDS_START 303650
<< end >>
