magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1302 -1364 41238 1680
<< metal1 >>
rect 78 0 114 395
rect 150 0 186 395
rect 222 79 258 420
rect 294 0 330 395
rect 366 0 402 395
rect 846 0 882 395
rect 918 0 954 395
rect 990 79 1026 420
rect 1062 0 1098 395
rect 1134 0 1170 395
rect 1326 0 1362 395
rect 1398 0 1434 395
rect 1470 79 1506 420
rect 1542 0 1578 395
rect 1614 0 1650 395
rect 2094 0 2130 395
rect 2166 0 2202 395
rect 2238 79 2274 420
rect 2310 0 2346 395
rect 2382 0 2418 395
rect 2574 0 2610 395
rect 2646 0 2682 395
rect 2718 79 2754 420
rect 2790 0 2826 395
rect 2862 0 2898 395
rect 3342 0 3378 395
rect 3414 0 3450 395
rect 3486 79 3522 420
rect 3558 0 3594 395
rect 3630 0 3666 395
rect 3822 0 3858 395
rect 3894 0 3930 395
rect 3966 79 4002 420
rect 4038 0 4074 395
rect 4110 0 4146 395
rect 4590 0 4626 395
rect 4662 0 4698 395
rect 4734 79 4770 420
rect 4806 0 4842 395
rect 4878 0 4914 395
rect 5070 0 5106 395
rect 5142 0 5178 395
rect 5214 79 5250 420
rect 5286 0 5322 395
rect 5358 0 5394 395
rect 5838 0 5874 395
rect 5910 0 5946 395
rect 5982 79 6018 420
rect 6054 0 6090 395
rect 6126 0 6162 395
rect 6318 0 6354 395
rect 6390 0 6426 395
rect 6462 79 6498 420
rect 6534 0 6570 395
rect 6606 0 6642 395
rect 7086 0 7122 395
rect 7158 0 7194 395
rect 7230 79 7266 420
rect 7302 0 7338 395
rect 7374 0 7410 395
rect 7566 0 7602 395
rect 7638 0 7674 395
rect 7710 79 7746 420
rect 7782 0 7818 395
rect 7854 0 7890 395
rect 8334 0 8370 395
rect 8406 0 8442 395
rect 8478 79 8514 420
rect 8550 0 8586 395
rect 8622 0 8658 395
rect 8814 0 8850 395
rect 8886 0 8922 395
rect 8958 79 8994 420
rect 9030 0 9066 395
rect 9102 0 9138 395
rect 9582 0 9618 395
rect 9654 0 9690 395
rect 9726 79 9762 420
rect 9798 0 9834 395
rect 9870 0 9906 395
rect 10062 0 10098 395
rect 10134 0 10170 395
rect 10206 79 10242 420
rect 10278 0 10314 395
rect 10350 0 10386 395
rect 10830 0 10866 395
rect 10902 0 10938 395
rect 10974 79 11010 420
rect 11046 0 11082 395
rect 11118 0 11154 395
rect 11310 0 11346 395
rect 11382 0 11418 395
rect 11454 79 11490 420
rect 11526 0 11562 395
rect 11598 0 11634 395
rect 12078 0 12114 395
rect 12150 0 12186 395
rect 12222 79 12258 420
rect 12294 0 12330 395
rect 12366 0 12402 395
rect 12558 0 12594 395
rect 12630 0 12666 395
rect 12702 79 12738 420
rect 12774 0 12810 395
rect 12846 0 12882 395
rect 13326 0 13362 395
rect 13398 0 13434 395
rect 13470 79 13506 420
rect 13542 0 13578 395
rect 13614 0 13650 395
rect 13806 0 13842 395
rect 13878 0 13914 395
rect 13950 79 13986 420
rect 14022 0 14058 395
rect 14094 0 14130 395
rect 14574 0 14610 395
rect 14646 0 14682 395
rect 14718 79 14754 420
rect 14790 0 14826 395
rect 14862 0 14898 395
rect 15054 0 15090 395
rect 15126 0 15162 395
rect 15198 79 15234 420
rect 15270 0 15306 395
rect 15342 0 15378 395
rect 15822 0 15858 395
rect 15894 0 15930 395
rect 15966 79 16002 420
rect 16038 0 16074 395
rect 16110 0 16146 395
rect 16302 0 16338 395
rect 16374 0 16410 395
rect 16446 79 16482 420
rect 16518 0 16554 395
rect 16590 0 16626 395
rect 17070 0 17106 395
rect 17142 0 17178 395
rect 17214 79 17250 420
rect 17286 0 17322 395
rect 17358 0 17394 395
rect 17550 0 17586 395
rect 17622 0 17658 395
rect 17694 79 17730 420
rect 17766 0 17802 395
rect 17838 0 17874 395
rect 18318 0 18354 395
rect 18390 0 18426 395
rect 18462 79 18498 420
rect 18534 0 18570 395
rect 18606 0 18642 395
rect 18798 0 18834 395
rect 18870 0 18906 395
rect 18942 79 18978 420
rect 19014 0 19050 395
rect 19086 0 19122 395
rect 19566 0 19602 395
rect 19638 0 19674 395
rect 19710 79 19746 420
rect 19782 0 19818 395
rect 19854 0 19890 395
rect 20046 0 20082 395
rect 20118 0 20154 395
rect 20190 79 20226 420
rect 20262 0 20298 395
rect 20334 0 20370 395
rect 20814 0 20850 395
rect 20886 0 20922 395
rect 20958 79 20994 420
rect 21030 0 21066 395
rect 21102 0 21138 395
rect 21294 0 21330 395
rect 21366 0 21402 395
rect 21438 79 21474 420
rect 21510 0 21546 395
rect 21582 0 21618 395
rect 22062 0 22098 395
rect 22134 0 22170 395
rect 22206 79 22242 420
rect 22278 0 22314 395
rect 22350 0 22386 395
rect 22542 0 22578 395
rect 22614 0 22650 395
rect 22686 79 22722 420
rect 22758 0 22794 395
rect 22830 0 22866 395
rect 23310 0 23346 395
rect 23382 0 23418 395
rect 23454 79 23490 420
rect 23526 0 23562 395
rect 23598 0 23634 395
rect 23790 0 23826 395
rect 23862 0 23898 395
rect 23934 79 23970 420
rect 24006 0 24042 395
rect 24078 0 24114 395
rect 24558 0 24594 395
rect 24630 0 24666 395
rect 24702 79 24738 420
rect 24774 0 24810 395
rect 24846 0 24882 395
rect 25038 0 25074 395
rect 25110 0 25146 395
rect 25182 79 25218 420
rect 25254 0 25290 395
rect 25326 0 25362 395
rect 25806 0 25842 395
rect 25878 0 25914 395
rect 25950 79 25986 420
rect 26022 0 26058 395
rect 26094 0 26130 395
rect 26286 0 26322 395
rect 26358 0 26394 395
rect 26430 79 26466 420
rect 26502 0 26538 395
rect 26574 0 26610 395
rect 27054 0 27090 395
rect 27126 0 27162 395
rect 27198 79 27234 420
rect 27270 0 27306 395
rect 27342 0 27378 395
rect 27534 0 27570 395
rect 27606 0 27642 395
rect 27678 79 27714 420
rect 27750 0 27786 395
rect 27822 0 27858 395
rect 28302 0 28338 395
rect 28374 0 28410 395
rect 28446 79 28482 420
rect 28518 0 28554 395
rect 28590 0 28626 395
rect 28782 0 28818 395
rect 28854 0 28890 395
rect 28926 79 28962 420
rect 28998 0 29034 395
rect 29070 0 29106 395
rect 29550 0 29586 395
rect 29622 0 29658 395
rect 29694 79 29730 420
rect 29766 0 29802 395
rect 29838 0 29874 395
rect 30030 0 30066 395
rect 30102 0 30138 395
rect 30174 79 30210 420
rect 30246 0 30282 395
rect 30318 0 30354 395
rect 30798 0 30834 395
rect 30870 0 30906 395
rect 30942 79 30978 420
rect 31014 0 31050 395
rect 31086 0 31122 395
rect 31278 0 31314 395
rect 31350 0 31386 395
rect 31422 79 31458 420
rect 31494 0 31530 395
rect 31566 0 31602 395
rect 32046 0 32082 395
rect 32118 0 32154 395
rect 32190 79 32226 420
rect 32262 0 32298 395
rect 32334 0 32370 395
rect 32526 0 32562 395
rect 32598 0 32634 395
rect 32670 79 32706 420
rect 32742 0 32778 395
rect 32814 0 32850 395
rect 33294 0 33330 395
rect 33366 0 33402 395
rect 33438 79 33474 420
rect 33510 0 33546 395
rect 33582 0 33618 395
rect 33774 0 33810 395
rect 33846 0 33882 395
rect 33918 79 33954 420
rect 33990 0 34026 395
rect 34062 0 34098 395
rect 34542 0 34578 395
rect 34614 0 34650 395
rect 34686 79 34722 420
rect 34758 0 34794 395
rect 34830 0 34866 395
rect 35022 0 35058 395
rect 35094 0 35130 395
rect 35166 79 35202 420
rect 35238 0 35274 395
rect 35310 0 35346 395
rect 35790 0 35826 395
rect 35862 0 35898 395
rect 35934 79 35970 420
rect 36006 0 36042 395
rect 36078 0 36114 395
rect 36270 0 36306 395
rect 36342 0 36378 395
rect 36414 79 36450 420
rect 36486 0 36522 395
rect 36558 0 36594 395
rect 37038 0 37074 395
rect 37110 0 37146 395
rect 37182 79 37218 420
rect 37254 0 37290 395
rect 37326 0 37362 395
rect 37518 0 37554 395
rect 37590 0 37626 395
rect 37662 79 37698 420
rect 37734 0 37770 395
rect 37806 0 37842 395
rect 38286 0 38322 395
rect 38358 0 38394 395
rect 38430 79 38466 420
rect 38502 0 38538 395
rect 38574 0 38610 395
rect 38766 0 38802 395
rect 38838 0 38874 395
rect 38910 79 38946 420
rect 38982 0 39018 395
rect 39054 0 39090 395
rect 39534 0 39570 395
rect 39606 0 39642 395
rect 39678 79 39714 420
rect 39750 0 39786 395
rect 39822 0 39858 395
<< metal2 >>
rect 0 323 39936 371
rect 186 199 294 275
rect 954 199 1062 275
rect 1434 199 1542 275
rect 2202 199 2310 275
rect 2682 199 2790 275
rect 3450 199 3558 275
rect 3930 199 4038 275
rect 4698 199 4806 275
rect 5178 199 5286 275
rect 5946 199 6054 275
rect 6426 199 6534 275
rect 7194 199 7302 275
rect 7674 199 7782 275
rect 8442 199 8550 275
rect 8922 199 9030 275
rect 9690 199 9798 275
rect 10170 199 10278 275
rect 10938 199 11046 275
rect 11418 199 11526 275
rect 12186 199 12294 275
rect 12666 199 12774 275
rect 13434 199 13542 275
rect 13914 199 14022 275
rect 14682 199 14790 275
rect 15162 199 15270 275
rect 15930 199 16038 275
rect 16410 199 16518 275
rect 17178 199 17286 275
rect 17658 199 17766 275
rect 18426 199 18534 275
rect 18906 199 19014 275
rect 19674 199 19782 275
rect 20154 199 20262 275
rect 20922 199 21030 275
rect 21402 199 21510 275
rect 22170 199 22278 275
rect 22650 199 22758 275
rect 23418 199 23526 275
rect 23898 199 24006 275
rect 24666 199 24774 275
rect 25146 199 25254 275
rect 25914 199 26022 275
rect 26394 199 26502 275
rect 27162 199 27270 275
rect 27642 199 27750 275
rect 28410 199 28518 275
rect 28890 199 28998 275
rect 29658 199 29766 275
rect 30138 199 30246 275
rect 30906 199 31014 275
rect 31386 199 31494 275
rect 32154 199 32262 275
rect 32634 199 32742 275
rect 33402 199 33510 275
rect 33882 199 33990 275
rect 34650 199 34758 275
rect 35130 199 35238 275
rect 35898 199 36006 275
rect 36378 199 36486 275
rect 37146 199 37254 275
rect 37626 199 37734 275
rect 38394 199 38502 275
rect 38874 199 38982 275
rect 39642 199 39750 275
rect 0 103 39936 151
rect 186 -55 294 55
rect 954 -55 1062 55
rect 1434 -55 1542 55
rect 2202 -55 2310 55
rect 2682 -55 2790 55
rect 3450 -55 3558 55
rect 3930 -55 4038 55
rect 4698 -55 4806 55
rect 5178 -55 5286 55
rect 5946 -55 6054 55
rect 6426 -55 6534 55
rect 7194 -55 7302 55
rect 7674 -55 7782 55
rect 8442 -55 8550 55
rect 8922 -55 9030 55
rect 9690 -55 9798 55
rect 10170 -55 10278 55
rect 10938 -55 11046 55
rect 11418 -55 11526 55
rect 12186 -55 12294 55
rect 12666 -55 12774 55
rect 13434 -55 13542 55
rect 13914 -55 14022 55
rect 14682 -55 14790 55
rect 15162 -55 15270 55
rect 15930 -55 16038 55
rect 16410 -55 16518 55
rect 17178 -55 17286 55
rect 17658 -55 17766 55
rect 18426 -55 18534 55
rect 18906 -55 19014 55
rect 19674 -55 19782 55
rect 20154 -55 20262 55
rect 20922 -55 21030 55
rect 21402 -55 21510 55
rect 22170 -55 22278 55
rect 22650 -55 22758 55
rect 23418 -55 23526 55
rect 23898 -55 24006 55
rect 24666 -55 24774 55
rect 25146 -55 25254 55
rect 25914 -55 26022 55
rect 26394 -55 26502 55
rect 27162 -55 27270 55
rect 27642 -55 27750 55
rect 28410 -55 28518 55
rect 28890 -55 28998 55
rect 29658 -55 29766 55
rect 30138 -55 30246 55
rect 30906 -55 31014 55
rect 31386 -55 31494 55
rect 32154 -55 32262 55
rect 32634 -55 32742 55
rect 33402 -55 33510 55
rect 33882 -55 33990 55
rect 34650 -55 34758 55
rect 35130 -55 35238 55
rect 35898 -55 36006 55
rect 36378 -55 36486 55
rect 37146 -55 37254 55
rect 37626 -55 37734 55
rect 38394 -55 38502 55
rect 38874 -55 38982 55
rect 39642 -55 39750 55
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_63
timestamp 1624857261
transform 1 0 0 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_62
timestamp 1624857261
transform -1 0 1248 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_61
timestamp 1624857261
transform 1 0 1248 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_60
timestamp 1624857261
transform -1 0 2496 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_59
timestamp 1624857261
transform 1 0 2496 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_58
timestamp 1624857261
transform -1 0 3744 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_57
timestamp 1624857261
transform 1 0 3744 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_56
timestamp 1624857261
transform -1 0 4992 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_55
timestamp 1624857261
transform 1 0 4992 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_54
timestamp 1624857261
transform -1 0 6240 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_53
timestamp 1624857261
transform 1 0 6240 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_52
timestamp 1624857261
transform -1 0 7488 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_51
timestamp 1624857261
transform 1 0 7488 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_50
timestamp 1624857261
transform -1 0 8736 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_49
timestamp 1624857261
transform 1 0 8736 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_48
timestamp 1624857261
transform -1 0 9984 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_47
timestamp 1624857261
transform 1 0 9984 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_46
timestamp 1624857261
transform -1 0 11232 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_45
timestamp 1624857261
transform 1 0 11232 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_44
timestamp 1624857261
transform -1 0 12480 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_43
timestamp 1624857261
transform 1 0 12480 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_42
timestamp 1624857261
transform -1 0 13728 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_41
timestamp 1624857261
transform 1 0 13728 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_40
timestamp 1624857261
transform -1 0 14976 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_39
timestamp 1624857261
transform 1 0 14976 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_38
timestamp 1624857261
transform -1 0 16224 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_37
timestamp 1624857261
transform 1 0 16224 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_36
timestamp 1624857261
transform -1 0 17472 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_35
timestamp 1624857261
transform 1 0 17472 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_34
timestamp 1624857261
transform -1 0 18720 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_33
timestamp 1624857261
transform 1 0 18720 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_32
timestamp 1624857261
transform -1 0 19968 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_31
timestamp 1624857261
transform 1 0 19968 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_30
timestamp 1624857261
transform -1 0 21216 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_29
timestamp 1624857261
transform 1 0 21216 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_28
timestamp 1624857261
transform -1 0 22464 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_27
timestamp 1624857261
transform 1 0 22464 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_26
timestamp 1624857261
transform -1 0 23712 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_25
timestamp 1624857261
transform 1 0 23712 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_24
timestamp 1624857261
transform -1 0 24960 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_23
timestamp 1624857261
transform 1 0 24960 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_22
timestamp 1624857261
transform -1 0 26208 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_21
timestamp 1624857261
transform 1 0 26208 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_20
timestamp 1624857261
transform -1 0 27456 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_19
timestamp 1624857261
transform 1 0 27456 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_18
timestamp 1624857261
transform -1 0 28704 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_17
timestamp 1624857261
transform 1 0 28704 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_16
timestamp 1624857261
transform -1 0 29952 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_15
timestamp 1624857261
transform 1 0 29952 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_14
timestamp 1624857261
transform -1 0 31200 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_13
timestamp 1624857261
transform 1 0 31200 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_12
timestamp 1624857261
transform -1 0 32448 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_11
timestamp 1624857261
transform 1 0 32448 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_10
timestamp 1624857261
transform -1 0 33696 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_9
timestamp 1624857261
transform 1 0 33696 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_8
timestamp 1624857261
transform -1 0 34944 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_7
timestamp 1624857261
transform 1 0 34944 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_6
timestamp 1624857261
transform -1 0 36192 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_5
timestamp 1624857261
transform 1 0 36192 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_4
timestamp 1624857261
transform -1 0 37440 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_3
timestamp 1624857261
transform 1 0 37440 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_2
timestamp 1624857261
transform -1 0 38688 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_1
timestamp 1624857261
transform 1 0 38688 0 1 0
box -42 -104 624 420
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1624857261
transform -1 0 39936 0 1 0
box -42 -104 624 420
<< labels >>
rlabel metal1 s 78 0 114 395 4 bl_0_0
port 261 se
rlabel metal1 s 150 0 186 395 4 br_0_0
port 263 se
rlabel metal1 s 294 0 330 395 4 bl_1_0
port 262 se
rlabel metal1 s 366 0 402 395 4 br_1_0
port 264 se
rlabel metal1 s 1134 0 1170 395 4 bl_0_1
port 265 se
rlabel metal1 s 1062 0 1098 395 4 br_0_1
port 267 se
rlabel metal1 s 918 0 954 395 4 bl_1_1
port 266 se
rlabel metal1 s 846 0 882 395 4 br_1_1
port 268 se
rlabel metal1 s 1326 0 1362 395 4 bl_0_2
port 269 se
rlabel metal1 s 1398 0 1434 395 4 br_0_2
port 271 se
rlabel metal1 s 1542 0 1578 395 4 bl_1_2
port 270 se
rlabel metal1 s 1614 0 1650 395 4 br_1_2
port 272 se
rlabel metal1 s 2382 0 2418 395 4 bl_0_3
port 273 se
rlabel metal1 s 2310 0 2346 395 4 br_0_3
port 275 se
rlabel metal1 s 2166 0 2202 395 4 bl_1_3
port 274 se
rlabel metal1 s 2094 0 2130 395 4 br_1_3
port 276 se
rlabel metal1 s 2574 0 2610 395 4 bl_0_4
port 277 se
rlabel metal1 s 2646 0 2682 395 4 br_0_4
port 279 se
rlabel metal1 s 2790 0 2826 395 4 bl_1_4
port 278 se
rlabel metal1 s 2862 0 2898 395 4 br_1_4
port 280 se
rlabel metal1 s 3630 0 3666 395 4 bl_0_5
port 281 se
rlabel metal1 s 3558 0 3594 395 4 br_0_5
port 283 se
rlabel metal1 s 3414 0 3450 395 4 bl_1_5
port 282 se
rlabel metal1 s 3342 0 3378 395 4 br_1_5
port 284 se
rlabel metal1 s 3822 0 3858 395 4 bl_0_6
port 285 se
rlabel metal1 s 3894 0 3930 395 4 br_0_6
port 287 se
rlabel metal1 s 4038 0 4074 395 4 bl_1_6
port 286 se
rlabel metal1 s 4110 0 4146 395 4 br_1_6
port 288 se
rlabel metal1 s 4878 0 4914 395 4 bl_0_7
port 289 se
rlabel metal1 s 4806 0 4842 395 4 br_0_7
port 291 se
rlabel metal1 s 4662 0 4698 395 4 bl_1_7
port 290 se
rlabel metal1 s 4590 0 4626 395 4 br_1_7
port 292 se
rlabel metal1 s 5070 0 5106 395 4 bl_0_8
port 293 se
rlabel metal1 s 5142 0 5178 395 4 br_0_8
port 295 se
rlabel metal1 s 5286 0 5322 395 4 bl_1_8
port 294 se
rlabel metal1 s 5358 0 5394 395 4 br_1_8
port 296 se
rlabel metal1 s 6126 0 6162 395 4 bl_0_9
port 297 se
rlabel metal1 s 6054 0 6090 395 4 br_0_9
port 299 se
rlabel metal1 s 5910 0 5946 395 4 bl_1_9
port 298 se
rlabel metal1 s 5838 0 5874 395 4 br_1_9
port 300 se
rlabel metal1 s 6318 0 6354 395 4 bl_0_10
port 301 se
rlabel metal1 s 6390 0 6426 395 4 br_0_10
port 303 se
rlabel metal1 s 6534 0 6570 395 4 bl_1_10
port 302 se
rlabel metal1 s 6606 0 6642 395 4 br_1_10
port 304 se
rlabel metal1 s 7374 0 7410 395 4 bl_0_11
port 305 se
rlabel metal1 s 7302 0 7338 395 4 br_0_11
port 307 se
rlabel metal1 s 7158 0 7194 395 4 bl_1_11
port 306 se
rlabel metal1 s 7086 0 7122 395 4 br_1_11
port 308 se
rlabel metal1 s 7566 0 7602 395 4 bl_0_12
port 309 se
rlabel metal1 s 7638 0 7674 395 4 br_0_12
port 311 se
rlabel metal1 s 7782 0 7818 395 4 bl_1_12
port 310 se
rlabel metal1 s 7854 0 7890 395 4 br_1_12
port 312 se
rlabel metal1 s 8622 0 8658 395 4 bl_0_13
port 313 se
rlabel metal1 s 8550 0 8586 395 4 br_0_13
port 315 se
rlabel metal1 s 8406 0 8442 395 4 bl_1_13
port 314 se
rlabel metal1 s 8334 0 8370 395 4 br_1_13
port 316 se
rlabel metal1 s 8814 0 8850 395 4 bl_0_14
port 317 se
rlabel metal1 s 8886 0 8922 395 4 br_0_14
port 319 se
rlabel metal1 s 9030 0 9066 395 4 bl_1_14
port 318 se
rlabel metal1 s 9102 0 9138 395 4 br_1_14
port 320 se
rlabel metal1 s 9870 0 9906 395 4 bl_0_15
port 321 se
rlabel metal1 s 9798 0 9834 395 4 br_0_15
port 323 se
rlabel metal1 s 9654 0 9690 395 4 bl_1_15
port 322 se
rlabel metal1 s 9582 0 9618 395 4 br_1_15
port 324 se
rlabel metal1 s 10062 0 10098 395 4 bl_0_16
port 325 se
rlabel metal1 s 10134 0 10170 395 4 br_0_16
port 327 se
rlabel metal1 s 10278 0 10314 395 4 bl_1_16
port 326 se
rlabel metal1 s 10350 0 10386 395 4 br_1_16
port 328 se
rlabel metal1 s 11118 0 11154 395 4 bl_0_17
port 329 se
rlabel metal1 s 11046 0 11082 395 4 br_0_17
port 331 se
rlabel metal1 s 10902 0 10938 395 4 bl_1_17
port 330 se
rlabel metal1 s 10830 0 10866 395 4 br_1_17
port 332 se
rlabel metal1 s 11310 0 11346 395 4 bl_0_18
port 333 se
rlabel metal1 s 11382 0 11418 395 4 br_0_18
port 335 se
rlabel metal1 s 11526 0 11562 395 4 bl_1_18
port 334 se
rlabel metal1 s 11598 0 11634 395 4 br_1_18
port 336 se
rlabel metal1 s 12366 0 12402 395 4 bl_0_19
port 337 se
rlabel metal1 s 12294 0 12330 395 4 br_0_19
port 339 se
rlabel metal1 s 12150 0 12186 395 4 bl_1_19
port 338 se
rlabel metal1 s 12078 0 12114 395 4 br_1_19
port 340 se
rlabel metal1 s 12558 0 12594 395 4 bl_0_20
port 341 se
rlabel metal1 s 12630 0 12666 395 4 br_0_20
port 343 se
rlabel metal1 s 12774 0 12810 395 4 bl_1_20
port 342 se
rlabel metal1 s 12846 0 12882 395 4 br_1_20
port 344 se
rlabel metal1 s 13614 0 13650 395 4 bl_0_21
port 345 se
rlabel metal1 s 13542 0 13578 395 4 br_0_21
port 347 se
rlabel metal1 s 13398 0 13434 395 4 bl_1_21
port 346 se
rlabel metal1 s 13326 0 13362 395 4 br_1_21
port 348 se
rlabel metal1 s 13806 0 13842 395 4 bl_0_22
port 349 se
rlabel metal1 s 13878 0 13914 395 4 br_0_22
port 351 se
rlabel metal1 s 14022 0 14058 395 4 bl_1_22
port 350 se
rlabel metal1 s 14094 0 14130 395 4 br_1_22
port 352 se
rlabel metal1 s 14862 0 14898 395 4 bl_0_23
port 353 se
rlabel metal1 s 14790 0 14826 395 4 br_0_23
port 355 se
rlabel metal1 s 14646 0 14682 395 4 bl_1_23
port 354 se
rlabel metal1 s 14574 0 14610 395 4 br_1_23
port 356 se
rlabel metal1 s 15054 0 15090 395 4 bl_0_24
port 357 se
rlabel metal1 s 15126 0 15162 395 4 br_0_24
port 359 se
rlabel metal1 s 15270 0 15306 395 4 bl_1_24
port 358 se
rlabel metal1 s 15342 0 15378 395 4 br_1_24
port 360 se
rlabel metal1 s 16110 0 16146 395 4 bl_0_25
port 361 se
rlabel metal1 s 16038 0 16074 395 4 br_0_25
port 363 se
rlabel metal1 s 15894 0 15930 395 4 bl_1_25
port 362 se
rlabel metal1 s 15822 0 15858 395 4 br_1_25
port 364 se
rlabel metal1 s 16302 0 16338 395 4 bl_0_26
port 365 se
rlabel metal1 s 16374 0 16410 395 4 br_0_26
port 367 se
rlabel metal1 s 16518 0 16554 395 4 bl_1_26
port 366 se
rlabel metal1 s 16590 0 16626 395 4 br_1_26
port 368 se
rlabel metal1 s 17358 0 17394 395 4 bl_0_27
port 369 se
rlabel metal1 s 17286 0 17322 395 4 br_0_27
port 371 se
rlabel metal1 s 17142 0 17178 395 4 bl_1_27
port 370 se
rlabel metal1 s 17070 0 17106 395 4 br_1_27
port 372 se
rlabel metal1 s 17550 0 17586 395 4 bl_0_28
port 373 se
rlabel metal1 s 17622 0 17658 395 4 br_0_28
port 375 se
rlabel metal1 s 17766 0 17802 395 4 bl_1_28
port 374 se
rlabel metal1 s 17838 0 17874 395 4 br_1_28
port 376 se
rlabel metal1 s 18606 0 18642 395 4 bl_0_29
port 377 se
rlabel metal1 s 18534 0 18570 395 4 br_0_29
port 379 se
rlabel metal1 s 18390 0 18426 395 4 bl_1_29
port 378 se
rlabel metal1 s 18318 0 18354 395 4 br_1_29
port 380 se
rlabel metal1 s 18798 0 18834 395 4 bl_0_30
port 381 se
rlabel metal1 s 18870 0 18906 395 4 br_0_30
port 383 se
rlabel metal1 s 19014 0 19050 395 4 bl_1_30
port 382 se
rlabel metal1 s 19086 0 19122 395 4 br_1_30
port 384 se
rlabel metal1 s 19854 0 19890 395 4 bl_0_31
port 385 se
rlabel metal1 s 19782 0 19818 395 4 br_0_31
port 387 se
rlabel metal1 s 19638 0 19674 395 4 bl_1_31
port 386 se
rlabel metal1 s 19566 0 19602 395 4 br_1_31
port 388 se
rlabel metal1 s 20046 0 20082 395 4 bl_0_32
port 389 se
rlabel metal1 s 20118 0 20154 395 4 br_0_32
port 391 se
rlabel metal1 s 20262 0 20298 395 4 bl_1_32
port 390 se
rlabel metal1 s 20334 0 20370 395 4 br_1_32
port 392 se
rlabel metal1 s 21102 0 21138 395 4 bl_0_33
port 393 se
rlabel metal1 s 21030 0 21066 395 4 br_0_33
port 395 se
rlabel metal1 s 20886 0 20922 395 4 bl_1_33
port 394 se
rlabel metal1 s 20814 0 20850 395 4 br_1_33
port 396 se
rlabel metal1 s 21294 0 21330 395 4 bl_0_34
port 397 se
rlabel metal1 s 21366 0 21402 395 4 br_0_34
port 399 se
rlabel metal1 s 21510 0 21546 395 4 bl_1_34
port 398 se
rlabel metal1 s 21582 0 21618 395 4 br_1_34
port 400 se
rlabel metal1 s 22350 0 22386 395 4 bl_0_35
port 401 se
rlabel metal1 s 22278 0 22314 395 4 br_0_35
port 403 se
rlabel metal1 s 22134 0 22170 395 4 bl_1_35
port 402 se
rlabel metal1 s 22062 0 22098 395 4 br_1_35
port 404 se
rlabel metal1 s 22542 0 22578 395 4 bl_0_36
port 405 se
rlabel metal1 s 22614 0 22650 395 4 br_0_36
port 407 se
rlabel metal1 s 22758 0 22794 395 4 bl_1_36
port 406 se
rlabel metal1 s 22830 0 22866 395 4 br_1_36
port 408 se
rlabel metal1 s 23598 0 23634 395 4 bl_0_37
port 409 se
rlabel metal1 s 23526 0 23562 395 4 br_0_37
port 411 se
rlabel metal1 s 23382 0 23418 395 4 bl_1_37
port 410 se
rlabel metal1 s 23310 0 23346 395 4 br_1_37
port 412 se
rlabel metal1 s 23790 0 23826 395 4 bl_0_38
port 413 se
rlabel metal1 s 23862 0 23898 395 4 br_0_38
port 415 se
rlabel metal1 s 24006 0 24042 395 4 bl_1_38
port 414 se
rlabel metal1 s 24078 0 24114 395 4 br_1_38
port 416 se
rlabel metal1 s 24846 0 24882 395 4 bl_0_39
port 417 se
rlabel metal1 s 24774 0 24810 395 4 br_0_39
port 419 se
rlabel metal1 s 24630 0 24666 395 4 bl_1_39
port 418 se
rlabel metal1 s 24558 0 24594 395 4 br_1_39
port 420 se
rlabel metal1 s 25038 0 25074 395 4 bl_0_40
port 421 se
rlabel metal1 s 25110 0 25146 395 4 br_0_40
port 423 se
rlabel metal1 s 25254 0 25290 395 4 bl_1_40
port 422 se
rlabel metal1 s 25326 0 25362 395 4 br_1_40
port 424 se
rlabel metal1 s 26094 0 26130 395 4 bl_0_41
port 425 se
rlabel metal1 s 26022 0 26058 395 4 br_0_41
port 427 se
rlabel metal1 s 25878 0 25914 395 4 bl_1_41
port 426 se
rlabel metal1 s 25806 0 25842 395 4 br_1_41
port 428 se
rlabel metal1 s 26286 0 26322 395 4 bl_0_42
port 429 se
rlabel metal1 s 26358 0 26394 395 4 br_0_42
port 431 se
rlabel metal1 s 26502 0 26538 395 4 bl_1_42
port 430 se
rlabel metal1 s 26574 0 26610 395 4 br_1_42
port 432 se
rlabel metal1 s 27342 0 27378 395 4 bl_0_43
port 433 se
rlabel metal1 s 27270 0 27306 395 4 br_0_43
port 435 se
rlabel metal1 s 27126 0 27162 395 4 bl_1_43
port 434 se
rlabel metal1 s 27054 0 27090 395 4 br_1_43
port 436 se
rlabel metal1 s 27534 0 27570 395 4 bl_0_44
port 437 se
rlabel metal1 s 27606 0 27642 395 4 br_0_44
port 439 se
rlabel metal1 s 27750 0 27786 395 4 bl_1_44
port 438 se
rlabel metal1 s 27822 0 27858 395 4 br_1_44
port 440 se
rlabel metal1 s 28590 0 28626 395 4 bl_0_45
port 441 se
rlabel metal1 s 28518 0 28554 395 4 br_0_45
port 443 se
rlabel metal1 s 28374 0 28410 395 4 bl_1_45
port 442 se
rlabel metal1 s 28302 0 28338 395 4 br_1_45
port 444 se
rlabel metal1 s 28782 0 28818 395 4 bl_0_46
port 445 se
rlabel metal1 s 28854 0 28890 395 4 br_0_46
port 447 se
rlabel metal1 s 28998 0 29034 395 4 bl_1_46
port 446 se
rlabel metal1 s 29070 0 29106 395 4 br_1_46
port 448 se
rlabel metal1 s 29838 0 29874 395 4 bl_0_47
port 449 se
rlabel metal1 s 29766 0 29802 395 4 br_0_47
port 451 se
rlabel metal1 s 29622 0 29658 395 4 bl_1_47
port 450 se
rlabel metal1 s 29550 0 29586 395 4 br_1_47
port 452 se
rlabel metal1 s 30030 0 30066 395 4 bl_0_48
port 453 se
rlabel metal1 s 30102 0 30138 395 4 br_0_48
port 455 se
rlabel metal1 s 30246 0 30282 395 4 bl_1_48
port 454 se
rlabel metal1 s 30318 0 30354 395 4 br_1_48
port 456 se
rlabel metal1 s 31086 0 31122 395 4 bl_0_49
port 457 se
rlabel metal1 s 31014 0 31050 395 4 br_0_49
port 459 se
rlabel metal1 s 30870 0 30906 395 4 bl_1_49
port 458 se
rlabel metal1 s 30798 0 30834 395 4 br_1_49
port 460 se
rlabel metal1 s 31278 0 31314 395 4 bl_0_50
port 461 se
rlabel metal1 s 31350 0 31386 395 4 br_0_50
port 463 se
rlabel metal1 s 31494 0 31530 395 4 bl_1_50
port 462 se
rlabel metal1 s 31566 0 31602 395 4 br_1_50
port 464 se
rlabel metal1 s 32334 0 32370 395 4 bl_0_51
port 465 se
rlabel metal1 s 32262 0 32298 395 4 br_0_51
port 467 se
rlabel metal1 s 32118 0 32154 395 4 bl_1_51
port 466 se
rlabel metal1 s 32046 0 32082 395 4 br_1_51
port 468 se
rlabel metal1 s 32526 0 32562 395 4 bl_0_52
port 469 se
rlabel metal1 s 32598 0 32634 395 4 br_0_52
port 471 se
rlabel metal1 s 32742 0 32778 395 4 bl_1_52
port 470 se
rlabel metal1 s 32814 0 32850 395 4 br_1_52
port 472 se
rlabel metal1 s 33582 0 33618 395 4 bl_0_53
port 473 se
rlabel metal1 s 33510 0 33546 395 4 br_0_53
port 475 se
rlabel metal1 s 33366 0 33402 395 4 bl_1_53
port 474 se
rlabel metal1 s 33294 0 33330 395 4 br_1_53
port 476 se
rlabel metal1 s 33774 0 33810 395 4 bl_0_54
port 477 se
rlabel metal1 s 33846 0 33882 395 4 br_0_54
port 479 se
rlabel metal1 s 33990 0 34026 395 4 bl_1_54
port 478 se
rlabel metal1 s 34062 0 34098 395 4 br_1_54
port 480 se
rlabel metal1 s 34830 0 34866 395 4 bl_0_55
port 481 se
rlabel metal1 s 34758 0 34794 395 4 br_0_55
port 483 se
rlabel metal1 s 34614 0 34650 395 4 bl_1_55
port 482 se
rlabel metal1 s 34542 0 34578 395 4 br_1_55
port 484 se
rlabel metal1 s 35022 0 35058 395 4 bl_0_56
port 485 se
rlabel metal1 s 35094 0 35130 395 4 br_0_56
port 487 se
rlabel metal1 s 35238 0 35274 395 4 bl_1_56
port 486 se
rlabel metal1 s 35310 0 35346 395 4 br_1_56
port 488 se
rlabel metal1 s 36078 0 36114 395 4 bl_0_57
port 489 se
rlabel metal1 s 36006 0 36042 395 4 br_0_57
port 491 se
rlabel metal1 s 35862 0 35898 395 4 bl_1_57
port 490 se
rlabel metal1 s 35790 0 35826 395 4 br_1_57
port 492 se
rlabel metal1 s 36270 0 36306 395 4 bl_0_58
port 493 se
rlabel metal1 s 36342 0 36378 395 4 br_0_58
port 495 se
rlabel metal1 s 36486 0 36522 395 4 bl_1_58
port 494 se
rlabel metal1 s 36558 0 36594 395 4 br_1_58
port 496 se
rlabel metal1 s 37326 0 37362 395 4 bl_0_59
port 497 se
rlabel metal1 s 37254 0 37290 395 4 br_0_59
port 499 se
rlabel metal1 s 37110 0 37146 395 4 bl_1_59
port 498 se
rlabel metal1 s 37038 0 37074 395 4 br_1_59
port 500 se
rlabel metal1 s 37518 0 37554 395 4 bl_0_60
port 501 se
rlabel metal1 s 37590 0 37626 395 4 br_0_60
port 503 se
rlabel metal1 s 37734 0 37770 395 4 bl_1_60
port 502 se
rlabel metal1 s 37806 0 37842 395 4 br_1_60
port 504 se
rlabel metal1 s 38574 0 38610 395 4 bl_0_61
port 505 se
rlabel metal1 s 38502 0 38538 395 4 br_0_61
port 507 se
rlabel metal1 s 38358 0 38394 395 4 bl_1_61
port 506 se
rlabel metal1 s 38286 0 38322 395 4 br_1_61
port 508 se
rlabel metal1 s 38766 0 38802 395 4 bl_0_62
port 509 se
rlabel metal1 s 38838 0 38874 395 4 br_0_62
port 511 se
rlabel metal1 s 38982 0 39018 395 4 bl_1_62
port 510 se
rlabel metal1 s 39054 0 39090 395 4 br_1_62
port 512 se
rlabel metal1 s 39822 0 39858 395 4 bl_0_63
port 513 se
rlabel metal1 s 39750 0 39786 395 4 br_0_63
port 515 se
rlabel metal1 s 39606 0 39642 395 4 bl_1_63
port 514 se
rlabel metal1 s 39534 0 39570 395 4 br_1_63
port 516 se
rlabel metal2 s 0 323 39936 371 4 wl_0_0
port 517 se
rlabel metal2 s 0 103 39936 151 4 wl_1_0
port 518 se
rlabel metal1 s 26430 79 26466 420 4 vdd
rlabel metal1 s 12702 79 12738 420 4 vdd
rlabel metal1 s 1470 79 1506 420 4 vdd
rlabel metal1 s 2718 79 2754 420 4 vdd
rlabel metal1 s 22206 79 22242 420 4 vdd
rlabel metal1 s 23934 79 23970 420 4 vdd
rlabel metal1 s 35934 79 35970 420 4 vdd
rlabel metal1 s 37662 79 37698 420 4 vdd
rlabel metal1 s 38430 79 38466 420 4 vdd
rlabel metal1 s 3486 79 3522 420 4 vdd
rlabel metal1 s 22686 79 22722 420 4 vdd
rlabel metal1 s 5982 79 6018 420 4 vdd
rlabel metal1 s 10206 79 10242 420 4 vdd
rlabel metal1 s 13950 79 13986 420 4 vdd
rlabel metal1 s 4734 79 4770 420 4 vdd
rlabel metal1 s 20958 79 20994 420 4 vdd
rlabel metal1 s 30174 79 30210 420 4 vdd
rlabel metal1 s 10974 79 11010 420 4 vdd
rlabel metal1 s 16446 79 16482 420 4 vdd
rlabel metal1 s 17694 79 17730 420 4 vdd
rlabel metal1 s 6462 79 6498 420 4 vdd
rlabel metal1 s 29694 79 29730 420 4 vdd
rlabel metal1 s 21438 79 21474 420 4 vdd
rlabel metal1 s 27198 79 27234 420 4 vdd
rlabel metal1 s 7710 79 7746 420 4 vdd
rlabel metal1 s 38910 79 38946 420 4 vdd
rlabel metal1 s 24702 79 24738 420 4 vdd
rlabel metal1 s 39678 79 39714 420 4 vdd
rlabel metal1 s 14718 79 14754 420 4 vdd
rlabel metal1 s 12222 79 12258 420 4 vdd
rlabel metal1 s 8958 79 8994 420 4 vdd
rlabel metal1 s 8478 79 8514 420 4 vdd
rlabel metal1 s 18462 79 18498 420 4 vdd
rlabel metal1 s 37182 79 37218 420 4 vdd
rlabel metal1 s 15198 79 15234 420 4 vdd
rlabel metal1 s 36414 79 36450 420 4 vdd
rlabel metal1 s 19710 79 19746 420 4 vdd
rlabel metal1 s 33438 79 33474 420 4 vdd
rlabel metal1 s 17214 79 17250 420 4 vdd
rlabel metal1 s 30942 79 30978 420 4 vdd
rlabel metal1 s 28446 79 28482 420 4 vdd
rlabel metal1 s 13470 79 13506 420 4 vdd
rlabel metal1 s 27678 79 27714 420 4 vdd
rlabel metal1 s 32190 79 32226 420 4 vdd
rlabel metal1 s 34686 79 34722 420 4 vdd
rlabel metal1 s 25950 79 25986 420 4 vdd
rlabel metal1 s 5214 79 5250 420 4 vdd
rlabel metal1 s 32670 79 32706 420 4 vdd
rlabel metal1 s 2238 79 2274 420 4 vdd
rlabel metal1 s 20190 79 20226 420 4 vdd
rlabel metal1 s 3966 79 4002 420 4 vdd
rlabel metal1 s 990 79 1026 420 4 vdd
rlabel metal1 s 31422 79 31458 420 4 vdd
rlabel metal1 s 33918 79 33954 420 4 vdd
rlabel metal1 s 11454 79 11490 420 4 vdd
rlabel metal1 s 18942 79 18978 420 4 vdd
rlabel metal1 s 25182 79 25218 420 4 vdd
rlabel metal1 s 9726 79 9762 420 4 vdd
rlabel metal1 s 15966 79 16002 420 4 vdd
rlabel metal1 s 7230 79 7266 420 4 vdd
rlabel metal1 s 28926 79 28962 420 4 vdd
rlabel metal1 s 23454 79 23490 420 4 vdd
rlabel metal1 s 35166 79 35202 420 4 vdd
rlabel metal1 s 222 79 258 420 4 vdd
port 1 se
rlabel metal2 s 954 -55 1062 55 4 gnd
rlabel metal2 s 1434 199 1542 275 4 gnd
rlabel metal2 s 7194 199 7302 275 4 gnd
rlabel metal2 s 22650 199 22758 275 4 gnd
rlabel metal2 s 6426 199 6534 275 4 gnd
rlabel metal2 s 9690 199 9798 275 4 gnd
rlabel metal2 s 37626 -55 37734 55 4 gnd
rlabel metal2 s 33882 -55 33990 55 4 gnd
rlabel metal2 s 10938 -55 11046 55 4 gnd
rlabel metal2 s 15162 199 15270 275 4 gnd
rlabel metal2 s 4698 199 4806 275 4 gnd
rlabel metal2 s 31386 -55 31494 55 4 gnd
rlabel metal2 s 10170 199 10278 275 4 gnd
rlabel metal2 s 20154 -55 20262 55 4 gnd
rlabel metal2 s 22170 -55 22278 55 4 gnd
rlabel metal2 s 25914 199 26022 275 4 gnd
rlabel metal2 s 5946 -55 6054 55 4 gnd
rlabel metal2 s 30906 199 31014 275 4 gnd
rlabel metal2 s 2202 -55 2310 55 4 gnd
rlabel metal2 s 26394 199 26502 275 4 gnd
rlabel metal2 s 28890 199 28998 275 4 gnd
rlabel metal2 s 8442 199 8550 275 4 gnd
rlabel metal2 s 4698 -55 4806 55 4 gnd
rlabel metal2 s 12186 -55 12294 55 4 gnd
rlabel metal2 s 20922 -55 21030 55 4 gnd
rlabel metal2 s 20922 199 21030 275 4 gnd
rlabel metal2 s 27642 199 27750 275 4 gnd
rlabel metal2 s 23418 199 23526 275 4 gnd
rlabel metal2 s 7194 -55 7302 55 4 gnd
rlabel metal2 s 28410 199 28518 275 4 gnd
rlabel metal2 s 15930 -55 16038 55 4 gnd
rlabel metal2 s 36378 199 36486 275 4 gnd
rlabel metal2 s 39642 199 39750 275 4 gnd
rlabel metal2 s 10938 199 11046 275 4 gnd
rlabel metal2 s 25146 199 25254 275 4 gnd
rlabel metal2 s 35898 199 36006 275 4 gnd
rlabel metal2 s 12186 199 12294 275 4 gnd
rlabel metal2 s 23898 -55 24006 55 4 gnd
rlabel metal2 s 8922 -55 9030 55 4 gnd
rlabel metal2 s 15930 199 16038 275 4 gnd
rlabel metal2 s 32154 -55 32262 55 4 gnd
rlabel metal2 s 33882 199 33990 275 4 gnd
rlabel metal2 s 6426 -55 6534 55 4 gnd
rlabel metal2 s 2682 199 2790 275 4 gnd
rlabel metal2 s 33402 -55 33510 55 4 gnd
rlabel metal2 s 11418 199 11526 275 4 gnd
rlabel metal2 s 32154 199 32262 275 4 gnd
rlabel metal2 s 38394 -55 38502 55 4 gnd
rlabel metal2 s 5178 -55 5286 55 4 gnd
rlabel metal2 s 8922 199 9030 275 4 gnd
rlabel metal2 s 186 -55 294 55 4 gnd
rlabel metal2 s 17658 -55 17766 55 4 gnd
rlabel metal2 s 38394 199 38502 275 4 gnd
rlabel metal2 s 38874 199 38982 275 4 gnd
rlabel metal2 s 15162 -55 15270 55 4 gnd
rlabel metal2 s 39642 -55 39750 55 4 gnd
rlabel metal2 s 25146 -55 25254 55 4 gnd
rlabel metal2 s 13914 199 14022 275 4 gnd
rlabel metal2 s 31386 199 31494 275 4 gnd
rlabel metal2 s 21402 199 21510 275 4 gnd
rlabel metal2 s 186 199 294 275 4 gnd
rlabel metal2 s 29658 199 29766 275 4 gnd
rlabel metal2 s 37146 -55 37254 55 4 gnd
rlabel metal2 s 2682 -55 2790 55 4 gnd
rlabel metal2 s 25914 -55 26022 55 4 gnd
rlabel metal2 s 36378 -55 36486 55 4 gnd
rlabel metal2 s 8442 -55 8550 55 4 gnd
rlabel metal2 s 35130 199 35238 275 4 gnd
rlabel metal2 s 32634 199 32742 275 4 gnd
rlabel metal2 s 2202 199 2310 275 4 gnd
rlabel metal2 s 37626 199 37734 275 4 gnd
rlabel metal2 s 5178 199 5286 275 4 gnd
rlabel metal2 s 35130 -55 35238 55 4 gnd
rlabel metal2 s 3450 -55 3558 55 4 gnd
rlabel metal2 s 32634 -55 32742 55 4 gnd
rlabel metal2 s 12666 -55 12774 55 4 gnd
rlabel metal2 s 18906 199 19014 275 4 gnd
rlabel metal2 s 18426 -55 18534 55 4 gnd
rlabel metal2 s 19674 199 19782 275 4 gnd
rlabel metal2 s 30138 -55 30246 55 4 gnd
rlabel metal2 s 9690 -55 9798 55 4 gnd
rlabel metal2 s 17178 -55 17286 55 4 gnd
rlabel metal2 s 24666 -55 24774 55 4 gnd
rlabel metal2 s 23418 -55 23526 55 4 gnd
rlabel metal2 s 14682 -55 14790 55 4 gnd
rlabel metal2 s 7674 199 7782 275 4 gnd
rlabel metal2 s 10170 -55 10278 55 4 gnd
rlabel metal2 s 13914 -55 14022 55 4 gnd
rlabel metal2 s 5946 199 6054 275 4 gnd
rlabel metal2 s 27642 -55 27750 55 4 gnd
rlabel metal2 s 27162 199 27270 275 4 gnd
rlabel metal2 s 22170 199 22278 275 4 gnd
rlabel metal2 s 3930 199 4038 275 4 gnd
rlabel metal2 s 19674 -55 19782 55 4 gnd
rlabel metal2 s 17658 199 17766 275 4 gnd
rlabel metal2 s 7674 -55 7782 55 4 gnd
rlabel metal2 s 12666 199 12774 275 4 gnd
rlabel metal2 s 33402 199 33510 275 4 gnd
rlabel metal2 s 16410 199 16518 275 4 gnd
rlabel metal2 s 13434 199 13542 275 4 gnd
rlabel metal2 s 29658 -55 29766 55 4 gnd
rlabel metal2 s 11418 -55 11526 55 4 gnd
rlabel metal2 s 35898 -55 36006 55 4 gnd
rlabel metal2 s 23898 199 24006 275 4 gnd
rlabel metal2 s 17178 199 17286 275 4 gnd
rlabel metal2 s 18426 199 18534 275 4 gnd
rlabel metal2 s 22650 -55 22758 55 4 gnd
rlabel metal2 s 30138 199 30246 275 4 gnd
rlabel metal2 s 3450 199 3558 275 4 gnd
rlabel metal2 s 16410 -55 16518 55 4 gnd
rlabel metal2 s 30906 -55 31014 55 4 gnd
rlabel metal2 s 1434 -55 1542 55 4 gnd
rlabel metal2 s 26394 -55 26502 55 4 gnd
rlabel metal2 s 18906 -55 19014 55 4 gnd
rlabel metal2 s 13434 -55 13542 55 4 gnd
rlabel metal2 s 28410 -55 28518 55 4 gnd
rlabel metal2 s 27162 -55 27270 55 4 gnd
rlabel metal2 s 28890 -55 28998 55 4 gnd
rlabel metal2 s 34650 199 34758 275 4 gnd
rlabel metal2 s 3930 -55 4038 55 4 gnd
rlabel metal2 s 21402 -55 21510 55 4 gnd
rlabel metal2 s 34650 -55 34758 55 4 gnd
rlabel metal2 s 38874 -55 38982 55 4 gnd
rlabel metal2 s 14682 199 14790 275 4 gnd
rlabel metal2 s 954 199 1062 275 4 gnd
rlabel metal2 s 20154 199 20262 275 4 gnd
rlabel metal2 s 37146 199 37254 275 4 gnd
rlabel metal2 s 24666 199 24774 275 4 gnd
port 2 se
<< properties >>
string FIXED_BBOX 0 0 39936 395
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 7140940
string GDS_START 7056696
<< end >>
