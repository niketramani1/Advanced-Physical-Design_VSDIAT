magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1288 -1260 2176 1357
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_0
timestamp 1624855509
transform 1 0 180 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_1
timestamp 1624855509
transform 1 0 416 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_2
timestamp 1624855509
transform 1 0 652 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180815  sky130_fd_pr__dfl1sd__example_5595914180815_0
timestamp 1624855509
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180815  sky130_fd_pr__dfl1sd__example_5595914180815_1
timestamp 1624855509
transform 1 0 888 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 916 97 916 97 0 FreeSans 300 0 0 0 D
flabel comment s 680 97 680 97 0 FreeSans 300 0 0 0 S
flabel comment s 444 97 444 97 0 FreeSans 300 0 0 0 D
flabel comment s 208 97 208 97 0 FreeSans 300 0 0 0 S
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 1653326
string GDS_START 1650798
<< end >>
