magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1310 -1503 1211 1274
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1624855509
transform 1 0 -50 0 1 13
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1624855509
transform 1 0 -50 0 1 -243
box 0 0 1 1
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 3504064
string GDS_START 3503280
<< end >>
