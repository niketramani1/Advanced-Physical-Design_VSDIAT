magic
tech sky130A
magscale 1 2
timestamp 1624855514
<< obsm3 >>
rect 100 7918 14940 8846
<< metal4 >>
rect 0 10225 15000 10821
rect 0 9273 15000 9869
rect 106 8780 170 8844
rect 187 8780 251 8844
rect 268 8780 332 8844
rect 349 8780 413 8844
rect 430 8780 494 8844
rect 510 8780 574 8844
rect 590 8780 654 8844
rect 670 8780 734 8844
rect 750 8780 814 8844
rect 830 8780 894 8844
rect 910 8780 974 8844
rect 990 8780 1054 8844
rect 1070 8780 1134 8844
rect 1150 8780 1214 8844
rect 1230 8780 1294 8844
rect 1310 8780 1374 8844
rect 1390 8780 1454 8844
rect 1470 8780 1534 8844
rect 1550 8780 1614 8844
rect 1630 8780 1694 8844
rect 1710 8780 1774 8844
rect 1790 8780 1854 8844
rect 1870 8780 1934 8844
rect 1950 8780 2014 8844
rect 2030 8780 2094 8844
rect 2110 8780 2174 8844
rect 2190 8780 2254 8844
rect 2270 8780 2334 8844
rect 2350 8780 2414 8844
rect 2430 8780 2494 8844
rect 2510 8780 2574 8844
rect 2590 8780 2654 8844
rect 2670 8780 2734 8844
rect 2750 8780 2814 8844
rect 2830 8780 2894 8844
rect 2910 8780 2974 8844
rect 2990 8780 3054 8844
rect 3070 8780 3134 8844
rect 3150 8780 3214 8844
rect 3230 8780 3294 8844
rect 3310 8780 3374 8844
rect 3390 8780 3454 8844
rect 3470 8780 3534 8844
rect 3550 8780 3614 8844
rect 3630 8780 3694 8844
rect 3710 8780 3774 8844
rect 3790 8780 3854 8844
rect 3870 8780 3934 8844
rect 3950 8780 4014 8844
rect 4030 8780 4094 8844
rect 4110 8780 4174 8844
rect 4190 8780 4254 8844
rect 4270 8780 4334 8844
rect 4350 8780 4414 8844
rect 4430 8780 4494 8844
rect 4510 8780 4574 8844
rect 4590 8780 4654 8844
rect 4670 8780 4734 8844
rect 4750 8780 4814 8844
rect 4830 8780 4894 8844
rect 10157 8780 10221 8844
rect 10239 8780 10303 8844
rect 10321 8780 10385 8844
rect 10403 8780 10467 8844
rect 10485 8780 10549 8844
rect 10567 8780 10631 8844
rect 10649 8780 10713 8844
rect 10731 8780 10795 8844
rect 10813 8780 10877 8844
rect 10895 8780 10959 8844
rect 10977 8780 11041 8844
rect 11059 8780 11123 8844
rect 11141 8780 11205 8844
rect 11223 8780 11287 8844
rect 11305 8780 11369 8844
rect 11387 8780 11451 8844
rect 11468 8780 11532 8844
rect 11549 8780 11613 8844
rect 11630 8780 11694 8844
rect 11711 8780 11775 8844
rect 11792 8780 11856 8844
rect 11873 8780 11937 8844
rect 11954 8780 12018 8844
rect 12035 8780 12099 8844
rect 12116 8780 12180 8844
rect 12197 8780 12261 8844
rect 12278 8780 12342 8844
rect 12359 8780 12423 8844
rect 12440 8780 12504 8844
rect 12521 8780 12585 8844
rect 12602 8780 12666 8844
rect 12683 8780 12747 8844
rect 12764 8780 12828 8844
rect 12845 8780 12909 8844
rect 12926 8780 12990 8844
rect 13007 8780 13071 8844
rect 13088 8780 13152 8844
rect 13169 8780 13233 8844
rect 13250 8780 13314 8844
rect 13331 8780 13395 8844
rect 13412 8780 13476 8844
rect 13493 8780 13557 8844
rect 13574 8780 13638 8844
rect 13655 8780 13719 8844
rect 13736 8780 13800 8844
rect 13817 8780 13881 8844
rect 13898 8780 13962 8844
rect 13979 8780 14043 8844
rect 14060 8780 14124 8844
rect 14141 8780 14205 8844
rect 14222 8780 14286 8844
rect 14303 8780 14367 8844
rect 14384 8780 14448 8844
rect 14465 8780 14529 8844
rect 14546 8780 14610 8844
rect 14627 8780 14691 8844
rect 14708 8780 14772 8844
rect 14789 8780 14853 8844
rect 14870 8780 14934 8844
rect 106 8694 170 8758
rect 187 8694 251 8758
rect 268 8694 332 8758
rect 349 8694 413 8758
rect 430 8694 494 8758
rect 510 8694 574 8758
rect 590 8694 654 8758
rect 670 8694 734 8758
rect 750 8694 814 8758
rect 830 8694 894 8758
rect 910 8694 974 8758
rect 990 8694 1054 8758
rect 1070 8694 1134 8758
rect 1150 8694 1214 8758
rect 1230 8694 1294 8758
rect 1310 8694 1374 8758
rect 1390 8694 1454 8758
rect 1470 8694 1534 8758
rect 1550 8694 1614 8758
rect 1630 8694 1694 8758
rect 1710 8694 1774 8758
rect 1790 8694 1854 8758
rect 1870 8694 1934 8758
rect 1950 8694 2014 8758
rect 2030 8694 2094 8758
rect 2110 8694 2174 8758
rect 2190 8694 2254 8758
rect 2270 8694 2334 8758
rect 2350 8694 2414 8758
rect 2430 8694 2494 8758
rect 2510 8694 2574 8758
rect 2590 8694 2654 8758
rect 2670 8694 2734 8758
rect 2750 8694 2814 8758
rect 2830 8694 2894 8758
rect 2910 8694 2974 8758
rect 2990 8694 3054 8758
rect 3070 8694 3134 8758
rect 3150 8694 3214 8758
rect 3230 8694 3294 8758
rect 3310 8694 3374 8758
rect 3390 8694 3454 8758
rect 3470 8694 3534 8758
rect 3550 8694 3614 8758
rect 3630 8694 3694 8758
rect 3710 8694 3774 8758
rect 3790 8694 3854 8758
rect 3870 8694 3934 8758
rect 3950 8694 4014 8758
rect 4030 8694 4094 8758
rect 4110 8694 4174 8758
rect 4190 8694 4254 8758
rect 4270 8694 4334 8758
rect 4350 8694 4414 8758
rect 4430 8694 4494 8758
rect 4510 8694 4574 8758
rect 4590 8694 4654 8758
rect 4670 8694 4734 8758
rect 4750 8694 4814 8758
rect 4830 8694 4894 8758
rect 10157 8694 10221 8758
rect 10239 8694 10303 8758
rect 10321 8694 10385 8758
rect 10403 8694 10467 8758
rect 10485 8694 10549 8758
rect 10567 8694 10631 8758
rect 10649 8694 10713 8758
rect 10731 8694 10795 8758
rect 10813 8694 10877 8758
rect 10895 8694 10959 8758
rect 10977 8694 11041 8758
rect 11059 8694 11123 8758
rect 11141 8694 11205 8758
rect 11223 8694 11287 8758
rect 11305 8694 11369 8758
rect 11387 8694 11451 8758
rect 11468 8694 11532 8758
rect 11549 8694 11613 8758
rect 11630 8694 11694 8758
rect 11711 8694 11775 8758
rect 11792 8694 11856 8758
rect 11873 8694 11937 8758
rect 11954 8694 12018 8758
rect 12035 8694 12099 8758
rect 12116 8694 12180 8758
rect 12197 8694 12261 8758
rect 12278 8694 12342 8758
rect 12359 8694 12423 8758
rect 12440 8694 12504 8758
rect 12521 8694 12585 8758
rect 12602 8694 12666 8758
rect 12683 8694 12747 8758
rect 12764 8694 12828 8758
rect 12845 8694 12909 8758
rect 12926 8694 12990 8758
rect 13007 8694 13071 8758
rect 13088 8694 13152 8758
rect 13169 8694 13233 8758
rect 13250 8694 13314 8758
rect 13331 8694 13395 8758
rect 13412 8694 13476 8758
rect 13493 8694 13557 8758
rect 13574 8694 13638 8758
rect 13655 8694 13719 8758
rect 13736 8694 13800 8758
rect 13817 8694 13881 8758
rect 13898 8694 13962 8758
rect 13979 8694 14043 8758
rect 14060 8694 14124 8758
rect 14141 8694 14205 8758
rect 14222 8694 14286 8758
rect 14303 8694 14367 8758
rect 14384 8694 14448 8758
rect 14465 8694 14529 8758
rect 14546 8694 14610 8758
rect 14627 8694 14691 8758
rect 14708 8694 14772 8758
rect 14789 8694 14853 8758
rect 14870 8694 14934 8758
rect 106 8608 170 8672
rect 187 8608 251 8672
rect 268 8608 332 8672
rect 349 8608 413 8672
rect 430 8608 494 8672
rect 510 8608 574 8672
rect 590 8608 654 8672
rect 670 8608 734 8672
rect 750 8608 814 8672
rect 830 8608 894 8672
rect 910 8608 974 8672
rect 990 8608 1054 8672
rect 1070 8608 1134 8672
rect 1150 8608 1214 8672
rect 1230 8608 1294 8672
rect 1310 8608 1374 8672
rect 1390 8608 1454 8672
rect 1470 8608 1534 8672
rect 1550 8608 1614 8672
rect 1630 8608 1694 8672
rect 1710 8608 1774 8672
rect 1790 8608 1854 8672
rect 1870 8608 1934 8672
rect 1950 8608 2014 8672
rect 2030 8608 2094 8672
rect 2110 8608 2174 8672
rect 2190 8608 2254 8672
rect 2270 8608 2334 8672
rect 2350 8608 2414 8672
rect 2430 8608 2494 8672
rect 2510 8608 2574 8672
rect 2590 8608 2654 8672
rect 2670 8608 2734 8672
rect 2750 8608 2814 8672
rect 2830 8608 2894 8672
rect 2910 8608 2974 8672
rect 2990 8608 3054 8672
rect 3070 8608 3134 8672
rect 3150 8608 3214 8672
rect 3230 8608 3294 8672
rect 3310 8608 3374 8672
rect 3390 8608 3454 8672
rect 3470 8608 3534 8672
rect 3550 8608 3614 8672
rect 3630 8608 3694 8672
rect 3710 8608 3774 8672
rect 3790 8608 3854 8672
rect 3870 8608 3934 8672
rect 3950 8608 4014 8672
rect 4030 8608 4094 8672
rect 4110 8608 4174 8672
rect 4190 8608 4254 8672
rect 4270 8608 4334 8672
rect 4350 8608 4414 8672
rect 4430 8608 4494 8672
rect 4510 8608 4574 8672
rect 4590 8608 4654 8672
rect 4670 8608 4734 8672
rect 4750 8608 4814 8672
rect 4830 8608 4894 8672
rect 10157 8608 10221 8672
rect 10239 8608 10303 8672
rect 10321 8608 10385 8672
rect 10403 8608 10467 8672
rect 10485 8608 10549 8672
rect 10567 8608 10631 8672
rect 10649 8608 10713 8672
rect 10731 8608 10795 8672
rect 10813 8608 10877 8672
rect 10895 8608 10959 8672
rect 10977 8608 11041 8672
rect 11059 8608 11123 8672
rect 11141 8608 11205 8672
rect 11223 8608 11287 8672
rect 11305 8608 11369 8672
rect 11387 8608 11451 8672
rect 11468 8608 11532 8672
rect 11549 8608 11613 8672
rect 11630 8608 11694 8672
rect 11711 8608 11775 8672
rect 11792 8608 11856 8672
rect 11873 8608 11937 8672
rect 11954 8608 12018 8672
rect 12035 8608 12099 8672
rect 12116 8608 12180 8672
rect 12197 8608 12261 8672
rect 12278 8608 12342 8672
rect 12359 8608 12423 8672
rect 12440 8608 12504 8672
rect 12521 8608 12585 8672
rect 12602 8608 12666 8672
rect 12683 8608 12747 8672
rect 12764 8608 12828 8672
rect 12845 8608 12909 8672
rect 12926 8608 12990 8672
rect 13007 8608 13071 8672
rect 13088 8608 13152 8672
rect 13169 8608 13233 8672
rect 13250 8608 13314 8672
rect 13331 8608 13395 8672
rect 13412 8608 13476 8672
rect 13493 8608 13557 8672
rect 13574 8608 13638 8672
rect 13655 8608 13719 8672
rect 13736 8608 13800 8672
rect 13817 8608 13881 8672
rect 13898 8608 13962 8672
rect 13979 8608 14043 8672
rect 14060 8608 14124 8672
rect 14141 8608 14205 8672
rect 14222 8608 14286 8672
rect 14303 8608 14367 8672
rect 14384 8608 14448 8672
rect 14465 8608 14529 8672
rect 14546 8608 14610 8672
rect 14627 8608 14691 8672
rect 14708 8608 14772 8672
rect 14789 8608 14853 8672
rect 14870 8608 14934 8672
rect 106 8522 170 8586
rect 187 8522 251 8586
rect 268 8522 332 8586
rect 349 8522 413 8586
rect 430 8522 494 8586
rect 510 8522 574 8586
rect 590 8522 654 8586
rect 670 8522 734 8586
rect 750 8522 814 8586
rect 830 8522 894 8586
rect 910 8522 974 8586
rect 990 8522 1054 8586
rect 1070 8522 1134 8586
rect 1150 8522 1214 8586
rect 1230 8522 1294 8586
rect 1310 8522 1374 8586
rect 1390 8522 1454 8586
rect 1470 8522 1534 8586
rect 1550 8522 1614 8586
rect 1630 8522 1694 8586
rect 1710 8522 1774 8586
rect 1790 8522 1854 8586
rect 1870 8522 1934 8586
rect 1950 8522 2014 8586
rect 2030 8522 2094 8586
rect 2110 8522 2174 8586
rect 2190 8522 2254 8586
rect 2270 8522 2334 8586
rect 2350 8522 2414 8586
rect 2430 8522 2494 8586
rect 2510 8522 2574 8586
rect 2590 8522 2654 8586
rect 2670 8522 2734 8586
rect 2750 8522 2814 8586
rect 2830 8522 2894 8586
rect 2910 8522 2974 8586
rect 2990 8522 3054 8586
rect 3070 8522 3134 8586
rect 3150 8522 3214 8586
rect 3230 8522 3294 8586
rect 3310 8522 3374 8586
rect 3390 8522 3454 8586
rect 3470 8522 3534 8586
rect 3550 8522 3614 8586
rect 3630 8522 3694 8586
rect 3710 8522 3774 8586
rect 3790 8522 3854 8586
rect 3870 8522 3934 8586
rect 3950 8522 4014 8586
rect 4030 8522 4094 8586
rect 4110 8522 4174 8586
rect 4190 8522 4254 8586
rect 4270 8522 4334 8586
rect 4350 8522 4414 8586
rect 4430 8522 4494 8586
rect 4510 8522 4574 8586
rect 4590 8522 4654 8586
rect 4670 8522 4734 8586
rect 4750 8522 4814 8586
rect 4830 8522 4894 8586
rect 10157 8522 10221 8586
rect 10239 8522 10303 8586
rect 10321 8522 10385 8586
rect 10403 8522 10467 8586
rect 10485 8522 10549 8586
rect 10567 8522 10631 8586
rect 10649 8522 10713 8586
rect 10731 8522 10795 8586
rect 10813 8522 10877 8586
rect 10895 8522 10959 8586
rect 10977 8522 11041 8586
rect 11059 8522 11123 8586
rect 11141 8522 11205 8586
rect 11223 8522 11287 8586
rect 11305 8522 11369 8586
rect 11387 8522 11451 8586
rect 11468 8522 11532 8586
rect 11549 8522 11613 8586
rect 11630 8522 11694 8586
rect 11711 8522 11775 8586
rect 11792 8522 11856 8586
rect 11873 8522 11937 8586
rect 11954 8522 12018 8586
rect 12035 8522 12099 8586
rect 12116 8522 12180 8586
rect 12197 8522 12261 8586
rect 12278 8522 12342 8586
rect 12359 8522 12423 8586
rect 12440 8522 12504 8586
rect 12521 8522 12585 8586
rect 12602 8522 12666 8586
rect 12683 8522 12747 8586
rect 12764 8522 12828 8586
rect 12845 8522 12909 8586
rect 12926 8522 12990 8586
rect 13007 8522 13071 8586
rect 13088 8522 13152 8586
rect 13169 8522 13233 8586
rect 13250 8522 13314 8586
rect 13331 8522 13395 8586
rect 13412 8522 13476 8586
rect 13493 8522 13557 8586
rect 13574 8522 13638 8586
rect 13655 8522 13719 8586
rect 13736 8522 13800 8586
rect 13817 8522 13881 8586
rect 13898 8522 13962 8586
rect 13979 8522 14043 8586
rect 14060 8522 14124 8586
rect 14141 8522 14205 8586
rect 14222 8522 14286 8586
rect 14303 8522 14367 8586
rect 14384 8522 14448 8586
rect 14465 8522 14529 8586
rect 14546 8522 14610 8586
rect 14627 8522 14691 8586
rect 14708 8522 14772 8586
rect 14789 8522 14853 8586
rect 14870 8522 14934 8586
rect 106 8436 170 8500
rect 187 8436 251 8500
rect 268 8436 332 8500
rect 349 8436 413 8500
rect 430 8436 494 8500
rect 510 8436 574 8500
rect 590 8436 654 8500
rect 670 8436 734 8500
rect 750 8436 814 8500
rect 830 8436 894 8500
rect 910 8436 974 8500
rect 990 8436 1054 8500
rect 1070 8436 1134 8500
rect 1150 8436 1214 8500
rect 1230 8436 1294 8500
rect 1310 8436 1374 8500
rect 1390 8436 1454 8500
rect 1470 8436 1534 8500
rect 1550 8436 1614 8500
rect 1630 8436 1694 8500
rect 1710 8436 1774 8500
rect 1790 8436 1854 8500
rect 1870 8436 1934 8500
rect 1950 8436 2014 8500
rect 2030 8436 2094 8500
rect 2110 8436 2174 8500
rect 2190 8436 2254 8500
rect 2270 8436 2334 8500
rect 2350 8436 2414 8500
rect 2430 8436 2494 8500
rect 2510 8436 2574 8500
rect 2590 8436 2654 8500
rect 2670 8436 2734 8500
rect 2750 8436 2814 8500
rect 2830 8436 2894 8500
rect 2910 8436 2974 8500
rect 2990 8436 3054 8500
rect 3070 8436 3134 8500
rect 3150 8436 3214 8500
rect 3230 8436 3294 8500
rect 3310 8436 3374 8500
rect 3390 8436 3454 8500
rect 3470 8436 3534 8500
rect 3550 8436 3614 8500
rect 3630 8436 3694 8500
rect 3710 8436 3774 8500
rect 3790 8436 3854 8500
rect 3870 8436 3934 8500
rect 3950 8436 4014 8500
rect 4030 8436 4094 8500
rect 4110 8436 4174 8500
rect 4190 8436 4254 8500
rect 4270 8436 4334 8500
rect 4350 8436 4414 8500
rect 4430 8436 4494 8500
rect 4510 8436 4574 8500
rect 4590 8436 4654 8500
rect 4670 8436 4734 8500
rect 4750 8436 4814 8500
rect 4830 8436 4894 8500
rect 10157 8436 10221 8500
rect 10239 8436 10303 8500
rect 10321 8436 10385 8500
rect 10403 8436 10467 8500
rect 10485 8436 10549 8500
rect 10567 8436 10631 8500
rect 10649 8436 10713 8500
rect 10731 8436 10795 8500
rect 10813 8436 10877 8500
rect 10895 8436 10959 8500
rect 10977 8436 11041 8500
rect 11059 8436 11123 8500
rect 11141 8436 11205 8500
rect 11223 8436 11287 8500
rect 11305 8436 11369 8500
rect 11387 8436 11451 8500
rect 11468 8436 11532 8500
rect 11549 8436 11613 8500
rect 11630 8436 11694 8500
rect 11711 8436 11775 8500
rect 11792 8436 11856 8500
rect 11873 8436 11937 8500
rect 11954 8436 12018 8500
rect 12035 8436 12099 8500
rect 12116 8436 12180 8500
rect 12197 8436 12261 8500
rect 12278 8436 12342 8500
rect 12359 8436 12423 8500
rect 12440 8436 12504 8500
rect 12521 8436 12585 8500
rect 12602 8436 12666 8500
rect 12683 8436 12747 8500
rect 12764 8436 12828 8500
rect 12845 8436 12909 8500
rect 12926 8436 12990 8500
rect 13007 8436 13071 8500
rect 13088 8436 13152 8500
rect 13169 8436 13233 8500
rect 13250 8436 13314 8500
rect 13331 8436 13395 8500
rect 13412 8436 13476 8500
rect 13493 8436 13557 8500
rect 13574 8436 13638 8500
rect 13655 8436 13719 8500
rect 13736 8436 13800 8500
rect 13817 8436 13881 8500
rect 13898 8436 13962 8500
rect 13979 8436 14043 8500
rect 14060 8436 14124 8500
rect 14141 8436 14205 8500
rect 14222 8436 14286 8500
rect 14303 8436 14367 8500
rect 14384 8436 14448 8500
rect 14465 8436 14529 8500
rect 14546 8436 14610 8500
rect 14627 8436 14691 8500
rect 14708 8436 14772 8500
rect 14789 8436 14853 8500
rect 14870 8436 14934 8500
rect 106 8350 170 8414
rect 187 8350 251 8414
rect 268 8350 332 8414
rect 349 8350 413 8414
rect 430 8350 494 8414
rect 510 8350 574 8414
rect 590 8350 654 8414
rect 670 8350 734 8414
rect 750 8350 814 8414
rect 830 8350 894 8414
rect 910 8350 974 8414
rect 990 8350 1054 8414
rect 1070 8350 1134 8414
rect 1150 8350 1214 8414
rect 1230 8350 1294 8414
rect 1310 8350 1374 8414
rect 1390 8350 1454 8414
rect 1470 8350 1534 8414
rect 1550 8350 1614 8414
rect 1630 8350 1694 8414
rect 1710 8350 1774 8414
rect 1790 8350 1854 8414
rect 1870 8350 1934 8414
rect 1950 8350 2014 8414
rect 2030 8350 2094 8414
rect 2110 8350 2174 8414
rect 2190 8350 2254 8414
rect 2270 8350 2334 8414
rect 2350 8350 2414 8414
rect 2430 8350 2494 8414
rect 2510 8350 2574 8414
rect 2590 8350 2654 8414
rect 2670 8350 2734 8414
rect 2750 8350 2814 8414
rect 2830 8350 2894 8414
rect 2910 8350 2974 8414
rect 2990 8350 3054 8414
rect 3070 8350 3134 8414
rect 3150 8350 3214 8414
rect 3230 8350 3294 8414
rect 3310 8350 3374 8414
rect 3390 8350 3454 8414
rect 3470 8350 3534 8414
rect 3550 8350 3614 8414
rect 3630 8350 3694 8414
rect 3710 8350 3774 8414
rect 3790 8350 3854 8414
rect 3870 8350 3934 8414
rect 3950 8350 4014 8414
rect 4030 8350 4094 8414
rect 4110 8350 4174 8414
rect 4190 8350 4254 8414
rect 4270 8350 4334 8414
rect 4350 8350 4414 8414
rect 4430 8350 4494 8414
rect 4510 8350 4574 8414
rect 4590 8350 4654 8414
rect 4670 8350 4734 8414
rect 4750 8350 4814 8414
rect 4830 8350 4894 8414
rect 10157 8350 10221 8414
rect 10239 8350 10303 8414
rect 10321 8350 10385 8414
rect 10403 8350 10467 8414
rect 10485 8350 10549 8414
rect 10567 8350 10631 8414
rect 10649 8350 10713 8414
rect 10731 8350 10795 8414
rect 10813 8350 10877 8414
rect 10895 8350 10959 8414
rect 10977 8350 11041 8414
rect 11059 8350 11123 8414
rect 11141 8350 11205 8414
rect 11223 8350 11287 8414
rect 11305 8350 11369 8414
rect 11387 8350 11451 8414
rect 11468 8350 11532 8414
rect 11549 8350 11613 8414
rect 11630 8350 11694 8414
rect 11711 8350 11775 8414
rect 11792 8350 11856 8414
rect 11873 8350 11937 8414
rect 11954 8350 12018 8414
rect 12035 8350 12099 8414
rect 12116 8350 12180 8414
rect 12197 8350 12261 8414
rect 12278 8350 12342 8414
rect 12359 8350 12423 8414
rect 12440 8350 12504 8414
rect 12521 8350 12585 8414
rect 12602 8350 12666 8414
rect 12683 8350 12747 8414
rect 12764 8350 12828 8414
rect 12845 8350 12909 8414
rect 12926 8350 12990 8414
rect 13007 8350 13071 8414
rect 13088 8350 13152 8414
rect 13169 8350 13233 8414
rect 13250 8350 13314 8414
rect 13331 8350 13395 8414
rect 13412 8350 13476 8414
rect 13493 8350 13557 8414
rect 13574 8350 13638 8414
rect 13655 8350 13719 8414
rect 13736 8350 13800 8414
rect 13817 8350 13881 8414
rect 13898 8350 13962 8414
rect 13979 8350 14043 8414
rect 14060 8350 14124 8414
rect 14141 8350 14205 8414
rect 14222 8350 14286 8414
rect 14303 8350 14367 8414
rect 14384 8350 14448 8414
rect 14465 8350 14529 8414
rect 14546 8350 14610 8414
rect 14627 8350 14691 8414
rect 14708 8350 14772 8414
rect 14789 8350 14853 8414
rect 14870 8350 14934 8414
rect 106 8264 170 8328
rect 187 8264 251 8328
rect 268 8264 332 8328
rect 349 8264 413 8328
rect 430 8264 494 8328
rect 510 8264 574 8328
rect 590 8264 654 8328
rect 670 8264 734 8328
rect 750 8264 814 8328
rect 830 8264 894 8328
rect 910 8264 974 8328
rect 990 8264 1054 8328
rect 1070 8264 1134 8328
rect 1150 8264 1214 8328
rect 1230 8264 1294 8328
rect 1310 8264 1374 8328
rect 1390 8264 1454 8328
rect 1470 8264 1534 8328
rect 1550 8264 1614 8328
rect 1630 8264 1694 8328
rect 1710 8264 1774 8328
rect 1790 8264 1854 8328
rect 1870 8264 1934 8328
rect 1950 8264 2014 8328
rect 2030 8264 2094 8328
rect 2110 8264 2174 8328
rect 2190 8264 2254 8328
rect 2270 8264 2334 8328
rect 2350 8264 2414 8328
rect 2430 8264 2494 8328
rect 2510 8264 2574 8328
rect 2590 8264 2654 8328
rect 2670 8264 2734 8328
rect 2750 8264 2814 8328
rect 2830 8264 2894 8328
rect 2910 8264 2974 8328
rect 2990 8264 3054 8328
rect 3070 8264 3134 8328
rect 3150 8264 3214 8328
rect 3230 8264 3294 8328
rect 3310 8264 3374 8328
rect 3390 8264 3454 8328
rect 3470 8264 3534 8328
rect 3550 8264 3614 8328
rect 3630 8264 3694 8328
rect 3710 8264 3774 8328
rect 3790 8264 3854 8328
rect 3870 8264 3934 8328
rect 3950 8264 4014 8328
rect 4030 8264 4094 8328
rect 4110 8264 4174 8328
rect 4190 8264 4254 8328
rect 4270 8264 4334 8328
rect 4350 8264 4414 8328
rect 4430 8264 4494 8328
rect 4510 8264 4574 8328
rect 4590 8264 4654 8328
rect 4670 8264 4734 8328
rect 4750 8264 4814 8328
rect 4830 8264 4894 8328
rect 10157 8264 10221 8328
rect 10239 8264 10303 8328
rect 10321 8264 10385 8328
rect 10403 8264 10467 8328
rect 10485 8264 10549 8328
rect 10567 8264 10631 8328
rect 10649 8264 10713 8328
rect 10731 8264 10795 8328
rect 10813 8264 10877 8328
rect 10895 8264 10959 8328
rect 10977 8264 11041 8328
rect 11059 8264 11123 8328
rect 11141 8264 11205 8328
rect 11223 8264 11287 8328
rect 11305 8264 11369 8328
rect 11387 8264 11451 8328
rect 11468 8264 11532 8328
rect 11549 8264 11613 8328
rect 11630 8264 11694 8328
rect 11711 8264 11775 8328
rect 11792 8264 11856 8328
rect 11873 8264 11937 8328
rect 11954 8264 12018 8328
rect 12035 8264 12099 8328
rect 12116 8264 12180 8328
rect 12197 8264 12261 8328
rect 12278 8264 12342 8328
rect 12359 8264 12423 8328
rect 12440 8264 12504 8328
rect 12521 8264 12585 8328
rect 12602 8264 12666 8328
rect 12683 8264 12747 8328
rect 12764 8264 12828 8328
rect 12845 8264 12909 8328
rect 12926 8264 12990 8328
rect 13007 8264 13071 8328
rect 13088 8264 13152 8328
rect 13169 8264 13233 8328
rect 13250 8264 13314 8328
rect 13331 8264 13395 8328
rect 13412 8264 13476 8328
rect 13493 8264 13557 8328
rect 13574 8264 13638 8328
rect 13655 8264 13719 8328
rect 13736 8264 13800 8328
rect 13817 8264 13881 8328
rect 13898 8264 13962 8328
rect 13979 8264 14043 8328
rect 14060 8264 14124 8328
rect 14141 8264 14205 8328
rect 14222 8264 14286 8328
rect 14303 8264 14367 8328
rect 14384 8264 14448 8328
rect 14465 8264 14529 8328
rect 14546 8264 14610 8328
rect 14627 8264 14691 8328
rect 14708 8264 14772 8328
rect 14789 8264 14853 8328
rect 14870 8264 14934 8328
rect 106 8178 170 8242
rect 187 8178 251 8242
rect 268 8178 332 8242
rect 349 8178 413 8242
rect 430 8178 494 8242
rect 510 8178 574 8242
rect 590 8178 654 8242
rect 670 8178 734 8242
rect 750 8178 814 8242
rect 830 8178 894 8242
rect 910 8178 974 8242
rect 990 8178 1054 8242
rect 1070 8178 1134 8242
rect 1150 8178 1214 8242
rect 1230 8178 1294 8242
rect 1310 8178 1374 8242
rect 1390 8178 1454 8242
rect 1470 8178 1534 8242
rect 1550 8178 1614 8242
rect 1630 8178 1694 8242
rect 1710 8178 1774 8242
rect 1790 8178 1854 8242
rect 1870 8178 1934 8242
rect 1950 8178 2014 8242
rect 2030 8178 2094 8242
rect 2110 8178 2174 8242
rect 2190 8178 2254 8242
rect 2270 8178 2334 8242
rect 2350 8178 2414 8242
rect 2430 8178 2494 8242
rect 2510 8178 2574 8242
rect 2590 8178 2654 8242
rect 2670 8178 2734 8242
rect 2750 8178 2814 8242
rect 2830 8178 2894 8242
rect 2910 8178 2974 8242
rect 2990 8178 3054 8242
rect 3070 8178 3134 8242
rect 3150 8178 3214 8242
rect 3230 8178 3294 8242
rect 3310 8178 3374 8242
rect 3390 8178 3454 8242
rect 3470 8178 3534 8242
rect 3550 8178 3614 8242
rect 3630 8178 3694 8242
rect 3710 8178 3774 8242
rect 3790 8178 3854 8242
rect 3870 8178 3934 8242
rect 3950 8178 4014 8242
rect 4030 8178 4094 8242
rect 4110 8178 4174 8242
rect 4190 8178 4254 8242
rect 4270 8178 4334 8242
rect 4350 8178 4414 8242
rect 4430 8178 4494 8242
rect 4510 8178 4574 8242
rect 4590 8178 4654 8242
rect 4670 8178 4734 8242
rect 4750 8178 4814 8242
rect 4830 8178 4894 8242
rect 10157 8178 10221 8242
rect 10239 8178 10303 8242
rect 10321 8178 10385 8242
rect 10403 8178 10467 8242
rect 10485 8178 10549 8242
rect 10567 8178 10631 8242
rect 10649 8178 10713 8242
rect 10731 8178 10795 8242
rect 10813 8178 10877 8242
rect 10895 8178 10959 8242
rect 10977 8178 11041 8242
rect 11059 8178 11123 8242
rect 11141 8178 11205 8242
rect 11223 8178 11287 8242
rect 11305 8178 11369 8242
rect 11387 8178 11451 8242
rect 11468 8178 11532 8242
rect 11549 8178 11613 8242
rect 11630 8178 11694 8242
rect 11711 8178 11775 8242
rect 11792 8178 11856 8242
rect 11873 8178 11937 8242
rect 11954 8178 12018 8242
rect 12035 8178 12099 8242
rect 12116 8178 12180 8242
rect 12197 8178 12261 8242
rect 12278 8178 12342 8242
rect 12359 8178 12423 8242
rect 12440 8178 12504 8242
rect 12521 8178 12585 8242
rect 12602 8178 12666 8242
rect 12683 8178 12747 8242
rect 12764 8178 12828 8242
rect 12845 8178 12909 8242
rect 12926 8178 12990 8242
rect 13007 8178 13071 8242
rect 13088 8178 13152 8242
rect 13169 8178 13233 8242
rect 13250 8178 13314 8242
rect 13331 8178 13395 8242
rect 13412 8178 13476 8242
rect 13493 8178 13557 8242
rect 13574 8178 13638 8242
rect 13655 8178 13719 8242
rect 13736 8178 13800 8242
rect 13817 8178 13881 8242
rect 13898 8178 13962 8242
rect 13979 8178 14043 8242
rect 14060 8178 14124 8242
rect 14141 8178 14205 8242
rect 14222 8178 14286 8242
rect 14303 8178 14367 8242
rect 14384 8178 14448 8242
rect 14465 8178 14529 8242
rect 14546 8178 14610 8242
rect 14627 8178 14691 8242
rect 14708 8178 14772 8242
rect 14789 8178 14853 8242
rect 14870 8178 14934 8242
rect 106 8092 170 8156
rect 187 8092 251 8156
rect 268 8092 332 8156
rect 349 8092 413 8156
rect 430 8092 494 8156
rect 510 8092 574 8156
rect 590 8092 654 8156
rect 670 8092 734 8156
rect 750 8092 814 8156
rect 830 8092 894 8156
rect 910 8092 974 8156
rect 990 8092 1054 8156
rect 1070 8092 1134 8156
rect 1150 8092 1214 8156
rect 1230 8092 1294 8156
rect 1310 8092 1374 8156
rect 1390 8092 1454 8156
rect 1470 8092 1534 8156
rect 1550 8092 1614 8156
rect 1630 8092 1694 8156
rect 1710 8092 1774 8156
rect 1790 8092 1854 8156
rect 1870 8092 1934 8156
rect 1950 8092 2014 8156
rect 2030 8092 2094 8156
rect 2110 8092 2174 8156
rect 2190 8092 2254 8156
rect 2270 8092 2334 8156
rect 2350 8092 2414 8156
rect 2430 8092 2494 8156
rect 2510 8092 2574 8156
rect 2590 8092 2654 8156
rect 2670 8092 2734 8156
rect 2750 8092 2814 8156
rect 2830 8092 2894 8156
rect 2910 8092 2974 8156
rect 2990 8092 3054 8156
rect 3070 8092 3134 8156
rect 3150 8092 3214 8156
rect 3230 8092 3294 8156
rect 3310 8092 3374 8156
rect 3390 8092 3454 8156
rect 3470 8092 3534 8156
rect 3550 8092 3614 8156
rect 3630 8092 3694 8156
rect 3710 8092 3774 8156
rect 3790 8092 3854 8156
rect 3870 8092 3934 8156
rect 3950 8092 4014 8156
rect 4030 8092 4094 8156
rect 4110 8092 4174 8156
rect 4190 8092 4254 8156
rect 4270 8092 4334 8156
rect 4350 8092 4414 8156
rect 4430 8092 4494 8156
rect 4510 8092 4574 8156
rect 4590 8092 4654 8156
rect 4670 8092 4734 8156
rect 4750 8092 4814 8156
rect 4830 8092 4894 8156
rect 10157 8092 10221 8156
rect 10239 8092 10303 8156
rect 10321 8092 10385 8156
rect 10403 8092 10467 8156
rect 10485 8092 10549 8156
rect 10567 8092 10631 8156
rect 10649 8092 10713 8156
rect 10731 8092 10795 8156
rect 10813 8092 10877 8156
rect 10895 8092 10959 8156
rect 10977 8092 11041 8156
rect 11059 8092 11123 8156
rect 11141 8092 11205 8156
rect 11223 8092 11287 8156
rect 11305 8092 11369 8156
rect 11387 8092 11451 8156
rect 11468 8092 11532 8156
rect 11549 8092 11613 8156
rect 11630 8092 11694 8156
rect 11711 8092 11775 8156
rect 11792 8092 11856 8156
rect 11873 8092 11937 8156
rect 11954 8092 12018 8156
rect 12035 8092 12099 8156
rect 12116 8092 12180 8156
rect 12197 8092 12261 8156
rect 12278 8092 12342 8156
rect 12359 8092 12423 8156
rect 12440 8092 12504 8156
rect 12521 8092 12585 8156
rect 12602 8092 12666 8156
rect 12683 8092 12747 8156
rect 12764 8092 12828 8156
rect 12845 8092 12909 8156
rect 12926 8092 12990 8156
rect 13007 8092 13071 8156
rect 13088 8092 13152 8156
rect 13169 8092 13233 8156
rect 13250 8092 13314 8156
rect 13331 8092 13395 8156
rect 13412 8092 13476 8156
rect 13493 8092 13557 8156
rect 13574 8092 13638 8156
rect 13655 8092 13719 8156
rect 13736 8092 13800 8156
rect 13817 8092 13881 8156
rect 13898 8092 13962 8156
rect 13979 8092 14043 8156
rect 14060 8092 14124 8156
rect 14141 8092 14205 8156
rect 14222 8092 14286 8156
rect 14303 8092 14367 8156
rect 14384 8092 14448 8156
rect 14465 8092 14529 8156
rect 14546 8092 14610 8156
rect 14627 8092 14691 8156
rect 14708 8092 14772 8156
rect 14789 8092 14853 8156
rect 14870 8092 14934 8156
rect 106 8006 170 8070
rect 187 8006 251 8070
rect 268 8006 332 8070
rect 349 8006 413 8070
rect 430 8006 494 8070
rect 510 8006 574 8070
rect 590 8006 654 8070
rect 670 8006 734 8070
rect 750 8006 814 8070
rect 830 8006 894 8070
rect 910 8006 974 8070
rect 990 8006 1054 8070
rect 1070 8006 1134 8070
rect 1150 8006 1214 8070
rect 1230 8006 1294 8070
rect 1310 8006 1374 8070
rect 1390 8006 1454 8070
rect 1470 8006 1534 8070
rect 1550 8006 1614 8070
rect 1630 8006 1694 8070
rect 1710 8006 1774 8070
rect 1790 8006 1854 8070
rect 1870 8006 1934 8070
rect 1950 8006 2014 8070
rect 2030 8006 2094 8070
rect 2110 8006 2174 8070
rect 2190 8006 2254 8070
rect 2270 8006 2334 8070
rect 2350 8006 2414 8070
rect 2430 8006 2494 8070
rect 2510 8006 2574 8070
rect 2590 8006 2654 8070
rect 2670 8006 2734 8070
rect 2750 8006 2814 8070
rect 2830 8006 2894 8070
rect 2910 8006 2974 8070
rect 2990 8006 3054 8070
rect 3070 8006 3134 8070
rect 3150 8006 3214 8070
rect 3230 8006 3294 8070
rect 3310 8006 3374 8070
rect 3390 8006 3454 8070
rect 3470 8006 3534 8070
rect 3550 8006 3614 8070
rect 3630 8006 3694 8070
rect 3710 8006 3774 8070
rect 3790 8006 3854 8070
rect 3870 8006 3934 8070
rect 3950 8006 4014 8070
rect 4030 8006 4094 8070
rect 4110 8006 4174 8070
rect 4190 8006 4254 8070
rect 4270 8006 4334 8070
rect 4350 8006 4414 8070
rect 4430 8006 4494 8070
rect 4510 8006 4574 8070
rect 4590 8006 4654 8070
rect 4670 8006 4734 8070
rect 4750 8006 4814 8070
rect 4830 8006 4894 8070
rect 10157 8006 10221 8070
rect 10239 8006 10303 8070
rect 10321 8006 10385 8070
rect 10403 8006 10467 8070
rect 10485 8006 10549 8070
rect 10567 8006 10631 8070
rect 10649 8006 10713 8070
rect 10731 8006 10795 8070
rect 10813 8006 10877 8070
rect 10895 8006 10959 8070
rect 10977 8006 11041 8070
rect 11059 8006 11123 8070
rect 11141 8006 11205 8070
rect 11223 8006 11287 8070
rect 11305 8006 11369 8070
rect 11387 8006 11451 8070
rect 11468 8006 11532 8070
rect 11549 8006 11613 8070
rect 11630 8006 11694 8070
rect 11711 8006 11775 8070
rect 11792 8006 11856 8070
rect 11873 8006 11937 8070
rect 11954 8006 12018 8070
rect 12035 8006 12099 8070
rect 12116 8006 12180 8070
rect 12197 8006 12261 8070
rect 12278 8006 12342 8070
rect 12359 8006 12423 8070
rect 12440 8006 12504 8070
rect 12521 8006 12585 8070
rect 12602 8006 12666 8070
rect 12683 8006 12747 8070
rect 12764 8006 12828 8070
rect 12845 8006 12909 8070
rect 12926 8006 12990 8070
rect 13007 8006 13071 8070
rect 13088 8006 13152 8070
rect 13169 8006 13233 8070
rect 13250 8006 13314 8070
rect 13331 8006 13395 8070
rect 13412 8006 13476 8070
rect 13493 8006 13557 8070
rect 13574 8006 13638 8070
rect 13655 8006 13719 8070
rect 13736 8006 13800 8070
rect 13817 8006 13881 8070
rect 13898 8006 13962 8070
rect 13979 8006 14043 8070
rect 14060 8006 14124 8070
rect 14141 8006 14205 8070
rect 14222 8006 14286 8070
rect 14303 8006 14367 8070
rect 14384 8006 14448 8070
rect 14465 8006 14529 8070
rect 14546 8006 14610 8070
rect 14627 8006 14691 8070
rect 14708 8006 14772 8070
rect 14789 8006 14853 8070
rect 14870 8006 14934 8070
rect 106 7920 170 7984
rect 187 7920 251 7984
rect 268 7920 332 7984
rect 349 7920 413 7984
rect 430 7920 494 7984
rect 510 7920 574 7984
rect 590 7920 654 7984
rect 670 7920 734 7984
rect 750 7920 814 7984
rect 830 7920 894 7984
rect 910 7920 974 7984
rect 990 7920 1054 7984
rect 1070 7920 1134 7984
rect 1150 7920 1214 7984
rect 1230 7920 1294 7984
rect 1310 7920 1374 7984
rect 1390 7920 1454 7984
rect 1470 7920 1534 7984
rect 1550 7920 1614 7984
rect 1630 7920 1694 7984
rect 1710 7920 1774 7984
rect 1790 7920 1854 7984
rect 1870 7920 1934 7984
rect 1950 7920 2014 7984
rect 2030 7920 2094 7984
rect 2110 7920 2174 7984
rect 2190 7920 2254 7984
rect 2270 7920 2334 7984
rect 2350 7920 2414 7984
rect 2430 7920 2494 7984
rect 2510 7920 2574 7984
rect 2590 7920 2654 7984
rect 2670 7920 2734 7984
rect 2750 7920 2814 7984
rect 2830 7920 2894 7984
rect 2910 7920 2974 7984
rect 2990 7920 3054 7984
rect 3070 7920 3134 7984
rect 3150 7920 3214 7984
rect 3230 7920 3294 7984
rect 3310 7920 3374 7984
rect 3390 7920 3454 7984
rect 3470 7920 3534 7984
rect 3550 7920 3614 7984
rect 3630 7920 3694 7984
rect 3710 7920 3774 7984
rect 3790 7920 3854 7984
rect 3870 7920 3934 7984
rect 3950 7920 4014 7984
rect 4030 7920 4094 7984
rect 4110 7920 4174 7984
rect 4190 7920 4254 7984
rect 4270 7920 4334 7984
rect 4350 7920 4414 7984
rect 4430 7920 4494 7984
rect 4510 7920 4574 7984
rect 4590 7920 4654 7984
rect 4670 7920 4734 7984
rect 4750 7920 4814 7984
rect 4830 7920 4894 7984
rect 10157 7920 10221 7984
rect 10239 7920 10303 7984
rect 10321 7920 10385 7984
rect 10403 7920 10467 7984
rect 10485 7920 10549 7984
rect 10567 7920 10631 7984
rect 10649 7920 10713 7984
rect 10731 7920 10795 7984
rect 10813 7920 10877 7984
rect 10895 7920 10959 7984
rect 10977 7920 11041 7984
rect 11059 7920 11123 7984
rect 11141 7920 11205 7984
rect 11223 7920 11287 7984
rect 11305 7920 11369 7984
rect 11387 7920 11451 7984
rect 11468 7920 11532 7984
rect 11549 7920 11613 7984
rect 11630 7920 11694 7984
rect 11711 7920 11775 7984
rect 11792 7920 11856 7984
rect 11873 7920 11937 7984
rect 11954 7920 12018 7984
rect 12035 7920 12099 7984
rect 12116 7920 12180 7984
rect 12197 7920 12261 7984
rect 12278 7920 12342 7984
rect 12359 7920 12423 7984
rect 12440 7920 12504 7984
rect 12521 7920 12585 7984
rect 12602 7920 12666 7984
rect 12683 7920 12747 7984
rect 12764 7920 12828 7984
rect 12845 7920 12909 7984
rect 12926 7920 12990 7984
rect 13007 7920 13071 7984
rect 13088 7920 13152 7984
rect 13169 7920 13233 7984
rect 13250 7920 13314 7984
rect 13331 7920 13395 7984
rect 13412 7920 13476 7984
rect 13493 7920 13557 7984
rect 13574 7920 13638 7984
rect 13655 7920 13719 7984
rect 13736 7920 13800 7984
rect 13817 7920 13881 7984
rect 13898 7920 13962 7984
rect 13979 7920 14043 7984
rect 14060 7920 14124 7984
rect 14141 7920 14205 7984
rect 14222 7920 14286 7984
rect 14303 7920 14367 7984
rect 14384 7920 14448 7984
rect 14465 7920 14529 7984
rect 14546 7920 14610 7984
rect 14627 7920 14691 7984
rect 14708 7920 14772 7984
rect 14789 7920 14853 7984
rect 14870 7920 14934 7984
<< obsm4 >>
rect 0 10901 15000 39600
rect 0 9949 15000 10145
rect 0 8844 15000 9193
rect 0 8780 106 8844
rect 170 8780 187 8844
rect 251 8780 268 8844
rect 332 8780 349 8844
rect 413 8780 430 8844
rect 494 8780 510 8844
rect 574 8780 590 8844
rect 654 8780 670 8844
rect 734 8780 750 8844
rect 814 8780 830 8844
rect 894 8780 910 8844
rect 974 8780 990 8844
rect 1054 8780 1070 8844
rect 1134 8780 1150 8844
rect 1214 8780 1230 8844
rect 1294 8780 1310 8844
rect 1374 8780 1390 8844
rect 1454 8780 1470 8844
rect 1534 8780 1550 8844
rect 1614 8780 1630 8844
rect 1694 8780 1710 8844
rect 1774 8780 1790 8844
rect 1854 8780 1870 8844
rect 1934 8780 1950 8844
rect 2014 8780 2030 8844
rect 2094 8780 2110 8844
rect 2174 8780 2190 8844
rect 2254 8780 2270 8844
rect 2334 8780 2350 8844
rect 2414 8780 2430 8844
rect 2494 8780 2510 8844
rect 2574 8780 2590 8844
rect 2654 8780 2670 8844
rect 2734 8780 2750 8844
rect 2814 8780 2830 8844
rect 2894 8780 2910 8844
rect 2974 8780 2990 8844
rect 3054 8780 3070 8844
rect 3134 8780 3150 8844
rect 3214 8780 3230 8844
rect 3294 8780 3310 8844
rect 3374 8780 3390 8844
rect 3454 8780 3470 8844
rect 3534 8780 3550 8844
rect 3614 8780 3630 8844
rect 3694 8780 3710 8844
rect 3774 8780 3790 8844
rect 3854 8780 3870 8844
rect 3934 8780 3950 8844
rect 4014 8780 4030 8844
rect 4094 8780 4110 8844
rect 4174 8780 4190 8844
rect 4254 8780 4270 8844
rect 4334 8780 4350 8844
rect 4414 8780 4430 8844
rect 4494 8780 4510 8844
rect 4574 8780 4590 8844
rect 4654 8780 4670 8844
rect 4734 8780 4750 8844
rect 4814 8780 4830 8844
rect 4894 8780 10157 8844
rect 10221 8780 10239 8844
rect 10303 8780 10321 8844
rect 10385 8780 10403 8844
rect 10467 8780 10485 8844
rect 10549 8780 10567 8844
rect 10631 8780 10649 8844
rect 10713 8780 10731 8844
rect 10795 8780 10813 8844
rect 10877 8780 10895 8844
rect 10959 8780 10977 8844
rect 11041 8780 11059 8844
rect 11123 8780 11141 8844
rect 11205 8780 11223 8844
rect 11287 8780 11305 8844
rect 11369 8780 11387 8844
rect 11451 8780 11468 8844
rect 11532 8780 11549 8844
rect 11613 8780 11630 8844
rect 11694 8780 11711 8844
rect 11775 8780 11792 8844
rect 11856 8780 11873 8844
rect 11937 8780 11954 8844
rect 12018 8780 12035 8844
rect 12099 8780 12116 8844
rect 12180 8780 12197 8844
rect 12261 8780 12278 8844
rect 12342 8780 12359 8844
rect 12423 8780 12440 8844
rect 12504 8780 12521 8844
rect 12585 8780 12602 8844
rect 12666 8780 12683 8844
rect 12747 8780 12764 8844
rect 12828 8780 12845 8844
rect 12909 8780 12926 8844
rect 12990 8780 13007 8844
rect 13071 8780 13088 8844
rect 13152 8780 13169 8844
rect 13233 8780 13250 8844
rect 13314 8780 13331 8844
rect 13395 8780 13412 8844
rect 13476 8780 13493 8844
rect 13557 8780 13574 8844
rect 13638 8780 13655 8844
rect 13719 8780 13736 8844
rect 13800 8780 13817 8844
rect 13881 8780 13898 8844
rect 13962 8780 13979 8844
rect 14043 8780 14060 8844
rect 14124 8780 14141 8844
rect 14205 8780 14222 8844
rect 14286 8780 14303 8844
rect 14367 8780 14384 8844
rect 14448 8780 14465 8844
rect 14529 8780 14546 8844
rect 14610 8780 14627 8844
rect 14691 8780 14708 8844
rect 14772 8780 14789 8844
rect 14853 8780 14870 8844
rect 14934 8780 15000 8844
rect 0 8758 15000 8780
rect 0 8694 106 8758
rect 170 8694 187 8758
rect 251 8694 268 8758
rect 332 8694 349 8758
rect 413 8694 430 8758
rect 494 8694 510 8758
rect 574 8694 590 8758
rect 654 8694 670 8758
rect 734 8694 750 8758
rect 814 8694 830 8758
rect 894 8694 910 8758
rect 974 8694 990 8758
rect 1054 8694 1070 8758
rect 1134 8694 1150 8758
rect 1214 8694 1230 8758
rect 1294 8694 1310 8758
rect 1374 8694 1390 8758
rect 1454 8694 1470 8758
rect 1534 8694 1550 8758
rect 1614 8694 1630 8758
rect 1694 8694 1710 8758
rect 1774 8694 1790 8758
rect 1854 8694 1870 8758
rect 1934 8694 1950 8758
rect 2014 8694 2030 8758
rect 2094 8694 2110 8758
rect 2174 8694 2190 8758
rect 2254 8694 2270 8758
rect 2334 8694 2350 8758
rect 2414 8694 2430 8758
rect 2494 8694 2510 8758
rect 2574 8694 2590 8758
rect 2654 8694 2670 8758
rect 2734 8694 2750 8758
rect 2814 8694 2830 8758
rect 2894 8694 2910 8758
rect 2974 8694 2990 8758
rect 3054 8694 3070 8758
rect 3134 8694 3150 8758
rect 3214 8694 3230 8758
rect 3294 8694 3310 8758
rect 3374 8694 3390 8758
rect 3454 8694 3470 8758
rect 3534 8694 3550 8758
rect 3614 8694 3630 8758
rect 3694 8694 3710 8758
rect 3774 8694 3790 8758
rect 3854 8694 3870 8758
rect 3934 8694 3950 8758
rect 4014 8694 4030 8758
rect 4094 8694 4110 8758
rect 4174 8694 4190 8758
rect 4254 8694 4270 8758
rect 4334 8694 4350 8758
rect 4414 8694 4430 8758
rect 4494 8694 4510 8758
rect 4574 8694 4590 8758
rect 4654 8694 4670 8758
rect 4734 8694 4750 8758
rect 4814 8694 4830 8758
rect 4894 8694 10157 8758
rect 10221 8694 10239 8758
rect 10303 8694 10321 8758
rect 10385 8694 10403 8758
rect 10467 8694 10485 8758
rect 10549 8694 10567 8758
rect 10631 8694 10649 8758
rect 10713 8694 10731 8758
rect 10795 8694 10813 8758
rect 10877 8694 10895 8758
rect 10959 8694 10977 8758
rect 11041 8694 11059 8758
rect 11123 8694 11141 8758
rect 11205 8694 11223 8758
rect 11287 8694 11305 8758
rect 11369 8694 11387 8758
rect 11451 8694 11468 8758
rect 11532 8694 11549 8758
rect 11613 8694 11630 8758
rect 11694 8694 11711 8758
rect 11775 8694 11792 8758
rect 11856 8694 11873 8758
rect 11937 8694 11954 8758
rect 12018 8694 12035 8758
rect 12099 8694 12116 8758
rect 12180 8694 12197 8758
rect 12261 8694 12278 8758
rect 12342 8694 12359 8758
rect 12423 8694 12440 8758
rect 12504 8694 12521 8758
rect 12585 8694 12602 8758
rect 12666 8694 12683 8758
rect 12747 8694 12764 8758
rect 12828 8694 12845 8758
rect 12909 8694 12926 8758
rect 12990 8694 13007 8758
rect 13071 8694 13088 8758
rect 13152 8694 13169 8758
rect 13233 8694 13250 8758
rect 13314 8694 13331 8758
rect 13395 8694 13412 8758
rect 13476 8694 13493 8758
rect 13557 8694 13574 8758
rect 13638 8694 13655 8758
rect 13719 8694 13736 8758
rect 13800 8694 13817 8758
rect 13881 8694 13898 8758
rect 13962 8694 13979 8758
rect 14043 8694 14060 8758
rect 14124 8694 14141 8758
rect 14205 8694 14222 8758
rect 14286 8694 14303 8758
rect 14367 8694 14384 8758
rect 14448 8694 14465 8758
rect 14529 8694 14546 8758
rect 14610 8694 14627 8758
rect 14691 8694 14708 8758
rect 14772 8694 14789 8758
rect 14853 8694 14870 8758
rect 14934 8694 15000 8758
rect 0 8672 15000 8694
rect 0 8608 106 8672
rect 170 8608 187 8672
rect 251 8608 268 8672
rect 332 8608 349 8672
rect 413 8608 430 8672
rect 494 8608 510 8672
rect 574 8608 590 8672
rect 654 8608 670 8672
rect 734 8608 750 8672
rect 814 8608 830 8672
rect 894 8608 910 8672
rect 974 8608 990 8672
rect 1054 8608 1070 8672
rect 1134 8608 1150 8672
rect 1214 8608 1230 8672
rect 1294 8608 1310 8672
rect 1374 8608 1390 8672
rect 1454 8608 1470 8672
rect 1534 8608 1550 8672
rect 1614 8608 1630 8672
rect 1694 8608 1710 8672
rect 1774 8608 1790 8672
rect 1854 8608 1870 8672
rect 1934 8608 1950 8672
rect 2014 8608 2030 8672
rect 2094 8608 2110 8672
rect 2174 8608 2190 8672
rect 2254 8608 2270 8672
rect 2334 8608 2350 8672
rect 2414 8608 2430 8672
rect 2494 8608 2510 8672
rect 2574 8608 2590 8672
rect 2654 8608 2670 8672
rect 2734 8608 2750 8672
rect 2814 8608 2830 8672
rect 2894 8608 2910 8672
rect 2974 8608 2990 8672
rect 3054 8608 3070 8672
rect 3134 8608 3150 8672
rect 3214 8608 3230 8672
rect 3294 8608 3310 8672
rect 3374 8608 3390 8672
rect 3454 8608 3470 8672
rect 3534 8608 3550 8672
rect 3614 8608 3630 8672
rect 3694 8608 3710 8672
rect 3774 8608 3790 8672
rect 3854 8608 3870 8672
rect 3934 8608 3950 8672
rect 4014 8608 4030 8672
rect 4094 8608 4110 8672
rect 4174 8608 4190 8672
rect 4254 8608 4270 8672
rect 4334 8608 4350 8672
rect 4414 8608 4430 8672
rect 4494 8608 4510 8672
rect 4574 8608 4590 8672
rect 4654 8608 4670 8672
rect 4734 8608 4750 8672
rect 4814 8608 4830 8672
rect 4894 8608 10157 8672
rect 10221 8608 10239 8672
rect 10303 8608 10321 8672
rect 10385 8608 10403 8672
rect 10467 8608 10485 8672
rect 10549 8608 10567 8672
rect 10631 8608 10649 8672
rect 10713 8608 10731 8672
rect 10795 8608 10813 8672
rect 10877 8608 10895 8672
rect 10959 8608 10977 8672
rect 11041 8608 11059 8672
rect 11123 8608 11141 8672
rect 11205 8608 11223 8672
rect 11287 8608 11305 8672
rect 11369 8608 11387 8672
rect 11451 8608 11468 8672
rect 11532 8608 11549 8672
rect 11613 8608 11630 8672
rect 11694 8608 11711 8672
rect 11775 8608 11792 8672
rect 11856 8608 11873 8672
rect 11937 8608 11954 8672
rect 12018 8608 12035 8672
rect 12099 8608 12116 8672
rect 12180 8608 12197 8672
rect 12261 8608 12278 8672
rect 12342 8608 12359 8672
rect 12423 8608 12440 8672
rect 12504 8608 12521 8672
rect 12585 8608 12602 8672
rect 12666 8608 12683 8672
rect 12747 8608 12764 8672
rect 12828 8608 12845 8672
rect 12909 8608 12926 8672
rect 12990 8608 13007 8672
rect 13071 8608 13088 8672
rect 13152 8608 13169 8672
rect 13233 8608 13250 8672
rect 13314 8608 13331 8672
rect 13395 8608 13412 8672
rect 13476 8608 13493 8672
rect 13557 8608 13574 8672
rect 13638 8608 13655 8672
rect 13719 8608 13736 8672
rect 13800 8608 13817 8672
rect 13881 8608 13898 8672
rect 13962 8608 13979 8672
rect 14043 8608 14060 8672
rect 14124 8608 14141 8672
rect 14205 8608 14222 8672
rect 14286 8608 14303 8672
rect 14367 8608 14384 8672
rect 14448 8608 14465 8672
rect 14529 8608 14546 8672
rect 14610 8608 14627 8672
rect 14691 8608 14708 8672
rect 14772 8608 14789 8672
rect 14853 8608 14870 8672
rect 14934 8608 15000 8672
rect 0 8586 15000 8608
rect 0 8522 106 8586
rect 170 8522 187 8586
rect 251 8522 268 8586
rect 332 8522 349 8586
rect 413 8522 430 8586
rect 494 8522 510 8586
rect 574 8522 590 8586
rect 654 8522 670 8586
rect 734 8522 750 8586
rect 814 8522 830 8586
rect 894 8522 910 8586
rect 974 8522 990 8586
rect 1054 8522 1070 8586
rect 1134 8522 1150 8586
rect 1214 8522 1230 8586
rect 1294 8522 1310 8586
rect 1374 8522 1390 8586
rect 1454 8522 1470 8586
rect 1534 8522 1550 8586
rect 1614 8522 1630 8586
rect 1694 8522 1710 8586
rect 1774 8522 1790 8586
rect 1854 8522 1870 8586
rect 1934 8522 1950 8586
rect 2014 8522 2030 8586
rect 2094 8522 2110 8586
rect 2174 8522 2190 8586
rect 2254 8522 2270 8586
rect 2334 8522 2350 8586
rect 2414 8522 2430 8586
rect 2494 8522 2510 8586
rect 2574 8522 2590 8586
rect 2654 8522 2670 8586
rect 2734 8522 2750 8586
rect 2814 8522 2830 8586
rect 2894 8522 2910 8586
rect 2974 8522 2990 8586
rect 3054 8522 3070 8586
rect 3134 8522 3150 8586
rect 3214 8522 3230 8586
rect 3294 8522 3310 8586
rect 3374 8522 3390 8586
rect 3454 8522 3470 8586
rect 3534 8522 3550 8586
rect 3614 8522 3630 8586
rect 3694 8522 3710 8586
rect 3774 8522 3790 8586
rect 3854 8522 3870 8586
rect 3934 8522 3950 8586
rect 4014 8522 4030 8586
rect 4094 8522 4110 8586
rect 4174 8522 4190 8586
rect 4254 8522 4270 8586
rect 4334 8522 4350 8586
rect 4414 8522 4430 8586
rect 4494 8522 4510 8586
rect 4574 8522 4590 8586
rect 4654 8522 4670 8586
rect 4734 8522 4750 8586
rect 4814 8522 4830 8586
rect 4894 8522 10157 8586
rect 10221 8522 10239 8586
rect 10303 8522 10321 8586
rect 10385 8522 10403 8586
rect 10467 8522 10485 8586
rect 10549 8522 10567 8586
rect 10631 8522 10649 8586
rect 10713 8522 10731 8586
rect 10795 8522 10813 8586
rect 10877 8522 10895 8586
rect 10959 8522 10977 8586
rect 11041 8522 11059 8586
rect 11123 8522 11141 8586
rect 11205 8522 11223 8586
rect 11287 8522 11305 8586
rect 11369 8522 11387 8586
rect 11451 8522 11468 8586
rect 11532 8522 11549 8586
rect 11613 8522 11630 8586
rect 11694 8522 11711 8586
rect 11775 8522 11792 8586
rect 11856 8522 11873 8586
rect 11937 8522 11954 8586
rect 12018 8522 12035 8586
rect 12099 8522 12116 8586
rect 12180 8522 12197 8586
rect 12261 8522 12278 8586
rect 12342 8522 12359 8586
rect 12423 8522 12440 8586
rect 12504 8522 12521 8586
rect 12585 8522 12602 8586
rect 12666 8522 12683 8586
rect 12747 8522 12764 8586
rect 12828 8522 12845 8586
rect 12909 8522 12926 8586
rect 12990 8522 13007 8586
rect 13071 8522 13088 8586
rect 13152 8522 13169 8586
rect 13233 8522 13250 8586
rect 13314 8522 13331 8586
rect 13395 8522 13412 8586
rect 13476 8522 13493 8586
rect 13557 8522 13574 8586
rect 13638 8522 13655 8586
rect 13719 8522 13736 8586
rect 13800 8522 13817 8586
rect 13881 8522 13898 8586
rect 13962 8522 13979 8586
rect 14043 8522 14060 8586
rect 14124 8522 14141 8586
rect 14205 8522 14222 8586
rect 14286 8522 14303 8586
rect 14367 8522 14384 8586
rect 14448 8522 14465 8586
rect 14529 8522 14546 8586
rect 14610 8522 14627 8586
rect 14691 8522 14708 8586
rect 14772 8522 14789 8586
rect 14853 8522 14870 8586
rect 14934 8522 15000 8586
rect 0 8500 15000 8522
rect 0 8436 106 8500
rect 170 8436 187 8500
rect 251 8436 268 8500
rect 332 8436 349 8500
rect 413 8436 430 8500
rect 494 8436 510 8500
rect 574 8436 590 8500
rect 654 8436 670 8500
rect 734 8436 750 8500
rect 814 8436 830 8500
rect 894 8436 910 8500
rect 974 8436 990 8500
rect 1054 8436 1070 8500
rect 1134 8436 1150 8500
rect 1214 8436 1230 8500
rect 1294 8436 1310 8500
rect 1374 8436 1390 8500
rect 1454 8436 1470 8500
rect 1534 8436 1550 8500
rect 1614 8436 1630 8500
rect 1694 8436 1710 8500
rect 1774 8436 1790 8500
rect 1854 8436 1870 8500
rect 1934 8436 1950 8500
rect 2014 8436 2030 8500
rect 2094 8436 2110 8500
rect 2174 8436 2190 8500
rect 2254 8436 2270 8500
rect 2334 8436 2350 8500
rect 2414 8436 2430 8500
rect 2494 8436 2510 8500
rect 2574 8436 2590 8500
rect 2654 8436 2670 8500
rect 2734 8436 2750 8500
rect 2814 8436 2830 8500
rect 2894 8436 2910 8500
rect 2974 8436 2990 8500
rect 3054 8436 3070 8500
rect 3134 8436 3150 8500
rect 3214 8436 3230 8500
rect 3294 8436 3310 8500
rect 3374 8436 3390 8500
rect 3454 8436 3470 8500
rect 3534 8436 3550 8500
rect 3614 8436 3630 8500
rect 3694 8436 3710 8500
rect 3774 8436 3790 8500
rect 3854 8436 3870 8500
rect 3934 8436 3950 8500
rect 4014 8436 4030 8500
rect 4094 8436 4110 8500
rect 4174 8436 4190 8500
rect 4254 8436 4270 8500
rect 4334 8436 4350 8500
rect 4414 8436 4430 8500
rect 4494 8436 4510 8500
rect 4574 8436 4590 8500
rect 4654 8436 4670 8500
rect 4734 8436 4750 8500
rect 4814 8436 4830 8500
rect 4894 8436 10157 8500
rect 10221 8436 10239 8500
rect 10303 8436 10321 8500
rect 10385 8436 10403 8500
rect 10467 8436 10485 8500
rect 10549 8436 10567 8500
rect 10631 8436 10649 8500
rect 10713 8436 10731 8500
rect 10795 8436 10813 8500
rect 10877 8436 10895 8500
rect 10959 8436 10977 8500
rect 11041 8436 11059 8500
rect 11123 8436 11141 8500
rect 11205 8436 11223 8500
rect 11287 8436 11305 8500
rect 11369 8436 11387 8500
rect 11451 8436 11468 8500
rect 11532 8436 11549 8500
rect 11613 8436 11630 8500
rect 11694 8436 11711 8500
rect 11775 8436 11792 8500
rect 11856 8436 11873 8500
rect 11937 8436 11954 8500
rect 12018 8436 12035 8500
rect 12099 8436 12116 8500
rect 12180 8436 12197 8500
rect 12261 8436 12278 8500
rect 12342 8436 12359 8500
rect 12423 8436 12440 8500
rect 12504 8436 12521 8500
rect 12585 8436 12602 8500
rect 12666 8436 12683 8500
rect 12747 8436 12764 8500
rect 12828 8436 12845 8500
rect 12909 8436 12926 8500
rect 12990 8436 13007 8500
rect 13071 8436 13088 8500
rect 13152 8436 13169 8500
rect 13233 8436 13250 8500
rect 13314 8436 13331 8500
rect 13395 8436 13412 8500
rect 13476 8436 13493 8500
rect 13557 8436 13574 8500
rect 13638 8436 13655 8500
rect 13719 8436 13736 8500
rect 13800 8436 13817 8500
rect 13881 8436 13898 8500
rect 13962 8436 13979 8500
rect 14043 8436 14060 8500
rect 14124 8436 14141 8500
rect 14205 8436 14222 8500
rect 14286 8436 14303 8500
rect 14367 8436 14384 8500
rect 14448 8436 14465 8500
rect 14529 8436 14546 8500
rect 14610 8436 14627 8500
rect 14691 8436 14708 8500
rect 14772 8436 14789 8500
rect 14853 8436 14870 8500
rect 14934 8436 15000 8500
rect 0 8414 15000 8436
rect 0 8350 106 8414
rect 170 8350 187 8414
rect 251 8350 268 8414
rect 332 8350 349 8414
rect 413 8350 430 8414
rect 494 8350 510 8414
rect 574 8350 590 8414
rect 654 8350 670 8414
rect 734 8350 750 8414
rect 814 8350 830 8414
rect 894 8350 910 8414
rect 974 8350 990 8414
rect 1054 8350 1070 8414
rect 1134 8350 1150 8414
rect 1214 8350 1230 8414
rect 1294 8350 1310 8414
rect 1374 8350 1390 8414
rect 1454 8350 1470 8414
rect 1534 8350 1550 8414
rect 1614 8350 1630 8414
rect 1694 8350 1710 8414
rect 1774 8350 1790 8414
rect 1854 8350 1870 8414
rect 1934 8350 1950 8414
rect 2014 8350 2030 8414
rect 2094 8350 2110 8414
rect 2174 8350 2190 8414
rect 2254 8350 2270 8414
rect 2334 8350 2350 8414
rect 2414 8350 2430 8414
rect 2494 8350 2510 8414
rect 2574 8350 2590 8414
rect 2654 8350 2670 8414
rect 2734 8350 2750 8414
rect 2814 8350 2830 8414
rect 2894 8350 2910 8414
rect 2974 8350 2990 8414
rect 3054 8350 3070 8414
rect 3134 8350 3150 8414
rect 3214 8350 3230 8414
rect 3294 8350 3310 8414
rect 3374 8350 3390 8414
rect 3454 8350 3470 8414
rect 3534 8350 3550 8414
rect 3614 8350 3630 8414
rect 3694 8350 3710 8414
rect 3774 8350 3790 8414
rect 3854 8350 3870 8414
rect 3934 8350 3950 8414
rect 4014 8350 4030 8414
rect 4094 8350 4110 8414
rect 4174 8350 4190 8414
rect 4254 8350 4270 8414
rect 4334 8350 4350 8414
rect 4414 8350 4430 8414
rect 4494 8350 4510 8414
rect 4574 8350 4590 8414
rect 4654 8350 4670 8414
rect 4734 8350 4750 8414
rect 4814 8350 4830 8414
rect 4894 8350 10157 8414
rect 10221 8350 10239 8414
rect 10303 8350 10321 8414
rect 10385 8350 10403 8414
rect 10467 8350 10485 8414
rect 10549 8350 10567 8414
rect 10631 8350 10649 8414
rect 10713 8350 10731 8414
rect 10795 8350 10813 8414
rect 10877 8350 10895 8414
rect 10959 8350 10977 8414
rect 11041 8350 11059 8414
rect 11123 8350 11141 8414
rect 11205 8350 11223 8414
rect 11287 8350 11305 8414
rect 11369 8350 11387 8414
rect 11451 8350 11468 8414
rect 11532 8350 11549 8414
rect 11613 8350 11630 8414
rect 11694 8350 11711 8414
rect 11775 8350 11792 8414
rect 11856 8350 11873 8414
rect 11937 8350 11954 8414
rect 12018 8350 12035 8414
rect 12099 8350 12116 8414
rect 12180 8350 12197 8414
rect 12261 8350 12278 8414
rect 12342 8350 12359 8414
rect 12423 8350 12440 8414
rect 12504 8350 12521 8414
rect 12585 8350 12602 8414
rect 12666 8350 12683 8414
rect 12747 8350 12764 8414
rect 12828 8350 12845 8414
rect 12909 8350 12926 8414
rect 12990 8350 13007 8414
rect 13071 8350 13088 8414
rect 13152 8350 13169 8414
rect 13233 8350 13250 8414
rect 13314 8350 13331 8414
rect 13395 8350 13412 8414
rect 13476 8350 13493 8414
rect 13557 8350 13574 8414
rect 13638 8350 13655 8414
rect 13719 8350 13736 8414
rect 13800 8350 13817 8414
rect 13881 8350 13898 8414
rect 13962 8350 13979 8414
rect 14043 8350 14060 8414
rect 14124 8350 14141 8414
rect 14205 8350 14222 8414
rect 14286 8350 14303 8414
rect 14367 8350 14384 8414
rect 14448 8350 14465 8414
rect 14529 8350 14546 8414
rect 14610 8350 14627 8414
rect 14691 8350 14708 8414
rect 14772 8350 14789 8414
rect 14853 8350 14870 8414
rect 14934 8350 15000 8414
rect 0 8328 15000 8350
rect 0 8264 106 8328
rect 170 8264 187 8328
rect 251 8264 268 8328
rect 332 8264 349 8328
rect 413 8264 430 8328
rect 494 8264 510 8328
rect 574 8264 590 8328
rect 654 8264 670 8328
rect 734 8264 750 8328
rect 814 8264 830 8328
rect 894 8264 910 8328
rect 974 8264 990 8328
rect 1054 8264 1070 8328
rect 1134 8264 1150 8328
rect 1214 8264 1230 8328
rect 1294 8264 1310 8328
rect 1374 8264 1390 8328
rect 1454 8264 1470 8328
rect 1534 8264 1550 8328
rect 1614 8264 1630 8328
rect 1694 8264 1710 8328
rect 1774 8264 1790 8328
rect 1854 8264 1870 8328
rect 1934 8264 1950 8328
rect 2014 8264 2030 8328
rect 2094 8264 2110 8328
rect 2174 8264 2190 8328
rect 2254 8264 2270 8328
rect 2334 8264 2350 8328
rect 2414 8264 2430 8328
rect 2494 8264 2510 8328
rect 2574 8264 2590 8328
rect 2654 8264 2670 8328
rect 2734 8264 2750 8328
rect 2814 8264 2830 8328
rect 2894 8264 2910 8328
rect 2974 8264 2990 8328
rect 3054 8264 3070 8328
rect 3134 8264 3150 8328
rect 3214 8264 3230 8328
rect 3294 8264 3310 8328
rect 3374 8264 3390 8328
rect 3454 8264 3470 8328
rect 3534 8264 3550 8328
rect 3614 8264 3630 8328
rect 3694 8264 3710 8328
rect 3774 8264 3790 8328
rect 3854 8264 3870 8328
rect 3934 8264 3950 8328
rect 4014 8264 4030 8328
rect 4094 8264 4110 8328
rect 4174 8264 4190 8328
rect 4254 8264 4270 8328
rect 4334 8264 4350 8328
rect 4414 8264 4430 8328
rect 4494 8264 4510 8328
rect 4574 8264 4590 8328
rect 4654 8264 4670 8328
rect 4734 8264 4750 8328
rect 4814 8264 4830 8328
rect 4894 8264 10157 8328
rect 10221 8264 10239 8328
rect 10303 8264 10321 8328
rect 10385 8264 10403 8328
rect 10467 8264 10485 8328
rect 10549 8264 10567 8328
rect 10631 8264 10649 8328
rect 10713 8264 10731 8328
rect 10795 8264 10813 8328
rect 10877 8264 10895 8328
rect 10959 8264 10977 8328
rect 11041 8264 11059 8328
rect 11123 8264 11141 8328
rect 11205 8264 11223 8328
rect 11287 8264 11305 8328
rect 11369 8264 11387 8328
rect 11451 8264 11468 8328
rect 11532 8264 11549 8328
rect 11613 8264 11630 8328
rect 11694 8264 11711 8328
rect 11775 8264 11792 8328
rect 11856 8264 11873 8328
rect 11937 8264 11954 8328
rect 12018 8264 12035 8328
rect 12099 8264 12116 8328
rect 12180 8264 12197 8328
rect 12261 8264 12278 8328
rect 12342 8264 12359 8328
rect 12423 8264 12440 8328
rect 12504 8264 12521 8328
rect 12585 8264 12602 8328
rect 12666 8264 12683 8328
rect 12747 8264 12764 8328
rect 12828 8264 12845 8328
rect 12909 8264 12926 8328
rect 12990 8264 13007 8328
rect 13071 8264 13088 8328
rect 13152 8264 13169 8328
rect 13233 8264 13250 8328
rect 13314 8264 13331 8328
rect 13395 8264 13412 8328
rect 13476 8264 13493 8328
rect 13557 8264 13574 8328
rect 13638 8264 13655 8328
rect 13719 8264 13736 8328
rect 13800 8264 13817 8328
rect 13881 8264 13898 8328
rect 13962 8264 13979 8328
rect 14043 8264 14060 8328
rect 14124 8264 14141 8328
rect 14205 8264 14222 8328
rect 14286 8264 14303 8328
rect 14367 8264 14384 8328
rect 14448 8264 14465 8328
rect 14529 8264 14546 8328
rect 14610 8264 14627 8328
rect 14691 8264 14708 8328
rect 14772 8264 14789 8328
rect 14853 8264 14870 8328
rect 14934 8264 15000 8328
rect 0 8242 15000 8264
rect 0 8178 106 8242
rect 170 8178 187 8242
rect 251 8178 268 8242
rect 332 8178 349 8242
rect 413 8178 430 8242
rect 494 8178 510 8242
rect 574 8178 590 8242
rect 654 8178 670 8242
rect 734 8178 750 8242
rect 814 8178 830 8242
rect 894 8178 910 8242
rect 974 8178 990 8242
rect 1054 8178 1070 8242
rect 1134 8178 1150 8242
rect 1214 8178 1230 8242
rect 1294 8178 1310 8242
rect 1374 8178 1390 8242
rect 1454 8178 1470 8242
rect 1534 8178 1550 8242
rect 1614 8178 1630 8242
rect 1694 8178 1710 8242
rect 1774 8178 1790 8242
rect 1854 8178 1870 8242
rect 1934 8178 1950 8242
rect 2014 8178 2030 8242
rect 2094 8178 2110 8242
rect 2174 8178 2190 8242
rect 2254 8178 2270 8242
rect 2334 8178 2350 8242
rect 2414 8178 2430 8242
rect 2494 8178 2510 8242
rect 2574 8178 2590 8242
rect 2654 8178 2670 8242
rect 2734 8178 2750 8242
rect 2814 8178 2830 8242
rect 2894 8178 2910 8242
rect 2974 8178 2990 8242
rect 3054 8178 3070 8242
rect 3134 8178 3150 8242
rect 3214 8178 3230 8242
rect 3294 8178 3310 8242
rect 3374 8178 3390 8242
rect 3454 8178 3470 8242
rect 3534 8178 3550 8242
rect 3614 8178 3630 8242
rect 3694 8178 3710 8242
rect 3774 8178 3790 8242
rect 3854 8178 3870 8242
rect 3934 8178 3950 8242
rect 4014 8178 4030 8242
rect 4094 8178 4110 8242
rect 4174 8178 4190 8242
rect 4254 8178 4270 8242
rect 4334 8178 4350 8242
rect 4414 8178 4430 8242
rect 4494 8178 4510 8242
rect 4574 8178 4590 8242
rect 4654 8178 4670 8242
rect 4734 8178 4750 8242
rect 4814 8178 4830 8242
rect 4894 8178 10157 8242
rect 10221 8178 10239 8242
rect 10303 8178 10321 8242
rect 10385 8178 10403 8242
rect 10467 8178 10485 8242
rect 10549 8178 10567 8242
rect 10631 8178 10649 8242
rect 10713 8178 10731 8242
rect 10795 8178 10813 8242
rect 10877 8178 10895 8242
rect 10959 8178 10977 8242
rect 11041 8178 11059 8242
rect 11123 8178 11141 8242
rect 11205 8178 11223 8242
rect 11287 8178 11305 8242
rect 11369 8178 11387 8242
rect 11451 8178 11468 8242
rect 11532 8178 11549 8242
rect 11613 8178 11630 8242
rect 11694 8178 11711 8242
rect 11775 8178 11792 8242
rect 11856 8178 11873 8242
rect 11937 8178 11954 8242
rect 12018 8178 12035 8242
rect 12099 8178 12116 8242
rect 12180 8178 12197 8242
rect 12261 8178 12278 8242
rect 12342 8178 12359 8242
rect 12423 8178 12440 8242
rect 12504 8178 12521 8242
rect 12585 8178 12602 8242
rect 12666 8178 12683 8242
rect 12747 8178 12764 8242
rect 12828 8178 12845 8242
rect 12909 8178 12926 8242
rect 12990 8178 13007 8242
rect 13071 8178 13088 8242
rect 13152 8178 13169 8242
rect 13233 8178 13250 8242
rect 13314 8178 13331 8242
rect 13395 8178 13412 8242
rect 13476 8178 13493 8242
rect 13557 8178 13574 8242
rect 13638 8178 13655 8242
rect 13719 8178 13736 8242
rect 13800 8178 13817 8242
rect 13881 8178 13898 8242
rect 13962 8178 13979 8242
rect 14043 8178 14060 8242
rect 14124 8178 14141 8242
rect 14205 8178 14222 8242
rect 14286 8178 14303 8242
rect 14367 8178 14384 8242
rect 14448 8178 14465 8242
rect 14529 8178 14546 8242
rect 14610 8178 14627 8242
rect 14691 8178 14708 8242
rect 14772 8178 14789 8242
rect 14853 8178 14870 8242
rect 14934 8178 15000 8242
rect 0 8156 15000 8178
rect 0 8092 106 8156
rect 170 8092 187 8156
rect 251 8092 268 8156
rect 332 8092 349 8156
rect 413 8092 430 8156
rect 494 8092 510 8156
rect 574 8092 590 8156
rect 654 8092 670 8156
rect 734 8092 750 8156
rect 814 8092 830 8156
rect 894 8092 910 8156
rect 974 8092 990 8156
rect 1054 8092 1070 8156
rect 1134 8092 1150 8156
rect 1214 8092 1230 8156
rect 1294 8092 1310 8156
rect 1374 8092 1390 8156
rect 1454 8092 1470 8156
rect 1534 8092 1550 8156
rect 1614 8092 1630 8156
rect 1694 8092 1710 8156
rect 1774 8092 1790 8156
rect 1854 8092 1870 8156
rect 1934 8092 1950 8156
rect 2014 8092 2030 8156
rect 2094 8092 2110 8156
rect 2174 8092 2190 8156
rect 2254 8092 2270 8156
rect 2334 8092 2350 8156
rect 2414 8092 2430 8156
rect 2494 8092 2510 8156
rect 2574 8092 2590 8156
rect 2654 8092 2670 8156
rect 2734 8092 2750 8156
rect 2814 8092 2830 8156
rect 2894 8092 2910 8156
rect 2974 8092 2990 8156
rect 3054 8092 3070 8156
rect 3134 8092 3150 8156
rect 3214 8092 3230 8156
rect 3294 8092 3310 8156
rect 3374 8092 3390 8156
rect 3454 8092 3470 8156
rect 3534 8092 3550 8156
rect 3614 8092 3630 8156
rect 3694 8092 3710 8156
rect 3774 8092 3790 8156
rect 3854 8092 3870 8156
rect 3934 8092 3950 8156
rect 4014 8092 4030 8156
rect 4094 8092 4110 8156
rect 4174 8092 4190 8156
rect 4254 8092 4270 8156
rect 4334 8092 4350 8156
rect 4414 8092 4430 8156
rect 4494 8092 4510 8156
rect 4574 8092 4590 8156
rect 4654 8092 4670 8156
rect 4734 8092 4750 8156
rect 4814 8092 4830 8156
rect 4894 8092 10157 8156
rect 10221 8092 10239 8156
rect 10303 8092 10321 8156
rect 10385 8092 10403 8156
rect 10467 8092 10485 8156
rect 10549 8092 10567 8156
rect 10631 8092 10649 8156
rect 10713 8092 10731 8156
rect 10795 8092 10813 8156
rect 10877 8092 10895 8156
rect 10959 8092 10977 8156
rect 11041 8092 11059 8156
rect 11123 8092 11141 8156
rect 11205 8092 11223 8156
rect 11287 8092 11305 8156
rect 11369 8092 11387 8156
rect 11451 8092 11468 8156
rect 11532 8092 11549 8156
rect 11613 8092 11630 8156
rect 11694 8092 11711 8156
rect 11775 8092 11792 8156
rect 11856 8092 11873 8156
rect 11937 8092 11954 8156
rect 12018 8092 12035 8156
rect 12099 8092 12116 8156
rect 12180 8092 12197 8156
rect 12261 8092 12278 8156
rect 12342 8092 12359 8156
rect 12423 8092 12440 8156
rect 12504 8092 12521 8156
rect 12585 8092 12602 8156
rect 12666 8092 12683 8156
rect 12747 8092 12764 8156
rect 12828 8092 12845 8156
rect 12909 8092 12926 8156
rect 12990 8092 13007 8156
rect 13071 8092 13088 8156
rect 13152 8092 13169 8156
rect 13233 8092 13250 8156
rect 13314 8092 13331 8156
rect 13395 8092 13412 8156
rect 13476 8092 13493 8156
rect 13557 8092 13574 8156
rect 13638 8092 13655 8156
rect 13719 8092 13736 8156
rect 13800 8092 13817 8156
rect 13881 8092 13898 8156
rect 13962 8092 13979 8156
rect 14043 8092 14060 8156
rect 14124 8092 14141 8156
rect 14205 8092 14222 8156
rect 14286 8092 14303 8156
rect 14367 8092 14384 8156
rect 14448 8092 14465 8156
rect 14529 8092 14546 8156
rect 14610 8092 14627 8156
rect 14691 8092 14708 8156
rect 14772 8092 14789 8156
rect 14853 8092 14870 8156
rect 14934 8092 15000 8156
rect 0 8070 15000 8092
rect 0 8006 106 8070
rect 170 8006 187 8070
rect 251 8006 268 8070
rect 332 8006 349 8070
rect 413 8006 430 8070
rect 494 8006 510 8070
rect 574 8006 590 8070
rect 654 8006 670 8070
rect 734 8006 750 8070
rect 814 8006 830 8070
rect 894 8006 910 8070
rect 974 8006 990 8070
rect 1054 8006 1070 8070
rect 1134 8006 1150 8070
rect 1214 8006 1230 8070
rect 1294 8006 1310 8070
rect 1374 8006 1390 8070
rect 1454 8006 1470 8070
rect 1534 8006 1550 8070
rect 1614 8006 1630 8070
rect 1694 8006 1710 8070
rect 1774 8006 1790 8070
rect 1854 8006 1870 8070
rect 1934 8006 1950 8070
rect 2014 8006 2030 8070
rect 2094 8006 2110 8070
rect 2174 8006 2190 8070
rect 2254 8006 2270 8070
rect 2334 8006 2350 8070
rect 2414 8006 2430 8070
rect 2494 8006 2510 8070
rect 2574 8006 2590 8070
rect 2654 8006 2670 8070
rect 2734 8006 2750 8070
rect 2814 8006 2830 8070
rect 2894 8006 2910 8070
rect 2974 8006 2990 8070
rect 3054 8006 3070 8070
rect 3134 8006 3150 8070
rect 3214 8006 3230 8070
rect 3294 8006 3310 8070
rect 3374 8006 3390 8070
rect 3454 8006 3470 8070
rect 3534 8006 3550 8070
rect 3614 8006 3630 8070
rect 3694 8006 3710 8070
rect 3774 8006 3790 8070
rect 3854 8006 3870 8070
rect 3934 8006 3950 8070
rect 4014 8006 4030 8070
rect 4094 8006 4110 8070
rect 4174 8006 4190 8070
rect 4254 8006 4270 8070
rect 4334 8006 4350 8070
rect 4414 8006 4430 8070
rect 4494 8006 4510 8070
rect 4574 8006 4590 8070
rect 4654 8006 4670 8070
rect 4734 8006 4750 8070
rect 4814 8006 4830 8070
rect 4894 8006 10157 8070
rect 10221 8006 10239 8070
rect 10303 8006 10321 8070
rect 10385 8006 10403 8070
rect 10467 8006 10485 8070
rect 10549 8006 10567 8070
rect 10631 8006 10649 8070
rect 10713 8006 10731 8070
rect 10795 8006 10813 8070
rect 10877 8006 10895 8070
rect 10959 8006 10977 8070
rect 11041 8006 11059 8070
rect 11123 8006 11141 8070
rect 11205 8006 11223 8070
rect 11287 8006 11305 8070
rect 11369 8006 11387 8070
rect 11451 8006 11468 8070
rect 11532 8006 11549 8070
rect 11613 8006 11630 8070
rect 11694 8006 11711 8070
rect 11775 8006 11792 8070
rect 11856 8006 11873 8070
rect 11937 8006 11954 8070
rect 12018 8006 12035 8070
rect 12099 8006 12116 8070
rect 12180 8006 12197 8070
rect 12261 8006 12278 8070
rect 12342 8006 12359 8070
rect 12423 8006 12440 8070
rect 12504 8006 12521 8070
rect 12585 8006 12602 8070
rect 12666 8006 12683 8070
rect 12747 8006 12764 8070
rect 12828 8006 12845 8070
rect 12909 8006 12926 8070
rect 12990 8006 13007 8070
rect 13071 8006 13088 8070
rect 13152 8006 13169 8070
rect 13233 8006 13250 8070
rect 13314 8006 13331 8070
rect 13395 8006 13412 8070
rect 13476 8006 13493 8070
rect 13557 8006 13574 8070
rect 13638 8006 13655 8070
rect 13719 8006 13736 8070
rect 13800 8006 13817 8070
rect 13881 8006 13898 8070
rect 13962 8006 13979 8070
rect 14043 8006 14060 8070
rect 14124 8006 14141 8070
rect 14205 8006 14222 8070
rect 14286 8006 14303 8070
rect 14367 8006 14384 8070
rect 14448 8006 14465 8070
rect 14529 8006 14546 8070
rect 14610 8006 14627 8070
rect 14691 8006 14708 8070
rect 14772 8006 14789 8070
rect 14853 8006 14870 8070
rect 14934 8006 15000 8070
rect 0 7984 15000 8006
rect 0 7920 106 7984
rect 170 7920 187 7984
rect 251 7920 268 7984
rect 332 7920 349 7984
rect 413 7920 430 7984
rect 494 7920 510 7984
rect 574 7920 590 7984
rect 654 7920 670 7984
rect 734 7920 750 7984
rect 814 7920 830 7984
rect 894 7920 910 7984
rect 974 7920 990 7984
rect 1054 7920 1070 7984
rect 1134 7920 1150 7984
rect 1214 7920 1230 7984
rect 1294 7920 1310 7984
rect 1374 7920 1390 7984
rect 1454 7920 1470 7984
rect 1534 7920 1550 7984
rect 1614 7920 1630 7984
rect 1694 7920 1710 7984
rect 1774 7920 1790 7984
rect 1854 7920 1870 7984
rect 1934 7920 1950 7984
rect 2014 7920 2030 7984
rect 2094 7920 2110 7984
rect 2174 7920 2190 7984
rect 2254 7920 2270 7984
rect 2334 7920 2350 7984
rect 2414 7920 2430 7984
rect 2494 7920 2510 7984
rect 2574 7920 2590 7984
rect 2654 7920 2670 7984
rect 2734 7920 2750 7984
rect 2814 7920 2830 7984
rect 2894 7920 2910 7984
rect 2974 7920 2990 7984
rect 3054 7920 3070 7984
rect 3134 7920 3150 7984
rect 3214 7920 3230 7984
rect 3294 7920 3310 7984
rect 3374 7920 3390 7984
rect 3454 7920 3470 7984
rect 3534 7920 3550 7984
rect 3614 7920 3630 7984
rect 3694 7920 3710 7984
rect 3774 7920 3790 7984
rect 3854 7920 3870 7984
rect 3934 7920 3950 7984
rect 4014 7920 4030 7984
rect 4094 7920 4110 7984
rect 4174 7920 4190 7984
rect 4254 7920 4270 7984
rect 4334 7920 4350 7984
rect 4414 7920 4430 7984
rect 4494 7920 4510 7984
rect 4574 7920 4590 7984
rect 4654 7920 4670 7984
rect 4734 7920 4750 7984
rect 4814 7920 4830 7984
rect 4894 7920 10157 7984
rect 10221 7920 10239 7984
rect 10303 7920 10321 7984
rect 10385 7920 10403 7984
rect 10467 7920 10485 7984
rect 10549 7920 10567 7984
rect 10631 7920 10649 7984
rect 10713 7920 10731 7984
rect 10795 7920 10813 7984
rect 10877 7920 10895 7984
rect 10959 7920 10977 7984
rect 11041 7920 11059 7984
rect 11123 7920 11141 7984
rect 11205 7920 11223 7984
rect 11287 7920 11305 7984
rect 11369 7920 11387 7984
rect 11451 7920 11468 7984
rect 11532 7920 11549 7984
rect 11613 7920 11630 7984
rect 11694 7920 11711 7984
rect 11775 7920 11792 7984
rect 11856 7920 11873 7984
rect 11937 7920 11954 7984
rect 12018 7920 12035 7984
rect 12099 7920 12116 7984
rect 12180 7920 12197 7984
rect 12261 7920 12278 7984
rect 12342 7920 12359 7984
rect 12423 7920 12440 7984
rect 12504 7920 12521 7984
rect 12585 7920 12602 7984
rect 12666 7920 12683 7984
rect 12747 7920 12764 7984
rect 12828 7920 12845 7984
rect 12909 7920 12926 7984
rect 12990 7920 13007 7984
rect 13071 7920 13088 7984
rect 13152 7920 13169 7984
rect 13233 7920 13250 7984
rect 13314 7920 13331 7984
rect 13395 7920 13412 7984
rect 13476 7920 13493 7984
rect 13557 7920 13574 7984
rect 13638 7920 13655 7984
rect 13719 7920 13736 7984
rect 13800 7920 13817 7984
rect 13881 7920 13898 7984
rect 13962 7920 13979 7984
rect 14043 7920 14060 7984
rect 14124 7920 14141 7984
rect 14205 7920 14222 7984
rect 14286 7920 14303 7984
rect 14367 7920 14384 7984
rect 14448 7920 14465 7984
rect 14529 7920 14546 7984
rect 14610 7920 14627 7984
rect 14691 7920 14708 7984
rect 14772 7920 14789 7984
rect 14853 7920 14870 7984
rect 14934 7920 15000 7984
rect 0 7 15000 7920
<< metal5 >>
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14807 2607 15000 3257
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 0 18917 15000 39600
rect 0 8827 14426 18917
rect 0 6967 15000 8827
rect 0 4467 14426 6967
rect 0 3577 15000 4467
rect 0 2607 14487 3577
rect 0 27 14426 2607
<< labels >>
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 3 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 106 7920 170 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 7920 170 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8006 170 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8006 170 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8092 170 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8092 170 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8178 170 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8178 170 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8264 170 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8264 170 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8350 170 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8350 170 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8436 170 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8436 170 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8522 170 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8522 170 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8608 170 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8608 170 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8694 170 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8694 170 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 106 8780 170 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 106 8780 170 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 7920 251 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 7920 251 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8006 251 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8006 251 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8092 251 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8092 251 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8178 251 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8178 251 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8264 251 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8264 251 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8350 251 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8350 251 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8436 251 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8436 251 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8522 251 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8522 251 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8608 251 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8608 251 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8694 251 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8694 251 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 187 8780 251 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 187 8780 251 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 7920 332 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 7920 332 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8006 332 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8006 332 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8092 332 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8092 332 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8178 332 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8178 332 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8264 332 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8264 332 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8350 332 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8350 332 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8436 332 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8436 332 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8522 332 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8522 332 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8608 332 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8608 332 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8694 332 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8694 332 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 268 8780 332 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 268 8780 332 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 7920 413 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 7920 413 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8006 413 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8006 413 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8092 413 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8092 413 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8178 413 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8178 413 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8264 413 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8264 413 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8350 413 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8350 413 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8436 413 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8436 413 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8522 413 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8522 413 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8608 413 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8608 413 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8694 413 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8694 413 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 349 8780 413 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 349 8780 413 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 7920 2094 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 7920 2094 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8006 2094 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8006 2094 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8092 2094 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8092 2094 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8178 2094 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8178 2094 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8264 2094 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8264 2094 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8350 2094 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8350 2094 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8436 2094 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8436 2094 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8522 2094 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8522 2094 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8608 2094 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8608 2094 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8694 2094 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8694 2094 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2030 8780 2094 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2030 8780 2094 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 7920 2174 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 7920 2174 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8006 2174 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8006 2174 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8092 2174 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8092 2174 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8178 2174 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8178 2174 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8264 2174 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8264 2174 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8350 2174 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8350 2174 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8436 2174 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8436 2174 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8522 2174 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8522 2174 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8608 2174 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8608 2174 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8694 2174 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8694 2174 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2110 8780 2174 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2110 8780 2174 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 7920 2254 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 7920 2254 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8006 2254 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8006 2254 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8092 2254 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8092 2254 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8178 2254 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8178 2254 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8264 2254 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8264 2254 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8350 2254 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8350 2254 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8436 2254 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8436 2254 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8522 2254 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8522 2254 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8608 2254 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8608 2254 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8694 2254 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8694 2254 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2190 8780 2254 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2190 8780 2254 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 7920 2334 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 7920 2334 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8006 2334 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8006 2334 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8092 2334 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8092 2334 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8178 2334 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8178 2334 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8264 2334 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8264 2334 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8350 2334 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8350 2334 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8436 2334 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8436 2334 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8522 2334 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8522 2334 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8608 2334 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8608 2334 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8694 2334 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8694 2334 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2270 8780 2334 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2270 8780 2334 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 7920 2414 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 7920 2414 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8006 2414 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8006 2414 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8092 2414 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8092 2414 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8178 2414 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8178 2414 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8264 2414 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8264 2414 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8350 2414 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8350 2414 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8436 2414 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8436 2414 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8522 2414 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8522 2414 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8608 2414 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8608 2414 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8694 2414 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8694 2414 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2350 8780 2414 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2350 8780 2414 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 7920 2494 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 7920 2494 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8006 2494 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8006 2494 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8092 2494 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8092 2494 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8178 2494 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8178 2494 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8264 2494 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8264 2494 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8350 2494 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8350 2494 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8436 2494 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8436 2494 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8522 2494 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8522 2494 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8608 2494 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8608 2494 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8694 2494 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8694 2494 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2430 8780 2494 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2430 8780 2494 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 7920 2574 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 7920 2574 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8006 2574 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8006 2574 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8092 2574 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8092 2574 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8178 2574 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8178 2574 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8264 2574 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8264 2574 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8350 2574 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8350 2574 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8436 2574 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8436 2574 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8522 2574 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8522 2574 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8608 2574 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8608 2574 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8694 2574 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8694 2574 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2510 8780 2574 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2510 8780 2574 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 7920 2654 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 7920 2654 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8006 2654 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8006 2654 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8092 2654 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8092 2654 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8178 2654 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8178 2654 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8264 2654 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8264 2654 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8350 2654 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8350 2654 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8436 2654 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8436 2654 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8522 2654 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8522 2654 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8608 2654 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8608 2654 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8694 2654 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8694 2654 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2590 8780 2654 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2590 8780 2654 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 7920 2734 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 7920 2734 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8006 2734 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8006 2734 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8092 2734 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8092 2734 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8178 2734 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8178 2734 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8264 2734 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8264 2734 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8350 2734 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8350 2734 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8436 2734 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8436 2734 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8522 2734 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8522 2734 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8608 2734 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8608 2734 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8694 2734 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8694 2734 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2670 8780 2734 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2670 8780 2734 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 7920 2814 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 7920 2814 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8006 2814 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8006 2814 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8092 2814 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8092 2814 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8178 2814 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8178 2814 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8264 2814 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8264 2814 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8350 2814 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8350 2814 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8436 2814 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8436 2814 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8522 2814 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8522 2814 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8608 2814 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8608 2814 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8694 2814 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8694 2814 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2750 8780 2814 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2750 8780 2814 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 7920 2894 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 7920 2894 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8006 2894 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8006 2894 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8092 2894 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8092 2894 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8178 2894 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8178 2894 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8264 2894 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8264 2894 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8350 2894 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8350 2894 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8436 2894 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8436 2894 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8522 2894 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8522 2894 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8608 2894 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8608 2894 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8694 2894 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8694 2894 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2830 8780 2894 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2830 8780 2894 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 7920 2974 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 7920 2974 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8006 2974 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8006 2974 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8092 2974 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8092 2974 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8178 2974 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8178 2974 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8264 2974 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8264 2974 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8350 2974 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8350 2974 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8436 2974 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8436 2974 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8522 2974 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8522 2974 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8608 2974 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8608 2974 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8694 2974 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8694 2974 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2910 8780 2974 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2910 8780 2974 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 7920 3054 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 7920 3054 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8006 3054 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8006 3054 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8092 3054 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8092 3054 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8178 3054 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8178 3054 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8264 3054 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8264 3054 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8350 3054 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8350 3054 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8436 3054 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8436 3054 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8522 3054 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8522 3054 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8608 3054 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8608 3054 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8694 3054 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8694 3054 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 2990 8780 3054 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 2990 8780 3054 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 7920 3134 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 7920 3134 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8006 3134 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8006 3134 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8092 3134 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8092 3134 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8178 3134 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8178 3134 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8264 3134 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8264 3134 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8350 3134 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8350 3134 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8436 3134 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8436 3134 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8522 3134 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8522 3134 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8608 3134 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8608 3134 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8694 3134 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8694 3134 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3070 8780 3134 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3070 8780 3134 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 7920 3214 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 7920 3214 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8006 3214 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8006 3214 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8092 3214 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8092 3214 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8178 3214 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8178 3214 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8264 3214 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8264 3214 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8350 3214 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8350 3214 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8436 3214 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8436 3214 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8522 3214 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8522 3214 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8608 3214 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8608 3214 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8694 3214 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8694 3214 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3150 8780 3214 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3150 8780 3214 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 7920 3294 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 7920 3294 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8006 3294 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8006 3294 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8092 3294 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8092 3294 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8178 3294 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8178 3294 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8264 3294 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8264 3294 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8350 3294 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8350 3294 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8436 3294 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8436 3294 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8522 3294 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8522 3294 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8608 3294 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8608 3294 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8694 3294 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8694 3294 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3230 8780 3294 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3230 8780 3294 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 7920 3374 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 7920 3374 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8006 3374 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8006 3374 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8092 3374 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8092 3374 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8178 3374 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8178 3374 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8264 3374 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8264 3374 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8350 3374 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8350 3374 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8436 3374 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8436 3374 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8522 3374 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8522 3374 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8608 3374 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8608 3374 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8694 3374 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8694 3374 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3310 8780 3374 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3310 8780 3374 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 7920 3454 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 7920 3454 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8006 3454 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8006 3454 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8092 3454 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8092 3454 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8178 3454 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8178 3454 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8264 3454 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8264 3454 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8350 3454 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8350 3454 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8436 3454 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8436 3454 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8522 3454 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8522 3454 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8608 3454 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8608 3454 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8694 3454 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8694 3454 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3390 8780 3454 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3390 8780 3454 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 7920 3534 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 7920 3534 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8006 3534 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8006 3534 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8092 3534 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8092 3534 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8178 3534 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8178 3534 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8264 3534 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8264 3534 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8350 3534 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8350 3534 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8436 3534 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8436 3534 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8522 3534 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8522 3534 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8608 3534 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8608 3534 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8694 3534 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8694 3534 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3470 8780 3534 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3470 8780 3534 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 7920 3614 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 7920 3614 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8006 3614 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8006 3614 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8092 3614 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8092 3614 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8178 3614 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8178 3614 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8264 3614 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8264 3614 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8350 3614 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8350 3614 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8436 3614 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8436 3614 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8522 3614 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8522 3614 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8608 3614 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8608 3614 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8694 3614 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8694 3614 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3550 8780 3614 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3550 8780 3614 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 7920 3694 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 7920 3694 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8006 3694 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8006 3694 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8092 3694 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8092 3694 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8178 3694 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8178 3694 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8264 3694 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8264 3694 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8350 3694 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8350 3694 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8436 3694 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8436 3694 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8522 3694 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8522 3694 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8608 3694 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8608 3694 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8694 3694 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8694 3694 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3630 8780 3694 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3630 8780 3694 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 7920 3774 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 7920 3774 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8006 3774 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8006 3774 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8092 3774 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8092 3774 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8178 3774 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8178 3774 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8264 3774 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8264 3774 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8350 3774 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8350 3774 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8436 3774 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8436 3774 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8522 3774 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8522 3774 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8608 3774 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8608 3774 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8694 3774 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8694 3774 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3710 8780 3774 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3710 8780 3774 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 7920 3854 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 7920 3854 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8006 3854 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8006 3854 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8092 3854 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8092 3854 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8178 3854 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8178 3854 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8264 3854 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8264 3854 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8350 3854 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8350 3854 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8436 3854 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8436 3854 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8522 3854 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8522 3854 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8608 3854 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8608 3854 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8694 3854 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8694 3854 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3790 8780 3854 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3790 8780 3854 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 7920 3934 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 7920 3934 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8006 3934 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8006 3934 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8092 3934 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8092 3934 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8178 3934 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8178 3934 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8264 3934 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8264 3934 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8350 3934 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8350 3934 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8436 3934 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8436 3934 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8522 3934 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8522 3934 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8608 3934 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8608 3934 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8694 3934 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8694 3934 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3870 8780 3934 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3870 8780 3934 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 7920 4014 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 7920 4014 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8006 4014 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8006 4014 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8092 4014 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8092 4014 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8178 4014 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8178 4014 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8264 4014 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8264 4014 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8350 4014 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8350 4014 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8436 4014 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8436 4014 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8522 4014 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8522 4014 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8608 4014 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8608 4014 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8694 4014 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8694 4014 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 3950 8780 4014 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 3950 8780 4014 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 7920 494 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 7920 494 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8006 494 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8006 494 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8092 494 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8092 494 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8178 494 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8178 494 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8264 494 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8264 494 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8350 494 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8350 494 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8436 494 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8436 494 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8522 494 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8522 494 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8608 494 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8608 494 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8694 494 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8694 494 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 430 8780 494 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 430 8780 494 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 7920 574 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 7920 574 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8006 574 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8006 574 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8092 574 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8092 574 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8178 574 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8178 574 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8264 574 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8264 574 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8350 574 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8350 574 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8436 574 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8436 574 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8522 574 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8522 574 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8608 574 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8608 574 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8694 574 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8694 574 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 510 8780 574 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 510 8780 574 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 7920 654 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 7920 654 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8006 654 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8006 654 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8092 654 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8092 654 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8178 654 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8178 654 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8264 654 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8264 654 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8350 654 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8350 654 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8436 654 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8436 654 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8522 654 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8522 654 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8608 654 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8608 654 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8694 654 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8694 654 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 590 8780 654 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 590 8780 654 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 7920 4094 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 7920 4094 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8006 4094 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8006 4094 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8092 4094 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8092 4094 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8178 4094 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8178 4094 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8264 4094 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8264 4094 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8350 4094 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8350 4094 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8436 4094 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8436 4094 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8522 4094 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8522 4094 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8608 4094 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8608 4094 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8694 4094 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8694 4094 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4030 8780 4094 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4030 8780 4094 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 7920 4174 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 7920 4174 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8006 4174 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8006 4174 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8092 4174 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8092 4174 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8178 4174 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8178 4174 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8264 4174 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8264 4174 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8350 4174 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8350 4174 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8436 4174 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8436 4174 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8522 4174 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8522 4174 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8608 4174 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8608 4174 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8694 4174 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8694 4174 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4110 8780 4174 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4110 8780 4174 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 7920 4254 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 7920 4254 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8006 4254 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8006 4254 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8092 4254 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8092 4254 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8178 4254 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8178 4254 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8264 4254 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8264 4254 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8350 4254 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8350 4254 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8436 4254 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8436 4254 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8522 4254 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8522 4254 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8608 4254 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8608 4254 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8694 4254 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8694 4254 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4190 8780 4254 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4190 8780 4254 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 7920 4334 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 7920 4334 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8006 4334 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8006 4334 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8092 4334 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8092 4334 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8178 4334 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8178 4334 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8264 4334 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8264 4334 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8350 4334 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8350 4334 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8436 4334 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8436 4334 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8522 4334 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8522 4334 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8608 4334 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8608 4334 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8694 4334 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8694 4334 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4270 8780 4334 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4270 8780 4334 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 7920 4414 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 7920 4414 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8006 4414 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8006 4414 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8092 4414 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8092 4414 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8178 4414 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8178 4414 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8264 4414 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8264 4414 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8350 4414 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8350 4414 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8436 4414 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8436 4414 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8522 4414 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8522 4414 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8608 4414 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8608 4414 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8694 4414 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8694 4414 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4350 8780 4414 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4350 8780 4414 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 7920 4494 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 7920 4494 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8006 4494 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8006 4494 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8092 4494 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8092 4494 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8178 4494 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8178 4494 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8264 4494 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8264 4494 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8350 4494 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8350 4494 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8436 4494 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8436 4494 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8522 4494 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8522 4494 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8608 4494 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8608 4494 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8694 4494 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8694 4494 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4430 8780 4494 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4430 8780 4494 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 7920 4574 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 7920 4574 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8006 4574 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8006 4574 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8092 4574 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8092 4574 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8178 4574 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8178 4574 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8264 4574 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8264 4574 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8350 4574 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8350 4574 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8436 4574 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8436 4574 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8522 4574 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8522 4574 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8608 4574 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8608 4574 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8694 4574 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8694 4574 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4510 8780 4574 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4510 8780 4574 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 7920 4654 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 7920 4654 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8006 4654 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8006 4654 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8092 4654 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8092 4654 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8178 4654 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8178 4654 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8264 4654 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8264 4654 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8350 4654 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8350 4654 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8436 4654 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8436 4654 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8522 4654 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8522 4654 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8608 4654 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8608 4654 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8694 4654 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8694 4654 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4590 8780 4654 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4590 8780 4654 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 7920 4734 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 7920 4734 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8006 4734 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8006 4734 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8092 4734 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8092 4734 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8178 4734 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8178 4734 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8264 4734 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8264 4734 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8350 4734 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8350 4734 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8436 4734 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8436 4734 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8522 4734 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8522 4734 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8608 4734 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8608 4734 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8694 4734 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8694 4734 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4670 8780 4734 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4670 8780 4734 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 7920 4814 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 7920 4814 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8006 4814 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8006 4814 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8092 4814 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8092 4814 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8178 4814 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8178 4814 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8264 4814 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8264 4814 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8350 4814 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8350 4814 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8436 4814 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8436 4814 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8522 4814 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8522 4814 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8608 4814 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8608 4814 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8694 4814 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8694 4814 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4750 8780 4814 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4750 8780 4814 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 7920 4894 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 7920 4894 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8006 4894 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8006 4894 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8092 4894 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8092 4894 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8178 4894 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8178 4894 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8264 4894 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8264 4894 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8350 4894 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8350 4894 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8436 4894 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8436 4894 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8522 4894 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8522 4894 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8608 4894 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8608 4894 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8694 4894 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8694 4894 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 4830 8780 4894 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 4830 8780 4894 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 7920 734 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 7920 734 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8006 734 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8006 734 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8092 734 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8092 734 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8178 734 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8178 734 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8264 734 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8264 734 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8350 734 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8350 734 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8436 734 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8436 734 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8522 734 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8522 734 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8608 734 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8608 734 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8694 734 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8694 734 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 670 8780 734 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 670 8780 734 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 7920 814 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 7920 814 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8006 814 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8006 814 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8092 814 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8092 814 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8178 814 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8178 814 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8264 814 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8264 814 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8350 814 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8350 814 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8436 814 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8436 814 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8522 814 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8522 814 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8608 814 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8608 814 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8694 814 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8694 814 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 750 8780 814 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 750 8780 814 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 7920 894 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 7920 894 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8006 894 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8006 894 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8092 894 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8092 894 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8178 894 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8178 894 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8264 894 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8264 894 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8350 894 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8350 894 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8436 894 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8436 894 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8522 894 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8522 894 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8608 894 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8608 894 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8694 894 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8694 894 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 830 8780 894 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 830 8780 894 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 7920 974 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 7920 974 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8006 974 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8006 974 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8092 974 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8092 974 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8178 974 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8178 974 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8264 974 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8264 974 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8350 974 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8350 974 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8436 974 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8436 974 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8522 974 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8522 974 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8608 974 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8608 974 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8694 974 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8694 974 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 910 8780 974 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 910 8780 974 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 7920 1054 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 7920 1054 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8006 1054 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8006 1054 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8092 1054 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8092 1054 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8178 1054 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8178 1054 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8264 1054 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8264 1054 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8350 1054 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8350 1054 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8436 1054 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8436 1054 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8522 1054 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8522 1054 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8608 1054 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8608 1054 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8694 1054 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8694 1054 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 990 8780 1054 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 990 8780 1054 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 7920 1134 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 7920 1134 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8006 1134 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8006 1134 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8092 1134 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8092 1134 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8178 1134 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8178 1134 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8264 1134 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8264 1134 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8350 1134 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8350 1134 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8436 1134 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8436 1134 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8522 1134 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8522 1134 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8608 1134 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8608 1134 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8694 1134 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8694 1134 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1070 8780 1134 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1070 8780 1134 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 7920 1214 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 7920 1214 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8006 1214 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8006 1214 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8092 1214 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8092 1214 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8178 1214 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8178 1214 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8264 1214 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8264 1214 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8350 1214 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8350 1214 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8436 1214 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8436 1214 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8522 1214 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8522 1214 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8608 1214 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8608 1214 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8694 1214 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8694 1214 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1150 8780 1214 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1150 8780 1214 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 7920 10221 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 7920 10221 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8006 10221 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8006 10221 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8092 10221 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8092 10221 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8178 10221 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8178 10221 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8264 10221 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8264 10221 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8350 10221 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8350 10221 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8436 10221 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8436 10221 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8522 10221 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8522 10221 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8608 10221 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8608 10221 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8694 10221 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8694 10221 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10157 8780 10221 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10157 8780 10221 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 7920 10303 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 7920 10303 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8006 10303 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8006 10303 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8092 10303 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8092 10303 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8178 10303 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8178 10303 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8264 10303 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8264 10303 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8350 10303 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8350 10303 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8436 10303 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8436 10303 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8522 10303 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8522 10303 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8608 10303 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8608 10303 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8694 10303 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8694 10303 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10239 8780 10303 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10239 8780 10303 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 7920 10385 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 7920 10385 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8006 10385 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8006 10385 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8092 10385 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8092 10385 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8178 10385 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8178 10385 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8264 10385 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8264 10385 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8350 10385 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8350 10385 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8436 10385 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8436 10385 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8522 10385 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8522 10385 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8608 10385 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8608 10385 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8694 10385 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8694 10385 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10321 8780 10385 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10321 8780 10385 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 7920 10467 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 7920 10467 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8006 10467 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8006 10467 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8092 10467 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8092 10467 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8178 10467 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8178 10467 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8264 10467 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8264 10467 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8350 10467 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8350 10467 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8436 10467 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8436 10467 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8522 10467 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8522 10467 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8608 10467 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8608 10467 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8694 10467 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8694 10467 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10403 8780 10467 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10403 8780 10467 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 7920 10549 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 7920 10549 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8006 10549 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8006 10549 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8092 10549 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8092 10549 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8178 10549 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8178 10549 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8264 10549 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8264 10549 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8350 10549 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8350 10549 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8436 10549 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8436 10549 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8522 10549 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8522 10549 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8608 10549 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8608 10549 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8694 10549 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8694 10549 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10485 8780 10549 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10485 8780 10549 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 7920 10631 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 7920 10631 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8006 10631 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8006 10631 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8092 10631 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8092 10631 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8178 10631 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8178 10631 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8264 10631 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8264 10631 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8350 10631 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8350 10631 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8436 10631 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8436 10631 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8522 10631 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8522 10631 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8608 10631 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8608 10631 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8694 10631 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8694 10631 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10567 8780 10631 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10567 8780 10631 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 7920 10713 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 7920 10713 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8006 10713 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8006 10713 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8092 10713 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8092 10713 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8178 10713 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8178 10713 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8264 10713 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8264 10713 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8350 10713 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8350 10713 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8436 10713 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8436 10713 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8522 10713 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8522 10713 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8608 10713 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8608 10713 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8694 10713 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8694 10713 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10649 8780 10713 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10649 8780 10713 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 7920 10795 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 7920 10795 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8006 10795 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8006 10795 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8092 10795 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8092 10795 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8178 10795 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8178 10795 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8264 10795 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8264 10795 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8350 10795 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8350 10795 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8436 10795 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8436 10795 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8522 10795 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8522 10795 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8608 10795 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8608 10795 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8694 10795 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8694 10795 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10731 8780 10795 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10731 8780 10795 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 7920 10877 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 7920 10877 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8006 10877 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8006 10877 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8092 10877 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8092 10877 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8178 10877 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8178 10877 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8264 10877 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8264 10877 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8350 10877 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8350 10877 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8436 10877 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8436 10877 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8522 10877 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8522 10877 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8608 10877 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8608 10877 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8694 10877 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8694 10877 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10813 8780 10877 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10813 8780 10877 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 7920 10959 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 7920 10959 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8006 10959 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8006 10959 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8092 10959 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8092 10959 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8178 10959 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8178 10959 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8264 10959 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8264 10959 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8350 10959 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8350 10959 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8436 10959 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8436 10959 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8522 10959 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8522 10959 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8608 10959 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8608 10959 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8694 10959 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8694 10959 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10895 8780 10959 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10895 8780 10959 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 7920 11041 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 7920 11041 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8006 11041 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8006 11041 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8092 11041 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8092 11041 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8178 11041 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8178 11041 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8264 11041 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8264 11041 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8350 11041 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8350 11041 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8436 11041 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8436 11041 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8522 11041 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8522 11041 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8608 11041 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8608 11041 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8694 11041 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8694 11041 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 10977 8780 11041 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10977 8780 11041 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 7920 11123 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 7920 11123 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8006 11123 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8006 11123 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8092 11123 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8092 11123 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8178 11123 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8178 11123 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8264 11123 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8264 11123 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8350 11123 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8350 11123 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8436 11123 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8436 11123 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8522 11123 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8522 11123 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8608 11123 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8608 11123 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8694 11123 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8694 11123 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11059 8780 11123 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11059 8780 11123 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 7920 11205 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 7920 11205 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8006 11205 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8006 11205 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8092 11205 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8092 11205 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8178 11205 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8178 11205 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8264 11205 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8264 11205 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8350 11205 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8350 11205 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8436 11205 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8436 11205 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8522 11205 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8522 11205 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8608 11205 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8608 11205 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8694 11205 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8694 11205 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11141 8780 11205 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11141 8780 11205 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 7920 11287 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 7920 11287 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8006 11287 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8006 11287 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8092 11287 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8092 11287 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8178 11287 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8178 11287 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8264 11287 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8264 11287 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8350 11287 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8350 11287 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8436 11287 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8436 11287 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8522 11287 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8522 11287 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8608 11287 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8608 11287 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8694 11287 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8694 11287 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11223 8780 11287 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11223 8780 11287 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 7920 11369 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 7920 11369 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8006 11369 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8006 11369 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8092 11369 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8092 11369 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8178 11369 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8178 11369 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8264 11369 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8264 11369 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8350 11369 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8350 11369 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8436 11369 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8436 11369 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8522 11369 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8522 11369 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8608 11369 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8608 11369 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8694 11369 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8694 11369 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11305 8780 11369 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11305 8780 11369 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 7920 11451 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 7920 11451 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8006 11451 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8006 11451 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8092 11451 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8092 11451 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8178 11451 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8178 11451 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8264 11451 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8264 11451 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8350 11451 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8350 11451 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8436 11451 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8436 11451 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8522 11451 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8522 11451 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8608 11451 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8608 11451 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8694 11451 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8694 11451 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11387 8780 11451 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11387 8780 11451 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 7920 11532 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 7920 11532 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8006 11532 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8006 11532 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8092 11532 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8092 11532 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8178 11532 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8178 11532 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8264 11532 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8264 11532 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8350 11532 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8350 11532 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8436 11532 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8436 11532 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8522 11532 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8522 11532 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8608 11532 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8608 11532 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8694 11532 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8694 11532 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11468 8780 11532 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11468 8780 11532 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 7920 11613 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 7920 11613 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8006 11613 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8006 11613 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8092 11613 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8092 11613 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8178 11613 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8178 11613 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8264 11613 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8264 11613 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8350 11613 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8350 11613 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8436 11613 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8436 11613 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8522 11613 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8522 11613 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8608 11613 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8608 11613 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8694 11613 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8694 11613 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11549 8780 11613 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11549 8780 11613 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 7920 11694 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 7920 11694 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8006 11694 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8006 11694 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8092 11694 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8092 11694 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8178 11694 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8178 11694 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8264 11694 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8264 11694 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8350 11694 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8350 11694 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8436 11694 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8436 11694 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8522 11694 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8522 11694 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8608 11694 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8608 11694 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8694 11694 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8694 11694 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11630 8780 11694 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11630 8780 11694 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 7920 11775 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 7920 11775 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8006 11775 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8006 11775 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8092 11775 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8092 11775 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8178 11775 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8178 11775 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8264 11775 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8264 11775 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8350 11775 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8350 11775 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8436 11775 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8436 11775 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8522 11775 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8522 11775 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8608 11775 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8608 11775 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8694 11775 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8694 11775 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11711 8780 11775 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11711 8780 11775 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 7920 11856 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 7920 11856 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8006 11856 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8006 11856 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8092 11856 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8092 11856 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8178 11856 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8178 11856 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8264 11856 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8264 11856 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8350 11856 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8350 11856 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8436 11856 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8436 11856 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8522 11856 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8522 11856 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8608 11856 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8608 11856 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8694 11856 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8694 11856 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11792 8780 11856 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11792 8780 11856 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 7920 11937 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 7920 11937 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8006 11937 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8006 11937 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8092 11937 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8092 11937 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8178 11937 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8178 11937 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8264 11937 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8264 11937 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8350 11937 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8350 11937 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8436 11937 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8436 11937 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8522 11937 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8522 11937 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8608 11937 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8608 11937 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8694 11937 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8694 11937 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11873 8780 11937 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11873 8780 11937 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 7920 12018 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 7920 12018 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8006 12018 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8006 12018 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8092 12018 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8092 12018 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8178 12018 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8178 12018 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8264 12018 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8264 12018 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8350 12018 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8350 12018 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8436 12018 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8436 12018 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8522 12018 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8522 12018 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8608 12018 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8608 12018 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8694 12018 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8694 12018 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 11954 8780 12018 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 11954 8780 12018 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 7920 1294 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 7920 1294 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8006 1294 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8006 1294 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8092 1294 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8092 1294 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8178 1294 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8178 1294 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8264 1294 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8264 1294 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8350 1294 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8350 1294 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8436 1294 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8436 1294 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8522 1294 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8522 1294 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8608 1294 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8608 1294 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8694 1294 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8694 1294 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1230 8780 1294 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1230 8780 1294 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 7920 1374 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 7920 1374 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8006 1374 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8006 1374 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8092 1374 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8092 1374 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8178 1374 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8178 1374 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8264 1374 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8264 1374 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8350 1374 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8350 1374 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8436 1374 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8436 1374 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8522 1374 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8522 1374 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8608 1374 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8608 1374 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8694 1374 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8694 1374 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1310 8780 1374 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1310 8780 1374 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 7920 1454 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 7920 1454 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8006 1454 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8006 1454 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8092 1454 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8092 1454 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8178 1454 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8178 1454 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8264 1454 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8264 1454 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8350 1454 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8350 1454 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8436 1454 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8436 1454 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8522 1454 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8522 1454 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8608 1454 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8608 1454 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8694 1454 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8694 1454 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1390 8780 1454 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1390 8780 1454 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 7920 12099 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 7920 12099 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8006 12099 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8006 12099 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8092 12099 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8092 12099 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8178 12099 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8178 12099 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8264 12099 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8264 12099 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8350 12099 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8350 12099 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8436 12099 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8436 12099 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8522 12099 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8522 12099 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8608 12099 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8608 12099 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8694 12099 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8694 12099 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12035 8780 12099 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12035 8780 12099 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 7920 12180 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 7920 12180 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8006 12180 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8006 12180 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8092 12180 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8092 12180 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8178 12180 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8178 12180 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8264 12180 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8264 12180 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8350 12180 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8350 12180 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8436 12180 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8436 12180 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8522 12180 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8522 12180 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8608 12180 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8608 12180 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8694 12180 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8694 12180 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12116 8780 12180 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12116 8780 12180 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 7920 12261 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 7920 12261 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8006 12261 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8006 12261 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8092 12261 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8092 12261 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8178 12261 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8178 12261 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8264 12261 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8264 12261 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8350 12261 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8350 12261 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8436 12261 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8436 12261 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8522 12261 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8522 12261 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8608 12261 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8608 12261 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8694 12261 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8694 12261 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12197 8780 12261 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12197 8780 12261 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 7920 12342 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 7920 12342 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8006 12342 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8006 12342 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8092 12342 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8092 12342 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8178 12342 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8178 12342 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8264 12342 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8264 12342 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8350 12342 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8350 12342 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8436 12342 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8436 12342 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8522 12342 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8522 12342 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8608 12342 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8608 12342 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8694 12342 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8694 12342 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12278 8780 12342 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12278 8780 12342 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 7920 12423 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 7920 12423 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8006 12423 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8006 12423 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8092 12423 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8092 12423 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8178 12423 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8178 12423 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8264 12423 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8264 12423 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8350 12423 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8350 12423 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8436 12423 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8436 12423 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8522 12423 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8522 12423 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8608 12423 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8608 12423 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8694 12423 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8694 12423 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12359 8780 12423 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12359 8780 12423 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 7920 12504 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 7920 12504 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8006 12504 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8006 12504 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8092 12504 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8092 12504 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8178 12504 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8178 12504 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8264 12504 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8264 12504 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8350 12504 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8350 12504 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8436 12504 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8436 12504 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8522 12504 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8522 12504 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8608 12504 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8608 12504 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8694 12504 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8694 12504 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12440 8780 12504 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12440 8780 12504 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 7920 12585 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 7920 12585 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8006 12585 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8006 12585 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8092 12585 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8092 12585 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8178 12585 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8178 12585 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8264 12585 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8264 12585 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8350 12585 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8350 12585 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8436 12585 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8436 12585 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8522 12585 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8522 12585 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8608 12585 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8608 12585 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8694 12585 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8694 12585 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12521 8780 12585 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12521 8780 12585 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 7920 12666 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 7920 12666 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8006 12666 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8006 12666 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8092 12666 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8092 12666 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8178 12666 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8178 12666 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8264 12666 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8264 12666 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8350 12666 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8350 12666 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8436 12666 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8436 12666 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8522 12666 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8522 12666 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8608 12666 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8608 12666 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8694 12666 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8694 12666 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12602 8780 12666 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12602 8780 12666 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 7920 12747 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 7920 12747 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8006 12747 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8006 12747 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8092 12747 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8092 12747 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8178 12747 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8178 12747 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8264 12747 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8264 12747 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8350 12747 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8350 12747 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8436 12747 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8436 12747 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8522 12747 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8522 12747 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8608 12747 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8608 12747 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8694 12747 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8694 12747 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12683 8780 12747 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12683 8780 12747 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 7920 12828 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 7920 12828 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8006 12828 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8006 12828 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8092 12828 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8092 12828 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8178 12828 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8178 12828 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8264 12828 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8264 12828 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8350 12828 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8350 12828 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8436 12828 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8436 12828 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8522 12828 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8522 12828 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8608 12828 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8608 12828 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8694 12828 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8694 12828 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12764 8780 12828 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12764 8780 12828 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 7920 12909 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 7920 12909 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8006 12909 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8006 12909 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8092 12909 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8092 12909 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8178 12909 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8178 12909 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8264 12909 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8264 12909 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8350 12909 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8350 12909 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8436 12909 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8436 12909 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8522 12909 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8522 12909 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8608 12909 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8608 12909 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8694 12909 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8694 12909 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12845 8780 12909 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12845 8780 12909 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 7920 12990 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 7920 12990 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8006 12990 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8006 12990 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8092 12990 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8092 12990 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8178 12990 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8178 12990 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8264 12990 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8264 12990 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8350 12990 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8350 12990 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8436 12990 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8436 12990 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8522 12990 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8522 12990 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8608 12990 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8608 12990 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8694 12990 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8694 12990 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 12926 8780 12990 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 12926 8780 12990 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 7920 13071 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 7920 13071 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8006 13071 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8006 13071 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8092 13071 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8092 13071 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8178 13071 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8178 13071 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8264 13071 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8264 13071 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8350 13071 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8350 13071 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8436 13071 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8436 13071 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8522 13071 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8522 13071 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8608 13071 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8608 13071 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8694 13071 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8694 13071 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13007 8780 13071 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13007 8780 13071 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 7920 13152 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 7920 13152 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8006 13152 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8006 13152 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8092 13152 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8092 13152 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8178 13152 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8178 13152 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8264 13152 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8264 13152 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8350 13152 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8350 13152 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8436 13152 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8436 13152 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8522 13152 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8522 13152 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8608 13152 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8608 13152 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8694 13152 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8694 13152 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13088 8780 13152 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13088 8780 13152 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 7920 13233 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 7920 13233 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8006 13233 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8006 13233 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8092 13233 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8092 13233 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8178 13233 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8178 13233 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8264 13233 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8264 13233 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8350 13233 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8350 13233 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8436 13233 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8436 13233 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8522 13233 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8522 13233 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8608 13233 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8608 13233 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8694 13233 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8694 13233 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13169 8780 13233 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13169 8780 13233 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 7920 13314 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 7920 13314 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8006 13314 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8006 13314 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8092 13314 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8092 13314 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8178 13314 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8178 13314 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8264 13314 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8264 13314 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8350 13314 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8350 13314 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8436 13314 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8436 13314 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8522 13314 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8522 13314 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8608 13314 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8608 13314 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8694 13314 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8694 13314 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13250 8780 13314 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13250 8780 13314 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 7920 13395 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 7920 13395 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8006 13395 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8006 13395 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8092 13395 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8092 13395 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8178 13395 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8178 13395 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8264 13395 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8264 13395 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8350 13395 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8350 13395 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8436 13395 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8436 13395 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8522 13395 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8522 13395 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8608 13395 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8608 13395 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8694 13395 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8694 13395 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13331 8780 13395 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13331 8780 13395 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 7920 13476 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 7920 13476 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8006 13476 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8006 13476 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8092 13476 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8092 13476 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8178 13476 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8178 13476 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8264 13476 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8264 13476 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8350 13476 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8350 13476 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8436 13476 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8436 13476 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8522 13476 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8522 13476 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8608 13476 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8608 13476 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8694 13476 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8694 13476 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13412 8780 13476 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13412 8780 13476 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 7920 13557 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 7920 13557 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8006 13557 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8006 13557 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8092 13557 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8092 13557 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8178 13557 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8178 13557 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8264 13557 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8264 13557 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8350 13557 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8350 13557 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8436 13557 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8436 13557 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8522 13557 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8522 13557 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8608 13557 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8608 13557 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8694 13557 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8694 13557 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13493 8780 13557 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13493 8780 13557 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 7920 13638 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 7920 13638 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8006 13638 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8006 13638 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8092 13638 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8092 13638 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8178 13638 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8178 13638 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8264 13638 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8264 13638 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8350 13638 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8350 13638 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8436 13638 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8436 13638 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8522 13638 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8522 13638 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8608 13638 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8608 13638 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8694 13638 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8694 13638 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13574 8780 13638 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13574 8780 13638 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 7920 13719 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 7920 13719 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8006 13719 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8006 13719 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8092 13719 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8092 13719 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8178 13719 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8178 13719 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8264 13719 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8264 13719 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8350 13719 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8350 13719 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8436 13719 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8436 13719 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8522 13719 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8522 13719 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8608 13719 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8608 13719 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8694 13719 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8694 13719 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13655 8780 13719 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13655 8780 13719 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 7920 13800 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 7920 13800 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8006 13800 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8006 13800 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8092 13800 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8092 13800 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8178 13800 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8178 13800 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8264 13800 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8264 13800 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8350 13800 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8350 13800 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8436 13800 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8436 13800 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8522 13800 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8522 13800 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8608 13800 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8608 13800 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8694 13800 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8694 13800 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13736 8780 13800 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13736 8780 13800 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 7920 13881 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 7920 13881 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8006 13881 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8006 13881 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8092 13881 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8092 13881 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8178 13881 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8178 13881 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8264 13881 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8264 13881 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8350 13881 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8350 13881 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8436 13881 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8436 13881 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8522 13881 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8522 13881 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8608 13881 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8608 13881 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8694 13881 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8694 13881 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13817 8780 13881 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13817 8780 13881 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 7920 13962 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 7920 13962 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8006 13962 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8006 13962 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8092 13962 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8092 13962 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8178 13962 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8178 13962 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8264 13962 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8264 13962 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8350 13962 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8350 13962 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8436 13962 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8436 13962 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8522 13962 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8522 13962 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8608 13962 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8608 13962 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8694 13962 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8694 13962 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13898 8780 13962 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13898 8780 13962 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 7920 14043 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 7920 14043 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8006 14043 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8006 14043 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8092 14043 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8092 14043 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8178 14043 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8178 14043 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8264 14043 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8264 14043 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8350 14043 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8350 14043 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8436 14043 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8436 14043 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8522 14043 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8522 14043 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8608 14043 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8608 14043 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8694 14043 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8694 14043 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 13979 8780 14043 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 13979 8780 14043 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 7920 1534 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 7920 1534 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8006 1534 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8006 1534 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8092 1534 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8092 1534 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8178 1534 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8178 1534 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8264 1534 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8264 1534 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8350 1534 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8350 1534 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8436 1534 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8436 1534 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8522 1534 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8522 1534 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8608 1534 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8608 1534 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8694 1534 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8694 1534 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1470 8780 1534 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1470 8780 1534 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 7920 1614 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 7920 1614 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8006 1614 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8006 1614 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8092 1614 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8092 1614 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8178 1614 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8178 1614 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8264 1614 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8264 1614 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8350 1614 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8350 1614 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8436 1614 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8436 1614 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8522 1614 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8522 1614 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8608 1614 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8608 1614 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8694 1614 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8694 1614 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1550 8780 1614 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1550 8780 1614 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 7920 14124 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 7920 14124 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8006 14124 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8006 14124 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8092 14124 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8092 14124 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8178 14124 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8178 14124 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8264 14124 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8264 14124 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8350 14124 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8350 14124 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8436 14124 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8436 14124 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8522 14124 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8522 14124 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8608 14124 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8608 14124 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8694 14124 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8694 14124 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14060 8780 14124 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14060 8780 14124 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 7920 14205 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 7920 14205 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8006 14205 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8006 14205 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8092 14205 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8092 14205 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8178 14205 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8178 14205 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8264 14205 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8264 14205 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8350 14205 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8350 14205 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8436 14205 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8436 14205 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8522 14205 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8522 14205 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8608 14205 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8608 14205 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8694 14205 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8694 14205 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14141 8780 14205 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14141 8780 14205 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 7920 14286 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 7920 14286 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8006 14286 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8006 14286 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8092 14286 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8092 14286 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8178 14286 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8178 14286 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8264 14286 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8264 14286 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8350 14286 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8350 14286 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8436 14286 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8436 14286 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8522 14286 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8522 14286 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8608 14286 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8608 14286 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8694 14286 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8694 14286 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14222 8780 14286 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14222 8780 14286 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 7920 14367 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 7920 14367 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8006 14367 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8006 14367 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8092 14367 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8092 14367 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8178 14367 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8178 14367 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8264 14367 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8264 14367 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8350 14367 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8350 14367 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8436 14367 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8436 14367 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8522 14367 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8522 14367 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8608 14367 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8608 14367 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8694 14367 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8694 14367 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14303 8780 14367 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14303 8780 14367 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 7920 14448 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 7920 14448 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8006 14448 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8006 14448 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8092 14448 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8092 14448 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8178 14448 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8178 14448 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8264 14448 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8264 14448 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8350 14448 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8350 14448 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8436 14448 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8436 14448 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8522 14448 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8522 14448 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8608 14448 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8608 14448 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8694 14448 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8694 14448 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14384 8780 14448 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14384 8780 14448 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 7920 14529 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 7920 14529 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8006 14529 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8006 14529 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8092 14529 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8092 14529 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8178 14529 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8178 14529 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8264 14529 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8264 14529 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8350 14529 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8350 14529 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8436 14529 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8436 14529 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8522 14529 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8522 14529 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8608 14529 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8608 14529 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8694 14529 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8694 14529 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14465 8780 14529 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14465 8780 14529 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 7920 14610 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 7920 14610 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8006 14610 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8006 14610 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8092 14610 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8092 14610 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8178 14610 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8178 14610 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8264 14610 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8264 14610 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8350 14610 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8350 14610 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8436 14610 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8436 14610 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8522 14610 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8522 14610 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8608 14610 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8608 14610 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8694 14610 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8694 14610 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14546 8780 14610 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14546 8780 14610 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 7920 14691 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 7920 14691 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8006 14691 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8006 14691 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8092 14691 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8092 14691 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8178 14691 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8178 14691 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8264 14691 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8264 14691 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8350 14691 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8350 14691 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8436 14691 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8436 14691 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8522 14691 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8522 14691 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8608 14691 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8608 14691 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8694 14691 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8694 14691 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14627 8780 14691 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14627 8780 14691 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 7920 14772 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 7920 14772 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8006 14772 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8006 14772 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8092 14772 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8092 14772 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8178 14772 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8178 14772 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8264 14772 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8264 14772 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8350 14772 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8350 14772 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8436 14772 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8436 14772 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8522 14772 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8522 14772 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8608 14772 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8608 14772 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8694 14772 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8694 14772 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14708 8780 14772 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14708 8780 14772 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 7920 14853 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 7920 14853 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8006 14853 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8006 14853 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8092 14853 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8092 14853 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8178 14853 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8178 14853 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8264 14853 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8264 14853 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8350 14853 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8350 14853 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8436 14853 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8436 14853 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8522 14853 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8522 14853 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8608 14853 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8608 14853 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8694 14853 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8694 14853 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14789 8780 14853 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14789 8780 14853 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 7920 14934 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 7920 14934 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8006 14934 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8006 14934 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8092 14934 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8092 14934 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8178 14934 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8178 14934 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8264 14934 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8264 14934 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8350 14934 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8350 14934 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8436 14934 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8436 14934 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8522 14934 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8522 14934 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8608 14934 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8608 14934 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8694 14934 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8694 14934 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 14870 8780 14934 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 14870 8780 14934 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 7920 1694 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 7920 1694 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8006 1694 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8006 1694 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8092 1694 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8092 1694 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8178 1694 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8178 1694 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8264 1694 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8264 1694 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8350 1694 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8350 1694 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8436 1694 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8436 1694 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8522 1694 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8522 1694 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8608 1694 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8608 1694 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8694 1694 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8694 1694 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1630 8780 1694 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1630 8780 1694 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 7920 1774 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 7920 1774 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8006 1774 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8006 1774 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8092 1774 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8092 1774 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8178 1774 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8178 1774 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8264 1774 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8264 1774 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8350 1774 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8350 1774 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8436 1774 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8436 1774 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8522 1774 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8522 1774 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8608 1774 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8608 1774 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8694 1774 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8694 1774 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1710 8780 1774 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1710 8780 1774 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 7920 1854 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 7920 1854 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8006 1854 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8006 1854 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8092 1854 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8092 1854 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8178 1854 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8178 1854 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8264 1854 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8264 1854 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8350 1854 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8350 1854 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8436 1854 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8436 1854 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8522 1854 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8522 1854 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8608 1854 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8608 1854 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8694 1854 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8694 1854 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1790 8780 1854 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1790 8780 1854 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 7920 1934 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 7920 1934 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8006 1934 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8006 1934 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8092 1934 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8092 1934 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8178 1934 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8178 1934 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8264 1934 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8264 1934 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8350 1934 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8350 1934 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8436 1934 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8436 1934 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8522 1934 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8522 1934 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8608 1934 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8608 1934 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8694 1934 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8694 1934 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1870 8780 1934 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1870 8780 1934 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 7920 2014 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 7920 2014 7984 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8006 2014 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8006 2014 8070 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8092 2014 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8092 2014 8156 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8178 2014 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8178 2014 8242 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8264 2014 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8264 2014 8328 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8350 2014 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8350 2014 8414 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8436 2014 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8436 2014 8500 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8522 2014 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8522 2014 8586 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8608 2014 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8608 2014 8672 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8694 2014 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8694 2014 8758 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 1950 8780 2014 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 1950 8780 2014 8844 6 VSSD
port 9 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 39600
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 35319472
string GDS_START 35226960
<< end >>
