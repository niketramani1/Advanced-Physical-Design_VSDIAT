magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1296 -1277 3500 2731
<< nwell >>
rect -36 679 2240 1471
<< locali >>
rect 0 1397 2204 1431
rect 64 674 98 740
rect 1047 690 1081 724
rect 0 -17 2204 17
use pinv_16  pinv_16_0
timestamp 1624857261
transform 1 0 0 0 1 0
box -36 -17 2240 1471
<< labels >>
rlabel locali s 1064 707 1064 707 4 Z
port 2 se
rlabel locali s 81 707 81 707 4 A
port 1 se
rlabel locali s 1102 0 1102 0 4 gnd
port 4 se
rlabel locali s 1102 1414 1102 1414 4 vdd
port 3 se
<< properties >>
string FIXED_BBOX 0 0 2204 1414
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 9213084
string GDS_START 9212286
<< end >>
