magic
tech sky130A
magscale 1 2
timestamp 1624855602
<< nwell >>
rect -66 377 6786 897
<< pwell >>
rect 0 -17 6720 17
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4063 831
rect 4097 797 4159 831
rect 4193 797 4255 831
rect 4289 797 4351 831
rect 4385 797 4447 831
rect 4481 797 4543 831
rect 4577 797 4639 831
rect 4673 797 4735 831
rect 4769 797 4831 831
rect 4865 797 4927 831
rect 4961 797 5023 831
rect 5057 797 5119 831
rect 5153 797 5215 831
rect 5249 797 5311 831
rect 5345 797 5407 831
rect 5441 797 5503 831
rect 5537 797 5599 831
rect 5633 797 5695 831
rect 5729 797 5791 831
rect 5825 797 5887 831
rect 5921 797 5983 831
rect 6017 797 6079 831
rect 6113 797 6175 831
rect 6209 797 6271 831
rect 6305 797 6367 831
rect 6401 797 6463 831
rect 6497 797 6559 831
rect 6593 797 6655 831
rect 6689 797 6720 831
rect 44 316 926 363
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 5023 17
rect 5057 -17 5119 17
rect 5153 -17 5215 17
rect 5249 -17 5311 17
rect 5345 -17 5407 17
rect 5441 -17 5503 17
rect 5537 -17 5599 17
rect 5633 -17 5695 17
rect 5729 -17 5791 17
rect 5825 -17 5887 17
rect 5921 -17 5983 17
rect 6017 -17 6079 17
rect 6113 -17 6175 17
rect 6209 -17 6271 17
rect 6305 -17 6367 17
rect 6401 -17 6463 17
rect 6497 -17 6559 17
rect 6593 -17 6655 17
rect 6689 -17 6720 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
rect 4063 797 4097 831
rect 4159 797 4193 831
rect 4255 797 4289 831
rect 4351 797 4385 831
rect 4447 797 4481 831
rect 4543 797 4577 831
rect 4639 797 4673 831
rect 4735 797 4769 831
rect 4831 797 4865 831
rect 4927 797 4961 831
rect 5023 797 5057 831
rect 5119 797 5153 831
rect 5215 797 5249 831
rect 5311 797 5345 831
rect 5407 797 5441 831
rect 5503 797 5537 831
rect 5599 797 5633 831
rect 5695 797 5729 831
rect 5791 797 5825 831
rect 5887 797 5921 831
rect 5983 797 6017 831
rect 6079 797 6113 831
rect 6175 797 6209 831
rect 6271 797 6305 831
rect 6367 797 6401 831
rect 6463 797 6497 831
rect 6559 797 6593 831
rect 6655 797 6689 831
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
rect 4735 -17 4769 17
rect 4831 -17 4865 17
rect 4927 -17 4961 17
rect 5023 -17 5057 17
rect 5119 -17 5153 17
rect 5215 -17 5249 17
rect 5311 -17 5345 17
rect 5407 -17 5441 17
rect 5503 -17 5537 17
rect 5599 -17 5633 17
rect 5695 -17 5729 17
rect 5791 -17 5825 17
rect 5887 -17 5921 17
rect 5983 -17 6017 17
rect 6079 -17 6113 17
rect 6175 -17 6209 17
rect 6271 -17 6305 17
rect 6367 -17 6401 17
rect 6463 -17 6497 17
rect 6559 -17 6593 17
rect 6655 -17 6689 17
<< obsli1 >>
rect 22 729 136 751
rect 22 695 30 729
rect 64 695 102 729
rect 22 435 136 695
rect 170 453 232 751
rect 268 729 446 735
rect 302 695 340 729
rect 374 695 412 729
rect 268 489 446 695
rect 480 453 542 751
rect 576 729 754 735
rect 610 695 648 729
rect 682 695 720 729
rect 576 489 754 695
rect 788 453 858 751
rect 892 729 1070 735
rect 926 695 964 729
rect 998 695 1036 729
rect 892 489 1070 695
rect 1104 453 1166 751
rect 1200 729 1378 735
rect 1234 695 1272 729
rect 1306 695 1344 729
rect 1200 489 1378 695
rect 1412 453 1482 751
rect 170 397 1482 453
rect 1516 729 1696 735
rect 1550 695 1588 729
rect 1622 695 1660 729
rect 1694 695 1696 729
rect 1516 447 1696 695
rect 1786 498 1852 751
rect 1786 464 1802 498
rect 1836 464 1852 498
rect 960 282 1482 397
rect 22 119 129 282
rect 163 239 1482 282
rect 163 151 234 239
rect 22 85 23 119
rect 57 85 95 119
rect 268 119 446 205
rect 480 146 558 239
rect 302 85 340 119
rect 374 85 412 119
rect 592 119 771 205
rect 805 146 854 239
rect 592 85 664 119
rect 698 85 736 119
rect 770 85 771 119
rect 888 119 1066 205
rect 1104 146 1182 239
rect 888 85 960 119
rect 994 85 1032 119
rect 1216 119 1395 205
rect 1429 146 1478 239
rect 1516 205 1696 279
rect 1216 85 1288 119
rect 1322 85 1360 119
rect 1394 85 1395 119
rect 1512 119 1696 205
rect 1786 158 1852 464
rect 1886 729 2064 751
rect 1920 695 1958 729
rect 1992 695 2030 729
rect 1886 435 2064 695
rect 2098 498 2164 751
rect 2098 464 2114 498
rect 2148 464 2164 498
rect 1904 313 2038 379
rect 1512 85 1584 119
rect 1618 85 1656 119
rect 1690 85 1696 119
rect 1886 119 2064 279
rect 2098 158 2164 464
rect 2198 729 2376 751
rect 2232 695 2270 729
rect 2304 695 2342 729
rect 2198 435 2376 695
rect 2410 498 2476 751
rect 2410 464 2426 498
rect 2460 464 2476 498
rect 2216 313 2350 379
rect 1886 85 1958 119
rect 1992 85 2030 119
rect 2198 119 2376 279
rect 2410 158 2476 464
rect 2510 729 2688 751
rect 2544 695 2582 729
rect 2616 695 2654 729
rect 2510 435 2688 695
rect 2722 498 2788 751
rect 2722 464 2738 498
rect 2772 464 2788 498
rect 2528 313 2662 379
rect 2198 85 2270 119
rect 2304 85 2342 119
rect 2510 119 2688 279
rect 2722 158 2788 464
rect 2822 729 3000 751
rect 2856 695 2894 729
rect 2928 695 2966 729
rect 2822 435 3000 695
rect 3034 498 3100 751
rect 3034 464 3050 498
rect 3084 464 3100 498
rect 2840 313 2974 379
rect 2510 85 2582 119
rect 2616 85 2654 119
rect 2822 119 3000 279
rect 3034 158 3100 464
rect 3134 729 3312 751
rect 3168 695 3206 729
rect 3240 695 3278 729
rect 3134 435 3312 695
rect 3346 498 3412 751
rect 3346 464 3362 498
rect 3396 464 3412 498
rect 3152 313 3286 379
rect 2822 85 2894 119
rect 2928 85 2966 119
rect 3134 119 3312 279
rect 3346 158 3412 464
rect 3446 729 3624 751
rect 3480 695 3518 729
rect 3552 695 3590 729
rect 3446 435 3624 695
rect 3658 498 3724 751
rect 3658 464 3674 498
rect 3708 464 3724 498
rect 3464 313 3598 379
rect 3134 85 3206 119
rect 3240 85 3278 119
rect 3446 119 3624 279
rect 3658 158 3724 464
rect 3758 729 3936 751
rect 3792 695 3830 729
rect 3864 695 3902 729
rect 3758 435 3936 695
rect 3970 498 4052 751
rect 3970 464 3986 498
rect 4020 464 4052 498
rect 3776 313 3910 379
rect 3446 85 3518 119
rect 3552 85 3590 119
rect 3758 119 3936 279
rect 3970 158 4052 464
rect 4086 729 4192 751
rect 4120 695 4158 729
rect 4086 435 4192 695
rect 4282 498 4348 751
rect 4282 464 4298 498
rect 4332 464 4348 498
rect 4086 313 4220 379
rect 3758 85 3830 119
rect 3864 85 3902 119
rect 4086 119 4192 279
rect 4282 158 4348 464
rect 4382 729 4560 751
rect 4416 695 4454 729
rect 4488 695 4526 729
rect 4382 435 4560 695
rect 4594 498 4660 751
rect 4594 464 4610 498
rect 4644 464 4660 498
rect 4400 313 4534 379
rect 4086 85 4158 119
rect 4382 119 4560 279
rect 4594 158 4660 464
rect 4694 729 4872 751
rect 4728 695 4766 729
rect 4800 695 4838 729
rect 4694 435 4872 695
rect 4906 498 4972 751
rect 4906 464 4922 498
rect 4956 464 4972 498
rect 4712 313 4846 379
rect 4382 85 4454 119
rect 4488 85 4526 119
rect 4694 119 4872 279
rect 4906 158 4972 464
rect 5006 729 5184 751
rect 5040 695 5078 729
rect 5112 695 5150 729
rect 5006 435 5184 695
rect 5218 498 5284 751
rect 5218 464 5234 498
rect 5268 464 5284 498
rect 5024 313 5158 379
rect 4694 85 4766 119
rect 4800 85 4838 119
rect 5006 119 5184 279
rect 5218 158 5284 464
rect 5318 729 5496 751
rect 5352 695 5390 729
rect 5424 695 5462 729
rect 5318 435 5496 695
rect 5530 498 5596 751
rect 5530 464 5546 498
rect 5580 464 5596 498
rect 5336 313 5470 379
rect 5006 85 5078 119
rect 5112 85 5150 119
rect 5318 119 5496 279
rect 5530 158 5596 464
rect 5630 729 5808 751
rect 5664 695 5702 729
rect 5736 695 5774 729
rect 5630 435 5808 695
rect 5842 498 5908 751
rect 5842 464 5858 498
rect 5892 464 5908 498
rect 5648 313 5782 379
rect 5318 85 5390 119
rect 5424 85 5462 119
rect 5630 119 5808 279
rect 5842 158 5908 464
rect 5942 729 6120 751
rect 5976 695 6014 729
rect 6048 695 6086 729
rect 5942 435 6120 695
rect 6154 498 6220 751
rect 6154 464 6170 498
rect 6204 464 6220 498
rect 5960 313 6094 379
rect 5630 85 5702 119
rect 5736 85 5774 119
rect 5942 119 6120 279
rect 6154 158 6220 464
rect 6254 729 6432 751
rect 6288 695 6326 729
rect 6360 695 6398 729
rect 6254 435 6432 695
rect 6466 498 6548 751
rect 6466 464 6482 498
rect 6516 464 6548 498
rect 6272 313 6406 379
rect 5942 85 6014 119
rect 6048 85 6086 119
rect 6254 119 6432 279
rect 6466 158 6548 464
rect 6582 729 6688 751
rect 6616 695 6654 729
rect 6582 435 6688 695
rect 6254 85 6326 119
rect 6360 85 6398 119
rect 6582 119 6688 299
rect 6582 85 6654 119
rect 268 83 446 85
<< obsli1c >>
rect 30 695 64 729
rect 102 695 136 729
rect 268 695 302 729
rect 340 695 374 729
rect 412 695 446 729
rect 576 695 610 729
rect 648 695 682 729
rect 720 695 754 729
rect 892 695 926 729
rect 964 695 998 729
rect 1036 695 1070 729
rect 1200 695 1234 729
rect 1272 695 1306 729
rect 1344 695 1378 729
rect 1516 695 1550 729
rect 1588 695 1622 729
rect 1660 695 1694 729
rect 1802 464 1836 498
rect 23 85 57 119
rect 95 85 129 119
rect 268 85 302 119
rect 340 85 374 119
rect 412 85 446 119
rect 664 85 698 119
rect 736 85 770 119
rect 960 85 994 119
rect 1032 85 1066 119
rect 1288 85 1322 119
rect 1360 85 1394 119
rect 1886 695 1920 729
rect 1958 695 1992 729
rect 2030 695 2064 729
rect 2114 464 2148 498
rect 1584 85 1618 119
rect 1656 85 1690 119
rect 2198 695 2232 729
rect 2270 695 2304 729
rect 2342 695 2376 729
rect 2426 464 2460 498
rect 1958 85 1992 119
rect 2030 85 2064 119
rect 2510 695 2544 729
rect 2582 695 2616 729
rect 2654 695 2688 729
rect 2738 464 2772 498
rect 2270 85 2304 119
rect 2342 85 2376 119
rect 2822 695 2856 729
rect 2894 695 2928 729
rect 2966 695 3000 729
rect 3050 464 3084 498
rect 2582 85 2616 119
rect 2654 85 2688 119
rect 3134 695 3168 729
rect 3206 695 3240 729
rect 3278 695 3312 729
rect 3362 464 3396 498
rect 2894 85 2928 119
rect 2966 85 3000 119
rect 3446 695 3480 729
rect 3518 695 3552 729
rect 3590 695 3624 729
rect 3674 464 3708 498
rect 3206 85 3240 119
rect 3278 85 3312 119
rect 3758 695 3792 729
rect 3830 695 3864 729
rect 3902 695 3936 729
rect 3986 464 4020 498
rect 3518 85 3552 119
rect 3590 85 3624 119
rect 4086 695 4120 729
rect 4158 695 4192 729
rect 4298 464 4332 498
rect 3830 85 3864 119
rect 3902 85 3936 119
rect 4382 695 4416 729
rect 4454 695 4488 729
rect 4526 695 4560 729
rect 4610 464 4644 498
rect 4158 85 4192 119
rect 4694 695 4728 729
rect 4766 695 4800 729
rect 4838 695 4872 729
rect 4922 464 4956 498
rect 4454 85 4488 119
rect 4526 85 4560 119
rect 5006 695 5040 729
rect 5078 695 5112 729
rect 5150 695 5184 729
rect 5234 464 5268 498
rect 4766 85 4800 119
rect 4838 85 4872 119
rect 5318 695 5352 729
rect 5390 695 5424 729
rect 5462 695 5496 729
rect 5546 464 5580 498
rect 5078 85 5112 119
rect 5150 85 5184 119
rect 5630 695 5664 729
rect 5702 695 5736 729
rect 5774 695 5808 729
rect 5858 464 5892 498
rect 5390 85 5424 119
rect 5462 85 5496 119
rect 5942 695 5976 729
rect 6014 695 6048 729
rect 6086 695 6120 729
rect 6170 464 6204 498
rect 5702 85 5736 119
rect 5774 85 5808 119
rect 6254 695 6288 729
rect 6326 695 6360 729
rect 6398 695 6432 729
rect 6482 464 6516 498
rect 6014 85 6048 119
rect 6086 85 6120 119
rect 6582 695 6616 729
rect 6654 695 6688 729
rect 6326 85 6360 119
rect 6398 85 6432 119
rect 6654 85 6688 119
<< metal1 >>
rect 0 831 6720 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4063 831
rect 4097 797 4159 831
rect 4193 797 4255 831
rect 4289 797 4351 831
rect 4385 797 4447 831
rect 4481 797 4543 831
rect 4577 797 4639 831
rect 4673 797 4735 831
rect 4769 797 4831 831
rect 4865 797 4927 831
rect 4961 797 5023 831
rect 5057 797 5119 831
rect 5153 797 5215 831
rect 5249 797 5311 831
rect 5345 797 5407 831
rect 5441 797 5503 831
rect 5537 797 5599 831
rect 5633 797 5695 831
rect 5729 797 5791 831
rect 5825 797 5887 831
rect 5921 797 5983 831
rect 6017 797 6079 831
rect 6113 797 6175 831
rect 6209 797 6271 831
rect 6305 797 6367 831
rect 6401 797 6463 831
rect 6497 797 6559 831
rect 6593 797 6655 831
rect 6689 797 6720 831
rect 0 791 6720 797
rect 0 729 6720 763
rect 0 695 30 729
rect 64 695 102 729
rect 136 695 268 729
rect 302 695 340 729
rect 374 695 412 729
rect 446 695 576 729
rect 610 695 648 729
rect 682 695 720 729
rect 754 695 892 729
rect 926 695 964 729
rect 998 695 1036 729
rect 1070 695 1200 729
rect 1234 695 1272 729
rect 1306 695 1344 729
rect 1378 695 1516 729
rect 1550 695 1588 729
rect 1622 695 1660 729
rect 1694 695 1886 729
rect 1920 695 1958 729
rect 1992 695 2030 729
rect 2064 695 2198 729
rect 2232 695 2270 729
rect 2304 695 2342 729
rect 2376 695 2510 729
rect 2544 695 2582 729
rect 2616 695 2654 729
rect 2688 695 2822 729
rect 2856 695 2894 729
rect 2928 695 2966 729
rect 3000 695 3134 729
rect 3168 695 3206 729
rect 3240 695 3278 729
rect 3312 695 3446 729
rect 3480 695 3518 729
rect 3552 695 3590 729
rect 3624 695 3758 729
rect 3792 695 3830 729
rect 3864 695 3902 729
rect 3936 695 4086 729
rect 4120 695 4158 729
rect 4192 695 4382 729
rect 4416 695 4454 729
rect 4488 695 4526 729
rect 4560 695 4694 729
rect 4728 695 4766 729
rect 4800 695 4838 729
rect 4872 695 5006 729
rect 5040 695 5078 729
rect 5112 695 5150 729
rect 5184 695 5318 729
rect 5352 695 5390 729
rect 5424 695 5462 729
rect 5496 695 5630 729
rect 5664 695 5702 729
rect 5736 695 5774 729
rect 5808 695 5942 729
rect 5976 695 6014 729
rect 6048 695 6086 729
rect 6120 695 6254 729
rect 6288 695 6326 729
rect 6360 695 6398 729
rect 6432 695 6582 729
rect 6616 695 6654 729
rect 6688 695 6720 729
rect 0 689 6720 695
rect 1790 498 6528 504
rect 1790 464 1802 498
rect 1836 464 2114 498
rect 2148 464 2426 498
rect 2460 464 2738 498
rect 2772 464 3050 498
rect 3084 464 3362 498
rect 3396 464 3674 498
rect 3708 464 3986 498
rect 4020 464 4298 498
rect 4332 464 4610 498
rect 4644 464 4922 498
rect 4956 464 5234 498
rect 5268 464 5546 498
rect 5580 464 5858 498
rect 5892 464 6170 498
rect 6204 464 6482 498
rect 6516 464 6528 498
rect 1790 458 6528 464
rect 0 119 6720 125
rect 0 85 23 119
rect 57 85 95 119
rect 129 85 268 119
rect 302 85 340 119
rect 374 85 412 119
rect 446 85 664 119
rect 698 85 736 119
rect 770 85 960 119
rect 994 85 1032 119
rect 1066 85 1288 119
rect 1322 85 1360 119
rect 1394 85 1584 119
rect 1618 85 1656 119
rect 1690 85 1958 119
rect 1992 85 2030 119
rect 2064 85 2270 119
rect 2304 85 2342 119
rect 2376 85 2582 119
rect 2616 85 2654 119
rect 2688 85 2894 119
rect 2928 85 2966 119
rect 3000 85 3206 119
rect 3240 85 3278 119
rect 3312 85 3518 119
rect 3552 85 3590 119
rect 3624 85 3830 119
rect 3864 85 3902 119
rect 3936 85 4158 119
rect 4192 85 4454 119
rect 4488 85 4526 119
rect 4560 85 4766 119
rect 4800 85 4838 119
rect 4872 85 5078 119
rect 5112 85 5150 119
rect 5184 85 5390 119
rect 5424 85 5462 119
rect 5496 85 5702 119
rect 5736 85 5774 119
rect 5808 85 6014 119
rect 6048 85 6086 119
rect 6120 85 6326 119
rect 6360 85 6398 119
rect 6432 85 6654 119
rect 6688 85 6720 119
rect 0 51 6720 85
rect 0 17 6720 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 5023 17
rect 5057 -17 5119 17
rect 5153 -17 5215 17
rect 5249 -17 5311 17
rect 5345 -17 5407 17
rect 5441 -17 5503 17
rect 5537 -17 5599 17
rect 5633 -17 5695 17
rect 5729 -17 5791 17
rect 5825 -17 5887 17
rect 5921 -17 5983 17
rect 6017 -17 6079 17
rect 6113 -17 6175 17
rect 6209 -17 6271 17
rect 6305 -17 6367 17
rect 6401 -17 6463 17
rect 6497 -17 6559 17
rect 6593 -17 6655 17
rect 6689 -17 6720 17
rect 0 -23 6720 -17
<< obsm1 >>
rect 992 310 6418 356
<< labels >>
rlabel locali s 44 316 926 363 6 A
port 1 nsew signal input
rlabel metal1 s 1790 458 6528 504 6 X
port 6 nsew signal output
rlabel metal1 s 0 51 6720 125 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 6655 -17 6689 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 6559 -17 6593 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 6463 -17 6497 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 6367 -17 6401 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 6271 -17 6305 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 6175 -17 6209 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 6079 -17 6113 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5983 -17 6017 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5887 -17 5921 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5791 -17 5825 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5695 -17 5729 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5599 -17 5633 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5503 -17 5537 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5407 -17 5441 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5311 -17 5345 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5215 -17 5249 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5119 -17 5153 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 5023 -17 5057 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4927 -17 4961 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4831 -17 4865 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4735 -17 4769 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4639 -17 4673 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4543 -17 4577 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4447 -17 4481 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4351 -17 4385 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4255 -17 4289 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4159 -17 4193 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 4063 -17 4097 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3967 -17 4001 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3871 -17 3905 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3775 -17 3809 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3679 -17 3713 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3583 -17 3617 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3487 -17 3521 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3391 -17 3425 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3295 -17 3329 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3199 -17 3233 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3103 -17 3137 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 3007 -17 3041 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2911 -17 2945 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2815 -17 2849 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2719 -17 2753 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2623 -17 2657 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2527 -17 2561 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2431 -17 2465 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2335 -17 2369 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2239 -17 2273 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2143 -17 2177 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 2047 -17 2081 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1951 -17 1985 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1855 -17 1889 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1759 -17 1793 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1663 -17 1697 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1567 -17 1601 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1471 -17 1505 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1375 -17 1409 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1279 -17 1313 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1183 -17 1217 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1087 -17 1121 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 991 -17 1025 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 895 -17 929 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 799 -17 833 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 703 -17 737 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 607 -17 641 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 511 -17 545 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 415 -17 449 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 319 -17 353 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 223 -17 257 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 127 -17 161 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 31 -17 65 17 8 VNB
port 3 nsew ground bidirectional
rlabel locali s 0 -17 6720 17 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 0 -17 6720 17 8 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 6720 23 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 6655 797 6689 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 6559 797 6593 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 6463 797 6497 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 6367 797 6401 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 6271 797 6305 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 6175 797 6209 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 6079 797 6113 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5983 797 6017 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5887 797 5921 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5791 797 5825 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5695 797 5729 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5599 797 5633 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5503 797 5537 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5407 797 5441 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5311 797 5345 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5215 797 5249 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5119 797 5153 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 5023 797 5057 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4927 797 4961 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4831 797 4865 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4735 797 4769 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4639 797 4673 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4543 797 4577 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4447 797 4481 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4351 797 4385 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4255 797 4289 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4159 797 4193 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 4063 797 4097 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3967 797 4001 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3871 797 3905 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3775 797 3809 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3679 797 3713 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3583 797 3617 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3487 797 3521 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3391 797 3425 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3295 797 3329 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3199 797 3233 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3103 797 3137 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 3007 797 3041 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2911 797 2945 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2815 797 2849 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2719 797 2753 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2623 797 2657 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2527 797 2561 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2431 797 2465 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2335 797 2369 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2239 797 2273 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2143 797 2177 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 2047 797 2081 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1951 797 1985 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1855 797 1889 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1759 797 1793 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1663 797 1697 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1567 797 1601 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1471 797 1505 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1375 797 1409 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1279 797 1313 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1183 797 1217 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1087 797 1121 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 991 797 1025 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 895 797 929 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 799 797 833 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 703 797 737 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 607 797 641 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 511 797 545 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 415 797 449 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 319 797 353 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 223 797 257 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 127 797 161 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 31 797 65 831 6 VPB
port 4 nsew power bidirectional
rlabel locali s 0 797 6720 831 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 6786 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 791 6720 837 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 6720 763 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 6720 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 1108086
string GDS_START 1048330
<< end >>
