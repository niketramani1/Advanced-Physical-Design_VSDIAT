magic
tech sky130A
magscale 1 2
timestamp 1624855596
<< checkpaint >>
rect -1326 -1283 1614 2157
<< nwell >>
rect -66 377 354 897
<< pwell >>
rect 0 -17 288 17
<< mvnmos >>
rect 101 107 201 257
<< mvpmos >>
rect 97 443 197 743
<< mvndiff >>
rect 44 249 101 257
rect 44 215 56 249
rect 90 215 101 249
rect 44 149 101 215
rect 44 115 56 149
rect 90 115 101 149
rect 44 107 101 115
rect 201 249 258 257
rect 201 215 212 249
rect 246 215 258 249
rect 201 149 258 215
rect 201 115 212 149
rect 246 115 258 149
rect 201 107 258 115
<< mvpdiff >>
rect 40 735 97 743
rect 40 701 52 735
rect 86 701 97 735
rect 40 652 97 701
rect 40 618 52 652
rect 86 618 97 652
rect 40 568 97 618
rect 40 534 52 568
rect 86 534 97 568
rect 40 485 97 534
rect 40 451 52 485
rect 86 451 97 485
rect 40 443 97 451
rect 197 735 254 743
rect 197 701 208 735
rect 242 701 254 735
rect 197 652 254 701
rect 197 618 208 652
rect 242 618 254 652
rect 197 568 254 618
rect 197 534 208 568
rect 242 534 254 568
rect 197 485 254 534
rect 197 451 208 485
rect 242 451 254 485
rect 197 443 254 451
<< mvndiffc >>
rect 56 215 90 249
rect 56 115 90 149
rect 212 215 246 249
rect 212 115 246 149
<< mvpdiffc >>
rect 52 701 86 735
rect 52 618 86 652
rect 52 534 86 568
rect 52 451 86 485
rect 208 701 242 735
rect 208 618 242 652
rect 208 534 242 568
rect 208 451 242 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 288 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
<< poly >>
rect 97 743 197 769
rect 97 417 197 443
rect 97 371 201 417
rect 97 337 117 371
rect 151 337 201 371
rect 97 283 201 337
rect 101 257 201 283
rect 101 81 201 107
<< polycont >>
rect 117 337 151 371
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 288 831
rect 18 735 136 751
rect 18 701 24 735
rect 86 701 96 735
rect 130 701 136 735
rect 18 652 136 701
rect 18 618 52 652
rect 86 618 136 652
rect 18 568 136 618
rect 18 534 52 568
rect 86 534 136 568
rect 18 485 136 534
rect 18 451 52 485
rect 86 451 136 485
rect 18 435 136 451
rect 192 735 269 751
rect 192 701 208 735
rect 242 701 269 735
rect 192 652 269 701
rect 192 618 208 652
rect 242 618 269 652
rect 192 568 269 618
rect 192 534 208 568
rect 242 534 269 568
rect 192 485 269 534
rect 192 451 208 485
rect 242 451 269 485
rect 192 435 269 451
rect 25 371 167 387
rect 25 337 117 371
rect 151 337 167 371
rect 25 310 167 337
rect 18 249 136 265
rect 18 215 56 249
rect 90 215 136 249
rect 18 149 136 215
rect 18 115 56 149
rect 90 115 136 149
rect 18 113 136 115
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 136 113
rect 203 249 269 435
rect 203 215 212 249
rect 246 215 269 249
rect 203 149 269 215
rect 203 115 212 149
rect 246 115 269 149
rect 203 99 269 115
rect 18 73 136 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 24 701 52 735
rect 52 701 58 735
rect 96 701 130 735
rect 24 79 58 113
rect 96 79 130 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< metal1 >>
rect 0 831 288 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 288 831
rect 0 791 288 797
rect 0 735 288 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 288 735
rect 0 689 288 701
rect 0 113 288 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 288 113
rect 0 51 288 79
rect 0 17 288 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
rect 0 -23 288 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_1
flabel metal1 s 0 51 288 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 0 288 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 689 288 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 288 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 612 257 646 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 288 814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string LEFsymmetry X Y
string GDS_END 217464
string GDS_START 211758
<< end >>
