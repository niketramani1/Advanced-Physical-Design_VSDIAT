magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1309 -1309 42619 2437
<< locali >>
rect -17 1137 17 1153
rect -17 1087 17 1103
rect 1784 1137 1818 1153
rect 1784 1087 1818 1103
rect 11768 1137 11802 1153
rect 11768 1087 11802 1103
rect 21752 1137 21786 1153
rect 21752 1087 21786 1103
rect 31736 1137 31770 1153
rect 31736 1087 31770 1103
rect 41293 1137 41327 1153
rect 41293 1087 41327 1103
rect 1586 535 1620 551
rect 1935 517 1969 551
rect 11570 535 11604 551
rect 1586 485 1620 501
rect 11919 517 11953 551
rect 21554 535 21588 551
rect 11570 485 11604 501
rect 21903 517 21937 551
rect 31538 535 31572 551
rect 21554 485 21588 501
rect 31887 517 31921 551
rect 31538 485 31572 501
rect 1357 287 1391 303
rect 11341 287 11375 303
rect 21325 287 21359 303
rect 31309 287 31343 303
rect 1391 253 1503 287
rect 11375 253 11487 287
rect 21359 253 21471 287
rect 31343 253 31455 287
rect 1357 237 1391 253
rect 11341 237 11375 253
rect 21325 237 21359 253
rect 31309 237 31343 253
rect -17 17 17 33
rect -17 -33 17 -17
rect 1784 17 1818 33
rect 1784 -33 1818 -17
rect 11768 17 11802 33
rect 11768 -33 11802 -17
rect 21752 17 21786 33
rect 21752 -33 21786 -17
rect 31736 17 31770 33
rect 31736 -33 31770 -17
rect 41293 17 41327 33
rect 41293 -33 41327 -17
<< viali >>
rect -17 1103 17 1137
rect 1784 1103 1818 1137
rect 11768 1103 11802 1137
rect 21752 1103 21786 1137
rect 31736 1103 31770 1137
rect 41293 1103 41327 1137
rect 1586 501 1620 535
rect 11570 501 11604 535
rect 21554 501 21588 535
rect 31538 501 31572 535
rect 1357 253 1391 287
rect 11341 253 11375 287
rect 21325 253 21359 287
rect 31309 253 31343 287
rect -17 -17 17 17
rect 1784 -17 1818 17
rect 11768 -17 11802 17
rect 21752 -17 21786 17
rect 31736 -17 31770 17
rect 41293 -17 41327 17
<< metal1 >>
rect -32 1094 -26 1146
rect 26 1134 32 1146
rect 1772 1137 1830 1143
rect 1772 1134 1784 1137
rect 26 1106 1784 1134
rect 26 1094 32 1106
rect 1772 1103 1784 1106
rect 1818 1134 1830 1137
rect 11756 1137 11814 1143
rect 11756 1134 11768 1137
rect 1818 1106 11768 1134
rect 1818 1103 1830 1106
rect 1772 1097 1830 1103
rect 11756 1103 11768 1106
rect 11802 1134 11814 1137
rect 21740 1137 21798 1143
rect 21740 1134 21752 1137
rect 11802 1106 21752 1134
rect 11802 1103 11814 1106
rect 11756 1097 11814 1103
rect 21740 1103 21752 1106
rect 21786 1134 21798 1137
rect 31724 1137 31782 1143
rect 31724 1134 31736 1137
rect 21786 1106 31736 1134
rect 21786 1103 21798 1106
rect 21740 1097 21798 1103
rect 31724 1103 31736 1106
rect 31770 1134 31782 1137
rect 41278 1134 41284 1146
rect 31770 1106 41284 1134
rect 31770 1103 31782 1106
rect 31724 1097 31782 1103
rect 41278 1094 41284 1106
rect 41336 1094 41342 1146
rect 1571 492 1577 544
rect 1629 492 1635 544
rect 11555 492 11561 544
rect 11613 492 11619 544
rect 21539 492 21545 544
rect 21597 492 21603 544
rect 31523 492 31529 544
rect 31581 492 31587 544
rect 1342 244 1348 296
rect 1400 244 1406 296
rect 11326 244 11332 296
rect 11384 244 11390 296
rect 21310 244 21316 296
rect 21368 244 21374 296
rect 31294 244 31300 296
rect 31352 244 31358 296
rect -32 -26 -26 26
rect 26 14 32 26
rect 1772 17 1830 23
rect 1772 14 1784 17
rect 26 -14 1784 14
rect 26 -26 32 -14
rect 1772 -17 1784 -14
rect 1818 14 1830 17
rect 11756 17 11814 23
rect 11756 14 11768 17
rect 1818 -14 11768 14
rect 1818 -17 1830 -14
rect 1772 -23 1830 -17
rect 11756 -17 11768 -14
rect 11802 14 11814 17
rect 21740 17 21798 23
rect 21740 14 21752 17
rect 11802 -14 21752 14
rect 11802 -17 11814 -14
rect 11756 -23 11814 -17
rect 21740 -17 21752 -14
rect 21786 14 21798 17
rect 31724 17 31782 23
rect 31724 14 31736 17
rect 21786 -14 31736 14
rect 21786 -17 21798 -14
rect 21740 -23 21798 -17
rect 31724 -17 31736 -14
rect 31770 14 31782 17
rect 41278 14 41284 26
rect 31770 -14 41284 14
rect 31770 -17 31782 -14
rect 31724 -23 31782 -17
rect 41278 -26 41284 -14
rect 41336 -26 41342 26
<< via1 >>
rect -26 1137 26 1146
rect -26 1103 -17 1137
rect -17 1103 17 1137
rect 17 1103 26 1137
rect -26 1094 26 1103
rect 41284 1137 41336 1146
rect 41284 1103 41293 1137
rect 41293 1103 41327 1137
rect 41327 1103 41336 1137
rect 41284 1094 41336 1103
rect 1577 535 1629 544
rect 1577 501 1586 535
rect 1586 501 1620 535
rect 1620 501 1629 535
rect 1577 492 1629 501
rect 11561 535 11613 544
rect 11561 501 11570 535
rect 11570 501 11604 535
rect 11604 501 11613 535
rect 11561 492 11613 501
rect 21545 535 21597 544
rect 21545 501 21554 535
rect 21554 501 21588 535
rect 21588 501 21597 535
rect 21545 492 21597 501
rect 31529 535 31581 544
rect 31529 501 31538 535
rect 31538 501 31572 535
rect 31572 501 31581 535
rect 31529 492 31581 501
rect 1348 287 1400 296
rect 1348 253 1357 287
rect 1357 253 1391 287
rect 1391 253 1400 287
rect 1348 244 1400 253
rect 11332 287 11384 296
rect 11332 253 11341 287
rect 11341 253 11375 287
rect 11375 253 11384 287
rect 11332 244 11384 253
rect 21316 287 21368 296
rect 21316 253 21325 287
rect 21325 253 21359 287
rect 21359 253 21368 287
rect 21316 244 21368 253
rect 31300 287 31352 296
rect 31300 253 31309 287
rect 31309 253 31343 287
rect 31343 253 31352 287
rect 31300 244 31352 253
rect -26 17 26 26
rect -26 -17 -17 17
rect -17 -17 17 17
rect 17 -17 26 17
rect -26 -26 26 -17
rect 41284 17 41336 26
rect 41284 -17 41293 17
rect 41293 -17 41327 17
rect 41327 -17 41336 17
rect 41284 -26 41336 -17
<< metal2 >>
rect -28 1148 28 1157
rect -28 1083 28 1092
rect 41282 1148 41338 1157
rect 41282 1083 41338 1092
rect 1575 546 1631 555
rect 1575 481 1631 490
rect 11559 546 11615 555
rect 11559 481 11615 490
rect 21543 546 21599 555
rect 21543 481 21599 490
rect 31527 546 31583 555
rect 31527 481 31583 490
rect 1348 296 1400 302
rect 1348 238 1400 244
rect 11332 296 11384 302
rect 11332 238 11384 244
rect 21316 296 21368 302
rect 21316 238 21368 244
rect 31300 296 31352 302
rect 31300 238 31352 244
rect -28 28 28 37
rect -28 -37 28 -28
rect 41282 28 41338 37
rect 41282 -37 41338 -28
<< via2 >>
rect -28 1146 28 1148
rect -28 1094 -26 1146
rect -26 1094 26 1146
rect 26 1094 28 1146
rect -28 1092 28 1094
rect 41282 1146 41338 1148
rect 41282 1094 41284 1146
rect 41284 1094 41336 1146
rect 41336 1094 41338 1146
rect 41282 1092 41338 1094
rect 1575 544 1631 546
rect 1575 492 1577 544
rect 1577 492 1629 544
rect 1629 492 1631 544
rect 1575 490 1631 492
rect 11559 544 11615 546
rect 11559 492 11561 544
rect 11561 492 11613 544
rect 11613 492 11615 544
rect 11559 490 11615 492
rect 21543 544 21599 546
rect 21543 492 21545 544
rect 21545 492 21597 544
rect 21597 492 21599 544
rect 21543 490 21599 492
rect 31527 544 31583 546
rect 31527 492 31529 544
rect 31529 492 31581 544
rect 31581 492 31583 544
rect 31527 490 31583 492
rect -28 26 28 28
rect -28 -26 -26 26
rect -26 -26 26 26
rect 26 -26 28 26
rect -28 -28 28 -26
rect 41282 26 41338 28
rect 41282 -26 41284 26
rect 41284 -26 41336 26
rect 41336 -26 41338 26
rect 41282 -28 41338 -26
<< metal3 >>
rect -49 1148 49 1169
rect -49 1092 -28 1148
rect 28 1092 49 1148
rect -49 1071 49 1092
rect 41261 1148 41359 1169
rect 41261 1092 41282 1148
rect 41338 1092 41359 1148
rect 41261 1071 41359 1092
rect 1570 548 1636 551
rect 11554 548 11620 551
rect 21538 548 21604 551
rect 31522 548 31588 551
rect 0 546 41310 548
rect 0 490 1575 546
rect 1631 490 11559 546
rect 11615 490 21543 546
rect 21599 490 31527 546
rect 31583 490 41310 546
rect 0 488 41310 490
rect 1570 485 1636 488
rect 11554 485 11620 488
rect 21538 485 21604 488
rect 31522 485 31588 488
rect -49 28 49 49
rect -49 -28 -28 28
rect 28 -28 49 28
rect -49 -49 49 -28
rect 41261 28 41359 49
rect 41261 -28 41282 28
rect 41338 -28 41359 28
rect 41261 -49 41359 -28
use contact_14  contact_14_7
timestamp 1624857261
transform 1 0 -29 0 1 -33
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1624857261
transform 1 0 -29 0 1 -33
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1624857261
transform 1 0 -32 0 1 -32
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1624857261
transform 1 0 -33 0 1 -37
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1624857261
transform 1 0 -29 0 1 1087
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1624857261
transform 1 0 -29 0 1 1087
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1624857261
transform 1 0 -32 0 1 1088
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1624857261
transform 1 0 -33 0 1 1083
box 0 0 1 1
use pand2  pand2_3
timestamp 1624857261
transform 1 0 1374 0 1 0
box -36 -17 890 1177
use contact_14  contact_14_23
timestamp 1624857261
transform 1 0 1345 0 1 237
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1624857261
transform 1 0 1342 0 1 238
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1624857261
transform 1 0 1574 0 1 485
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1624857261
transform 1 0 1571 0 1 486
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1624857261
transform 1 0 1570 0 1 481
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1624857261
transform 1 0 1772 0 1 -33
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1624857261
transform 1 0 1772 0 1 1087
box 0 0 1 1
use pand2  pand2_2
timestamp 1624857261
transform 1 0 11358 0 1 0
box -36 -17 890 1177
use contact_14  contact_14_19
timestamp 1624857261
transform 1 0 11329 0 1 237
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1624857261
transform 1 0 11326 0 1 238
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1624857261
transform 1 0 11558 0 1 485
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1624857261
transform 1 0 11555 0 1 486
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1624857261
transform 1 0 11554 0 1 481
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1624857261
transform 1 0 11756 0 1 -33
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1624857261
transform 1 0 11756 0 1 1087
box 0 0 1 1
use pand2  pand2_1
timestamp 1624857261
transform 1 0 21342 0 1 0
box -36 -17 890 1177
use contact_14  contact_14_15
timestamp 1624857261
transform 1 0 21313 0 1 237
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1624857261
transform 1 0 21310 0 1 238
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1624857261
transform 1 0 21542 0 1 485
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1624857261
transform 1 0 21539 0 1 486
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1624857261
transform 1 0 21538 0 1 481
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1624857261
transform 1 0 21740 0 1 -33
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1624857261
transform 1 0 21740 0 1 1087
box 0 0 1 1
use pand2  pand2_0
timestamp 1624857261
transform 1 0 31326 0 1 0
box -36 -17 890 1177
use contact_14  contact_14_11
timestamp 1624857261
transform 1 0 31297 0 1 237
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1624857261
transform 1 0 31294 0 1 238
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1624857261
transform 1 0 31526 0 1 485
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1624857261
transform 1 0 31523 0 1 486
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1624857261
transform 1 0 31522 0 1 481
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1624857261
transform 1 0 31724 0 1 -33
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1624857261
transform 1 0 31724 0 1 1087
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1624857261
transform 1 0 41281 0 1 -33
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1624857261
transform 1 0 41281 0 1 -33
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1624857261
transform 1 0 41278 0 1 -32
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1624857261
transform 1 0 41277 0 1 -37
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1624857261
transform 1 0 41281 0 1 1087
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1624857261
transform 1 0 41281 0 1 1087
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1624857261
transform 1 0 41278 0 1 1088
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1624857261
transform 1 0 41277 0 1 1083
box 0 0 1 1
<< labels >>
rlabel metal3 s 0 488 41310 548 4 en
port 5 se
rlabel metal2 s 1360 256 1388 284 4 wmask_in_0
port 1 se
rlabel locali s 1952 534 1952 534 4 wmask_out_0
port 6 se
rlabel metal2 s 11344 256 11372 284 4 wmask_in_1
port 2 se
rlabel locali s 11936 534 11936 534 4 wmask_out_1
port 7 se
rlabel metal2 s 21328 256 21356 284 4 wmask_in_2
port 3 se
rlabel locali s 21920 534 21920 534 4 wmask_out_2
port 8 se
rlabel metal2 s 31312 256 31340 284 4 wmask_in_3
port 4 se
rlabel locali s 31904 534 31904 534 4 wmask_out_3
port 9 se
rlabel metal3 s -49 -49 49 49 4 gnd
rlabel metal3 s 41261 -49 41359 49 4 gnd
port 11 se
rlabel metal3 s -49 1071 49 1169 4 vdd
rlabel metal3 s 41261 1071 41359 1169 4 vdd
port 10 se
<< properties >>
string FIXED_BBOX 41277 -37 41343 0
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 7874986
string GDS_START 7869226
<< end >>
