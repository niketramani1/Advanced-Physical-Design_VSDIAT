magic
tech sky130A
magscale 1 2
timestamp 1624855514
<< obsm3 >>
rect 99 1778 14858 2706
<< metal4 >>
rect 0 10625 15000 11221
rect 0 9673 15000 10269
rect 105 2640 169 2704
rect 187 2640 251 2704
rect 269 2640 333 2704
rect 351 2640 415 2704
rect 433 2640 497 2704
rect 515 2640 579 2704
rect 597 2640 661 2704
rect 678 2640 742 2704
rect 759 2640 823 2704
rect 840 2640 904 2704
rect 921 2640 985 2704
rect 1002 2640 1066 2704
rect 1083 2640 1147 2704
rect 1164 2640 1228 2704
rect 1245 2640 1309 2704
rect 1326 2640 1390 2704
rect 1407 2640 1471 2704
rect 1488 2640 1552 2704
rect 1569 2640 1633 2704
rect 1650 2640 1714 2704
rect 1731 2640 1795 2704
rect 1812 2640 1876 2704
rect 1893 2640 1957 2704
rect 1974 2640 2038 2704
rect 2055 2640 2119 2704
rect 2136 2640 2200 2704
rect 2217 2640 2281 2704
rect 2298 2640 2362 2704
rect 2379 2640 2443 2704
rect 2460 2640 2524 2704
rect 2541 2640 2605 2704
rect 2622 2640 2686 2704
rect 2703 2640 2767 2704
rect 2784 2640 2848 2704
rect 2865 2640 2929 2704
rect 2946 2640 3010 2704
rect 3027 2640 3091 2704
rect 3108 2640 3172 2704
rect 3189 2640 3253 2704
rect 3270 2640 3334 2704
rect 3351 2640 3415 2704
rect 3432 2640 3496 2704
rect 3513 2640 3577 2704
rect 3594 2640 3658 2704
rect 3675 2640 3739 2704
rect 3756 2640 3820 2704
rect 3837 2640 3901 2704
rect 3918 2640 3982 2704
rect 3999 2640 4063 2704
rect 4080 2640 4144 2704
rect 4161 2640 4225 2704
rect 4242 2640 4306 2704
rect 4323 2640 4387 2704
rect 4404 2640 4468 2704
rect 4485 2640 4549 2704
rect 4566 2640 4630 2704
rect 4647 2640 4711 2704
rect 4728 2640 4792 2704
rect 4809 2640 4873 2704
rect 10084 2640 10148 2704
rect 10166 2640 10230 2704
rect 10248 2640 10312 2704
rect 10330 2640 10394 2704
rect 10412 2640 10476 2704
rect 10494 2640 10558 2704
rect 10576 2640 10640 2704
rect 10657 2640 10721 2704
rect 10738 2640 10802 2704
rect 10819 2640 10883 2704
rect 10900 2640 10964 2704
rect 10981 2640 11045 2704
rect 11062 2640 11126 2704
rect 11143 2640 11207 2704
rect 11224 2640 11288 2704
rect 11305 2640 11369 2704
rect 11386 2640 11450 2704
rect 11467 2640 11531 2704
rect 11548 2640 11612 2704
rect 11629 2640 11693 2704
rect 11710 2640 11774 2704
rect 11791 2640 11855 2704
rect 11872 2640 11936 2704
rect 11953 2640 12017 2704
rect 12034 2640 12098 2704
rect 12115 2640 12179 2704
rect 12196 2640 12260 2704
rect 12277 2640 12341 2704
rect 12358 2640 12422 2704
rect 12439 2640 12503 2704
rect 12520 2640 12584 2704
rect 12601 2640 12665 2704
rect 12682 2640 12746 2704
rect 12763 2640 12827 2704
rect 12844 2640 12908 2704
rect 12925 2640 12989 2704
rect 13006 2640 13070 2704
rect 13087 2640 13151 2704
rect 13168 2640 13232 2704
rect 13249 2640 13313 2704
rect 13330 2640 13394 2704
rect 13411 2640 13475 2704
rect 13492 2640 13556 2704
rect 13573 2640 13637 2704
rect 13654 2640 13718 2704
rect 13735 2640 13799 2704
rect 13816 2640 13880 2704
rect 13897 2640 13961 2704
rect 13978 2640 14042 2704
rect 14059 2640 14123 2704
rect 14140 2640 14204 2704
rect 14221 2640 14285 2704
rect 14302 2640 14366 2704
rect 14383 2640 14447 2704
rect 14464 2640 14528 2704
rect 14545 2640 14609 2704
rect 14626 2640 14690 2704
rect 14707 2640 14771 2704
rect 14788 2640 14852 2704
rect 105 2554 169 2618
rect 187 2554 251 2618
rect 269 2554 333 2618
rect 351 2554 415 2618
rect 433 2554 497 2618
rect 515 2554 579 2618
rect 597 2554 661 2618
rect 678 2554 742 2618
rect 759 2554 823 2618
rect 840 2554 904 2618
rect 921 2554 985 2618
rect 1002 2554 1066 2618
rect 1083 2554 1147 2618
rect 1164 2554 1228 2618
rect 1245 2554 1309 2618
rect 1326 2554 1390 2618
rect 1407 2554 1471 2618
rect 1488 2554 1552 2618
rect 1569 2554 1633 2618
rect 1650 2554 1714 2618
rect 1731 2554 1795 2618
rect 1812 2554 1876 2618
rect 1893 2554 1957 2618
rect 1974 2554 2038 2618
rect 2055 2554 2119 2618
rect 2136 2554 2200 2618
rect 2217 2554 2281 2618
rect 2298 2554 2362 2618
rect 2379 2554 2443 2618
rect 2460 2554 2524 2618
rect 2541 2554 2605 2618
rect 2622 2554 2686 2618
rect 2703 2554 2767 2618
rect 2784 2554 2848 2618
rect 2865 2554 2929 2618
rect 2946 2554 3010 2618
rect 3027 2554 3091 2618
rect 3108 2554 3172 2618
rect 3189 2554 3253 2618
rect 3270 2554 3334 2618
rect 3351 2554 3415 2618
rect 3432 2554 3496 2618
rect 3513 2554 3577 2618
rect 3594 2554 3658 2618
rect 3675 2554 3739 2618
rect 3756 2554 3820 2618
rect 3837 2554 3901 2618
rect 3918 2554 3982 2618
rect 3999 2554 4063 2618
rect 4080 2554 4144 2618
rect 4161 2554 4225 2618
rect 4242 2554 4306 2618
rect 4323 2554 4387 2618
rect 4404 2554 4468 2618
rect 4485 2554 4549 2618
rect 4566 2554 4630 2618
rect 4647 2554 4711 2618
rect 4728 2554 4792 2618
rect 4809 2554 4873 2618
rect 10084 2554 10148 2618
rect 10166 2554 10230 2618
rect 10248 2554 10312 2618
rect 10330 2554 10394 2618
rect 10412 2554 10476 2618
rect 10494 2554 10558 2618
rect 10576 2554 10640 2618
rect 10657 2554 10721 2618
rect 10738 2554 10802 2618
rect 10819 2554 10883 2618
rect 10900 2554 10964 2618
rect 10981 2554 11045 2618
rect 11062 2554 11126 2618
rect 11143 2554 11207 2618
rect 11224 2554 11288 2618
rect 11305 2554 11369 2618
rect 11386 2554 11450 2618
rect 11467 2554 11531 2618
rect 11548 2554 11612 2618
rect 11629 2554 11693 2618
rect 11710 2554 11774 2618
rect 11791 2554 11855 2618
rect 11872 2554 11936 2618
rect 11953 2554 12017 2618
rect 12034 2554 12098 2618
rect 12115 2554 12179 2618
rect 12196 2554 12260 2618
rect 12277 2554 12341 2618
rect 12358 2554 12422 2618
rect 12439 2554 12503 2618
rect 12520 2554 12584 2618
rect 12601 2554 12665 2618
rect 12682 2554 12746 2618
rect 12763 2554 12827 2618
rect 12844 2554 12908 2618
rect 12925 2554 12989 2618
rect 13006 2554 13070 2618
rect 13087 2554 13151 2618
rect 13168 2554 13232 2618
rect 13249 2554 13313 2618
rect 13330 2554 13394 2618
rect 13411 2554 13475 2618
rect 13492 2554 13556 2618
rect 13573 2554 13637 2618
rect 13654 2554 13718 2618
rect 13735 2554 13799 2618
rect 13816 2554 13880 2618
rect 13897 2554 13961 2618
rect 13978 2554 14042 2618
rect 14059 2554 14123 2618
rect 14140 2554 14204 2618
rect 14221 2554 14285 2618
rect 14302 2554 14366 2618
rect 14383 2554 14447 2618
rect 14464 2554 14528 2618
rect 14545 2554 14609 2618
rect 14626 2554 14690 2618
rect 14707 2554 14771 2618
rect 14788 2554 14852 2618
rect 105 2468 169 2532
rect 187 2468 251 2532
rect 269 2468 333 2532
rect 351 2468 415 2532
rect 433 2468 497 2532
rect 515 2468 579 2532
rect 597 2468 661 2532
rect 678 2468 742 2532
rect 759 2468 823 2532
rect 840 2468 904 2532
rect 921 2468 985 2532
rect 1002 2468 1066 2532
rect 1083 2468 1147 2532
rect 1164 2468 1228 2532
rect 1245 2468 1309 2532
rect 1326 2468 1390 2532
rect 1407 2468 1471 2532
rect 1488 2468 1552 2532
rect 1569 2468 1633 2532
rect 1650 2468 1714 2532
rect 1731 2468 1795 2532
rect 1812 2468 1876 2532
rect 1893 2468 1957 2532
rect 1974 2468 2038 2532
rect 2055 2468 2119 2532
rect 2136 2468 2200 2532
rect 2217 2468 2281 2532
rect 2298 2468 2362 2532
rect 2379 2468 2443 2532
rect 2460 2468 2524 2532
rect 2541 2468 2605 2532
rect 2622 2468 2686 2532
rect 2703 2468 2767 2532
rect 2784 2468 2848 2532
rect 2865 2468 2929 2532
rect 2946 2468 3010 2532
rect 3027 2468 3091 2532
rect 3108 2468 3172 2532
rect 3189 2468 3253 2532
rect 3270 2468 3334 2532
rect 3351 2468 3415 2532
rect 3432 2468 3496 2532
rect 3513 2468 3577 2532
rect 3594 2468 3658 2532
rect 3675 2468 3739 2532
rect 3756 2468 3820 2532
rect 3837 2468 3901 2532
rect 3918 2468 3982 2532
rect 3999 2468 4063 2532
rect 4080 2468 4144 2532
rect 4161 2468 4225 2532
rect 4242 2468 4306 2532
rect 4323 2468 4387 2532
rect 4404 2468 4468 2532
rect 4485 2468 4549 2532
rect 4566 2468 4630 2532
rect 4647 2468 4711 2532
rect 4728 2468 4792 2532
rect 4809 2468 4873 2532
rect 10084 2468 10148 2532
rect 10166 2468 10230 2532
rect 10248 2468 10312 2532
rect 10330 2468 10394 2532
rect 10412 2468 10476 2532
rect 10494 2468 10558 2532
rect 10576 2468 10640 2532
rect 10657 2468 10721 2532
rect 10738 2468 10802 2532
rect 10819 2468 10883 2532
rect 10900 2468 10964 2532
rect 10981 2468 11045 2532
rect 11062 2468 11126 2532
rect 11143 2468 11207 2532
rect 11224 2468 11288 2532
rect 11305 2468 11369 2532
rect 11386 2468 11450 2532
rect 11467 2468 11531 2532
rect 11548 2468 11612 2532
rect 11629 2468 11693 2532
rect 11710 2468 11774 2532
rect 11791 2468 11855 2532
rect 11872 2468 11936 2532
rect 11953 2468 12017 2532
rect 12034 2468 12098 2532
rect 12115 2468 12179 2532
rect 12196 2468 12260 2532
rect 12277 2468 12341 2532
rect 12358 2468 12422 2532
rect 12439 2468 12503 2532
rect 12520 2468 12584 2532
rect 12601 2468 12665 2532
rect 12682 2468 12746 2532
rect 12763 2468 12827 2532
rect 12844 2468 12908 2532
rect 12925 2468 12989 2532
rect 13006 2468 13070 2532
rect 13087 2468 13151 2532
rect 13168 2468 13232 2532
rect 13249 2468 13313 2532
rect 13330 2468 13394 2532
rect 13411 2468 13475 2532
rect 13492 2468 13556 2532
rect 13573 2468 13637 2532
rect 13654 2468 13718 2532
rect 13735 2468 13799 2532
rect 13816 2468 13880 2532
rect 13897 2468 13961 2532
rect 13978 2468 14042 2532
rect 14059 2468 14123 2532
rect 14140 2468 14204 2532
rect 14221 2468 14285 2532
rect 14302 2468 14366 2532
rect 14383 2468 14447 2532
rect 14464 2468 14528 2532
rect 14545 2468 14609 2532
rect 14626 2468 14690 2532
rect 14707 2468 14771 2532
rect 14788 2468 14852 2532
rect 105 2382 169 2446
rect 187 2382 251 2446
rect 269 2382 333 2446
rect 351 2382 415 2446
rect 433 2382 497 2446
rect 515 2382 579 2446
rect 597 2382 661 2446
rect 678 2382 742 2446
rect 759 2382 823 2446
rect 840 2382 904 2446
rect 921 2382 985 2446
rect 1002 2382 1066 2446
rect 1083 2382 1147 2446
rect 1164 2382 1228 2446
rect 1245 2382 1309 2446
rect 1326 2382 1390 2446
rect 1407 2382 1471 2446
rect 1488 2382 1552 2446
rect 1569 2382 1633 2446
rect 1650 2382 1714 2446
rect 1731 2382 1795 2446
rect 1812 2382 1876 2446
rect 1893 2382 1957 2446
rect 1974 2382 2038 2446
rect 2055 2382 2119 2446
rect 2136 2382 2200 2446
rect 2217 2382 2281 2446
rect 2298 2382 2362 2446
rect 2379 2382 2443 2446
rect 2460 2382 2524 2446
rect 2541 2382 2605 2446
rect 2622 2382 2686 2446
rect 2703 2382 2767 2446
rect 2784 2382 2848 2446
rect 2865 2382 2929 2446
rect 2946 2382 3010 2446
rect 3027 2382 3091 2446
rect 3108 2382 3172 2446
rect 3189 2382 3253 2446
rect 3270 2382 3334 2446
rect 3351 2382 3415 2446
rect 3432 2382 3496 2446
rect 3513 2382 3577 2446
rect 3594 2382 3658 2446
rect 3675 2382 3739 2446
rect 3756 2382 3820 2446
rect 3837 2382 3901 2446
rect 3918 2382 3982 2446
rect 3999 2382 4063 2446
rect 4080 2382 4144 2446
rect 4161 2382 4225 2446
rect 4242 2382 4306 2446
rect 4323 2382 4387 2446
rect 4404 2382 4468 2446
rect 4485 2382 4549 2446
rect 4566 2382 4630 2446
rect 4647 2382 4711 2446
rect 4728 2382 4792 2446
rect 4809 2382 4873 2446
rect 10084 2382 10148 2446
rect 10166 2382 10230 2446
rect 10248 2382 10312 2446
rect 10330 2382 10394 2446
rect 10412 2382 10476 2446
rect 10494 2382 10558 2446
rect 10576 2382 10640 2446
rect 10657 2382 10721 2446
rect 10738 2382 10802 2446
rect 10819 2382 10883 2446
rect 10900 2382 10964 2446
rect 10981 2382 11045 2446
rect 11062 2382 11126 2446
rect 11143 2382 11207 2446
rect 11224 2382 11288 2446
rect 11305 2382 11369 2446
rect 11386 2382 11450 2446
rect 11467 2382 11531 2446
rect 11548 2382 11612 2446
rect 11629 2382 11693 2446
rect 11710 2382 11774 2446
rect 11791 2382 11855 2446
rect 11872 2382 11936 2446
rect 11953 2382 12017 2446
rect 12034 2382 12098 2446
rect 12115 2382 12179 2446
rect 12196 2382 12260 2446
rect 12277 2382 12341 2446
rect 12358 2382 12422 2446
rect 12439 2382 12503 2446
rect 12520 2382 12584 2446
rect 12601 2382 12665 2446
rect 12682 2382 12746 2446
rect 12763 2382 12827 2446
rect 12844 2382 12908 2446
rect 12925 2382 12989 2446
rect 13006 2382 13070 2446
rect 13087 2382 13151 2446
rect 13168 2382 13232 2446
rect 13249 2382 13313 2446
rect 13330 2382 13394 2446
rect 13411 2382 13475 2446
rect 13492 2382 13556 2446
rect 13573 2382 13637 2446
rect 13654 2382 13718 2446
rect 13735 2382 13799 2446
rect 13816 2382 13880 2446
rect 13897 2382 13961 2446
rect 13978 2382 14042 2446
rect 14059 2382 14123 2446
rect 14140 2382 14204 2446
rect 14221 2382 14285 2446
rect 14302 2382 14366 2446
rect 14383 2382 14447 2446
rect 14464 2382 14528 2446
rect 14545 2382 14609 2446
rect 14626 2382 14690 2446
rect 14707 2382 14771 2446
rect 14788 2382 14852 2446
rect 105 2296 169 2360
rect 187 2296 251 2360
rect 269 2296 333 2360
rect 351 2296 415 2360
rect 433 2296 497 2360
rect 515 2296 579 2360
rect 597 2296 661 2360
rect 678 2296 742 2360
rect 759 2296 823 2360
rect 840 2296 904 2360
rect 921 2296 985 2360
rect 1002 2296 1066 2360
rect 1083 2296 1147 2360
rect 1164 2296 1228 2360
rect 1245 2296 1309 2360
rect 1326 2296 1390 2360
rect 1407 2296 1471 2360
rect 1488 2296 1552 2360
rect 1569 2296 1633 2360
rect 1650 2296 1714 2360
rect 1731 2296 1795 2360
rect 1812 2296 1876 2360
rect 1893 2296 1957 2360
rect 1974 2296 2038 2360
rect 2055 2296 2119 2360
rect 2136 2296 2200 2360
rect 2217 2296 2281 2360
rect 2298 2296 2362 2360
rect 2379 2296 2443 2360
rect 2460 2296 2524 2360
rect 2541 2296 2605 2360
rect 2622 2296 2686 2360
rect 2703 2296 2767 2360
rect 2784 2296 2848 2360
rect 2865 2296 2929 2360
rect 2946 2296 3010 2360
rect 3027 2296 3091 2360
rect 3108 2296 3172 2360
rect 3189 2296 3253 2360
rect 3270 2296 3334 2360
rect 3351 2296 3415 2360
rect 3432 2296 3496 2360
rect 3513 2296 3577 2360
rect 3594 2296 3658 2360
rect 3675 2296 3739 2360
rect 3756 2296 3820 2360
rect 3837 2296 3901 2360
rect 3918 2296 3982 2360
rect 3999 2296 4063 2360
rect 4080 2296 4144 2360
rect 4161 2296 4225 2360
rect 4242 2296 4306 2360
rect 4323 2296 4387 2360
rect 4404 2296 4468 2360
rect 4485 2296 4549 2360
rect 4566 2296 4630 2360
rect 4647 2296 4711 2360
rect 4728 2296 4792 2360
rect 4809 2296 4873 2360
rect 10084 2296 10148 2360
rect 10166 2296 10230 2360
rect 10248 2296 10312 2360
rect 10330 2296 10394 2360
rect 10412 2296 10476 2360
rect 10494 2296 10558 2360
rect 10576 2296 10640 2360
rect 10657 2296 10721 2360
rect 10738 2296 10802 2360
rect 10819 2296 10883 2360
rect 10900 2296 10964 2360
rect 10981 2296 11045 2360
rect 11062 2296 11126 2360
rect 11143 2296 11207 2360
rect 11224 2296 11288 2360
rect 11305 2296 11369 2360
rect 11386 2296 11450 2360
rect 11467 2296 11531 2360
rect 11548 2296 11612 2360
rect 11629 2296 11693 2360
rect 11710 2296 11774 2360
rect 11791 2296 11855 2360
rect 11872 2296 11936 2360
rect 11953 2296 12017 2360
rect 12034 2296 12098 2360
rect 12115 2296 12179 2360
rect 12196 2296 12260 2360
rect 12277 2296 12341 2360
rect 12358 2296 12422 2360
rect 12439 2296 12503 2360
rect 12520 2296 12584 2360
rect 12601 2296 12665 2360
rect 12682 2296 12746 2360
rect 12763 2296 12827 2360
rect 12844 2296 12908 2360
rect 12925 2296 12989 2360
rect 13006 2296 13070 2360
rect 13087 2296 13151 2360
rect 13168 2296 13232 2360
rect 13249 2296 13313 2360
rect 13330 2296 13394 2360
rect 13411 2296 13475 2360
rect 13492 2296 13556 2360
rect 13573 2296 13637 2360
rect 13654 2296 13718 2360
rect 13735 2296 13799 2360
rect 13816 2296 13880 2360
rect 13897 2296 13961 2360
rect 13978 2296 14042 2360
rect 14059 2296 14123 2360
rect 14140 2296 14204 2360
rect 14221 2296 14285 2360
rect 14302 2296 14366 2360
rect 14383 2296 14447 2360
rect 14464 2296 14528 2360
rect 14545 2296 14609 2360
rect 14626 2296 14690 2360
rect 14707 2296 14771 2360
rect 14788 2296 14852 2360
rect 105 2210 169 2274
rect 187 2210 251 2274
rect 269 2210 333 2274
rect 351 2210 415 2274
rect 433 2210 497 2274
rect 515 2210 579 2274
rect 597 2210 661 2274
rect 678 2210 742 2274
rect 759 2210 823 2274
rect 840 2210 904 2274
rect 921 2210 985 2274
rect 1002 2210 1066 2274
rect 1083 2210 1147 2274
rect 1164 2210 1228 2274
rect 1245 2210 1309 2274
rect 1326 2210 1390 2274
rect 1407 2210 1471 2274
rect 1488 2210 1552 2274
rect 1569 2210 1633 2274
rect 1650 2210 1714 2274
rect 1731 2210 1795 2274
rect 1812 2210 1876 2274
rect 1893 2210 1957 2274
rect 1974 2210 2038 2274
rect 2055 2210 2119 2274
rect 2136 2210 2200 2274
rect 2217 2210 2281 2274
rect 2298 2210 2362 2274
rect 2379 2210 2443 2274
rect 2460 2210 2524 2274
rect 2541 2210 2605 2274
rect 2622 2210 2686 2274
rect 2703 2210 2767 2274
rect 2784 2210 2848 2274
rect 2865 2210 2929 2274
rect 2946 2210 3010 2274
rect 3027 2210 3091 2274
rect 3108 2210 3172 2274
rect 3189 2210 3253 2274
rect 3270 2210 3334 2274
rect 3351 2210 3415 2274
rect 3432 2210 3496 2274
rect 3513 2210 3577 2274
rect 3594 2210 3658 2274
rect 3675 2210 3739 2274
rect 3756 2210 3820 2274
rect 3837 2210 3901 2274
rect 3918 2210 3982 2274
rect 3999 2210 4063 2274
rect 4080 2210 4144 2274
rect 4161 2210 4225 2274
rect 4242 2210 4306 2274
rect 4323 2210 4387 2274
rect 4404 2210 4468 2274
rect 4485 2210 4549 2274
rect 4566 2210 4630 2274
rect 4647 2210 4711 2274
rect 4728 2210 4792 2274
rect 4809 2210 4873 2274
rect 10084 2210 10148 2274
rect 10166 2210 10230 2274
rect 10248 2210 10312 2274
rect 10330 2210 10394 2274
rect 10412 2210 10476 2274
rect 10494 2210 10558 2274
rect 10576 2210 10640 2274
rect 10657 2210 10721 2274
rect 10738 2210 10802 2274
rect 10819 2210 10883 2274
rect 10900 2210 10964 2274
rect 10981 2210 11045 2274
rect 11062 2210 11126 2274
rect 11143 2210 11207 2274
rect 11224 2210 11288 2274
rect 11305 2210 11369 2274
rect 11386 2210 11450 2274
rect 11467 2210 11531 2274
rect 11548 2210 11612 2274
rect 11629 2210 11693 2274
rect 11710 2210 11774 2274
rect 11791 2210 11855 2274
rect 11872 2210 11936 2274
rect 11953 2210 12017 2274
rect 12034 2210 12098 2274
rect 12115 2210 12179 2274
rect 12196 2210 12260 2274
rect 12277 2210 12341 2274
rect 12358 2210 12422 2274
rect 12439 2210 12503 2274
rect 12520 2210 12584 2274
rect 12601 2210 12665 2274
rect 12682 2210 12746 2274
rect 12763 2210 12827 2274
rect 12844 2210 12908 2274
rect 12925 2210 12989 2274
rect 13006 2210 13070 2274
rect 13087 2210 13151 2274
rect 13168 2210 13232 2274
rect 13249 2210 13313 2274
rect 13330 2210 13394 2274
rect 13411 2210 13475 2274
rect 13492 2210 13556 2274
rect 13573 2210 13637 2274
rect 13654 2210 13718 2274
rect 13735 2210 13799 2274
rect 13816 2210 13880 2274
rect 13897 2210 13961 2274
rect 13978 2210 14042 2274
rect 14059 2210 14123 2274
rect 14140 2210 14204 2274
rect 14221 2210 14285 2274
rect 14302 2210 14366 2274
rect 14383 2210 14447 2274
rect 14464 2210 14528 2274
rect 14545 2210 14609 2274
rect 14626 2210 14690 2274
rect 14707 2210 14771 2274
rect 14788 2210 14852 2274
rect 105 2124 169 2188
rect 187 2124 251 2188
rect 269 2124 333 2188
rect 351 2124 415 2188
rect 433 2124 497 2188
rect 515 2124 579 2188
rect 597 2124 661 2188
rect 678 2124 742 2188
rect 759 2124 823 2188
rect 840 2124 904 2188
rect 921 2124 985 2188
rect 1002 2124 1066 2188
rect 1083 2124 1147 2188
rect 1164 2124 1228 2188
rect 1245 2124 1309 2188
rect 1326 2124 1390 2188
rect 1407 2124 1471 2188
rect 1488 2124 1552 2188
rect 1569 2124 1633 2188
rect 1650 2124 1714 2188
rect 1731 2124 1795 2188
rect 1812 2124 1876 2188
rect 1893 2124 1957 2188
rect 1974 2124 2038 2188
rect 2055 2124 2119 2188
rect 2136 2124 2200 2188
rect 2217 2124 2281 2188
rect 2298 2124 2362 2188
rect 2379 2124 2443 2188
rect 2460 2124 2524 2188
rect 2541 2124 2605 2188
rect 2622 2124 2686 2188
rect 2703 2124 2767 2188
rect 2784 2124 2848 2188
rect 2865 2124 2929 2188
rect 2946 2124 3010 2188
rect 3027 2124 3091 2188
rect 3108 2124 3172 2188
rect 3189 2124 3253 2188
rect 3270 2124 3334 2188
rect 3351 2124 3415 2188
rect 3432 2124 3496 2188
rect 3513 2124 3577 2188
rect 3594 2124 3658 2188
rect 3675 2124 3739 2188
rect 3756 2124 3820 2188
rect 3837 2124 3901 2188
rect 3918 2124 3982 2188
rect 3999 2124 4063 2188
rect 4080 2124 4144 2188
rect 4161 2124 4225 2188
rect 4242 2124 4306 2188
rect 4323 2124 4387 2188
rect 4404 2124 4468 2188
rect 4485 2124 4549 2188
rect 4566 2124 4630 2188
rect 4647 2124 4711 2188
rect 4728 2124 4792 2188
rect 4809 2124 4873 2188
rect 10084 2124 10148 2188
rect 10166 2124 10230 2188
rect 10248 2124 10312 2188
rect 10330 2124 10394 2188
rect 10412 2124 10476 2188
rect 10494 2124 10558 2188
rect 10576 2124 10640 2188
rect 10657 2124 10721 2188
rect 10738 2124 10802 2188
rect 10819 2124 10883 2188
rect 10900 2124 10964 2188
rect 10981 2124 11045 2188
rect 11062 2124 11126 2188
rect 11143 2124 11207 2188
rect 11224 2124 11288 2188
rect 11305 2124 11369 2188
rect 11386 2124 11450 2188
rect 11467 2124 11531 2188
rect 11548 2124 11612 2188
rect 11629 2124 11693 2188
rect 11710 2124 11774 2188
rect 11791 2124 11855 2188
rect 11872 2124 11936 2188
rect 11953 2124 12017 2188
rect 12034 2124 12098 2188
rect 12115 2124 12179 2188
rect 12196 2124 12260 2188
rect 12277 2124 12341 2188
rect 12358 2124 12422 2188
rect 12439 2124 12503 2188
rect 12520 2124 12584 2188
rect 12601 2124 12665 2188
rect 12682 2124 12746 2188
rect 12763 2124 12827 2188
rect 12844 2124 12908 2188
rect 12925 2124 12989 2188
rect 13006 2124 13070 2188
rect 13087 2124 13151 2188
rect 13168 2124 13232 2188
rect 13249 2124 13313 2188
rect 13330 2124 13394 2188
rect 13411 2124 13475 2188
rect 13492 2124 13556 2188
rect 13573 2124 13637 2188
rect 13654 2124 13718 2188
rect 13735 2124 13799 2188
rect 13816 2124 13880 2188
rect 13897 2124 13961 2188
rect 13978 2124 14042 2188
rect 14059 2124 14123 2188
rect 14140 2124 14204 2188
rect 14221 2124 14285 2188
rect 14302 2124 14366 2188
rect 14383 2124 14447 2188
rect 14464 2124 14528 2188
rect 14545 2124 14609 2188
rect 14626 2124 14690 2188
rect 14707 2124 14771 2188
rect 14788 2124 14852 2188
rect 105 2038 169 2102
rect 187 2038 251 2102
rect 269 2038 333 2102
rect 351 2038 415 2102
rect 433 2038 497 2102
rect 515 2038 579 2102
rect 597 2038 661 2102
rect 678 2038 742 2102
rect 759 2038 823 2102
rect 840 2038 904 2102
rect 921 2038 985 2102
rect 1002 2038 1066 2102
rect 1083 2038 1147 2102
rect 1164 2038 1228 2102
rect 1245 2038 1309 2102
rect 1326 2038 1390 2102
rect 1407 2038 1471 2102
rect 1488 2038 1552 2102
rect 1569 2038 1633 2102
rect 1650 2038 1714 2102
rect 1731 2038 1795 2102
rect 1812 2038 1876 2102
rect 1893 2038 1957 2102
rect 1974 2038 2038 2102
rect 2055 2038 2119 2102
rect 2136 2038 2200 2102
rect 2217 2038 2281 2102
rect 2298 2038 2362 2102
rect 2379 2038 2443 2102
rect 2460 2038 2524 2102
rect 2541 2038 2605 2102
rect 2622 2038 2686 2102
rect 2703 2038 2767 2102
rect 2784 2038 2848 2102
rect 2865 2038 2929 2102
rect 2946 2038 3010 2102
rect 3027 2038 3091 2102
rect 3108 2038 3172 2102
rect 3189 2038 3253 2102
rect 3270 2038 3334 2102
rect 3351 2038 3415 2102
rect 3432 2038 3496 2102
rect 3513 2038 3577 2102
rect 3594 2038 3658 2102
rect 3675 2038 3739 2102
rect 3756 2038 3820 2102
rect 3837 2038 3901 2102
rect 3918 2038 3982 2102
rect 3999 2038 4063 2102
rect 4080 2038 4144 2102
rect 4161 2038 4225 2102
rect 4242 2038 4306 2102
rect 4323 2038 4387 2102
rect 4404 2038 4468 2102
rect 4485 2038 4549 2102
rect 4566 2038 4630 2102
rect 4647 2038 4711 2102
rect 4728 2038 4792 2102
rect 4809 2038 4873 2102
rect 10084 2038 10148 2102
rect 10166 2038 10230 2102
rect 10248 2038 10312 2102
rect 10330 2038 10394 2102
rect 10412 2038 10476 2102
rect 10494 2038 10558 2102
rect 10576 2038 10640 2102
rect 10657 2038 10721 2102
rect 10738 2038 10802 2102
rect 10819 2038 10883 2102
rect 10900 2038 10964 2102
rect 10981 2038 11045 2102
rect 11062 2038 11126 2102
rect 11143 2038 11207 2102
rect 11224 2038 11288 2102
rect 11305 2038 11369 2102
rect 11386 2038 11450 2102
rect 11467 2038 11531 2102
rect 11548 2038 11612 2102
rect 11629 2038 11693 2102
rect 11710 2038 11774 2102
rect 11791 2038 11855 2102
rect 11872 2038 11936 2102
rect 11953 2038 12017 2102
rect 12034 2038 12098 2102
rect 12115 2038 12179 2102
rect 12196 2038 12260 2102
rect 12277 2038 12341 2102
rect 12358 2038 12422 2102
rect 12439 2038 12503 2102
rect 12520 2038 12584 2102
rect 12601 2038 12665 2102
rect 12682 2038 12746 2102
rect 12763 2038 12827 2102
rect 12844 2038 12908 2102
rect 12925 2038 12989 2102
rect 13006 2038 13070 2102
rect 13087 2038 13151 2102
rect 13168 2038 13232 2102
rect 13249 2038 13313 2102
rect 13330 2038 13394 2102
rect 13411 2038 13475 2102
rect 13492 2038 13556 2102
rect 13573 2038 13637 2102
rect 13654 2038 13718 2102
rect 13735 2038 13799 2102
rect 13816 2038 13880 2102
rect 13897 2038 13961 2102
rect 13978 2038 14042 2102
rect 14059 2038 14123 2102
rect 14140 2038 14204 2102
rect 14221 2038 14285 2102
rect 14302 2038 14366 2102
rect 14383 2038 14447 2102
rect 14464 2038 14528 2102
rect 14545 2038 14609 2102
rect 14626 2038 14690 2102
rect 14707 2038 14771 2102
rect 14788 2038 14852 2102
rect 105 1952 169 2016
rect 187 1952 251 2016
rect 269 1952 333 2016
rect 351 1952 415 2016
rect 433 1952 497 2016
rect 515 1952 579 2016
rect 597 1952 661 2016
rect 678 1952 742 2016
rect 759 1952 823 2016
rect 840 1952 904 2016
rect 921 1952 985 2016
rect 1002 1952 1066 2016
rect 1083 1952 1147 2016
rect 1164 1952 1228 2016
rect 1245 1952 1309 2016
rect 1326 1952 1390 2016
rect 1407 1952 1471 2016
rect 1488 1952 1552 2016
rect 1569 1952 1633 2016
rect 1650 1952 1714 2016
rect 1731 1952 1795 2016
rect 1812 1952 1876 2016
rect 1893 1952 1957 2016
rect 1974 1952 2038 2016
rect 2055 1952 2119 2016
rect 2136 1952 2200 2016
rect 2217 1952 2281 2016
rect 2298 1952 2362 2016
rect 2379 1952 2443 2016
rect 2460 1952 2524 2016
rect 2541 1952 2605 2016
rect 2622 1952 2686 2016
rect 2703 1952 2767 2016
rect 2784 1952 2848 2016
rect 2865 1952 2929 2016
rect 2946 1952 3010 2016
rect 3027 1952 3091 2016
rect 3108 1952 3172 2016
rect 3189 1952 3253 2016
rect 3270 1952 3334 2016
rect 3351 1952 3415 2016
rect 3432 1952 3496 2016
rect 3513 1952 3577 2016
rect 3594 1952 3658 2016
rect 3675 1952 3739 2016
rect 3756 1952 3820 2016
rect 3837 1952 3901 2016
rect 3918 1952 3982 2016
rect 3999 1952 4063 2016
rect 4080 1952 4144 2016
rect 4161 1952 4225 2016
rect 4242 1952 4306 2016
rect 4323 1952 4387 2016
rect 4404 1952 4468 2016
rect 4485 1952 4549 2016
rect 4566 1952 4630 2016
rect 4647 1952 4711 2016
rect 4728 1952 4792 2016
rect 4809 1952 4873 2016
rect 10084 1952 10148 2016
rect 10166 1952 10230 2016
rect 10248 1952 10312 2016
rect 10330 1952 10394 2016
rect 10412 1952 10476 2016
rect 10494 1952 10558 2016
rect 10576 1952 10640 2016
rect 10657 1952 10721 2016
rect 10738 1952 10802 2016
rect 10819 1952 10883 2016
rect 10900 1952 10964 2016
rect 10981 1952 11045 2016
rect 11062 1952 11126 2016
rect 11143 1952 11207 2016
rect 11224 1952 11288 2016
rect 11305 1952 11369 2016
rect 11386 1952 11450 2016
rect 11467 1952 11531 2016
rect 11548 1952 11612 2016
rect 11629 1952 11693 2016
rect 11710 1952 11774 2016
rect 11791 1952 11855 2016
rect 11872 1952 11936 2016
rect 11953 1952 12017 2016
rect 12034 1952 12098 2016
rect 12115 1952 12179 2016
rect 12196 1952 12260 2016
rect 12277 1952 12341 2016
rect 12358 1952 12422 2016
rect 12439 1952 12503 2016
rect 12520 1952 12584 2016
rect 12601 1952 12665 2016
rect 12682 1952 12746 2016
rect 12763 1952 12827 2016
rect 12844 1952 12908 2016
rect 12925 1952 12989 2016
rect 13006 1952 13070 2016
rect 13087 1952 13151 2016
rect 13168 1952 13232 2016
rect 13249 1952 13313 2016
rect 13330 1952 13394 2016
rect 13411 1952 13475 2016
rect 13492 1952 13556 2016
rect 13573 1952 13637 2016
rect 13654 1952 13718 2016
rect 13735 1952 13799 2016
rect 13816 1952 13880 2016
rect 13897 1952 13961 2016
rect 13978 1952 14042 2016
rect 14059 1952 14123 2016
rect 14140 1952 14204 2016
rect 14221 1952 14285 2016
rect 14302 1952 14366 2016
rect 14383 1952 14447 2016
rect 14464 1952 14528 2016
rect 14545 1952 14609 2016
rect 14626 1952 14690 2016
rect 14707 1952 14771 2016
rect 14788 1952 14852 2016
rect 105 1866 169 1930
rect 187 1866 251 1930
rect 269 1866 333 1930
rect 351 1866 415 1930
rect 433 1866 497 1930
rect 515 1866 579 1930
rect 597 1866 661 1930
rect 678 1866 742 1930
rect 759 1866 823 1930
rect 840 1866 904 1930
rect 921 1866 985 1930
rect 1002 1866 1066 1930
rect 1083 1866 1147 1930
rect 1164 1866 1228 1930
rect 1245 1866 1309 1930
rect 1326 1866 1390 1930
rect 1407 1866 1471 1930
rect 1488 1866 1552 1930
rect 1569 1866 1633 1930
rect 1650 1866 1714 1930
rect 1731 1866 1795 1930
rect 1812 1866 1876 1930
rect 1893 1866 1957 1930
rect 1974 1866 2038 1930
rect 2055 1866 2119 1930
rect 2136 1866 2200 1930
rect 2217 1866 2281 1930
rect 2298 1866 2362 1930
rect 2379 1866 2443 1930
rect 2460 1866 2524 1930
rect 2541 1866 2605 1930
rect 2622 1866 2686 1930
rect 2703 1866 2767 1930
rect 2784 1866 2848 1930
rect 2865 1866 2929 1930
rect 2946 1866 3010 1930
rect 3027 1866 3091 1930
rect 3108 1866 3172 1930
rect 3189 1866 3253 1930
rect 3270 1866 3334 1930
rect 3351 1866 3415 1930
rect 3432 1866 3496 1930
rect 3513 1866 3577 1930
rect 3594 1866 3658 1930
rect 3675 1866 3739 1930
rect 3756 1866 3820 1930
rect 3837 1866 3901 1930
rect 3918 1866 3982 1930
rect 3999 1866 4063 1930
rect 4080 1866 4144 1930
rect 4161 1866 4225 1930
rect 4242 1866 4306 1930
rect 4323 1866 4387 1930
rect 4404 1866 4468 1930
rect 4485 1866 4549 1930
rect 4566 1866 4630 1930
rect 4647 1866 4711 1930
rect 4728 1866 4792 1930
rect 4809 1866 4873 1930
rect 10084 1866 10148 1930
rect 10166 1866 10230 1930
rect 10248 1866 10312 1930
rect 10330 1866 10394 1930
rect 10412 1866 10476 1930
rect 10494 1866 10558 1930
rect 10576 1866 10640 1930
rect 10657 1866 10721 1930
rect 10738 1866 10802 1930
rect 10819 1866 10883 1930
rect 10900 1866 10964 1930
rect 10981 1866 11045 1930
rect 11062 1866 11126 1930
rect 11143 1866 11207 1930
rect 11224 1866 11288 1930
rect 11305 1866 11369 1930
rect 11386 1866 11450 1930
rect 11467 1866 11531 1930
rect 11548 1866 11612 1930
rect 11629 1866 11693 1930
rect 11710 1866 11774 1930
rect 11791 1866 11855 1930
rect 11872 1866 11936 1930
rect 11953 1866 12017 1930
rect 12034 1866 12098 1930
rect 12115 1866 12179 1930
rect 12196 1866 12260 1930
rect 12277 1866 12341 1930
rect 12358 1866 12422 1930
rect 12439 1866 12503 1930
rect 12520 1866 12584 1930
rect 12601 1866 12665 1930
rect 12682 1866 12746 1930
rect 12763 1866 12827 1930
rect 12844 1866 12908 1930
rect 12925 1866 12989 1930
rect 13006 1866 13070 1930
rect 13087 1866 13151 1930
rect 13168 1866 13232 1930
rect 13249 1866 13313 1930
rect 13330 1866 13394 1930
rect 13411 1866 13475 1930
rect 13492 1866 13556 1930
rect 13573 1866 13637 1930
rect 13654 1866 13718 1930
rect 13735 1866 13799 1930
rect 13816 1866 13880 1930
rect 13897 1866 13961 1930
rect 13978 1866 14042 1930
rect 14059 1866 14123 1930
rect 14140 1866 14204 1930
rect 14221 1866 14285 1930
rect 14302 1866 14366 1930
rect 14383 1866 14447 1930
rect 14464 1866 14528 1930
rect 14545 1866 14609 1930
rect 14626 1866 14690 1930
rect 14707 1866 14771 1930
rect 14788 1866 14852 1930
rect 105 1780 169 1844
rect 187 1780 251 1844
rect 269 1780 333 1844
rect 351 1780 415 1844
rect 433 1780 497 1844
rect 515 1780 579 1844
rect 597 1780 661 1844
rect 678 1780 742 1844
rect 759 1780 823 1844
rect 840 1780 904 1844
rect 921 1780 985 1844
rect 1002 1780 1066 1844
rect 1083 1780 1147 1844
rect 1164 1780 1228 1844
rect 1245 1780 1309 1844
rect 1326 1780 1390 1844
rect 1407 1780 1471 1844
rect 1488 1780 1552 1844
rect 1569 1780 1633 1844
rect 1650 1780 1714 1844
rect 1731 1780 1795 1844
rect 1812 1780 1876 1844
rect 1893 1780 1957 1844
rect 1974 1780 2038 1844
rect 2055 1780 2119 1844
rect 2136 1780 2200 1844
rect 2217 1780 2281 1844
rect 2298 1780 2362 1844
rect 2379 1780 2443 1844
rect 2460 1780 2524 1844
rect 2541 1780 2605 1844
rect 2622 1780 2686 1844
rect 2703 1780 2767 1844
rect 2784 1780 2848 1844
rect 2865 1780 2929 1844
rect 2946 1780 3010 1844
rect 3027 1780 3091 1844
rect 3108 1780 3172 1844
rect 3189 1780 3253 1844
rect 3270 1780 3334 1844
rect 3351 1780 3415 1844
rect 3432 1780 3496 1844
rect 3513 1780 3577 1844
rect 3594 1780 3658 1844
rect 3675 1780 3739 1844
rect 3756 1780 3820 1844
rect 3837 1780 3901 1844
rect 3918 1780 3982 1844
rect 3999 1780 4063 1844
rect 4080 1780 4144 1844
rect 4161 1780 4225 1844
rect 4242 1780 4306 1844
rect 4323 1780 4387 1844
rect 4404 1780 4468 1844
rect 4485 1780 4549 1844
rect 4566 1780 4630 1844
rect 4647 1780 4711 1844
rect 4728 1780 4792 1844
rect 4809 1780 4873 1844
rect 10084 1780 10148 1844
rect 10166 1780 10230 1844
rect 10248 1780 10312 1844
rect 10330 1780 10394 1844
rect 10412 1780 10476 1844
rect 10494 1780 10558 1844
rect 10576 1780 10640 1844
rect 10657 1780 10721 1844
rect 10738 1780 10802 1844
rect 10819 1780 10883 1844
rect 10900 1780 10964 1844
rect 10981 1780 11045 1844
rect 11062 1780 11126 1844
rect 11143 1780 11207 1844
rect 11224 1780 11288 1844
rect 11305 1780 11369 1844
rect 11386 1780 11450 1844
rect 11467 1780 11531 1844
rect 11548 1780 11612 1844
rect 11629 1780 11693 1844
rect 11710 1780 11774 1844
rect 11791 1780 11855 1844
rect 11872 1780 11936 1844
rect 11953 1780 12017 1844
rect 12034 1780 12098 1844
rect 12115 1780 12179 1844
rect 12196 1780 12260 1844
rect 12277 1780 12341 1844
rect 12358 1780 12422 1844
rect 12439 1780 12503 1844
rect 12520 1780 12584 1844
rect 12601 1780 12665 1844
rect 12682 1780 12746 1844
rect 12763 1780 12827 1844
rect 12844 1780 12908 1844
rect 12925 1780 12989 1844
rect 13006 1780 13070 1844
rect 13087 1780 13151 1844
rect 13168 1780 13232 1844
rect 13249 1780 13313 1844
rect 13330 1780 13394 1844
rect 13411 1780 13475 1844
rect 13492 1780 13556 1844
rect 13573 1780 13637 1844
rect 13654 1780 13718 1844
rect 13735 1780 13799 1844
rect 13816 1780 13880 1844
rect 13897 1780 13961 1844
rect 13978 1780 14042 1844
rect 14059 1780 14123 1844
rect 14140 1780 14204 1844
rect 14221 1780 14285 1844
rect 14302 1780 14366 1844
rect 14383 1780 14447 1844
rect 14464 1780 14528 1844
rect 14545 1780 14609 1844
rect 14626 1780 14690 1844
rect 14707 1780 14771 1844
rect 14788 1780 14852 1844
<< obsm4 >>
rect 0 11301 15000 40000
rect 0 10349 15000 10545
rect 0 2704 15000 9593
rect 0 2640 105 2704
rect 169 2640 187 2704
rect 251 2640 269 2704
rect 333 2640 351 2704
rect 415 2640 433 2704
rect 497 2640 515 2704
rect 579 2640 597 2704
rect 661 2640 678 2704
rect 742 2640 759 2704
rect 823 2640 840 2704
rect 904 2640 921 2704
rect 985 2640 1002 2704
rect 1066 2640 1083 2704
rect 1147 2640 1164 2704
rect 1228 2640 1245 2704
rect 1309 2640 1326 2704
rect 1390 2640 1407 2704
rect 1471 2640 1488 2704
rect 1552 2640 1569 2704
rect 1633 2640 1650 2704
rect 1714 2640 1731 2704
rect 1795 2640 1812 2704
rect 1876 2640 1893 2704
rect 1957 2640 1974 2704
rect 2038 2640 2055 2704
rect 2119 2640 2136 2704
rect 2200 2640 2217 2704
rect 2281 2640 2298 2704
rect 2362 2640 2379 2704
rect 2443 2640 2460 2704
rect 2524 2640 2541 2704
rect 2605 2640 2622 2704
rect 2686 2640 2703 2704
rect 2767 2640 2784 2704
rect 2848 2640 2865 2704
rect 2929 2640 2946 2704
rect 3010 2640 3027 2704
rect 3091 2640 3108 2704
rect 3172 2640 3189 2704
rect 3253 2640 3270 2704
rect 3334 2640 3351 2704
rect 3415 2640 3432 2704
rect 3496 2640 3513 2704
rect 3577 2640 3594 2704
rect 3658 2640 3675 2704
rect 3739 2640 3756 2704
rect 3820 2640 3837 2704
rect 3901 2640 3918 2704
rect 3982 2640 3999 2704
rect 4063 2640 4080 2704
rect 4144 2640 4161 2704
rect 4225 2640 4242 2704
rect 4306 2640 4323 2704
rect 4387 2640 4404 2704
rect 4468 2640 4485 2704
rect 4549 2640 4566 2704
rect 4630 2640 4647 2704
rect 4711 2640 4728 2704
rect 4792 2640 4809 2704
rect 4873 2640 10084 2704
rect 10148 2640 10166 2704
rect 10230 2640 10248 2704
rect 10312 2640 10330 2704
rect 10394 2640 10412 2704
rect 10476 2640 10494 2704
rect 10558 2640 10576 2704
rect 10640 2640 10657 2704
rect 10721 2640 10738 2704
rect 10802 2640 10819 2704
rect 10883 2640 10900 2704
rect 10964 2640 10981 2704
rect 11045 2640 11062 2704
rect 11126 2640 11143 2704
rect 11207 2640 11224 2704
rect 11288 2640 11305 2704
rect 11369 2640 11386 2704
rect 11450 2640 11467 2704
rect 11531 2640 11548 2704
rect 11612 2640 11629 2704
rect 11693 2640 11710 2704
rect 11774 2640 11791 2704
rect 11855 2640 11872 2704
rect 11936 2640 11953 2704
rect 12017 2640 12034 2704
rect 12098 2640 12115 2704
rect 12179 2640 12196 2704
rect 12260 2640 12277 2704
rect 12341 2640 12358 2704
rect 12422 2640 12439 2704
rect 12503 2640 12520 2704
rect 12584 2640 12601 2704
rect 12665 2640 12682 2704
rect 12746 2640 12763 2704
rect 12827 2640 12844 2704
rect 12908 2640 12925 2704
rect 12989 2640 13006 2704
rect 13070 2640 13087 2704
rect 13151 2640 13168 2704
rect 13232 2640 13249 2704
rect 13313 2640 13330 2704
rect 13394 2640 13411 2704
rect 13475 2640 13492 2704
rect 13556 2640 13573 2704
rect 13637 2640 13654 2704
rect 13718 2640 13735 2704
rect 13799 2640 13816 2704
rect 13880 2640 13897 2704
rect 13961 2640 13978 2704
rect 14042 2640 14059 2704
rect 14123 2640 14140 2704
rect 14204 2640 14221 2704
rect 14285 2640 14302 2704
rect 14366 2640 14383 2704
rect 14447 2640 14464 2704
rect 14528 2640 14545 2704
rect 14609 2640 14626 2704
rect 14690 2640 14707 2704
rect 14771 2640 14788 2704
rect 14852 2640 15000 2704
rect 0 2618 15000 2640
rect 0 2554 105 2618
rect 169 2554 187 2618
rect 251 2554 269 2618
rect 333 2554 351 2618
rect 415 2554 433 2618
rect 497 2554 515 2618
rect 579 2554 597 2618
rect 661 2554 678 2618
rect 742 2554 759 2618
rect 823 2554 840 2618
rect 904 2554 921 2618
rect 985 2554 1002 2618
rect 1066 2554 1083 2618
rect 1147 2554 1164 2618
rect 1228 2554 1245 2618
rect 1309 2554 1326 2618
rect 1390 2554 1407 2618
rect 1471 2554 1488 2618
rect 1552 2554 1569 2618
rect 1633 2554 1650 2618
rect 1714 2554 1731 2618
rect 1795 2554 1812 2618
rect 1876 2554 1893 2618
rect 1957 2554 1974 2618
rect 2038 2554 2055 2618
rect 2119 2554 2136 2618
rect 2200 2554 2217 2618
rect 2281 2554 2298 2618
rect 2362 2554 2379 2618
rect 2443 2554 2460 2618
rect 2524 2554 2541 2618
rect 2605 2554 2622 2618
rect 2686 2554 2703 2618
rect 2767 2554 2784 2618
rect 2848 2554 2865 2618
rect 2929 2554 2946 2618
rect 3010 2554 3027 2618
rect 3091 2554 3108 2618
rect 3172 2554 3189 2618
rect 3253 2554 3270 2618
rect 3334 2554 3351 2618
rect 3415 2554 3432 2618
rect 3496 2554 3513 2618
rect 3577 2554 3594 2618
rect 3658 2554 3675 2618
rect 3739 2554 3756 2618
rect 3820 2554 3837 2618
rect 3901 2554 3918 2618
rect 3982 2554 3999 2618
rect 4063 2554 4080 2618
rect 4144 2554 4161 2618
rect 4225 2554 4242 2618
rect 4306 2554 4323 2618
rect 4387 2554 4404 2618
rect 4468 2554 4485 2618
rect 4549 2554 4566 2618
rect 4630 2554 4647 2618
rect 4711 2554 4728 2618
rect 4792 2554 4809 2618
rect 4873 2554 10084 2618
rect 10148 2554 10166 2618
rect 10230 2554 10248 2618
rect 10312 2554 10330 2618
rect 10394 2554 10412 2618
rect 10476 2554 10494 2618
rect 10558 2554 10576 2618
rect 10640 2554 10657 2618
rect 10721 2554 10738 2618
rect 10802 2554 10819 2618
rect 10883 2554 10900 2618
rect 10964 2554 10981 2618
rect 11045 2554 11062 2618
rect 11126 2554 11143 2618
rect 11207 2554 11224 2618
rect 11288 2554 11305 2618
rect 11369 2554 11386 2618
rect 11450 2554 11467 2618
rect 11531 2554 11548 2618
rect 11612 2554 11629 2618
rect 11693 2554 11710 2618
rect 11774 2554 11791 2618
rect 11855 2554 11872 2618
rect 11936 2554 11953 2618
rect 12017 2554 12034 2618
rect 12098 2554 12115 2618
rect 12179 2554 12196 2618
rect 12260 2554 12277 2618
rect 12341 2554 12358 2618
rect 12422 2554 12439 2618
rect 12503 2554 12520 2618
rect 12584 2554 12601 2618
rect 12665 2554 12682 2618
rect 12746 2554 12763 2618
rect 12827 2554 12844 2618
rect 12908 2554 12925 2618
rect 12989 2554 13006 2618
rect 13070 2554 13087 2618
rect 13151 2554 13168 2618
rect 13232 2554 13249 2618
rect 13313 2554 13330 2618
rect 13394 2554 13411 2618
rect 13475 2554 13492 2618
rect 13556 2554 13573 2618
rect 13637 2554 13654 2618
rect 13718 2554 13735 2618
rect 13799 2554 13816 2618
rect 13880 2554 13897 2618
rect 13961 2554 13978 2618
rect 14042 2554 14059 2618
rect 14123 2554 14140 2618
rect 14204 2554 14221 2618
rect 14285 2554 14302 2618
rect 14366 2554 14383 2618
rect 14447 2554 14464 2618
rect 14528 2554 14545 2618
rect 14609 2554 14626 2618
rect 14690 2554 14707 2618
rect 14771 2554 14788 2618
rect 14852 2554 15000 2618
rect 0 2532 15000 2554
rect 0 2468 105 2532
rect 169 2468 187 2532
rect 251 2468 269 2532
rect 333 2468 351 2532
rect 415 2468 433 2532
rect 497 2468 515 2532
rect 579 2468 597 2532
rect 661 2468 678 2532
rect 742 2468 759 2532
rect 823 2468 840 2532
rect 904 2468 921 2532
rect 985 2468 1002 2532
rect 1066 2468 1083 2532
rect 1147 2468 1164 2532
rect 1228 2468 1245 2532
rect 1309 2468 1326 2532
rect 1390 2468 1407 2532
rect 1471 2468 1488 2532
rect 1552 2468 1569 2532
rect 1633 2468 1650 2532
rect 1714 2468 1731 2532
rect 1795 2468 1812 2532
rect 1876 2468 1893 2532
rect 1957 2468 1974 2532
rect 2038 2468 2055 2532
rect 2119 2468 2136 2532
rect 2200 2468 2217 2532
rect 2281 2468 2298 2532
rect 2362 2468 2379 2532
rect 2443 2468 2460 2532
rect 2524 2468 2541 2532
rect 2605 2468 2622 2532
rect 2686 2468 2703 2532
rect 2767 2468 2784 2532
rect 2848 2468 2865 2532
rect 2929 2468 2946 2532
rect 3010 2468 3027 2532
rect 3091 2468 3108 2532
rect 3172 2468 3189 2532
rect 3253 2468 3270 2532
rect 3334 2468 3351 2532
rect 3415 2468 3432 2532
rect 3496 2468 3513 2532
rect 3577 2468 3594 2532
rect 3658 2468 3675 2532
rect 3739 2468 3756 2532
rect 3820 2468 3837 2532
rect 3901 2468 3918 2532
rect 3982 2468 3999 2532
rect 4063 2468 4080 2532
rect 4144 2468 4161 2532
rect 4225 2468 4242 2532
rect 4306 2468 4323 2532
rect 4387 2468 4404 2532
rect 4468 2468 4485 2532
rect 4549 2468 4566 2532
rect 4630 2468 4647 2532
rect 4711 2468 4728 2532
rect 4792 2468 4809 2532
rect 4873 2468 10084 2532
rect 10148 2468 10166 2532
rect 10230 2468 10248 2532
rect 10312 2468 10330 2532
rect 10394 2468 10412 2532
rect 10476 2468 10494 2532
rect 10558 2468 10576 2532
rect 10640 2468 10657 2532
rect 10721 2468 10738 2532
rect 10802 2468 10819 2532
rect 10883 2468 10900 2532
rect 10964 2468 10981 2532
rect 11045 2468 11062 2532
rect 11126 2468 11143 2532
rect 11207 2468 11224 2532
rect 11288 2468 11305 2532
rect 11369 2468 11386 2532
rect 11450 2468 11467 2532
rect 11531 2468 11548 2532
rect 11612 2468 11629 2532
rect 11693 2468 11710 2532
rect 11774 2468 11791 2532
rect 11855 2468 11872 2532
rect 11936 2468 11953 2532
rect 12017 2468 12034 2532
rect 12098 2468 12115 2532
rect 12179 2468 12196 2532
rect 12260 2468 12277 2532
rect 12341 2468 12358 2532
rect 12422 2468 12439 2532
rect 12503 2468 12520 2532
rect 12584 2468 12601 2532
rect 12665 2468 12682 2532
rect 12746 2468 12763 2532
rect 12827 2468 12844 2532
rect 12908 2468 12925 2532
rect 12989 2468 13006 2532
rect 13070 2468 13087 2532
rect 13151 2468 13168 2532
rect 13232 2468 13249 2532
rect 13313 2468 13330 2532
rect 13394 2468 13411 2532
rect 13475 2468 13492 2532
rect 13556 2468 13573 2532
rect 13637 2468 13654 2532
rect 13718 2468 13735 2532
rect 13799 2468 13816 2532
rect 13880 2468 13897 2532
rect 13961 2468 13978 2532
rect 14042 2468 14059 2532
rect 14123 2468 14140 2532
rect 14204 2468 14221 2532
rect 14285 2468 14302 2532
rect 14366 2468 14383 2532
rect 14447 2468 14464 2532
rect 14528 2468 14545 2532
rect 14609 2468 14626 2532
rect 14690 2468 14707 2532
rect 14771 2468 14788 2532
rect 14852 2468 15000 2532
rect 0 2446 15000 2468
rect 0 2382 105 2446
rect 169 2382 187 2446
rect 251 2382 269 2446
rect 333 2382 351 2446
rect 415 2382 433 2446
rect 497 2382 515 2446
rect 579 2382 597 2446
rect 661 2382 678 2446
rect 742 2382 759 2446
rect 823 2382 840 2446
rect 904 2382 921 2446
rect 985 2382 1002 2446
rect 1066 2382 1083 2446
rect 1147 2382 1164 2446
rect 1228 2382 1245 2446
rect 1309 2382 1326 2446
rect 1390 2382 1407 2446
rect 1471 2382 1488 2446
rect 1552 2382 1569 2446
rect 1633 2382 1650 2446
rect 1714 2382 1731 2446
rect 1795 2382 1812 2446
rect 1876 2382 1893 2446
rect 1957 2382 1974 2446
rect 2038 2382 2055 2446
rect 2119 2382 2136 2446
rect 2200 2382 2217 2446
rect 2281 2382 2298 2446
rect 2362 2382 2379 2446
rect 2443 2382 2460 2446
rect 2524 2382 2541 2446
rect 2605 2382 2622 2446
rect 2686 2382 2703 2446
rect 2767 2382 2784 2446
rect 2848 2382 2865 2446
rect 2929 2382 2946 2446
rect 3010 2382 3027 2446
rect 3091 2382 3108 2446
rect 3172 2382 3189 2446
rect 3253 2382 3270 2446
rect 3334 2382 3351 2446
rect 3415 2382 3432 2446
rect 3496 2382 3513 2446
rect 3577 2382 3594 2446
rect 3658 2382 3675 2446
rect 3739 2382 3756 2446
rect 3820 2382 3837 2446
rect 3901 2382 3918 2446
rect 3982 2382 3999 2446
rect 4063 2382 4080 2446
rect 4144 2382 4161 2446
rect 4225 2382 4242 2446
rect 4306 2382 4323 2446
rect 4387 2382 4404 2446
rect 4468 2382 4485 2446
rect 4549 2382 4566 2446
rect 4630 2382 4647 2446
rect 4711 2382 4728 2446
rect 4792 2382 4809 2446
rect 4873 2382 10084 2446
rect 10148 2382 10166 2446
rect 10230 2382 10248 2446
rect 10312 2382 10330 2446
rect 10394 2382 10412 2446
rect 10476 2382 10494 2446
rect 10558 2382 10576 2446
rect 10640 2382 10657 2446
rect 10721 2382 10738 2446
rect 10802 2382 10819 2446
rect 10883 2382 10900 2446
rect 10964 2382 10981 2446
rect 11045 2382 11062 2446
rect 11126 2382 11143 2446
rect 11207 2382 11224 2446
rect 11288 2382 11305 2446
rect 11369 2382 11386 2446
rect 11450 2382 11467 2446
rect 11531 2382 11548 2446
rect 11612 2382 11629 2446
rect 11693 2382 11710 2446
rect 11774 2382 11791 2446
rect 11855 2382 11872 2446
rect 11936 2382 11953 2446
rect 12017 2382 12034 2446
rect 12098 2382 12115 2446
rect 12179 2382 12196 2446
rect 12260 2382 12277 2446
rect 12341 2382 12358 2446
rect 12422 2382 12439 2446
rect 12503 2382 12520 2446
rect 12584 2382 12601 2446
rect 12665 2382 12682 2446
rect 12746 2382 12763 2446
rect 12827 2382 12844 2446
rect 12908 2382 12925 2446
rect 12989 2382 13006 2446
rect 13070 2382 13087 2446
rect 13151 2382 13168 2446
rect 13232 2382 13249 2446
rect 13313 2382 13330 2446
rect 13394 2382 13411 2446
rect 13475 2382 13492 2446
rect 13556 2382 13573 2446
rect 13637 2382 13654 2446
rect 13718 2382 13735 2446
rect 13799 2382 13816 2446
rect 13880 2382 13897 2446
rect 13961 2382 13978 2446
rect 14042 2382 14059 2446
rect 14123 2382 14140 2446
rect 14204 2382 14221 2446
rect 14285 2382 14302 2446
rect 14366 2382 14383 2446
rect 14447 2382 14464 2446
rect 14528 2382 14545 2446
rect 14609 2382 14626 2446
rect 14690 2382 14707 2446
rect 14771 2382 14788 2446
rect 14852 2382 15000 2446
rect 0 2360 15000 2382
rect 0 2296 105 2360
rect 169 2296 187 2360
rect 251 2296 269 2360
rect 333 2296 351 2360
rect 415 2296 433 2360
rect 497 2296 515 2360
rect 579 2296 597 2360
rect 661 2296 678 2360
rect 742 2296 759 2360
rect 823 2296 840 2360
rect 904 2296 921 2360
rect 985 2296 1002 2360
rect 1066 2296 1083 2360
rect 1147 2296 1164 2360
rect 1228 2296 1245 2360
rect 1309 2296 1326 2360
rect 1390 2296 1407 2360
rect 1471 2296 1488 2360
rect 1552 2296 1569 2360
rect 1633 2296 1650 2360
rect 1714 2296 1731 2360
rect 1795 2296 1812 2360
rect 1876 2296 1893 2360
rect 1957 2296 1974 2360
rect 2038 2296 2055 2360
rect 2119 2296 2136 2360
rect 2200 2296 2217 2360
rect 2281 2296 2298 2360
rect 2362 2296 2379 2360
rect 2443 2296 2460 2360
rect 2524 2296 2541 2360
rect 2605 2296 2622 2360
rect 2686 2296 2703 2360
rect 2767 2296 2784 2360
rect 2848 2296 2865 2360
rect 2929 2296 2946 2360
rect 3010 2296 3027 2360
rect 3091 2296 3108 2360
rect 3172 2296 3189 2360
rect 3253 2296 3270 2360
rect 3334 2296 3351 2360
rect 3415 2296 3432 2360
rect 3496 2296 3513 2360
rect 3577 2296 3594 2360
rect 3658 2296 3675 2360
rect 3739 2296 3756 2360
rect 3820 2296 3837 2360
rect 3901 2296 3918 2360
rect 3982 2296 3999 2360
rect 4063 2296 4080 2360
rect 4144 2296 4161 2360
rect 4225 2296 4242 2360
rect 4306 2296 4323 2360
rect 4387 2296 4404 2360
rect 4468 2296 4485 2360
rect 4549 2296 4566 2360
rect 4630 2296 4647 2360
rect 4711 2296 4728 2360
rect 4792 2296 4809 2360
rect 4873 2296 10084 2360
rect 10148 2296 10166 2360
rect 10230 2296 10248 2360
rect 10312 2296 10330 2360
rect 10394 2296 10412 2360
rect 10476 2296 10494 2360
rect 10558 2296 10576 2360
rect 10640 2296 10657 2360
rect 10721 2296 10738 2360
rect 10802 2296 10819 2360
rect 10883 2296 10900 2360
rect 10964 2296 10981 2360
rect 11045 2296 11062 2360
rect 11126 2296 11143 2360
rect 11207 2296 11224 2360
rect 11288 2296 11305 2360
rect 11369 2296 11386 2360
rect 11450 2296 11467 2360
rect 11531 2296 11548 2360
rect 11612 2296 11629 2360
rect 11693 2296 11710 2360
rect 11774 2296 11791 2360
rect 11855 2296 11872 2360
rect 11936 2296 11953 2360
rect 12017 2296 12034 2360
rect 12098 2296 12115 2360
rect 12179 2296 12196 2360
rect 12260 2296 12277 2360
rect 12341 2296 12358 2360
rect 12422 2296 12439 2360
rect 12503 2296 12520 2360
rect 12584 2296 12601 2360
rect 12665 2296 12682 2360
rect 12746 2296 12763 2360
rect 12827 2296 12844 2360
rect 12908 2296 12925 2360
rect 12989 2296 13006 2360
rect 13070 2296 13087 2360
rect 13151 2296 13168 2360
rect 13232 2296 13249 2360
rect 13313 2296 13330 2360
rect 13394 2296 13411 2360
rect 13475 2296 13492 2360
rect 13556 2296 13573 2360
rect 13637 2296 13654 2360
rect 13718 2296 13735 2360
rect 13799 2296 13816 2360
rect 13880 2296 13897 2360
rect 13961 2296 13978 2360
rect 14042 2296 14059 2360
rect 14123 2296 14140 2360
rect 14204 2296 14221 2360
rect 14285 2296 14302 2360
rect 14366 2296 14383 2360
rect 14447 2296 14464 2360
rect 14528 2296 14545 2360
rect 14609 2296 14626 2360
rect 14690 2296 14707 2360
rect 14771 2296 14788 2360
rect 14852 2296 15000 2360
rect 0 2274 15000 2296
rect 0 2210 105 2274
rect 169 2210 187 2274
rect 251 2210 269 2274
rect 333 2210 351 2274
rect 415 2210 433 2274
rect 497 2210 515 2274
rect 579 2210 597 2274
rect 661 2210 678 2274
rect 742 2210 759 2274
rect 823 2210 840 2274
rect 904 2210 921 2274
rect 985 2210 1002 2274
rect 1066 2210 1083 2274
rect 1147 2210 1164 2274
rect 1228 2210 1245 2274
rect 1309 2210 1326 2274
rect 1390 2210 1407 2274
rect 1471 2210 1488 2274
rect 1552 2210 1569 2274
rect 1633 2210 1650 2274
rect 1714 2210 1731 2274
rect 1795 2210 1812 2274
rect 1876 2210 1893 2274
rect 1957 2210 1974 2274
rect 2038 2210 2055 2274
rect 2119 2210 2136 2274
rect 2200 2210 2217 2274
rect 2281 2210 2298 2274
rect 2362 2210 2379 2274
rect 2443 2210 2460 2274
rect 2524 2210 2541 2274
rect 2605 2210 2622 2274
rect 2686 2210 2703 2274
rect 2767 2210 2784 2274
rect 2848 2210 2865 2274
rect 2929 2210 2946 2274
rect 3010 2210 3027 2274
rect 3091 2210 3108 2274
rect 3172 2210 3189 2274
rect 3253 2210 3270 2274
rect 3334 2210 3351 2274
rect 3415 2210 3432 2274
rect 3496 2210 3513 2274
rect 3577 2210 3594 2274
rect 3658 2210 3675 2274
rect 3739 2210 3756 2274
rect 3820 2210 3837 2274
rect 3901 2210 3918 2274
rect 3982 2210 3999 2274
rect 4063 2210 4080 2274
rect 4144 2210 4161 2274
rect 4225 2210 4242 2274
rect 4306 2210 4323 2274
rect 4387 2210 4404 2274
rect 4468 2210 4485 2274
rect 4549 2210 4566 2274
rect 4630 2210 4647 2274
rect 4711 2210 4728 2274
rect 4792 2210 4809 2274
rect 4873 2210 10084 2274
rect 10148 2210 10166 2274
rect 10230 2210 10248 2274
rect 10312 2210 10330 2274
rect 10394 2210 10412 2274
rect 10476 2210 10494 2274
rect 10558 2210 10576 2274
rect 10640 2210 10657 2274
rect 10721 2210 10738 2274
rect 10802 2210 10819 2274
rect 10883 2210 10900 2274
rect 10964 2210 10981 2274
rect 11045 2210 11062 2274
rect 11126 2210 11143 2274
rect 11207 2210 11224 2274
rect 11288 2210 11305 2274
rect 11369 2210 11386 2274
rect 11450 2210 11467 2274
rect 11531 2210 11548 2274
rect 11612 2210 11629 2274
rect 11693 2210 11710 2274
rect 11774 2210 11791 2274
rect 11855 2210 11872 2274
rect 11936 2210 11953 2274
rect 12017 2210 12034 2274
rect 12098 2210 12115 2274
rect 12179 2210 12196 2274
rect 12260 2210 12277 2274
rect 12341 2210 12358 2274
rect 12422 2210 12439 2274
rect 12503 2210 12520 2274
rect 12584 2210 12601 2274
rect 12665 2210 12682 2274
rect 12746 2210 12763 2274
rect 12827 2210 12844 2274
rect 12908 2210 12925 2274
rect 12989 2210 13006 2274
rect 13070 2210 13087 2274
rect 13151 2210 13168 2274
rect 13232 2210 13249 2274
rect 13313 2210 13330 2274
rect 13394 2210 13411 2274
rect 13475 2210 13492 2274
rect 13556 2210 13573 2274
rect 13637 2210 13654 2274
rect 13718 2210 13735 2274
rect 13799 2210 13816 2274
rect 13880 2210 13897 2274
rect 13961 2210 13978 2274
rect 14042 2210 14059 2274
rect 14123 2210 14140 2274
rect 14204 2210 14221 2274
rect 14285 2210 14302 2274
rect 14366 2210 14383 2274
rect 14447 2210 14464 2274
rect 14528 2210 14545 2274
rect 14609 2210 14626 2274
rect 14690 2210 14707 2274
rect 14771 2210 14788 2274
rect 14852 2210 15000 2274
rect 0 2188 15000 2210
rect 0 2124 105 2188
rect 169 2124 187 2188
rect 251 2124 269 2188
rect 333 2124 351 2188
rect 415 2124 433 2188
rect 497 2124 515 2188
rect 579 2124 597 2188
rect 661 2124 678 2188
rect 742 2124 759 2188
rect 823 2124 840 2188
rect 904 2124 921 2188
rect 985 2124 1002 2188
rect 1066 2124 1083 2188
rect 1147 2124 1164 2188
rect 1228 2124 1245 2188
rect 1309 2124 1326 2188
rect 1390 2124 1407 2188
rect 1471 2124 1488 2188
rect 1552 2124 1569 2188
rect 1633 2124 1650 2188
rect 1714 2124 1731 2188
rect 1795 2124 1812 2188
rect 1876 2124 1893 2188
rect 1957 2124 1974 2188
rect 2038 2124 2055 2188
rect 2119 2124 2136 2188
rect 2200 2124 2217 2188
rect 2281 2124 2298 2188
rect 2362 2124 2379 2188
rect 2443 2124 2460 2188
rect 2524 2124 2541 2188
rect 2605 2124 2622 2188
rect 2686 2124 2703 2188
rect 2767 2124 2784 2188
rect 2848 2124 2865 2188
rect 2929 2124 2946 2188
rect 3010 2124 3027 2188
rect 3091 2124 3108 2188
rect 3172 2124 3189 2188
rect 3253 2124 3270 2188
rect 3334 2124 3351 2188
rect 3415 2124 3432 2188
rect 3496 2124 3513 2188
rect 3577 2124 3594 2188
rect 3658 2124 3675 2188
rect 3739 2124 3756 2188
rect 3820 2124 3837 2188
rect 3901 2124 3918 2188
rect 3982 2124 3999 2188
rect 4063 2124 4080 2188
rect 4144 2124 4161 2188
rect 4225 2124 4242 2188
rect 4306 2124 4323 2188
rect 4387 2124 4404 2188
rect 4468 2124 4485 2188
rect 4549 2124 4566 2188
rect 4630 2124 4647 2188
rect 4711 2124 4728 2188
rect 4792 2124 4809 2188
rect 4873 2124 10084 2188
rect 10148 2124 10166 2188
rect 10230 2124 10248 2188
rect 10312 2124 10330 2188
rect 10394 2124 10412 2188
rect 10476 2124 10494 2188
rect 10558 2124 10576 2188
rect 10640 2124 10657 2188
rect 10721 2124 10738 2188
rect 10802 2124 10819 2188
rect 10883 2124 10900 2188
rect 10964 2124 10981 2188
rect 11045 2124 11062 2188
rect 11126 2124 11143 2188
rect 11207 2124 11224 2188
rect 11288 2124 11305 2188
rect 11369 2124 11386 2188
rect 11450 2124 11467 2188
rect 11531 2124 11548 2188
rect 11612 2124 11629 2188
rect 11693 2124 11710 2188
rect 11774 2124 11791 2188
rect 11855 2124 11872 2188
rect 11936 2124 11953 2188
rect 12017 2124 12034 2188
rect 12098 2124 12115 2188
rect 12179 2124 12196 2188
rect 12260 2124 12277 2188
rect 12341 2124 12358 2188
rect 12422 2124 12439 2188
rect 12503 2124 12520 2188
rect 12584 2124 12601 2188
rect 12665 2124 12682 2188
rect 12746 2124 12763 2188
rect 12827 2124 12844 2188
rect 12908 2124 12925 2188
rect 12989 2124 13006 2188
rect 13070 2124 13087 2188
rect 13151 2124 13168 2188
rect 13232 2124 13249 2188
rect 13313 2124 13330 2188
rect 13394 2124 13411 2188
rect 13475 2124 13492 2188
rect 13556 2124 13573 2188
rect 13637 2124 13654 2188
rect 13718 2124 13735 2188
rect 13799 2124 13816 2188
rect 13880 2124 13897 2188
rect 13961 2124 13978 2188
rect 14042 2124 14059 2188
rect 14123 2124 14140 2188
rect 14204 2124 14221 2188
rect 14285 2124 14302 2188
rect 14366 2124 14383 2188
rect 14447 2124 14464 2188
rect 14528 2124 14545 2188
rect 14609 2124 14626 2188
rect 14690 2124 14707 2188
rect 14771 2124 14788 2188
rect 14852 2124 15000 2188
rect 0 2102 15000 2124
rect 0 2038 105 2102
rect 169 2038 187 2102
rect 251 2038 269 2102
rect 333 2038 351 2102
rect 415 2038 433 2102
rect 497 2038 515 2102
rect 579 2038 597 2102
rect 661 2038 678 2102
rect 742 2038 759 2102
rect 823 2038 840 2102
rect 904 2038 921 2102
rect 985 2038 1002 2102
rect 1066 2038 1083 2102
rect 1147 2038 1164 2102
rect 1228 2038 1245 2102
rect 1309 2038 1326 2102
rect 1390 2038 1407 2102
rect 1471 2038 1488 2102
rect 1552 2038 1569 2102
rect 1633 2038 1650 2102
rect 1714 2038 1731 2102
rect 1795 2038 1812 2102
rect 1876 2038 1893 2102
rect 1957 2038 1974 2102
rect 2038 2038 2055 2102
rect 2119 2038 2136 2102
rect 2200 2038 2217 2102
rect 2281 2038 2298 2102
rect 2362 2038 2379 2102
rect 2443 2038 2460 2102
rect 2524 2038 2541 2102
rect 2605 2038 2622 2102
rect 2686 2038 2703 2102
rect 2767 2038 2784 2102
rect 2848 2038 2865 2102
rect 2929 2038 2946 2102
rect 3010 2038 3027 2102
rect 3091 2038 3108 2102
rect 3172 2038 3189 2102
rect 3253 2038 3270 2102
rect 3334 2038 3351 2102
rect 3415 2038 3432 2102
rect 3496 2038 3513 2102
rect 3577 2038 3594 2102
rect 3658 2038 3675 2102
rect 3739 2038 3756 2102
rect 3820 2038 3837 2102
rect 3901 2038 3918 2102
rect 3982 2038 3999 2102
rect 4063 2038 4080 2102
rect 4144 2038 4161 2102
rect 4225 2038 4242 2102
rect 4306 2038 4323 2102
rect 4387 2038 4404 2102
rect 4468 2038 4485 2102
rect 4549 2038 4566 2102
rect 4630 2038 4647 2102
rect 4711 2038 4728 2102
rect 4792 2038 4809 2102
rect 4873 2038 10084 2102
rect 10148 2038 10166 2102
rect 10230 2038 10248 2102
rect 10312 2038 10330 2102
rect 10394 2038 10412 2102
rect 10476 2038 10494 2102
rect 10558 2038 10576 2102
rect 10640 2038 10657 2102
rect 10721 2038 10738 2102
rect 10802 2038 10819 2102
rect 10883 2038 10900 2102
rect 10964 2038 10981 2102
rect 11045 2038 11062 2102
rect 11126 2038 11143 2102
rect 11207 2038 11224 2102
rect 11288 2038 11305 2102
rect 11369 2038 11386 2102
rect 11450 2038 11467 2102
rect 11531 2038 11548 2102
rect 11612 2038 11629 2102
rect 11693 2038 11710 2102
rect 11774 2038 11791 2102
rect 11855 2038 11872 2102
rect 11936 2038 11953 2102
rect 12017 2038 12034 2102
rect 12098 2038 12115 2102
rect 12179 2038 12196 2102
rect 12260 2038 12277 2102
rect 12341 2038 12358 2102
rect 12422 2038 12439 2102
rect 12503 2038 12520 2102
rect 12584 2038 12601 2102
rect 12665 2038 12682 2102
rect 12746 2038 12763 2102
rect 12827 2038 12844 2102
rect 12908 2038 12925 2102
rect 12989 2038 13006 2102
rect 13070 2038 13087 2102
rect 13151 2038 13168 2102
rect 13232 2038 13249 2102
rect 13313 2038 13330 2102
rect 13394 2038 13411 2102
rect 13475 2038 13492 2102
rect 13556 2038 13573 2102
rect 13637 2038 13654 2102
rect 13718 2038 13735 2102
rect 13799 2038 13816 2102
rect 13880 2038 13897 2102
rect 13961 2038 13978 2102
rect 14042 2038 14059 2102
rect 14123 2038 14140 2102
rect 14204 2038 14221 2102
rect 14285 2038 14302 2102
rect 14366 2038 14383 2102
rect 14447 2038 14464 2102
rect 14528 2038 14545 2102
rect 14609 2038 14626 2102
rect 14690 2038 14707 2102
rect 14771 2038 14788 2102
rect 14852 2038 15000 2102
rect 0 2016 15000 2038
rect 0 1952 105 2016
rect 169 1952 187 2016
rect 251 1952 269 2016
rect 333 1952 351 2016
rect 415 1952 433 2016
rect 497 1952 515 2016
rect 579 1952 597 2016
rect 661 1952 678 2016
rect 742 1952 759 2016
rect 823 1952 840 2016
rect 904 1952 921 2016
rect 985 1952 1002 2016
rect 1066 1952 1083 2016
rect 1147 1952 1164 2016
rect 1228 1952 1245 2016
rect 1309 1952 1326 2016
rect 1390 1952 1407 2016
rect 1471 1952 1488 2016
rect 1552 1952 1569 2016
rect 1633 1952 1650 2016
rect 1714 1952 1731 2016
rect 1795 1952 1812 2016
rect 1876 1952 1893 2016
rect 1957 1952 1974 2016
rect 2038 1952 2055 2016
rect 2119 1952 2136 2016
rect 2200 1952 2217 2016
rect 2281 1952 2298 2016
rect 2362 1952 2379 2016
rect 2443 1952 2460 2016
rect 2524 1952 2541 2016
rect 2605 1952 2622 2016
rect 2686 1952 2703 2016
rect 2767 1952 2784 2016
rect 2848 1952 2865 2016
rect 2929 1952 2946 2016
rect 3010 1952 3027 2016
rect 3091 1952 3108 2016
rect 3172 1952 3189 2016
rect 3253 1952 3270 2016
rect 3334 1952 3351 2016
rect 3415 1952 3432 2016
rect 3496 1952 3513 2016
rect 3577 1952 3594 2016
rect 3658 1952 3675 2016
rect 3739 1952 3756 2016
rect 3820 1952 3837 2016
rect 3901 1952 3918 2016
rect 3982 1952 3999 2016
rect 4063 1952 4080 2016
rect 4144 1952 4161 2016
rect 4225 1952 4242 2016
rect 4306 1952 4323 2016
rect 4387 1952 4404 2016
rect 4468 1952 4485 2016
rect 4549 1952 4566 2016
rect 4630 1952 4647 2016
rect 4711 1952 4728 2016
rect 4792 1952 4809 2016
rect 4873 1952 10084 2016
rect 10148 1952 10166 2016
rect 10230 1952 10248 2016
rect 10312 1952 10330 2016
rect 10394 1952 10412 2016
rect 10476 1952 10494 2016
rect 10558 1952 10576 2016
rect 10640 1952 10657 2016
rect 10721 1952 10738 2016
rect 10802 1952 10819 2016
rect 10883 1952 10900 2016
rect 10964 1952 10981 2016
rect 11045 1952 11062 2016
rect 11126 1952 11143 2016
rect 11207 1952 11224 2016
rect 11288 1952 11305 2016
rect 11369 1952 11386 2016
rect 11450 1952 11467 2016
rect 11531 1952 11548 2016
rect 11612 1952 11629 2016
rect 11693 1952 11710 2016
rect 11774 1952 11791 2016
rect 11855 1952 11872 2016
rect 11936 1952 11953 2016
rect 12017 1952 12034 2016
rect 12098 1952 12115 2016
rect 12179 1952 12196 2016
rect 12260 1952 12277 2016
rect 12341 1952 12358 2016
rect 12422 1952 12439 2016
rect 12503 1952 12520 2016
rect 12584 1952 12601 2016
rect 12665 1952 12682 2016
rect 12746 1952 12763 2016
rect 12827 1952 12844 2016
rect 12908 1952 12925 2016
rect 12989 1952 13006 2016
rect 13070 1952 13087 2016
rect 13151 1952 13168 2016
rect 13232 1952 13249 2016
rect 13313 1952 13330 2016
rect 13394 1952 13411 2016
rect 13475 1952 13492 2016
rect 13556 1952 13573 2016
rect 13637 1952 13654 2016
rect 13718 1952 13735 2016
rect 13799 1952 13816 2016
rect 13880 1952 13897 2016
rect 13961 1952 13978 2016
rect 14042 1952 14059 2016
rect 14123 1952 14140 2016
rect 14204 1952 14221 2016
rect 14285 1952 14302 2016
rect 14366 1952 14383 2016
rect 14447 1952 14464 2016
rect 14528 1952 14545 2016
rect 14609 1952 14626 2016
rect 14690 1952 14707 2016
rect 14771 1952 14788 2016
rect 14852 1952 15000 2016
rect 0 1930 15000 1952
rect 0 1866 105 1930
rect 169 1866 187 1930
rect 251 1866 269 1930
rect 333 1866 351 1930
rect 415 1866 433 1930
rect 497 1866 515 1930
rect 579 1866 597 1930
rect 661 1866 678 1930
rect 742 1866 759 1930
rect 823 1866 840 1930
rect 904 1866 921 1930
rect 985 1866 1002 1930
rect 1066 1866 1083 1930
rect 1147 1866 1164 1930
rect 1228 1866 1245 1930
rect 1309 1866 1326 1930
rect 1390 1866 1407 1930
rect 1471 1866 1488 1930
rect 1552 1866 1569 1930
rect 1633 1866 1650 1930
rect 1714 1866 1731 1930
rect 1795 1866 1812 1930
rect 1876 1866 1893 1930
rect 1957 1866 1974 1930
rect 2038 1866 2055 1930
rect 2119 1866 2136 1930
rect 2200 1866 2217 1930
rect 2281 1866 2298 1930
rect 2362 1866 2379 1930
rect 2443 1866 2460 1930
rect 2524 1866 2541 1930
rect 2605 1866 2622 1930
rect 2686 1866 2703 1930
rect 2767 1866 2784 1930
rect 2848 1866 2865 1930
rect 2929 1866 2946 1930
rect 3010 1866 3027 1930
rect 3091 1866 3108 1930
rect 3172 1866 3189 1930
rect 3253 1866 3270 1930
rect 3334 1866 3351 1930
rect 3415 1866 3432 1930
rect 3496 1866 3513 1930
rect 3577 1866 3594 1930
rect 3658 1866 3675 1930
rect 3739 1866 3756 1930
rect 3820 1866 3837 1930
rect 3901 1866 3918 1930
rect 3982 1866 3999 1930
rect 4063 1866 4080 1930
rect 4144 1866 4161 1930
rect 4225 1866 4242 1930
rect 4306 1866 4323 1930
rect 4387 1866 4404 1930
rect 4468 1866 4485 1930
rect 4549 1866 4566 1930
rect 4630 1866 4647 1930
rect 4711 1866 4728 1930
rect 4792 1866 4809 1930
rect 4873 1866 10084 1930
rect 10148 1866 10166 1930
rect 10230 1866 10248 1930
rect 10312 1866 10330 1930
rect 10394 1866 10412 1930
rect 10476 1866 10494 1930
rect 10558 1866 10576 1930
rect 10640 1866 10657 1930
rect 10721 1866 10738 1930
rect 10802 1866 10819 1930
rect 10883 1866 10900 1930
rect 10964 1866 10981 1930
rect 11045 1866 11062 1930
rect 11126 1866 11143 1930
rect 11207 1866 11224 1930
rect 11288 1866 11305 1930
rect 11369 1866 11386 1930
rect 11450 1866 11467 1930
rect 11531 1866 11548 1930
rect 11612 1866 11629 1930
rect 11693 1866 11710 1930
rect 11774 1866 11791 1930
rect 11855 1866 11872 1930
rect 11936 1866 11953 1930
rect 12017 1866 12034 1930
rect 12098 1866 12115 1930
rect 12179 1866 12196 1930
rect 12260 1866 12277 1930
rect 12341 1866 12358 1930
rect 12422 1866 12439 1930
rect 12503 1866 12520 1930
rect 12584 1866 12601 1930
rect 12665 1866 12682 1930
rect 12746 1866 12763 1930
rect 12827 1866 12844 1930
rect 12908 1866 12925 1930
rect 12989 1866 13006 1930
rect 13070 1866 13087 1930
rect 13151 1866 13168 1930
rect 13232 1866 13249 1930
rect 13313 1866 13330 1930
rect 13394 1866 13411 1930
rect 13475 1866 13492 1930
rect 13556 1866 13573 1930
rect 13637 1866 13654 1930
rect 13718 1866 13735 1930
rect 13799 1866 13816 1930
rect 13880 1866 13897 1930
rect 13961 1866 13978 1930
rect 14042 1866 14059 1930
rect 14123 1866 14140 1930
rect 14204 1866 14221 1930
rect 14285 1866 14302 1930
rect 14366 1866 14383 1930
rect 14447 1866 14464 1930
rect 14528 1866 14545 1930
rect 14609 1866 14626 1930
rect 14690 1866 14707 1930
rect 14771 1866 14788 1930
rect 14852 1866 15000 1930
rect 0 1844 15000 1866
rect 0 1780 105 1844
rect 169 1780 187 1844
rect 251 1780 269 1844
rect 333 1780 351 1844
rect 415 1780 433 1844
rect 497 1780 515 1844
rect 579 1780 597 1844
rect 661 1780 678 1844
rect 742 1780 759 1844
rect 823 1780 840 1844
rect 904 1780 921 1844
rect 985 1780 1002 1844
rect 1066 1780 1083 1844
rect 1147 1780 1164 1844
rect 1228 1780 1245 1844
rect 1309 1780 1326 1844
rect 1390 1780 1407 1844
rect 1471 1780 1488 1844
rect 1552 1780 1569 1844
rect 1633 1780 1650 1844
rect 1714 1780 1731 1844
rect 1795 1780 1812 1844
rect 1876 1780 1893 1844
rect 1957 1780 1974 1844
rect 2038 1780 2055 1844
rect 2119 1780 2136 1844
rect 2200 1780 2217 1844
rect 2281 1780 2298 1844
rect 2362 1780 2379 1844
rect 2443 1780 2460 1844
rect 2524 1780 2541 1844
rect 2605 1780 2622 1844
rect 2686 1780 2703 1844
rect 2767 1780 2784 1844
rect 2848 1780 2865 1844
rect 2929 1780 2946 1844
rect 3010 1780 3027 1844
rect 3091 1780 3108 1844
rect 3172 1780 3189 1844
rect 3253 1780 3270 1844
rect 3334 1780 3351 1844
rect 3415 1780 3432 1844
rect 3496 1780 3513 1844
rect 3577 1780 3594 1844
rect 3658 1780 3675 1844
rect 3739 1780 3756 1844
rect 3820 1780 3837 1844
rect 3901 1780 3918 1844
rect 3982 1780 3999 1844
rect 4063 1780 4080 1844
rect 4144 1780 4161 1844
rect 4225 1780 4242 1844
rect 4306 1780 4323 1844
rect 4387 1780 4404 1844
rect 4468 1780 4485 1844
rect 4549 1780 4566 1844
rect 4630 1780 4647 1844
rect 4711 1780 4728 1844
rect 4792 1780 4809 1844
rect 4873 1780 10084 1844
rect 10148 1780 10166 1844
rect 10230 1780 10248 1844
rect 10312 1780 10330 1844
rect 10394 1780 10412 1844
rect 10476 1780 10494 1844
rect 10558 1780 10576 1844
rect 10640 1780 10657 1844
rect 10721 1780 10738 1844
rect 10802 1780 10819 1844
rect 10883 1780 10900 1844
rect 10964 1780 10981 1844
rect 11045 1780 11062 1844
rect 11126 1780 11143 1844
rect 11207 1780 11224 1844
rect 11288 1780 11305 1844
rect 11369 1780 11386 1844
rect 11450 1780 11467 1844
rect 11531 1780 11548 1844
rect 11612 1780 11629 1844
rect 11693 1780 11710 1844
rect 11774 1780 11791 1844
rect 11855 1780 11872 1844
rect 11936 1780 11953 1844
rect 12017 1780 12034 1844
rect 12098 1780 12115 1844
rect 12179 1780 12196 1844
rect 12260 1780 12277 1844
rect 12341 1780 12358 1844
rect 12422 1780 12439 1844
rect 12503 1780 12520 1844
rect 12584 1780 12601 1844
rect 12665 1780 12682 1844
rect 12746 1780 12763 1844
rect 12827 1780 12844 1844
rect 12908 1780 12925 1844
rect 12989 1780 13006 1844
rect 13070 1780 13087 1844
rect 13151 1780 13168 1844
rect 13232 1780 13249 1844
rect 13313 1780 13330 1844
rect 13394 1780 13411 1844
rect 13475 1780 13492 1844
rect 13556 1780 13573 1844
rect 13637 1780 13654 1844
rect 13718 1780 13735 1844
rect 13799 1780 13816 1844
rect 13880 1780 13897 1844
rect 13961 1780 13978 1844
rect 14042 1780 14059 1844
rect 14123 1780 14140 1844
rect 14204 1780 14221 1844
rect 14285 1780 14302 1844
rect 14366 1780 14383 1844
rect 14447 1780 14464 1844
rect 14528 1780 14545 1844
rect 14609 1780 14626 1844
rect 14690 1780 14707 1844
rect 14771 1780 14788 1844
rect 14852 1780 15000 1844
rect 0 407 15000 1780
<< metal5 >>
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14807 3007 15000 3657
rect 14746 427 15000 1477
<< obsm5 >>
rect 0 19317 15000 40000
rect 0 8017 14426 19317
rect 0 7367 15000 8017
rect 0 4867 14426 7367
rect 0 3977 15000 4867
rect 0 2687 14487 3977
rect 0 1797 15000 2687
rect 0 427 14426 1797
<< labels >>
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal4 s 105 2038 169 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 2038 169 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 2124 169 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 2124 169 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 2210 169 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 2210 169 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 2296 169 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 2296 169 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 2382 169 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 2382 169 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 2468 169 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 2468 169 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 2554 169 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 2554 169 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 2640 169 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 2640 169 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 1780 169 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 1780 169 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 1866 169 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 1866 169 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 105 1952 169 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 105 1952 169 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 2038 251 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 2038 251 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 2124 251 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 2124 251 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 2210 251 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 2210 251 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 2296 251 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 2296 251 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 2382 251 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 2382 251 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 2468 251 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 2468 251 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 2554 251 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 2554 251 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 2640 251 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 2640 251 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 1780 251 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 1780 251 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 1866 251 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 1866 251 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 187 1952 251 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 187 1952 251 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 2038 333 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 2038 333 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 2124 333 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 2124 333 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 2210 333 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 2210 333 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 2296 333 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 2296 333 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 2382 333 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 2382 333 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 2468 333 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 2468 333 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 2554 333 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 2554 333 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 2640 333 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 2640 333 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 1780 333 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 1780 333 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 1866 333 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 1866 333 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 269 1952 333 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 269 1952 333 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 2038 415 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 2038 415 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 2124 415 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 2124 415 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 2210 415 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 2210 415 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 2296 415 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 2296 415 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 2382 415 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 2382 415 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 2468 415 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 2468 415 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 2554 415 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 2554 415 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 2640 415 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 2640 415 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 1780 415 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 1780 415 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 1866 415 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 1866 415 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 351 1952 415 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 351 1952 415 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 2038 2119 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 2038 2119 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 2124 2119 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 2124 2119 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 2210 2119 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 2210 2119 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 2296 2119 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 2296 2119 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 2382 2119 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 2382 2119 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 2468 2119 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 2468 2119 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 2554 2119 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 2554 2119 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 2640 2119 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 2640 2119 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 1780 2119 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 1780 2119 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 1866 2119 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 1866 2119 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2055 1952 2119 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2055 1952 2119 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 2038 2200 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 2038 2200 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 2124 2200 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 2124 2200 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 2210 2200 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 2210 2200 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 2296 2200 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 2296 2200 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 2382 2200 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 2382 2200 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 2468 2200 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 2468 2200 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 2554 2200 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 2554 2200 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 2640 2200 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 2640 2200 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 1780 2200 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 1780 2200 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 1866 2200 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 1866 2200 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2136 1952 2200 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2136 1952 2200 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 2038 2281 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 2038 2281 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 2124 2281 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 2124 2281 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 2210 2281 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 2210 2281 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 2296 2281 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 2296 2281 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 2382 2281 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 2382 2281 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 2468 2281 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 2468 2281 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 2554 2281 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 2554 2281 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 2640 2281 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 2640 2281 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 1780 2281 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 1780 2281 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 1866 2281 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 1866 2281 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2217 1952 2281 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2217 1952 2281 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 2038 2362 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 2038 2362 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 2124 2362 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 2124 2362 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 2210 2362 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 2210 2362 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 2296 2362 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 2296 2362 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 2382 2362 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 2382 2362 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 2468 2362 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 2468 2362 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 2554 2362 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 2554 2362 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 2640 2362 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 2640 2362 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 1780 2362 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 1780 2362 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 1866 2362 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 1866 2362 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2298 1952 2362 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2298 1952 2362 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 2038 2443 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 2038 2443 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 2124 2443 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 2124 2443 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 2210 2443 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 2210 2443 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 2296 2443 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 2296 2443 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 2382 2443 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 2382 2443 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 2468 2443 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 2468 2443 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 2554 2443 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 2554 2443 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 2640 2443 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 2640 2443 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 1780 2443 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 1780 2443 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 1866 2443 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 1866 2443 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2379 1952 2443 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2379 1952 2443 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 2038 2524 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 2038 2524 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 2124 2524 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 2124 2524 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 2210 2524 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 2210 2524 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 2296 2524 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 2296 2524 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 2382 2524 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 2382 2524 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 2468 2524 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 2468 2524 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 2554 2524 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 2554 2524 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 2640 2524 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 2640 2524 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 1780 2524 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 1780 2524 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 1866 2524 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 1866 2524 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2460 1952 2524 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2460 1952 2524 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 2038 2605 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 2038 2605 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 2124 2605 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 2124 2605 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 2210 2605 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 2210 2605 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 2296 2605 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 2296 2605 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 2382 2605 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 2382 2605 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 2468 2605 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 2468 2605 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 2554 2605 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 2554 2605 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 2640 2605 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 2640 2605 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 1780 2605 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 1780 2605 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 1866 2605 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 1866 2605 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2541 1952 2605 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2541 1952 2605 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 2038 2686 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 2038 2686 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 2124 2686 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 2124 2686 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 2210 2686 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 2210 2686 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 2296 2686 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 2296 2686 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 2382 2686 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 2382 2686 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 2468 2686 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 2468 2686 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 2554 2686 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 2554 2686 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 2640 2686 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 2640 2686 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 1780 2686 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 1780 2686 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 1866 2686 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 1866 2686 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2622 1952 2686 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2622 1952 2686 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 2038 2767 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 2038 2767 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 2124 2767 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 2124 2767 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 2210 2767 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 2210 2767 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 2296 2767 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 2296 2767 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 2382 2767 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 2382 2767 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 2468 2767 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 2468 2767 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 2554 2767 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 2554 2767 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 2640 2767 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 2640 2767 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 1780 2767 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 1780 2767 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 1866 2767 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 1866 2767 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2703 1952 2767 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2703 1952 2767 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 2038 2848 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 2038 2848 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 2124 2848 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 2124 2848 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 2210 2848 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 2210 2848 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 2296 2848 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 2296 2848 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 2382 2848 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 2382 2848 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 2468 2848 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 2468 2848 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 2554 2848 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 2554 2848 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 2640 2848 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 2640 2848 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 1780 2848 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 1780 2848 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 1866 2848 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 1866 2848 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2784 1952 2848 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2784 1952 2848 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 2038 2929 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 2038 2929 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 2124 2929 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 2124 2929 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 2210 2929 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 2210 2929 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 2296 2929 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 2296 2929 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 2382 2929 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 2382 2929 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 2468 2929 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 2468 2929 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 2554 2929 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 2554 2929 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 2640 2929 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 2640 2929 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 1780 2929 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 1780 2929 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 1866 2929 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 1866 2929 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2865 1952 2929 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2865 1952 2929 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 2038 3010 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 2038 3010 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 2124 3010 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 2124 3010 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 2210 3010 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 2210 3010 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 2296 3010 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 2296 3010 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 2382 3010 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 2382 3010 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 2468 3010 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 2468 3010 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 2554 3010 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 2554 3010 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 2640 3010 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 2640 3010 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 1780 3010 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 1780 3010 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 1866 3010 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 1866 3010 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 2946 1952 3010 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 2946 1952 3010 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 2038 3091 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 2038 3091 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 2124 3091 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 2124 3091 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 2210 3091 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 2210 3091 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 2296 3091 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 2296 3091 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 2382 3091 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 2382 3091 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 2468 3091 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 2468 3091 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 2554 3091 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 2554 3091 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 2640 3091 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 2640 3091 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 1780 3091 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 1780 3091 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 1866 3091 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 1866 3091 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3027 1952 3091 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3027 1952 3091 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 2038 3172 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 2038 3172 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 2124 3172 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 2124 3172 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 2210 3172 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 2210 3172 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 2296 3172 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 2296 3172 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 2382 3172 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 2382 3172 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 2468 3172 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 2468 3172 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 2554 3172 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 2554 3172 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 2640 3172 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 2640 3172 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 1780 3172 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 1780 3172 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 1866 3172 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 1866 3172 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3108 1952 3172 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3108 1952 3172 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 2038 3253 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 2038 3253 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 2124 3253 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 2124 3253 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 2210 3253 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 2210 3253 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 2296 3253 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 2296 3253 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 2382 3253 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 2382 3253 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 2468 3253 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 2468 3253 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 2554 3253 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 2554 3253 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 2640 3253 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 2640 3253 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 1780 3253 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 1780 3253 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 1866 3253 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 1866 3253 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3189 1952 3253 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3189 1952 3253 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 2038 3334 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 2038 3334 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 2124 3334 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 2124 3334 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 2210 3334 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 2210 3334 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 2296 3334 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 2296 3334 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 2382 3334 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 2382 3334 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 2468 3334 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 2468 3334 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 2554 3334 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 2554 3334 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 2640 3334 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 2640 3334 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 1780 3334 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 1780 3334 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 1866 3334 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 1866 3334 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3270 1952 3334 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3270 1952 3334 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 2038 3415 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 2038 3415 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 2124 3415 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 2124 3415 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 2210 3415 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 2210 3415 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 2296 3415 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 2296 3415 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 2382 3415 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 2382 3415 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 2468 3415 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 2468 3415 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 2554 3415 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 2554 3415 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 2640 3415 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 2640 3415 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 1780 3415 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 1780 3415 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 1866 3415 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 1866 3415 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3351 1952 3415 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3351 1952 3415 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 2038 3496 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 2038 3496 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 2124 3496 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 2124 3496 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 2210 3496 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 2210 3496 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 2296 3496 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 2296 3496 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 2382 3496 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 2382 3496 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 2468 3496 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 2468 3496 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 2554 3496 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 2554 3496 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 2640 3496 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 2640 3496 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 1780 3496 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 1780 3496 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 1866 3496 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 1866 3496 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3432 1952 3496 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3432 1952 3496 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 2038 3577 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 2038 3577 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 2124 3577 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 2124 3577 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 2210 3577 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 2210 3577 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 2296 3577 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 2296 3577 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 2382 3577 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 2382 3577 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 2468 3577 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 2468 3577 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 2554 3577 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 2554 3577 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 2640 3577 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 2640 3577 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 1780 3577 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 1780 3577 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 1866 3577 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 1866 3577 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3513 1952 3577 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3513 1952 3577 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 2038 3658 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 2038 3658 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 2124 3658 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 2124 3658 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 2210 3658 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 2210 3658 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 2296 3658 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 2296 3658 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 2382 3658 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 2382 3658 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 2468 3658 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 2468 3658 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 2554 3658 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 2554 3658 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 2640 3658 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 2640 3658 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 1780 3658 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 1780 3658 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 1866 3658 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 1866 3658 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3594 1952 3658 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3594 1952 3658 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 2038 3739 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 2038 3739 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 2124 3739 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 2124 3739 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 2210 3739 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 2210 3739 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 2296 3739 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 2296 3739 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 2382 3739 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 2382 3739 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 2468 3739 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 2468 3739 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 2554 3739 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 2554 3739 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 2640 3739 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 2640 3739 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 1780 3739 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 1780 3739 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 1866 3739 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 1866 3739 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3675 1952 3739 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3675 1952 3739 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 2038 3820 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 2038 3820 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 2124 3820 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 2124 3820 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 2210 3820 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 2210 3820 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 2296 3820 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 2296 3820 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 2382 3820 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 2382 3820 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 2468 3820 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 2468 3820 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 2554 3820 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 2554 3820 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 2640 3820 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 2640 3820 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 1780 3820 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 1780 3820 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 1866 3820 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 1866 3820 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3756 1952 3820 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3756 1952 3820 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 2038 3901 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 2038 3901 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 2124 3901 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 2124 3901 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 2210 3901 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 2210 3901 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 2296 3901 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 2296 3901 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 2382 3901 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 2382 3901 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 2468 3901 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 2468 3901 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 2554 3901 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 2554 3901 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 2640 3901 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 2640 3901 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 1780 3901 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 1780 3901 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 1866 3901 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 1866 3901 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3837 1952 3901 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3837 1952 3901 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 2038 3982 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 2038 3982 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 2124 3982 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 2124 3982 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 2210 3982 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 2210 3982 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 2296 3982 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 2296 3982 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 2382 3982 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 2382 3982 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 2468 3982 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 2468 3982 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 2554 3982 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 2554 3982 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 2640 3982 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 2640 3982 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 1780 3982 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 1780 3982 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 1866 3982 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 1866 3982 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3918 1952 3982 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3918 1952 3982 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 2038 4063 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 2038 4063 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 2124 4063 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 2124 4063 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 2210 4063 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 2210 4063 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 2296 4063 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 2296 4063 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 2382 4063 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 2382 4063 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 2468 4063 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 2468 4063 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 2554 4063 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 2554 4063 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 2640 4063 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 2640 4063 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 1780 4063 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 1780 4063 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 1866 4063 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 1866 4063 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 3999 1952 4063 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 3999 1952 4063 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 2038 497 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 2038 497 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 2124 497 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 2124 497 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 2210 497 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 2210 497 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 2296 497 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 2296 497 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 2382 497 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 2382 497 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 2468 497 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 2468 497 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 2554 497 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 2554 497 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 2640 497 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 2640 497 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 1780 497 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 1780 497 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 1866 497 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 1866 497 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 433 1952 497 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 433 1952 497 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 2038 579 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 2038 579 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 2124 579 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 2124 579 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 2210 579 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 2210 579 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 2296 579 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 2296 579 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 2382 579 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 2382 579 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 2468 579 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 2468 579 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 2554 579 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 2554 579 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 2640 579 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 2640 579 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 1780 579 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 1780 579 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 1866 579 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 1866 579 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 515 1952 579 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 515 1952 579 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 2038 661 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 2038 661 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 2124 661 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 2124 661 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 2210 661 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 2210 661 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 2296 661 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 2296 661 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 2382 661 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 2382 661 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 2468 661 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 2468 661 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 2554 661 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 2554 661 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 2640 661 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 2640 661 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 1780 661 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 1780 661 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 1866 661 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 1866 661 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 597 1952 661 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 597 1952 661 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 2038 4144 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 2038 4144 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 2124 4144 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 2124 4144 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 2210 4144 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 2210 4144 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 2296 4144 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 2296 4144 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 2382 4144 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 2382 4144 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 2468 4144 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 2468 4144 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 2554 4144 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 2554 4144 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 2640 4144 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 2640 4144 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 1780 4144 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 1780 4144 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 1866 4144 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 1866 4144 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4080 1952 4144 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4080 1952 4144 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 2038 4225 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 2038 4225 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 2124 4225 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 2124 4225 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 2210 4225 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 2210 4225 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 2296 4225 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 2296 4225 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 2382 4225 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 2382 4225 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 2468 4225 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 2468 4225 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 2554 4225 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 2554 4225 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 2640 4225 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 2640 4225 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 1780 4225 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 1780 4225 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 1866 4225 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 1866 4225 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4161 1952 4225 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4161 1952 4225 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 2038 4306 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 2038 4306 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 2124 4306 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 2124 4306 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 2210 4306 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 2210 4306 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 2296 4306 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 2296 4306 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 2382 4306 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 2382 4306 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 2468 4306 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 2468 4306 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 2554 4306 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 2554 4306 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 2640 4306 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 2640 4306 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 1780 4306 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 1780 4306 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 1866 4306 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 1866 4306 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4242 1952 4306 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4242 1952 4306 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 2038 4387 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 2038 4387 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 2124 4387 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 2124 4387 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 2210 4387 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 2210 4387 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 2296 4387 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 2296 4387 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 2382 4387 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 2382 4387 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 2468 4387 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 2468 4387 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 2554 4387 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 2554 4387 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 2640 4387 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 2640 4387 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 1780 4387 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 1780 4387 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 1866 4387 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 1866 4387 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4323 1952 4387 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4323 1952 4387 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 2038 4468 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 2038 4468 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 2124 4468 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 2124 4468 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 2210 4468 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 2210 4468 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 2296 4468 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 2296 4468 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 2382 4468 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 2382 4468 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 2468 4468 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 2468 4468 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 2554 4468 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 2554 4468 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 2640 4468 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 2640 4468 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 1780 4468 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 1780 4468 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 1866 4468 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 1866 4468 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4404 1952 4468 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4404 1952 4468 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 2038 4549 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 2038 4549 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 2124 4549 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 2124 4549 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 2210 4549 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 2210 4549 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 2296 4549 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 2296 4549 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 2382 4549 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 2382 4549 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 2468 4549 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 2468 4549 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 2554 4549 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 2554 4549 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 2640 4549 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 2640 4549 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 1780 4549 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 1780 4549 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 1866 4549 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 1866 4549 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4485 1952 4549 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4485 1952 4549 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 2038 4630 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 2038 4630 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 2124 4630 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 2124 4630 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 2210 4630 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 2210 4630 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 2296 4630 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 2296 4630 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 2382 4630 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 2382 4630 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 2468 4630 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 2468 4630 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 2554 4630 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 2554 4630 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 2640 4630 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 2640 4630 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 1780 4630 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 1780 4630 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 1866 4630 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 1866 4630 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4566 1952 4630 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4566 1952 4630 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 2038 4711 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 2038 4711 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 2124 4711 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 2124 4711 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 2210 4711 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 2210 4711 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 2296 4711 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 2296 4711 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 2382 4711 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 2382 4711 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 2468 4711 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 2468 4711 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 2554 4711 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 2554 4711 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 2640 4711 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 2640 4711 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 1780 4711 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 1780 4711 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 1866 4711 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 1866 4711 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4647 1952 4711 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4647 1952 4711 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 2038 4792 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 2038 4792 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 2124 4792 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 2124 4792 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 2210 4792 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 2210 4792 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 2296 4792 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 2296 4792 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 2382 4792 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 2382 4792 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 2468 4792 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 2468 4792 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 2554 4792 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 2554 4792 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 2640 4792 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 2640 4792 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 1780 4792 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 1780 4792 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 1866 4792 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 1866 4792 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4728 1952 4792 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4728 1952 4792 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 2038 4873 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 2038 4873 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 2124 4873 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 2124 4873 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 2210 4873 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 2210 4873 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 2296 4873 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 2296 4873 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 2382 4873 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 2382 4873 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 2468 4873 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 2468 4873 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 2554 4873 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 2554 4873 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 2640 4873 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 2640 4873 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 1780 4873 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 1780 4873 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 1866 4873 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 1866 4873 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 4809 1952 4873 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 4809 1952 4873 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 2038 742 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 2038 742 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 2124 742 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 2124 742 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 2210 742 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 2210 742 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 2296 742 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 2296 742 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 2382 742 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 2382 742 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 2468 742 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 2468 742 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 2554 742 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 2554 742 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 2640 742 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 2640 742 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 1780 742 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 1780 742 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 1866 742 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 1866 742 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 678 1952 742 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 678 1952 742 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 2038 823 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 2038 823 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 2124 823 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 2124 823 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 2210 823 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 2210 823 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 2296 823 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 2296 823 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 2382 823 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 2382 823 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 2468 823 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 2468 823 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 2554 823 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 2554 823 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 2640 823 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 2640 823 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 1780 823 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 1780 823 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 1866 823 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 1866 823 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 759 1952 823 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 759 1952 823 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 2038 904 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 2038 904 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 2124 904 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 2124 904 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 2210 904 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 2210 904 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 2296 904 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 2296 904 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 2382 904 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 2382 904 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 2468 904 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 2468 904 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 2554 904 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 2554 904 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 2640 904 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 2640 904 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 1780 904 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 1780 904 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 1866 904 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 1866 904 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 840 1952 904 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 840 1952 904 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 2038 985 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 2038 985 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 2124 985 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 2124 985 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 2210 985 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 2210 985 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 2296 985 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 2296 985 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 2382 985 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 2382 985 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 2468 985 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 2468 985 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 2554 985 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 2554 985 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 2640 985 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 2640 985 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 1780 985 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 1780 985 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 1866 985 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 1866 985 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 921 1952 985 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 921 1952 985 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 2038 1066 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 2038 1066 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 2124 1066 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 2124 1066 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 2210 1066 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 2210 1066 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 2296 1066 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 2296 1066 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 2382 1066 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 2382 1066 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 2468 1066 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 2468 1066 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 2554 1066 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 2554 1066 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 2640 1066 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 2640 1066 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 1780 1066 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 1780 1066 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 1866 1066 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 1866 1066 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1002 1952 1066 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1002 1952 1066 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 2038 1147 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 2038 1147 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 2124 1147 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 2124 1147 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 2210 1147 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 2210 1147 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 2296 1147 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 2296 1147 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 2382 1147 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 2382 1147 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 2468 1147 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 2468 1147 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 2554 1147 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 2554 1147 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 2640 1147 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 2640 1147 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 1780 1147 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 1780 1147 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 1866 1147 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 1866 1147 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1083 1952 1147 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1083 1952 1147 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 2038 1228 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 2038 1228 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 2124 1228 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 2124 1228 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 2210 1228 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 2210 1228 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 2296 1228 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 2296 1228 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 2382 1228 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 2382 1228 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 2468 1228 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 2468 1228 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 2554 1228 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 2554 1228 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 2640 1228 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 2640 1228 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 1780 1228 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 1780 1228 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 1866 1228 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 1866 1228 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1164 1952 1228 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1164 1952 1228 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 2038 10148 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 2038 10148 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 2124 10148 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 2124 10148 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 2210 10148 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 2210 10148 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 2296 10148 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 2296 10148 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 2382 10148 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 2382 10148 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 2468 10148 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 2468 10148 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 2554 10148 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 2554 10148 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 2640 10148 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 2640 10148 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 1780 10148 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 1780 10148 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 1866 10148 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 1866 10148 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10084 1952 10148 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10084 1952 10148 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 2038 10230 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 2038 10230 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 2124 10230 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 2124 10230 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 2210 10230 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 2210 10230 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 2296 10230 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 2296 10230 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 2382 10230 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 2382 10230 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 2468 10230 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 2468 10230 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 2554 10230 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 2554 10230 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 2640 10230 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 2640 10230 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 1780 10230 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 1780 10230 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 1866 10230 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 1866 10230 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10166 1952 10230 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10166 1952 10230 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 2038 10312 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 2038 10312 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 2124 10312 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 2124 10312 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 2210 10312 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 2210 10312 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 2296 10312 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 2296 10312 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 2382 10312 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 2382 10312 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 2468 10312 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 2468 10312 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 2554 10312 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 2554 10312 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 2640 10312 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 2640 10312 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 1780 10312 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 1780 10312 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 1866 10312 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 1866 10312 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10248 1952 10312 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10248 1952 10312 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 2038 10394 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 2038 10394 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 2124 10394 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 2124 10394 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 2210 10394 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 2210 10394 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 2296 10394 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 2296 10394 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 2382 10394 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 2382 10394 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 2468 10394 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 2468 10394 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 2554 10394 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 2554 10394 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 2640 10394 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 2640 10394 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 1780 10394 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 1780 10394 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 1866 10394 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 1866 10394 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10330 1952 10394 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10330 1952 10394 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 2038 10476 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 2038 10476 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 2124 10476 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 2124 10476 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 2210 10476 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 2210 10476 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 2296 10476 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 2296 10476 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 2382 10476 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 2382 10476 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 2468 10476 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 2468 10476 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 2554 10476 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 2554 10476 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 2640 10476 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 2640 10476 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 1780 10476 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 1780 10476 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 1866 10476 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 1866 10476 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10412 1952 10476 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10412 1952 10476 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 2038 10558 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 2038 10558 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 2124 10558 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 2124 10558 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 2210 10558 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 2210 10558 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 2296 10558 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 2296 10558 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 2382 10558 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 2382 10558 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 2468 10558 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 2468 10558 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 2554 10558 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 2554 10558 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 2640 10558 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 2640 10558 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 1780 10558 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 1780 10558 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 1866 10558 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 1866 10558 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10494 1952 10558 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10494 1952 10558 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 2038 10640 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 2038 10640 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 2124 10640 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 2124 10640 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 2210 10640 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 2210 10640 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 2296 10640 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 2296 10640 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 2382 10640 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 2382 10640 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 2468 10640 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 2468 10640 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 2554 10640 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 2554 10640 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 2640 10640 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 2640 10640 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 1780 10640 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 1780 10640 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 1866 10640 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 1866 10640 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10576 1952 10640 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10576 1952 10640 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 2038 10721 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 2038 10721 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 2124 10721 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 2124 10721 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 2210 10721 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 2210 10721 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 2296 10721 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 2296 10721 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 2382 10721 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 2382 10721 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 2468 10721 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 2468 10721 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 2554 10721 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 2554 10721 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 2640 10721 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 2640 10721 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 1780 10721 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 1780 10721 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 1866 10721 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 1866 10721 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10657 1952 10721 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10657 1952 10721 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 2038 10802 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 2038 10802 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 2124 10802 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 2124 10802 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 2210 10802 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 2210 10802 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 2296 10802 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 2296 10802 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 2382 10802 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 2382 10802 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 2468 10802 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 2468 10802 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 2554 10802 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 2554 10802 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 2640 10802 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 2640 10802 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 1780 10802 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 1780 10802 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 1866 10802 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 1866 10802 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10738 1952 10802 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10738 1952 10802 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 2038 10883 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 2038 10883 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 2124 10883 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 2124 10883 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 2210 10883 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 2210 10883 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 2296 10883 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 2296 10883 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 2382 10883 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 2382 10883 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 2468 10883 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 2468 10883 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 2554 10883 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 2554 10883 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 2640 10883 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 2640 10883 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 1780 10883 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 1780 10883 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 1866 10883 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 1866 10883 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10819 1952 10883 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10819 1952 10883 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 2038 10964 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 2038 10964 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 2124 10964 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 2124 10964 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 2210 10964 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 2210 10964 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 2296 10964 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 2296 10964 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 2382 10964 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 2382 10964 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 2468 10964 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 2468 10964 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 2554 10964 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 2554 10964 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 2640 10964 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 2640 10964 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 1780 10964 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 1780 10964 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 1866 10964 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 1866 10964 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10900 1952 10964 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10900 1952 10964 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 2038 11045 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 2038 11045 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 2124 11045 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 2124 11045 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 2210 11045 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 2210 11045 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 2296 11045 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 2296 11045 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 2382 11045 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 2382 11045 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 2468 11045 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 2468 11045 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 2554 11045 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 2554 11045 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 2640 11045 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 2640 11045 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 1780 11045 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 1780 11045 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 1866 11045 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 1866 11045 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 10981 1952 11045 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 10981 1952 11045 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 2038 11126 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 2038 11126 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 2124 11126 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 2124 11126 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 2210 11126 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 2210 11126 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 2296 11126 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 2296 11126 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 2382 11126 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 2382 11126 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 2468 11126 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 2468 11126 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 2554 11126 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 2554 11126 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 2640 11126 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 2640 11126 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 1780 11126 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 1780 11126 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 1866 11126 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 1866 11126 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11062 1952 11126 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11062 1952 11126 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 2038 11207 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 2038 11207 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 2124 11207 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 2124 11207 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 2210 11207 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 2210 11207 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 2296 11207 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 2296 11207 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 2382 11207 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 2382 11207 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 2468 11207 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 2468 11207 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 2554 11207 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 2554 11207 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 2640 11207 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 2640 11207 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 1780 11207 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 1780 11207 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 1866 11207 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 1866 11207 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11143 1952 11207 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11143 1952 11207 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 2038 11288 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 2038 11288 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 2124 11288 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 2124 11288 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 2210 11288 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 2210 11288 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 2296 11288 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 2296 11288 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 2382 11288 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 2382 11288 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 2468 11288 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 2468 11288 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 2554 11288 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 2554 11288 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 2640 11288 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 2640 11288 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 1780 11288 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 1780 11288 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 1866 11288 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 1866 11288 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11224 1952 11288 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11224 1952 11288 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 2038 11369 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 2038 11369 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 2124 11369 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 2124 11369 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 2210 11369 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 2210 11369 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 2296 11369 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 2296 11369 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 2382 11369 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 2382 11369 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 2468 11369 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 2468 11369 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 2554 11369 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 2554 11369 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 2640 11369 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 2640 11369 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 1780 11369 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 1780 11369 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 1866 11369 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 1866 11369 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11305 1952 11369 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11305 1952 11369 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 2038 11450 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 2038 11450 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 2124 11450 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 2124 11450 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 2210 11450 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 2210 11450 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 2296 11450 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 2296 11450 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 2382 11450 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 2382 11450 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 2468 11450 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 2468 11450 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 2554 11450 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 2554 11450 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 2640 11450 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 2640 11450 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 1780 11450 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 1780 11450 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 1866 11450 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 1866 11450 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11386 1952 11450 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11386 1952 11450 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 2038 11531 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 2038 11531 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 2124 11531 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 2124 11531 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 2210 11531 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 2210 11531 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 2296 11531 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 2296 11531 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 2382 11531 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 2382 11531 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 2468 11531 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 2468 11531 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 2554 11531 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 2554 11531 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 2640 11531 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 2640 11531 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 1780 11531 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 1780 11531 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 1866 11531 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 1866 11531 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11467 1952 11531 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11467 1952 11531 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 2038 11612 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 2038 11612 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 2124 11612 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 2124 11612 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 2210 11612 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 2210 11612 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 2296 11612 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 2296 11612 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 2382 11612 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 2382 11612 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 2468 11612 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 2468 11612 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 2554 11612 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 2554 11612 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 2640 11612 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 2640 11612 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 1780 11612 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 1780 11612 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 1866 11612 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 1866 11612 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11548 1952 11612 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11548 1952 11612 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 2038 11693 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 2038 11693 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 2124 11693 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 2124 11693 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 2210 11693 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 2210 11693 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 2296 11693 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 2296 11693 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 2382 11693 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 2382 11693 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 2468 11693 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 2468 11693 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 2554 11693 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 2554 11693 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 2640 11693 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 2640 11693 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 1780 11693 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 1780 11693 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 1866 11693 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 1866 11693 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11629 1952 11693 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11629 1952 11693 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 2038 11774 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 2038 11774 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 2124 11774 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 2124 11774 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 2210 11774 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 2210 11774 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 2296 11774 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 2296 11774 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 2382 11774 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 2382 11774 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 2468 11774 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 2468 11774 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 2554 11774 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 2554 11774 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 2640 11774 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 2640 11774 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 1780 11774 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 1780 11774 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 1866 11774 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 1866 11774 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11710 1952 11774 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11710 1952 11774 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 2038 11855 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 2038 11855 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 2124 11855 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 2124 11855 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 2210 11855 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 2210 11855 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 2296 11855 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 2296 11855 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 2382 11855 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 2382 11855 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 2468 11855 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 2468 11855 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 2554 11855 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 2554 11855 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 2640 11855 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 2640 11855 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 1780 11855 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 1780 11855 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 1866 11855 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 1866 11855 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11791 1952 11855 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11791 1952 11855 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 2038 11936 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 2038 11936 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 2124 11936 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 2124 11936 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 2210 11936 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 2210 11936 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 2296 11936 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 2296 11936 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 2382 11936 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 2382 11936 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 2468 11936 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 2468 11936 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 2554 11936 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 2554 11936 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 2640 11936 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 2640 11936 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 1780 11936 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 1780 11936 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 1866 11936 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 1866 11936 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11872 1952 11936 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11872 1952 11936 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 2038 12017 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 2038 12017 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 2124 12017 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 2124 12017 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 2210 12017 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 2210 12017 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 2296 12017 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 2296 12017 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 2382 12017 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 2382 12017 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 2468 12017 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 2468 12017 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 2554 12017 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 2554 12017 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 2640 12017 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 2640 12017 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 1780 12017 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 1780 12017 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 1866 12017 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 1866 12017 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 11953 1952 12017 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 11953 1952 12017 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 2038 1309 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 2038 1309 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 2124 1309 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 2124 1309 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 2210 1309 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 2210 1309 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 2296 1309 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 2296 1309 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 2382 1309 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 2382 1309 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 2468 1309 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 2468 1309 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 2554 1309 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 2554 1309 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 2640 1309 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 2640 1309 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 1780 1309 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 1780 1309 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 1866 1309 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 1866 1309 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1245 1952 1309 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1245 1952 1309 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 2038 1390 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 2038 1390 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 2124 1390 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 2124 1390 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 2210 1390 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 2210 1390 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 2296 1390 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 2296 1390 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 2382 1390 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 2382 1390 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 2468 1390 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 2468 1390 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 2554 1390 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 2554 1390 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 2640 1390 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 2640 1390 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 1780 1390 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 1780 1390 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 1866 1390 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 1866 1390 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1326 1952 1390 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1326 1952 1390 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 2038 12098 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 2038 12098 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 2124 12098 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 2124 12098 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 2210 12098 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 2210 12098 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 2296 12098 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 2296 12098 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 2382 12098 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 2382 12098 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 2468 12098 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 2468 12098 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 2554 12098 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 2554 12098 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 2640 12098 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 2640 12098 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 1780 12098 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 1780 12098 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 1866 12098 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 1866 12098 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12034 1952 12098 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12034 1952 12098 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 2038 12179 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 2038 12179 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 2124 12179 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 2124 12179 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 2210 12179 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 2210 12179 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 2296 12179 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 2296 12179 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 2382 12179 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 2382 12179 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 2468 12179 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 2468 12179 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 2554 12179 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 2554 12179 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 2640 12179 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 2640 12179 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 1780 12179 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 1780 12179 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 1866 12179 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 1866 12179 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12115 1952 12179 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12115 1952 12179 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 2038 12260 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 2038 12260 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 2124 12260 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 2124 12260 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 2210 12260 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 2210 12260 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 2296 12260 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 2296 12260 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 2382 12260 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 2382 12260 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 2468 12260 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 2468 12260 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 2554 12260 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 2554 12260 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 2640 12260 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 2640 12260 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 1780 12260 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 1780 12260 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 1866 12260 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 1866 12260 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12196 1952 12260 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12196 1952 12260 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 2038 12341 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 2038 12341 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 2124 12341 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 2124 12341 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 2210 12341 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 2210 12341 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 2296 12341 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 2296 12341 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 2382 12341 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 2382 12341 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 2468 12341 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 2468 12341 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 2554 12341 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 2554 12341 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 2640 12341 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 2640 12341 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 1780 12341 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 1780 12341 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 1866 12341 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 1866 12341 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12277 1952 12341 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12277 1952 12341 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 2038 12422 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 2038 12422 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 2124 12422 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 2124 12422 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 2210 12422 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 2210 12422 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 2296 12422 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 2296 12422 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 2382 12422 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 2382 12422 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 2468 12422 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 2468 12422 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 2554 12422 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 2554 12422 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 2640 12422 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 2640 12422 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 1780 12422 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 1780 12422 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 1866 12422 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 1866 12422 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12358 1952 12422 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12358 1952 12422 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 2038 12503 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 2038 12503 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 2124 12503 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 2124 12503 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 2210 12503 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 2210 12503 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 2296 12503 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 2296 12503 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 2382 12503 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 2382 12503 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 2468 12503 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 2468 12503 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 2554 12503 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 2554 12503 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 2640 12503 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 2640 12503 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 1780 12503 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 1780 12503 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 1866 12503 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 1866 12503 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12439 1952 12503 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12439 1952 12503 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 2038 12584 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 2038 12584 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 2124 12584 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 2124 12584 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 2210 12584 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 2210 12584 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 2296 12584 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 2296 12584 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 2382 12584 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 2382 12584 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 2468 12584 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 2468 12584 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 2554 12584 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 2554 12584 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 2640 12584 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 2640 12584 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 1780 12584 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 1780 12584 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 1866 12584 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 1866 12584 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12520 1952 12584 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12520 1952 12584 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 2038 12665 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 2038 12665 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 2124 12665 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 2124 12665 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 2210 12665 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 2210 12665 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 2296 12665 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 2296 12665 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 2382 12665 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 2382 12665 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 2468 12665 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 2468 12665 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 2554 12665 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 2554 12665 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 2640 12665 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 2640 12665 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 1780 12665 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 1780 12665 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 1866 12665 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 1866 12665 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12601 1952 12665 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12601 1952 12665 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 2038 12746 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 2038 12746 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 2124 12746 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 2124 12746 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 2210 12746 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 2210 12746 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 2296 12746 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 2296 12746 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 2382 12746 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 2382 12746 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 2468 12746 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 2468 12746 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 2554 12746 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 2554 12746 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 2640 12746 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 2640 12746 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 1780 12746 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 1780 12746 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 1866 12746 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 1866 12746 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12682 1952 12746 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12682 1952 12746 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 2038 12827 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 2038 12827 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 2124 12827 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 2124 12827 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 2210 12827 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 2210 12827 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 2296 12827 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 2296 12827 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 2382 12827 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 2382 12827 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 2468 12827 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 2468 12827 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 2554 12827 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 2554 12827 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 2640 12827 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 2640 12827 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 1780 12827 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 1780 12827 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 1866 12827 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 1866 12827 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12763 1952 12827 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12763 1952 12827 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 2038 12908 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 2038 12908 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 2124 12908 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 2124 12908 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 2210 12908 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 2210 12908 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 2296 12908 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 2296 12908 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 2382 12908 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 2382 12908 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 2468 12908 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 2468 12908 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 2554 12908 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 2554 12908 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 2640 12908 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 2640 12908 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 1780 12908 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 1780 12908 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 1866 12908 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 1866 12908 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12844 1952 12908 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12844 1952 12908 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 2038 12989 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 2038 12989 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 2124 12989 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 2124 12989 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 2210 12989 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 2210 12989 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 2296 12989 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 2296 12989 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 2382 12989 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 2382 12989 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 2468 12989 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 2468 12989 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 2554 12989 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 2554 12989 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 2640 12989 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 2640 12989 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 1780 12989 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 1780 12989 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 1866 12989 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 1866 12989 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 12925 1952 12989 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 12925 1952 12989 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 2038 13070 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 2038 13070 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 2124 13070 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 2124 13070 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 2210 13070 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 2210 13070 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 2296 13070 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 2296 13070 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 2382 13070 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 2382 13070 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 2468 13070 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 2468 13070 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 2554 13070 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 2554 13070 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 2640 13070 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 2640 13070 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 1780 13070 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 1780 13070 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 1866 13070 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 1866 13070 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13006 1952 13070 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13006 1952 13070 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 2038 13151 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 2038 13151 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 2124 13151 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 2124 13151 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 2210 13151 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 2210 13151 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 2296 13151 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 2296 13151 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 2382 13151 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 2382 13151 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 2468 13151 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 2468 13151 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 2554 13151 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 2554 13151 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 2640 13151 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 2640 13151 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 1780 13151 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 1780 13151 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 1866 13151 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 1866 13151 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13087 1952 13151 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13087 1952 13151 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 2038 13232 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 2038 13232 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 2124 13232 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 2124 13232 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 2210 13232 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 2210 13232 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 2296 13232 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 2296 13232 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 2382 13232 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 2382 13232 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 2468 13232 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 2468 13232 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 2554 13232 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 2554 13232 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 2640 13232 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 2640 13232 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 1780 13232 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 1780 13232 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 1866 13232 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 1866 13232 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13168 1952 13232 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13168 1952 13232 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 2038 13313 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 2038 13313 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 2124 13313 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 2124 13313 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 2210 13313 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 2210 13313 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 2296 13313 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 2296 13313 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 2382 13313 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 2382 13313 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 2468 13313 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 2468 13313 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 2554 13313 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 2554 13313 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 2640 13313 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 2640 13313 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 1780 13313 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 1780 13313 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 1866 13313 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 1866 13313 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13249 1952 13313 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13249 1952 13313 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 2038 13394 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 2038 13394 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 2124 13394 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 2124 13394 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 2210 13394 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 2210 13394 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 2296 13394 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 2296 13394 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 2382 13394 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 2382 13394 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 2468 13394 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 2468 13394 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 2554 13394 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 2554 13394 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 2640 13394 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 2640 13394 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 1780 13394 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 1780 13394 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 1866 13394 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 1866 13394 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13330 1952 13394 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13330 1952 13394 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 2038 13475 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 2038 13475 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 2124 13475 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 2124 13475 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 2210 13475 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 2210 13475 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 2296 13475 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 2296 13475 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 2382 13475 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 2382 13475 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 2468 13475 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 2468 13475 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 2554 13475 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 2554 13475 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 2640 13475 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 2640 13475 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 1780 13475 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 1780 13475 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 1866 13475 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 1866 13475 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13411 1952 13475 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13411 1952 13475 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 2038 13556 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 2038 13556 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 2124 13556 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 2124 13556 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 2210 13556 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 2210 13556 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 2296 13556 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 2296 13556 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 2382 13556 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 2382 13556 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 2468 13556 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 2468 13556 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 2554 13556 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 2554 13556 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 2640 13556 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 2640 13556 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 1780 13556 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 1780 13556 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 1866 13556 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 1866 13556 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13492 1952 13556 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13492 1952 13556 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 2038 13637 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 2038 13637 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 2124 13637 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 2124 13637 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 2210 13637 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 2210 13637 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 2296 13637 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 2296 13637 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 2382 13637 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 2382 13637 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 2468 13637 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 2468 13637 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 2554 13637 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 2554 13637 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 2640 13637 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 2640 13637 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 1780 13637 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 1780 13637 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 1866 13637 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 1866 13637 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13573 1952 13637 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13573 1952 13637 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 2038 13718 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 2038 13718 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 2124 13718 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 2124 13718 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 2210 13718 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 2210 13718 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 2296 13718 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 2296 13718 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 2382 13718 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 2382 13718 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 2468 13718 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 2468 13718 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 2554 13718 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 2554 13718 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 2640 13718 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 2640 13718 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 1780 13718 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 1780 13718 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 1866 13718 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 1866 13718 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13654 1952 13718 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13654 1952 13718 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 2038 13799 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 2038 13799 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 2124 13799 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 2124 13799 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 2210 13799 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 2210 13799 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 2296 13799 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 2296 13799 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 2382 13799 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 2382 13799 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 2468 13799 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 2468 13799 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 2554 13799 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 2554 13799 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 2640 13799 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 2640 13799 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 1780 13799 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 1780 13799 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 1866 13799 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 1866 13799 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13735 1952 13799 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13735 1952 13799 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 2038 13880 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 2038 13880 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 2124 13880 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 2124 13880 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 2210 13880 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 2210 13880 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 2296 13880 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 2296 13880 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 2382 13880 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 2382 13880 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 2468 13880 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 2468 13880 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 2554 13880 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 2554 13880 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 2640 13880 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 2640 13880 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 1780 13880 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 1780 13880 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 1866 13880 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 1866 13880 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13816 1952 13880 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13816 1952 13880 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 2038 13961 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 2038 13961 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 2124 13961 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 2124 13961 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 2210 13961 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 2210 13961 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 2296 13961 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 2296 13961 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 2382 13961 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 2382 13961 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 2468 13961 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 2468 13961 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 2554 13961 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 2554 13961 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 2640 13961 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 2640 13961 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 1780 13961 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 1780 13961 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 1866 13961 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 1866 13961 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13897 1952 13961 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13897 1952 13961 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 2038 14042 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 2038 14042 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 2124 14042 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 2124 14042 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 2210 14042 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 2210 14042 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 2296 14042 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 2296 14042 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 2382 14042 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 2382 14042 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 2468 14042 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 2468 14042 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 2554 14042 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 2554 14042 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 2640 14042 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 2640 14042 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 1780 14042 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 1780 14042 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 1866 14042 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 1866 14042 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 13978 1952 14042 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 13978 1952 14042 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 2038 1471 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 2038 1471 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 2124 1471 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 2124 1471 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 2210 1471 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 2210 1471 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 2296 1471 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 2296 1471 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 2382 1471 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 2382 1471 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 2468 1471 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 2468 1471 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 2554 1471 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 2554 1471 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 2640 1471 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 2640 1471 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 1780 1471 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 1780 1471 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 1866 1471 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 1866 1471 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1407 1952 1471 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1407 1952 1471 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 2038 1552 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 2038 1552 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 2124 1552 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 2124 1552 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 2210 1552 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 2210 1552 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 2296 1552 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 2296 1552 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 2382 1552 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 2382 1552 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 2468 1552 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 2468 1552 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 2554 1552 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 2554 1552 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 2640 1552 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 2640 1552 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 1780 1552 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 1780 1552 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 1866 1552 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 1866 1552 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1488 1952 1552 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1488 1952 1552 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 2038 1633 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 2038 1633 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 2124 1633 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 2124 1633 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 2210 1633 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 2210 1633 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 2296 1633 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 2296 1633 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 2382 1633 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 2382 1633 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 2468 1633 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 2468 1633 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 2554 1633 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 2554 1633 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 2640 1633 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 2640 1633 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 1780 1633 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 1780 1633 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 1866 1633 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 1866 1633 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1569 1952 1633 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1569 1952 1633 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 2038 14123 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 2038 14123 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 2124 14123 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 2124 14123 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 2210 14123 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 2210 14123 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 2296 14123 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 2296 14123 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 2382 14123 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 2382 14123 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 2468 14123 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 2468 14123 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 2554 14123 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 2554 14123 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 2640 14123 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 2640 14123 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 1780 14123 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 1780 14123 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 1866 14123 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 1866 14123 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14059 1952 14123 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14059 1952 14123 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 2038 14204 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 2038 14204 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 2124 14204 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 2124 14204 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 2210 14204 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 2210 14204 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 2296 14204 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 2296 14204 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 2382 14204 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 2382 14204 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 2468 14204 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 2468 14204 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 2554 14204 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 2554 14204 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 2640 14204 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 2640 14204 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 1780 14204 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 1780 14204 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 1866 14204 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 1866 14204 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14140 1952 14204 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14140 1952 14204 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 2038 14285 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 2038 14285 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 2124 14285 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 2124 14285 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 2210 14285 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 2210 14285 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 2296 14285 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 2296 14285 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 2382 14285 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 2382 14285 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 2468 14285 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 2468 14285 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 2554 14285 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 2554 14285 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 2640 14285 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 2640 14285 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 1780 14285 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 1780 14285 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 1866 14285 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 1866 14285 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14221 1952 14285 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14221 1952 14285 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 2038 14366 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 2038 14366 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 2124 14366 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 2124 14366 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 2210 14366 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 2210 14366 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 2296 14366 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 2296 14366 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 2382 14366 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 2382 14366 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 2468 14366 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 2468 14366 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 2554 14366 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 2554 14366 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 2640 14366 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 2640 14366 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 1780 14366 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 1780 14366 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 1866 14366 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 1866 14366 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14302 1952 14366 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14302 1952 14366 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 2038 14447 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 2038 14447 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 2124 14447 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 2124 14447 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 2210 14447 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 2210 14447 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 2296 14447 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 2296 14447 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 2382 14447 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 2382 14447 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 2468 14447 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 2468 14447 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 2554 14447 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 2554 14447 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 2640 14447 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 2640 14447 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 1780 14447 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 1780 14447 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 1866 14447 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 1866 14447 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14383 1952 14447 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14383 1952 14447 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 2038 14528 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 2038 14528 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 2124 14528 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 2124 14528 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 2210 14528 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 2210 14528 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 2296 14528 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 2296 14528 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 2382 14528 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 2382 14528 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 2468 14528 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 2468 14528 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 2554 14528 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 2554 14528 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 2640 14528 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 2640 14528 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 1780 14528 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 1780 14528 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 1866 14528 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 1866 14528 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14464 1952 14528 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14464 1952 14528 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 2038 14609 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 2038 14609 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 2124 14609 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 2124 14609 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 2210 14609 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 2210 14609 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 2296 14609 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 2296 14609 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 2382 14609 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 2382 14609 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 2468 14609 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 2468 14609 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 2554 14609 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 2554 14609 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 2640 14609 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 2640 14609 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 1780 14609 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 1780 14609 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 1866 14609 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 1866 14609 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14545 1952 14609 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14545 1952 14609 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 2038 14690 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 2038 14690 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 2124 14690 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 2124 14690 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 2210 14690 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 2210 14690 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 2296 14690 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 2296 14690 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 2382 14690 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 2382 14690 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 2468 14690 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 2468 14690 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 2554 14690 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 2554 14690 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 2640 14690 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 2640 14690 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 1780 14690 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 1780 14690 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 1866 14690 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 1866 14690 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14626 1952 14690 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14626 1952 14690 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 2038 14771 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 2038 14771 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 2124 14771 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 2124 14771 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 2210 14771 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 2210 14771 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 2296 14771 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 2296 14771 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 2382 14771 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 2382 14771 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 2468 14771 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 2468 14771 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 2554 14771 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 2554 14771 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 2640 14771 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 2640 14771 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 1780 14771 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 1780 14771 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 1866 14771 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 1866 14771 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14707 1952 14771 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14707 1952 14771 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 2038 14852 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 2038 14852 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 2124 14852 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 2124 14852 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 2210 14852 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 2210 14852 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 2296 14852 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 2296 14852 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 2382 14852 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 2382 14852 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 2468 14852 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 2468 14852 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 2554 14852 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 2554 14852 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 2640 14852 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 2640 14852 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 1780 14852 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 1780 14852 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 1866 14852 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 1866 14852 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14788 1952 14852 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 14788 1952 14852 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 2038 1714 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 2038 1714 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 2124 1714 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 2124 1714 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 2210 1714 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 2210 1714 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 2296 1714 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 2296 1714 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 2382 1714 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 2382 1714 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 2468 1714 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 2468 1714 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 2554 1714 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 2554 1714 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 2640 1714 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 2640 1714 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 1780 1714 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 1780 1714 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 1866 1714 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 1866 1714 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1650 1952 1714 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1650 1952 1714 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 2038 1795 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 2038 1795 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 2124 1795 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 2124 1795 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 2210 1795 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 2210 1795 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 2296 1795 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 2296 1795 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 2382 1795 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 2382 1795 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 2468 1795 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 2468 1795 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 2554 1795 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 2554 1795 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 2640 1795 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 2640 1795 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 1780 1795 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 1780 1795 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 1866 1795 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 1866 1795 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1731 1952 1795 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1731 1952 1795 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 2038 1876 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 2038 1876 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 2124 1876 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 2124 1876 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 2210 1876 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 2210 1876 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 2296 1876 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 2296 1876 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 2382 1876 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 2382 1876 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 2468 1876 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 2468 1876 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 2554 1876 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 2554 1876 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 2640 1876 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 2640 1876 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 1780 1876 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 1780 1876 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 1866 1876 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 1866 1876 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1812 1952 1876 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1812 1952 1876 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 2038 1957 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 2038 1957 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 2124 1957 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 2124 1957 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 2210 1957 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 2210 1957 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 2296 1957 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 2296 1957 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 2382 1957 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 2382 1957 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 2468 1957 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 2468 1957 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 2554 1957 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 2554 1957 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 2640 1957 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 2640 1957 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 1780 1957 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 1780 1957 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 1866 1957 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 1866 1957 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1893 1952 1957 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1893 1952 1957 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 2038 2038 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 2038 2038 2102 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 2124 2038 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 2124 2038 2188 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 2210 2038 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 2210 2038 2274 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 2296 2038 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 2296 2038 2360 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 2382 2038 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 2382 2038 2446 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 2468 2038 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 2468 2038 2532 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 2554 2038 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 2554 2038 2618 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 2640 2038 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 2640 2038 2704 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 1780 2038 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 1780 2038 1844 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 1866 2038 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 1866 2038 1930 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 1974 1952 2038 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal3 s 1974 1952 2038 2016 6 VCCD
port 3 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 9 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 40000
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 35411070
string GDS_START 35319534
<< end >>
