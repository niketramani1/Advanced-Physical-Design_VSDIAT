magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1285 -1110 1385 1411
<< labels >>
flabel comment s 125 150 125 150 0 FreeSans 300 0 0 0 D
flabel comment s -25 150 -25 150 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 2025948
string GDS_START 2025308
<< end >>
