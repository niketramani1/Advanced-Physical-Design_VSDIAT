magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1531 -1464 41260 42060
<< obsactive >>
tri 25423 26223 40000 40800 ne
<< metal4 >>
rect 0 35957 287 40800
rect 0 14807 529 19800
rect 0 13617 296 14507
rect 0 12447 325 13337
rect 0 12081 4635 12147
rect 0 11425 100 12021
rect 0 11129 4310 11365
rect 0 10473 116 11069
rect 0 10347 3915 10413
rect 0 9117 295 10047
rect 0 8147 267 8837
rect 0 7177 277 7867
rect 0 5967 254 6897
rect 0 4757 305 5687
rect 0 3787 294 4477
rect 0 2577 757 3507
rect 0 1207 470 2297
rect 407 0 1497 254
rect 1777 0 2707 254
rect 2987 0 3677 254
rect 3957 0 4887 254
rect 5167 0 6097 254
rect 6377 0 7067 254
rect 7347 0 8037 254
rect 8317 0 9247 254
rect 9547 0 9613 4715
rect 9673 0 10269 4175
rect 10329 0 10565 4311
rect 10625 0 11221 5382
rect 11281 0 11347 5435
rect 11647 0 12537 254
rect 12817 0 13707 254
rect 14007 0 19000 371
rect 35157 0 40000 254
<< metal5 >>
rect 0 35957 254 40800
rect 0 14807 254 19797
rect 0 13637 254 14487
rect 0 12467 254 13317
rect 0 10347 254 12147
rect 0 9137 254 10027
rect 0 8167 254 8817
rect 0 7197 254 7847
rect 0 5987 254 6877
rect 0 4777 305 5667
rect 0 3807 254 4457
rect 0 2597 254 3487
rect 0 1227 254 2277
rect 427 0 1477 254
rect 1797 0 2687 254
rect 3007 0 3657 254
rect 3977 0 4867 254
rect 5187 0 6077 254
rect 6397 0 7047 254
rect 7367 0 8017 254
rect 8337 0 9227 254
rect 9547 0 11347 5431
rect 11667 0 12517 254
rect 12837 0 13687 254
rect 14007 0 18997 371
rect 35157 0 40000 254
<< fillblock >>
tri 25423 26223 40000 40800 ne
use sky130_fd_io__corner_bus_overlay  sky130_fd_io__corner_bus_overlay_0
timestamp 1624855509
transform 1 0 0 0 1 67
box 0 0 40000 40733
<< labels >>
flabel metal4 s 0 11425 100 12021 3 FreeSans 650 0 0 0 AMUXBUS_A
port 1 nsew signal bidirectional
flabel metal4 s 10625 0 11221 100 3 FreeSans 650 90 0 0 AMUXBUS_A
port 1 nsew signal bidirectional
flabel metal4 s 0 10473 115 11069 3 FreeSans 650 0 0 0 AMUXBUS_B
port 2 nsew signal bidirectional
flabel metal4 s 9673 0 10269 115 3 FreeSans 650 90 0 0 AMUXBUS_B
port 2 nsew signal bidirectional
flabel metal5 s 0 10347 254 12147 3 FreeSans 650 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 127 11205 127 11205 3 FreeSans 650 180 0 0 VSSA
flabel metal5 s 0 8168 254 8817 3 FreeSans 650 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 10347 254 10413 3 FreeSans 650 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 8147 254 8837 3 FreeSans 650 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 11129 254 11365 3 FreeSans 650 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 12081 254 12147 3 FreeSans 650 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 7368 0 8017 254 3 FreeSans 650 270 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 9547 0 11347 254 3 FreeSans 650 270 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 10258 127 10258 127 3 FreeSans 650 90 0 0 VSSA
flabel metal4 s 11281 0 11347 254 3 FreeSans 650 90 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 10329 0 10565 254 3 FreeSans 650 90 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 7347 0 8037 254 3 FreeSans 650 270 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 9547 0 9613 254 3 FreeSans 650 90 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 0 3807 251 4457 3 FreeSans 650 180 0 0 VDDA
port 4 nsew power bidirectional
flabel metal4 s 0 3787 251 4477 3 FreeSans 650 180 0 0 VDDA
port 4 nsew power bidirectional
flabel metal5 s 3007 0 3657 251 3 FreeSans 650 270 0 0 VDDA
port 4 nsew power bidirectional
flabel metal4 s 2987 0 3677 251 3 FreeSans 650 270 0 0 VDDA
port 4 nsew power bidirectional
flabel metal5 s 0 7197 254 7847 3 FreeSans 650 180 0 0 VSWITCH
port 5 nsew power bidirectional
flabel metal4 s 0 7177 254 7867 3 FreeSans 650 180 0 0 VSWITCH
port 5 nsew power bidirectional
flabel metal5 s 6397 0 7047 254 3 FreeSans 650 270 0 0 VSWITCH
port 5 nsew power bidirectional
flabel metal4 s 6377 0 7067 254 3 FreeSans 650 270 0 0 VSWITCH
port 5 nsew power bidirectional
flabel metal5 s 0 13637 254 14487 3 FreeSans 650 180 0 0 VDDIO_Q
port 6 nsew power bidirectional
flabel metal4 s 0 13617 254 14507 3 FreeSans 650 180 0 0 VDDIO_Q
port 6 nsew power bidirectional
flabel metal5 s 12837 0 13687 254 3 FreeSans 650 270 0 0 VDDIO_Q
port 6 nsew power bidirectional
flabel metal4 s 12817 0 13707 254 3 FreeSans 650 270 0 0 VDDIO_Q
port 6 nsew power bidirectional
flabel metal5 s 0 1227 254 2277 3 FreeSans 650 180 0 0 VCCHIB
port 7 nsew power bidirectional
flabel metal4 s 0 1207 254 2297 3 FreeSans 650 180 0 0 VCCHIB
port 7 nsew power bidirectional
flabel metal5 s 427 0 1477 254 3 FreeSans 650 270 0 0 VCCHIB
port 7 nsew power bidirectional
flabel metal4 s 407 0 1497 254 3 FreeSans 650 270 0 0 VCCHIB
port 7 nsew power bidirectional
flabel metal5 s 0 14807 254 19797 3 FreeSans 650 180 0 0 VDDIO
port 8 nsew power bidirectional
flabel metal5 s 0 4777 254 5667 3 FreeSans 650 180 0 0 VDDIO
port 8 nsew power bidirectional
flabel metal4 s 0 4757 254 5687 3 FreeSans 650 180 0 0 VDDIO
port 8 nsew power bidirectional
flabel metal4 s 0 14808 254 19800 3 FreeSans 650 180 0 0 VDDIO
port 8 nsew power bidirectional
flabel metal5 s 3977 0 4867 254 3 FreeSans 650 270 0 0 VDDIO
port 8 nsew power bidirectional
flabel metal5 s 14007 0 18997 254 3 FreeSans 650 270 0 0 VDDIO
port 8 nsew power bidirectional
flabel metal4 s 14008 0 19000 254 3 FreeSans 650 270 0 0 VDDIO
port 8 nsew power bidirectional
flabel metal4 s 3957 0 4887 254 3 FreeSans 650 270 0 0 VDDIO
port 8 nsew power bidirectional
flabel metal5 s 0 2597 254 3487 3 FreeSans 650 180 0 0 VCCD
port 9 nsew power bidirectional
flabel metal4 s 0 2577 254 3507 3 FreeSans 650 180 0 0 VCCD
port 9 nsew power bidirectional
flabel metal5 s 1797 0 2687 254 3 FreeSans 650 270 0 0 VCCD
port 9 nsew power bidirectional
flabel metal4 s 1777 0 2707 254 3 FreeSans 650 270 0 0 VCCD
port 9 nsew power bidirectional
flabel metal5 s 0 5987 254 6877 3 FreeSans 650 180 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 0 5967 254 6897 3 FreeSans 650 180 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 0 35957 254 40800 3 FreeSans 650 180 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 127 38974 127 38974 3 FreeSans 650 180 0 0 VSSIO
flabel metal5 s 5187 0 6077 254 3 FreeSans 650 270 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 5167 0 6097 254 3 FreeSans 650 270 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 35157 0 40000 254 3 FreeSans 650 270 0 0 VSSIO
port 10 nsew ground bidirectional
flabel metal4 s 38174 127 38174 127 3 FreeSans 650 270 0 0 VSSIO
flabel metal5 s 0 9137 254 10027 3 FreeSans 650 180 0 0 VSSD
port 11 nsew ground bidirectional
flabel metal4 s 0 9117 254 10047 3 FreeSans 650 180 0 0 VSSD
port 11 nsew ground bidirectional
flabel metal5 s 8337 0 9227 254 3 FreeSans 650 270 0 0 VSSD
port 11 nsew ground bidirectional
flabel metal4 s 8317 0 9247 254 3 FreeSans 650 270 0 0 VSSD
port 11 nsew ground bidirectional
flabel metal5 s 0 12467 254 13317 3 FreeSans 650 180 0 0 VSSIO_Q
port 12 nsew ground bidirectional
flabel metal4 s 0 12447 254 13337 3 FreeSans 650 180 0 0 VSSIO_Q
port 12 nsew ground bidirectional
flabel metal5 s 11667 0 12517 254 3 FreeSans 650 270 0 0 VSSIO_Q
port 12 nsew ground bidirectional
flabel metal4 s 11647 0 12537 254 3 FreeSans 650 270 0 0 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 10625 0 11221 5382 1 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 9673 0 10269 4175 1 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal4 s 0 10347 3915 10413 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 8147 267 8837 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 11129 4310 11365 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 12081 4635 12147 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 7368 0 8017 254 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 9547 0 11347 5431 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 10257 126 10259 128 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 11281 0 11347 5435 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 10329 0 10565 4311 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 7347 0 8037 254 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 9547 0 9613 4715 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 3787 294 4477 1 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 3007 0 3657 251 1 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2987 0 3677 251 1 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 7177 277 7867 1 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 6397 0 7047 254 1 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 6377 0 7067 254 1 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 0 13617 296 14507 1 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 12837 0 13687 254 1 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 12817 0 13707 254 1 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 1207 470 2297 1 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 427 0 1477 254 1 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 407 0 1497 254 1 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 0 4777 305 5667 1 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 4757 305 5687 1 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 14807 529 19800 1 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 3977 0 4867 254 1 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14007 0 18997 371 1 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14007 0 19000 371 1 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 3957 0 4887 254 1 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 2577 757 3507 1 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 1797 0 2687 254 1 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 1777 0 2707 254 1 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 35957 287 40800 1 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 126 38973 128 38975 1 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 5187 0 6077 254 1 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 5167 0 6097 254 1 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 35157 0 40000 254 1 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 38173 126 38175 128 1 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 9117 295 10047 1 VSSD
port 11 nsew ground bidirectional
rlabel metal5 s 8337 0 9227 254 1 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 8317 0 9247 254 1 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 0 12447 325 13337 1 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal5 s 11667 0 12517 254 1 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 11647 0 12537 254 1 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string LEFclass ENDCAP TOPRIGHT
string FIXED_BBOX 0 0 40000 40800
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_END 1673972
string GDS_START 1661258
<< end >>
