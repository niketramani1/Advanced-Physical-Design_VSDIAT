magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1260 -1260 220024 145360
<< dnwell >>
rect 1730 1848 216936 142344
<< nwell >>
rect 1646 142260 217020 142428
rect 1646 1932 1814 142260
rect 216852 1932 217020 142260
rect 1646 1764 217020 1932
<< nsubdiff >>
rect 2041 142361 2091 142385
rect 2041 142327 2049 142361
rect 2083 142327 2091 142361
rect 2041 142303 2091 142327
rect 2377 142361 2427 142385
rect 2377 142327 2385 142361
rect 2419 142327 2427 142361
rect 2377 142303 2427 142327
rect 2713 142361 2763 142385
rect 2713 142327 2721 142361
rect 2755 142327 2763 142361
rect 2713 142303 2763 142327
rect 3049 142361 3099 142385
rect 3049 142327 3057 142361
rect 3091 142327 3099 142361
rect 3049 142303 3099 142327
rect 3385 142361 3435 142385
rect 3385 142327 3393 142361
rect 3427 142327 3435 142361
rect 3385 142303 3435 142327
rect 3721 142361 3771 142385
rect 3721 142327 3729 142361
rect 3763 142327 3771 142361
rect 3721 142303 3771 142327
rect 4057 142361 4107 142385
rect 4057 142327 4065 142361
rect 4099 142327 4107 142361
rect 4057 142303 4107 142327
rect 4393 142361 4443 142385
rect 4393 142327 4401 142361
rect 4435 142327 4443 142361
rect 4393 142303 4443 142327
rect 4729 142361 4779 142385
rect 4729 142327 4737 142361
rect 4771 142327 4779 142361
rect 4729 142303 4779 142327
rect 5065 142361 5115 142385
rect 5065 142327 5073 142361
rect 5107 142327 5115 142361
rect 5065 142303 5115 142327
rect 5401 142361 5451 142385
rect 5401 142327 5409 142361
rect 5443 142327 5451 142361
rect 5401 142303 5451 142327
rect 5737 142361 5787 142385
rect 5737 142327 5745 142361
rect 5779 142327 5787 142361
rect 5737 142303 5787 142327
rect 6073 142361 6123 142385
rect 6073 142327 6081 142361
rect 6115 142327 6123 142361
rect 6073 142303 6123 142327
rect 6409 142361 6459 142385
rect 6409 142327 6417 142361
rect 6451 142327 6459 142361
rect 6409 142303 6459 142327
rect 6745 142361 6795 142385
rect 6745 142327 6753 142361
rect 6787 142327 6795 142361
rect 6745 142303 6795 142327
rect 7081 142361 7131 142385
rect 7081 142327 7089 142361
rect 7123 142327 7131 142361
rect 7081 142303 7131 142327
rect 7417 142361 7467 142385
rect 7417 142327 7425 142361
rect 7459 142327 7467 142361
rect 7417 142303 7467 142327
rect 7753 142361 7803 142385
rect 7753 142327 7761 142361
rect 7795 142327 7803 142361
rect 7753 142303 7803 142327
rect 8089 142361 8139 142385
rect 8089 142327 8097 142361
rect 8131 142327 8139 142361
rect 8089 142303 8139 142327
rect 8425 142361 8475 142385
rect 8425 142327 8433 142361
rect 8467 142327 8475 142361
rect 8425 142303 8475 142327
rect 8761 142361 8811 142385
rect 8761 142327 8769 142361
rect 8803 142327 8811 142361
rect 8761 142303 8811 142327
rect 9097 142361 9147 142385
rect 9097 142327 9105 142361
rect 9139 142327 9147 142361
rect 9097 142303 9147 142327
rect 9433 142361 9483 142385
rect 9433 142327 9441 142361
rect 9475 142327 9483 142361
rect 9433 142303 9483 142327
rect 9769 142361 9819 142385
rect 9769 142327 9777 142361
rect 9811 142327 9819 142361
rect 9769 142303 9819 142327
rect 10105 142361 10155 142385
rect 10105 142327 10113 142361
rect 10147 142327 10155 142361
rect 10105 142303 10155 142327
rect 10441 142361 10491 142385
rect 10441 142327 10449 142361
rect 10483 142327 10491 142361
rect 10441 142303 10491 142327
rect 10777 142361 10827 142385
rect 10777 142327 10785 142361
rect 10819 142327 10827 142361
rect 10777 142303 10827 142327
rect 11113 142361 11163 142385
rect 11113 142327 11121 142361
rect 11155 142327 11163 142361
rect 11113 142303 11163 142327
rect 11449 142361 11499 142385
rect 11449 142327 11457 142361
rect 11491 142327 11499 142361
rect 11449 142303 11499 142327
rect 11785 142361 11835 142385
rect 11785 142327 11793 142361
rect 11827 142327 11835 142361
rect 11785 142303 11835 142327
rect 12121 142361 12171 142385
rect 12121 142327 12129 142361
rect 12163 142327 12171 142361
rect 12121 142303 12171 142327
rect 12457 142361 12507 142385
rect 12457 142327 12465 142361
rect 12499 142327 12507 142361
rect 12457 142303 12507 142327
rect 12793 142361 12843 142385
rect 12793 142327 12801 142361
rect 12835 142327 12843 142361
rect 12793 142303 12843 142327
rect 13129 142361 13179 142385
rect 13129 142327 13137 142361
rect 13171 142327 13179 142361
rect 13129 142303 13179 142327
rect 13465 142361 13515 142385
rect 13465 142327 13473 142361
rect 13507 142327 13515 142361
rect 13465 142303 13515 142327
rect 13801 142361 13851 142385
rect 13801 142327 13809 142361
rect 13843 142327 13851 142361
rect 13801 142303 13851 142327
rect 14137 142361 14187 142385
rect 14137 142327 14145 142361
rect 14179 142327 14187 142361
rect 14137 142303 14187 142327
rect 14473 142361 14523 142385
rect 14473 142327 14481 142361
rect 14515 142327 14523 142361
rect 14473 142303 14523 142327
rect 14809 142361 14859 142385
rect 14809 142327 14817 142361
rect 14851 142327 14859 142361
rect 14809 142303 14859 142327
rect 15145 142361 15195 142385
rect 15145 142327 15153 142361
rect 15187 142327 15195 142361
rect 15145 142303 15195 142327
rect 15481 142361 15531 142385
rect 15481 142327 15489 142361
rect 15523 142327 15531 142361
rect 15481 142303 15531 142327
rect 15817 142361 15867 142385
rect 15817 142327 15825 142361
rect 15859 142327 15867 142361
rect 15817 142303 15867 142327
rect 16153 142361 16203 142385
rect 16153 142327 16161 142361
rect 16195 142327 16203 142361
rect 16153 142303 16203 142327
rect 16489 142361 16539 142385
rect 16489 142327 16497 142361
rect 16531 142327 16539 142361
rect 16489 142303 16539 142327
rect 16825 142361 16875 142385
rect 16825 142327 16833 142361
rect 16867 142327 16875 142361
rect 16825 142303 16875 142327
rect 17161 142361 17211 142385
rect 17161 142327 17169 142361
rect 17203 142327 17211 142361
rect 17161 142303 17211 142327
rect 17497 142361 17547 142385
rect 17497 142327 17505 142361
rect 17539 142327 17547 142361
rect 17497 142303 17547 142327
rect 17833 142361 17883 142385
rect 17833 142327 17841 142361
rect 17875 142327 17883 142361
rect 17833 142303 17883 142327
rect 18169 142361 18219 142385
rect 18169 142327 18177 142361
rect 18211 142327 18219 142361
rect 18169 142303 18219 142327
rect 18505 142361 18555 142385
rect 18505 142327 18513 142361
rect 18547 142327 18555 142361
rect 18505 142303 18555 142327
rect 18841 142361 18891 142385
rect 18841 142327 18849 142361
rect 18883 142327 18891 142361
rect 18841 142303 18891 142327
rect 19177 142361 19227 142385
rect 19177 142327 19185 142361
rect 19219 142327 19227 142361
rect 19177 142303 19227 142327
rect 19513 142361 19563 142385
rect 19513 142327 19521 142361
rect 19555 142327 19563 142361
rect 19513 142303 19563 142327
rect 19849 142361 19899 142385
rect 19849 142327 19857 142361
rect 19891 142327 19899 142361
rect 19849 142303 19899 142327
rect 20185 142361 20235 142385
rect 20185 142327 20193 142361
rect 20227 142327 20235 142361
rect 20185 142303 20235 142327
rect 20521 142361 20571 142385
rect 20521 142327 20529 142361
rect 20563 142327 20571 142361
rect 20521 142303 20571 142327
rect 20857 142361 20907 142385
rect 20857 142327 20865 142361
rect 20899 142327 20907 142361
rect 20857 142303 20907 142327
rect 21193 142361 21243 142385
rect 21193 142327 21201 142361
rect 21235 142327 21243 142361
rect 21193 142303 21243 142327
rect 21529 142361 21579 142385
rect 21529 142327 21537 142361
rect 21571 142327 21579 142361
rect 21529 142303 21579 142327
rect 21865 142361 21915 142385
rect 21865 142327 21873 142361
rect 21907 142327 21915 142361
rect 21865 142303 21915 142327
rect 22201 142361 22251 142385
rect 22201 142327 22209 142361
rect 22243 142327 22251 142361
rect 22201 142303 22251 142327
rect 22537 142361 22587 142385
rect 22537 142327 22545 142361
rect 22579 142327 22587 142361
rect 22537 142303 22587 142327
rect 22873 142361 22923 142385
rect 22873 142327 22881 142361
rect 22915 142327 22923 142361
rect 22873 142303 22923 142327
rect 23209 142361 23259 142385
rect 23209 142327 23217 142361
rect 23251 142327 23259 142361
rect 23209 142303 23259 142327
rect 23545 142361 23595 142385
rect 23545 142327 23553 142361
rect 23587 142327 23595 142361
rect 23545 142303 23595 142327
rect 23881 142361 23931 142385
rect 23881 142327 23889 142361
rect 23923 142327 23931 142361
rect 23881 142303 23931 142327
rect 24217 142361 24267 142385
rect 24217 142327 24225 142361
rect 24259 142327 24267 142361
rect 24217 142303 24267 142327
rect 24553 142361 24603 142385
rect 24553 142327 24561 142361
rect 24595 142327 24603 142361
rect 24553 142303 24603 142327
rect 24889 142361 24939 142385
rect 24889 142327 24897 142361
rect 24931 142327 24939 142361
rect 24889 142303 24939 142327
rect 25225 142361 25275 142385
rect 25225 142327 25233 142361
rect 25267 142327 25275 142361
rect 25225 142303 25275 142327
rect 25561 142361 25611 142385
rect 25561 142327 25569 142361
rect 25603 142327 25611 142361
rect 25561 142303 25611 142327
rect 25897 142361 25947 142385
rect 25897 142327 25905 142361
rect 25939 142327 25947 142361
rect 25897 142303 25947 142327
rect 26233 142361 26283 142385
rect 26233 142327 26241 142361
rect 26275 142327 26283 142361
rect 26233 142303 26283 142327
rect 26569 142361 26619 142385
rect 26569 142327 26577 142361
rect 26611 142327 26619 142361
rect 26569 142303 26619 142327
rect 26905 142361 26955 142385
rect 26905 142327 26913 142361
rect 26947 142327 26955 142361
rect 26905 142303 26955 142327
rect 27241 142361 27291 142385
rect 27241 142327 27249 142361
rect 27283 142327 27291 142361
rect 27241 142303 27291 142327
rect 27577 142361 27627 142385
rect 27577 142327 27585 142361
rect 27619 142327 27627 142361
rect 27577 142303 27627 142327
rect 27913 142361 27963 142385
rect 27913 142327 27921 142361
rect 27955 142327 27963 142361
rect 27913 142303 27963 142327
rect 28249 142361 28299 142385
rect 28249 142327 28257 142361
rect 28291 142327 28299 142361
rect 28249 142303 28299 142327
rect 28585 142361 28635 142385
rect 28585 142327 28593 142361
rect 28627 142327 28635 142361
rect 28585 142303 28635 142327
rect 28921 142361 28971 142385
rect 28921 142327 28929 142361
rect 28963 142327 28971 142361
rect 28921 142303 28971 142327
rect 29257 142361 29307 142385
rect 29257 142327 29265 142361
rect 29299 142327 29307 142361
rect 29257 142303 29307 142327
rect 29593 142361 29643 142385
rect 29593 142327 29601 142361
rect 29635 142327 29643 142361
rect 29593 142303 29643 142327
rect 29929 142361 29979 142385
rect 29929 142327 29937 142361
rect 29971 142327 29979 142361
rect 29929 142303 29979 142327
rect 30265 142361 30315 142385
rect 30265 142327 30273 142361
rect 30307 142327 30315 142361
rect 30265 142303 30315 142327
rect 30601 142361 30651 142385
rect 30601 142327 30609 142361
rect 30643 142327 30651 142361
rect 30601 142303 30651 142327
rect 30937 142361 30987 142385
rect 30937 142327 30945 142361
rect 30979 142327 30987 142361
rect 30937 142303 30987 142327
rect 31273 142361 31323 142385
rect 31273 142327 31281 142361
rect 31315 142327 31323 142361
rect 31273 142303 31323 142327
rect 31609 142361 31659 142385
rect 31609 142327 31617 142361
rect 31651 142327 31659 142361
rect 31609 142303 31659 142327
rect 31945 142361 31995 142385
rect 31945 142327 31953 142361
rect 31987 142327 31995 142361
rect 31945 142303 31995 142327
rect 32281 142361 32331 142385
rect 32281 142327 32289 142361
rect 32323 142327 32331 142361
rect 32281 142303 32331 142327
rect 32617 142361 32667 142385
rect 32617 142327 32625 142361
rect 32659 142327 32667 142361
rect 32617 142303 32667 142327
rect 32953 142361 33003 142385
rect 32953 142327 32961 142361
rect 32995 142327 33003 142361
rect 32953 142303 33003 142327
rect 33289 142361 33339 142385
rect 33289 142327 33297 142361
rect 33331 142327 33339 142361
rect 33289 142303 33339 142327
rect 33625 142361 33675 142385
rect 33625 142327 33633 142361
rect 33667 142327 33675 142361
rect 33625 142303 33675 142327
rect 33961 142361 34011 142385
rect 33961 142327 33969 142361
rect 34003 142327 34011 142361
rect 33961 142303 34011 142327
rect 34297 142361 34347 142385
rect 34297 142327 34305 142361
rect 34339 142327 34347 142361
rect 34297 142303 34347 142327
rect 34633 142361 34683 142385
rect 34633 142327 34641 142361
rect 34675 142327 34683 142361
rect 34633 142303 34683 142327
rect 34969 142361 35019 142385
rect 34969 142327 34977 142361
rect 35011 142327 35019 142361
rect 34969 142303 35019 142327
rect 35305 142361 35355 142385
rect 35305 142327 35313 142361
rect 35347 142327 35355 142361
rect 35305 142303 35355 142327
rect 35641 142361 35691 142385
rect 35641 142327 35649 142361
rect 35683 142327 35691 142361
rect 35641 142303 35691 142327
rect 35977 142361 36027 142385
rect 35977 142327 35985 142361
rect 36019 142327 36027 142361
rect 35977 142303 36027 142327
rect 36313 142361 36363 142385
rect 36313 142327 36321 142361
rect 36355 142327 36363 142361
rect 36313 142303 36363 142327
rect 36649 142361 36699 142385
rect 36649 142327 36657 142361
rect 36691 142327 36699 142361
rect 36649 142303 36699 142327
rect 36985 142361 37035 142385
rect 36985 142327 36993 142361
rect 37027 142327 37035 142361
rect 36985 142303 37035 142327
rect 37321 142361 37371 142385
rect 37321 142327 37329 142361
rect 37363 142327 37371 142361
rect 37321 142303 37371 142327
rect 37657 142361 37707 142385
rect 37657 142327 37665 142361
rect 37699 142327 37707 142361
rect 37657 142303 37707 142327
rect 37993 142361 38043 142385
rect 37993 142327 38001 142361
rect 38035 142327 38043 142361
rect 37993 142303 38043 142327
rect 38329 142361 38379 142385
rect 38329 142327 38337 142361
rect 38371 142327 38379 142361
rect 38329 142303 38379 142327
rect 38665 142361 38715 142385
rect 38665 142327 38673 142361
rect 38707 142327 38715 142361
rect 38665 142303 38715 142327
rect 39001 142361 39051 142385
rect 39001 142327 39009 142361
rect 39043 142327 39051 142361
rect 39001 142303 39051 142327
rect 39337 142361 39387 142385
rect 39337 142327 39345 142361
rect 39379 142327 39387 142361
rect 39337 142303 39387 142327
rect 39673 142361 39723 142385
rect 39673 142327 39681 142361
rect 39715 142327 39723 142361
rect 39673 142303 39723 142327
rect 40009 142361 40059 142385
rect 40009 142327 40017 142361
rect 40051 142327 40059 142361
rect 40009 142303 40059 142327
rect 40345 142361 40395 142385
rect 40345 142327 40353 142361
rect 40387 142327 40395 142361
rect 40345 142303 40395 142327
rect 40681 142361 40731 142385
rect 40681 142327 40689 142361
rect 40723 142327 40731 142361
rect 40681 142303 40731 142327
rect 41017 142361 41067 142385
rect 41017 142327 41025 142361
rect 41059 142327 41067 142361
rect 41017 142303 41067 142327
rect 41353 142361 41403 142385
rect 41353 142327 41361 142361
rect 41395 142327 41403 142361
rect 41353 142303 41403 142327
rect 41689 142361 41739 142385
rect 41689 142327 41697 142361
rect 41731 142327 41739 142361
rect 41689 142303 41739 142327
rect 42025 142361 42075 142385
rect 42025 142327 42033 142361
rect 42067 142327 42075 142361
rect 42025 142303 42075 142327
rect 42361 142361 42411 142385
rect 42361 142327 42369 142361
rect 42403 142327 42411 142361
rect 42361 142303 42411 142327
rect 42697 142361 42747 142385
rect 42697 142327 42705 142361
rect 42739 142327 42747 142361
rect 42697 142303 42747 142327
rect 43033 142361 43083 142385
rect 43033 142327 43041 142361
rect 43075 142327 43083 142361
rect 43033 142303 43083 142327
rect 43369 142361 43419 142385
rect 43369 142327 43377 142361
rect 43411 142327 43419 142361
rect 43369 142303 43419 142327
rect 43705 142361 43755 142385
rect 43705 142327 43713 142361
rect 43747 142327 43755 142361
rect 43705 142303 43755 142327
rect 44041 142361 44091 142385
rect 44041 142327 44049 142361
rect 44083 142327 44091 142361
rect 44041 142303 44091 142327
rect 44377 142361 44427 142385
rect 44377 142327 44385 142361
rect 44419 142327 44427 142361
rect 44377 142303 44427 142327
rect 44713 142361 44763 142385
rect 44713 142327 44721 142361
rect 44755 142327 44763 142361
rect 44713 142303 44763 142327
rect 45049 142361 45099 142385
rect 45049 142327 45057 142361
rect 45091 142327 45099 142361
rect 45049 142303 45099 142327
rect 45385 142361 45435 142385
rect 45385 142327 45393 142361
rect 45427 142327 45435 142361
rect 45385 142303 45435 142327
rect 45721 142361 45771 142385
rect 45721 142327 45729 142361
rect 45763 142327 45771 142361
rect 45721 142303 45771 142327
rect 46057 142361 46107 142385
rect 46057 142327 46065 142361
rect 46099 142327 46107 142361
rect 46057 142303 46107 142327
rect 46393 142361 46443 142385
rect 46393 142327 46401 142361
rect 46435 142327 46443 142361
rect 46393 142303 46443 142327
rect 46729 142361 46779 142385
rect 46729 142327 46737 142361
rect 46771 142327 46779 142361
rect 46729 142303 46779 142327
rect 47065 142361 47115 142385
rect 47065 142327 47073 142361
rect 47107 142327 47115 142361
rect 47065 142303 47115 142327
rect 47401 142361 47451 142385
rect 47401 142327 47409 142361
rect 47443 142327 47451 142361
rect 47401 142303 47451 142327
rect 47737 142361 47787 142385
rect 47737 142327 47745 142361
rect 47779 142327 47787 142361
rect 47737 142303 47787 142327
rect 48073 142361 48123 142385
rect 48073 142327 48081 142361
rect 48115 142327 48123 142361
rect 48073 142303 48123 142327
rect 48409 142361 48459 142385
rect 48409 142327 48417 142361
rect 48451 142327 48459 142361
rect 48409 142303 48459 142327
rect 48745 142361 48795 142385
rect 48745 142327 48753 142361
rect 48787 142327 48795 142361
rect 48745 142303 48795 142327
rect 49081 142361 49131 142385
rect 49081 142327 49089 142361
rect 49123 142327 49131 142361
rect 49081 142303 49131 142327
rect 49417 142361 49467 142385
rect 49417 142327 49425 142361
rect 49459 142327 49467 142361
rect 49417 142303 49467 142327
rect 49753 142361 49803 142385
rect 49753 142327 49761 142361
rect 49795 142327 49803 142361
rect 49753 142303 49803 142327
rect 50089 142361 50139 142385
rect 50089 142327 50097 142361
rect 50131 142327 50139 142361
rect 50089 142303 50139 142327
rect 50425 142361 50475 142385
rect 50425 142327 50433 142361
rect 50467 142327 50475 142361
rect 50425 142303 50475 142327
rect 50761 142361 50811 142385
rect 50761 142327 50769 142361
rect 50803 142327 50811 142361
rect 50761 142303 50811 142327
rect 51097 142361 51147 142385
rect 51097 142327 51105 142361
rect 51139 142327 51147 142361
rect 51097 142303 51147 142327
rect 51433 142361 51483 142385
rect 51433 142327 51441 142361
rect 51475 142327 51483 142361
rect 51433 142303 51483 142327
rect 51769 142361 51819 142385
rect 51769 142327 51777 142361
rect 51811 142327 51819 142361
rect 51769 142303 51819 142327
rect 52105 142361 52155 142385
rect 52105 142327 52113 142361
rect 52147 142327 52155 142361
rect 52105 142303 52155 142327
rect 52441 142361 52491 142385
rect 52441 142327 52449 142361
rect 52483 142327 52491 142361
rect 52441 142303 52491 142327
rect 52777 142361 52827 142385
rect 52777 142327 52785 142361
rect 52819 142327 52827 142361
rect 52777 142303 52827 142327
rect 53113 142361 53163 142385
rect 53113 142327 53121 142361
rect 53155 142327 53163 142361
rect 53113 142303 53163 142327
rect 53449 142361 53499 142385
rect 53449 142327 53457 142361
rect 53491 142327 53499 142361
rect 53449 142303 53499 142327
rect 53785 142361 53835 142385
rect 53785 142327 53793 142361
rect 53827 142327 53835 142361
rect 53785 142303 53835 142327
rect 54121 142361 54171 142385
rect 54121 142327 54129 142361
rect 54163 142327 54171 142361
rect 54121 142303 54171 142327
rect 54457 142361 54507 142385
rect 54457 142327 54465 142361
rect 54499 142327 54507 142361
rect 54457 142303 54507 142327
rect 54793 142361 54843 142385
rect 54793 142327 54801 142361
rect 54835 142327 54843 142361
rect 54793 142303 54843 142327
rect 55129 142361 55179 142385
rect 55129 142327 55137 142361
rect 55171 142327 55179 142361
rect 55129 142303 55179 142327
rect 55465 142361 55515 142385
rect 55465 142327 55473 142361
rect 55507 142327 55515 142361
rect 55465 142303 55515 142327
rect 55801 142361 55851 142385
rect 55801 142327 55809 142361
rect 55843 142327 55851 142361
rect 55801 142303 55851 142327
rect 56137 142361 56187 142385
rect 56137 142327 56145 142361
rect 56179 142327 56187 142361
rect 56137 142303 56187 142327
rect 56473 142361 56523 142385
rect 56473 142327 56481 142361
rect 56515 142327 56523 142361
rect 56473 142303 56523 142327
rect 56809 142361 56859 142385
rect 56809 142327 56817 142361
rect 56851 142327 56859 142361
rect 56809 142303 56859 142327
rect 57145 142361 57195 142385
rect 57145 142327 57153 142361
rect 57187 142327 57195 142361
rect 57145 142303 57195 142327
rect 57481 142361 57531 142385
rect 57481 142327 57489 142361
rect 57523 142327 57531 142361
rect 57481 142303 57531 142327
rect 57817 142361 57867 142385
rect 57817 142327 57825 142361
rect 57859 142327 57867 142361
rect 57817 142303 57867 142327
rect 58153 142361 58203 142385
rect 58153 142327 58161 142361
rect 58195 142327 58203 142361
rect 58153 142303 58203 142327
rect 58489 142361 58539 142385
rect 58489 142327 58497 142361
rect 58531 142327 58539 142361
rect 58489 142303 58539 142327
rect 58825 142361 58875 142385
rect 58825 142327 58833 142361
rect 58867 142327 58875 142361
rect 58825 142303 58875 142327
rect 59161 142361 59211 142385
rect 59161 142327 59169 142361
rect 59203 142327 59211 142361
rect 59161 142303 59211 142327
rect 59497 142361 59547 142385
rect 59497 142327 59505 142361
rect 59539 142327 59547 142361
rect 59497 142303 59547 142327
rect 59833 142361 59883 142385
rect 59833 142327 59841 142361
rect 59875 142327 59883 142361
rect 59833 142303 59883 142327
rect 60169 142361 60219 142385
rect 60169 142327 60177 142361
rect 60211 142327 60219 142361
rect 60169 142303 60219 142327
rect 60505 142361 60555 142385
rect 60505 142327 60513 142361
rect 60547 142327 60555 142361
rect 60505 142303 60555 142327
rect 60841 142361 60891 142385
rect 60841 142327 60849 142361
rect 60883 142327 60891 142361
rect 60841 142303 60891 142327
rect 61177 142361 61227 142385
rect 61177 142327 61185 142361
rect 61219 142327 61227 142361
rect 61177 142303 61227 142327
rect 61513 142361 61563 142385
rect 61513 142327 61521 142361
rect 61555 142327 61563 142361
rect 61513 142303 61563 142327
rect 61849 142361 61899 142385
rect 61849 142327 61857 142361
rect 61891 142327 61899 142361
rect 61849 142303 61899 142327
rect 62185 142361 62235 142385
rect 62185 142327 62193 142361
rect 62227 142327 62235 142361
rect 62185 142303 62235 142327
rect 62521 142361 62571 142385
rect 62521 142327 62529 142361
rect 62563 142327 62571 142361
rect 62521 142303 62571 142327
rect 62857 142361 62907 142385
rect 62857 142327 62865 142361
rect 62899 142327 62907 142361
rect 62857 142303 62907 142327
rect 63193 142361 63243 142385
rect 63193 142327 63201 142361
rect 63235 142327 63243 142361
rect 63193 142303 63243 142327
rect 63529 142361 63579 142385
rect 63529 142327 63537 142361
rect 63571 142327 63579 142361
rect 63529 142303 63579 142327
rect 63865 142361 63915 142385
rect 63865 142327 63873 142361
rect 63907 142327 63915 142361
rect 63865 142303 63915 142327
rect 64201 142361 64251 142385
rect 64201 142327 64209 142361
rect 64243 142327 64251 142361
rect 64201 142303 64251 142327
rect 64537 142361 64587 142385
rect 64537 142327 64545 142361
rect 64579 142327 64587 142361
rect 64537 142303 64587 142327
rect 64873 142361 64923 142385
rect 64873 142327 64881 142361
rect 64915 142327 64923 142361
rect 64873 142303 64923 142327
rect 65209 142361 65259 142385
rect 65209 142327 65217 142361
rect 65251 142327 65259 142361
rect 65209 142303 65259 142327
rect 65545 142361 65595 142385
rect 65545 142327 65553 142361
rect 65587 142327 65595 142361
rect 65545 142303 65595 142327
rect 65881 142361 65931 142385
rect 65881 142327 65889 142361
rect 65923 142327 65931 142361
rect 65881 142303 65931 142327
rect 66217 142361 66267 142385
rect 66217 142327 66225 142361
rect 66259 142327 66267 142361
rect 66217 142303 66267 142327
rect 66553 142361 66603 142385
rect 66553 142327 66561 142361
rect 66595 142327 66603 142361
rect 66553 142303 66603 142327
rect 66889 142361 66939 142385
rect 66889 142327 66897 142361
rect 66931 142327 66939 142361
rect 66889 142303 66939 142327
rect 67225 142361 67275 142385
rect 67225 142327 67233 142361
rect 67267 142327 67275 142361
rect 67225 142303 67275 142327
rect 67561 142361 67611 142385
rect 67561 142327 67569 142361
rect 67603 142327 67611 142361
rect 67561 142303 67611 142327
rect 67897 142361 67947 142385
rect 67897 142327 67905 142361
rect 67939 142327 67947 142361
rect 67897 142303 67947 142327
rect 68233 142361 68283 142385
rect 68233 142327 68241 142361
rect 68275 142327 68283 142361
rect 68233 142303 68283 142327
rect 68569 142361 68619 142385
rect 68569 142327 68577 142361
rect 68611 142327 68619 142361
rect 68569 142303 68619 142327
rect 68905 142361 68955 142385
rect 68905 142327 68913 142361
rect 68947 142327 68955 142361
rect 68905 142303 68955 142327
rect 69241 142361 69291 142385
rect 69241 142327 69249 142361
rect 69283 142327 69291 142361
rect 69241 142303 69291 142327
rect 69577 142361 69627 142385
rect 69577 142327 69585 142361
rect 69619 142327 69627 142361
rect 69577 142303 69627 142327
rect 69913 142361 69963 142385
rect 69913 142327 69921 142361
rect 69955 142327 69963 142361
rect 69913 142303 69963 142327
rect 70249 142361 70299 142385
rect 70249 142327 70257 142361
rect 70291 142327 70299 142361
rect 70249 142303 70299 142327
rect 70585 142361 70635 142385
rect 70585 142327 70593 142361
rect 70627 142327 70635 142361
rect 70585 142303 70635 142327
rect 70921 142361 70971 142385
rect 70921 142327 70929 142361
rect 70963 142327 70971 142361
rect 70921 142303 70971 142327
rect 71257 142361 71307 142385
rect 71257 142327 71265 142361
rect 71299 142327 71307 142361
rect 71257 142303 71307 142327
rect 71593 142361 71643 142385
rect 71593 142327 71601 142361
rect 71635 142327 71643 142361
rect 71593 142303 71643 142327
rect 71929 142361 71979 142385
rect 71929 142327 71937 142361
rect 71971 142327 71979 142361
rect 71929 142303 71979 142327
rect 72265 142361 72315 142385
rect 72265 142327 72273 142361
rect 72307 142327 72315 142361
rect 72265 142303 72315 142327
rect 72601 142361 72651 142385
rect 72601 142327 72609 142361
rect 72643 142327 72651 142361
rect 72601 142303 72651 142327
rect 72937 142361 72987 142385
rect 72937 142327 72945 142361
rect 72979 142327 72987 142361
rect 72937 142303 72987 142327
rect 73273 142361 73323 142385
rect 73273 142327 73281 142361
rect 73315 142327 73323 142361
rect 73273 142303 73323 142327
rect 73609 142361 73659 142385
rect 73609 142327 73617 142361
rect 73651 142327 73659 142361
rect 73609 142303 73659 142327
rect 73945 142361 73995 142385
rect 73945 142327 73953 142361
rect 73987 142327 73995 142361
rect 73945 142303 73995 142327
rect 74281 142361 74331 142385
rect 74281 142327 74289 142361
rect 74323 142327 74331 142361
rect 74281 142303 74331 142327
rect 74617 142361 74667 142385
rect 74617 142327 74625 142361
rect 74659 142327 74667 142361
rect 74617 142303 74667 142327
rect 74953 142361 75003 142385
rect 74953 142327 74961 142361
rect 74995 142327 75003 142361
rect 74953 142303 75003 142327
rect 75289 142361 75339 142385
rect 75289 142327 75297 142361
rect 75331 142327 75339 142361
rect 75289 142303 75339 142327
rect 75625 142361 75675 142385
rect 75625 142327 75633 142361
rect 75667 142327 75675 142361
rect 75625 142303 75675 142327
rect 75961 142361 76011 142385
rect 75961 142327 75969 142361
rect 76003 142327 76011 142361
rect 75961 142303 76011 142327
rect 76297 142361 76347 142385
rect 76297 142327 76305 142361
rect 76339 142327 76347 142361
rect 76297 142303 76347 142327
rect 76633 142361 76683 142385
rect 76633 142327 76641 142361
rect 76675 142327 76683 142361
rect 76633 142303 76683 142327
rect 76969 142361 77019 142385
rect 76969 142327 76977 142361
rect 77011 142327 77019 142361
rect 76969 142303 77019 142327
rect 77305 142361 77355 142385
rect 77305 142327 77313 142361
rect 77347 142327 77355 142361
rect 77305 142303 77355 142327
rect 77641 142361 77691 142385
rect 77641 142327 77649 142361
rect 77683 142327 77691 142361
rect 77641 142303 77691 142327
rect 77977 142361 78027 142385
rect 77977 142327 77985 142361
rect 78019 142327 78027 142361
rect 77977 142303 78027 142327
rect 78313 142361 78363 142385
rect 78313 142327 78321 142361
rect 78355 142327 78363 142361
rect 78313 142303 78363 142327
rect 78649 142361 78699 142385
rect 78649 142327 78657 142361
rect 78691 142327 78699 142361
rect 78649 142303 78699 142327
rect 78985 142361 79035 142385
rect 78985 142327 78993 142361
rect 79027 142327 79035 142361
rect 78985 142303 79035 142327
rect 79321 142361 79371 142385
rect 79321 142327 79329 142361
rect 79363 142327 79371 142361
rect 79321 142303 79371 142327
rect 79657 142361 79707 142385
rect 79657 142327 79665 142361
rect 79699 142327 79707 142361
rect 79657 142303 79707 142327
rect 79993 142361 80043 142385
rect 79993 142327 80001 142361
rect 80035 142327 80043 142361
rect 79993 142303 80043 142327
rect 80329 142361 80379 142385
rect 80329 142327 80337 142361
rect 80371 142327 80379 142361
rect 80329 142303 80379 142327
rect 80665 142361 80715 142385
rect 80665 142327 80673 142361
rect 80707 142327 80715 142361
rect 80665 142303 80715 142327
rect 81001 142361 81051 142385
rect 81001 142327 81009 142361
rect 81043 142327 81051 142361
rect 81001 142303 81051 142327
rect 81337 142361 81387 142385
rect 81337 142327 81345 142361
rect 81379 142327 81387 142361
rect 81337 142303 81387 142327
rect 81673 142361 81723 142385
rect 81673 142327 81681 142361
rect 81715 142327 81723 142361
rect 81673 142303 81723 142327
rect 82009 142361 82059 142385
rect 82009 142327 82017 142361
rect 82051 142327 82059 142361
rect 82009 142303 82059 142327
rect 82345 142361 82395 142385
rect 82345 142327 82353 142361
rect 82387 142327 82395 142361
rect 82345 142303 82395 142327
rect 82681 142361 82731 142385
rect 82681 142327 82689 142361
rect 82723 142327 82731 142361
rect 82681 142303 82731 142327
rect 83017 142361 83067 142385
rect 83017 142327 83025 142361
rect 83059 142327 83067 142361
rect 83017 142303 83067 142327
rect 83353 142361 83403 142385
rect 83353 142327 83361 142361
rect 83395 142327 83403 142361
rect 83353 142303 83403 142327
rect 83689 142361 83739 142385
rect 83689 142327 83697 142361
rect 83731 142327 83739 142361
rect 83689 142303 83739 142327
rect 84025 142361 84075 142385
rect 84025 142327 84033 142361
rect 84067 142327 84075 142361
rect 84025 142303 84075 142327
rect 84361 142361 84411 142385
rect 84361 142327 84369 142361
rect 84403 142327 84411 142361
rect 84361 142303 84411 142327
rect 84697 142361 84747 142385
rect 84697 142327 84705 142361
rect 84739 142327 84747 142361
rect 84697 142303 84747 142327
rect 85033 142361 85083 142385
rect 85033 142327 85041 142361
rect 85075 142327 85083 142361
rect 85033 142303 85083 142327
rect 85369 142361 85419 142385
rect 85369 142327 85377 142361
rect 85411 142327 85419 142361
rect 85369 142303 85419 142327
rect 85705 142361 85755 142385
rect 85705 142327 85713 142361
rect 85747 142327 85755 142361
rect 85705 142303 85755 142327
rect 86041 142361 86091 142385
rect 86041 142327 86049 142361
rect 86083 142327 86091 142361
rect 86041 142303 86091 142327
rect 86377 142361 86427 142385
rect 86377 142327 86385 142361
rect 86419 142327 86427 142361
rect 86377 142303 86427 142327
rect 86713 142361 86763 142385
rect 86713 142327 86721 142361
rect 86755 142327 86763 142361
rect 86713 142303 86763 142327
rect 87049 142361 87099 142385
rect 87049 142327 87057 142361
rect 87091 142327 87099 142361
rect 87049 142303 87099 142327
rect 87385 142361 87435 142385
rect 87385 142327 87393 142361
rect 87427 142327 87435 142361
rect 87385 142303 87435 142327
rect 87721 142361 87771 142385
rect 87721 142327 87729 142361
rect 87763 142327 87771 142361
rect 87721 142303 87771 142327
rect 88057 142361 88107 142385
rect 88057 142327 88065 142361
rect 88099 142327 88107 142361
rect 88057 142303 88107 142327
rect 88393 142361 88443 142385
rect 88393 142327 88401 142361
rect 88435 142327 88443 142361
rect 88393 142303 88443 142327
rect 88729 142361 88779 142385
rect 88729 142327 88737 142361
rect 88771 142327 88779 142361
rect 88729 142303 88779 142327
rect 89065 142361 89115 142385
rect 89065 142327 89073 142361
rect 89107 142327 89115 142361
rect 89065 142303 89115 142327
rect 89401 142361 89451 142385
rect 89401 142327 89409 142361
rect 89443 142327 89451 142361
rect 89401 142303 89451 142327
rect 89737 142361 89787 142385
rect 89737 142327 89745 142361
rect 89779 142327 89787 142361
rect 89737 142303 89787 142327
rect 90073 142361 90123 142385
rect 90073 142327 90081 142361
rect 90115 142327 90123 142361
rect 90073 142303 90123 142327
rect 90409 142361 90459 142385
rect 90409 142327 90417 142361
rect 90451 142327 90459 142361
rect 90409 142303 90459 142327
rect 90745 142361 90795 142385
rect 90745 142327 90753 142361
rect 90787 142327 90795 142361
rect 90745 142303 90795 142327
rect 91081 142361 91131 142385
rect 91081 142327 91089 142361
rect 91123 142327 91131 142361
rect 91081 142303 91131 142327
rect 91417 142361 91467 142385
rect 91417 142327 91425 142361
rect 91459 142327 91467 142361
rect 91417 142303 91467 142327
rect 91753 142361 91803 142385
rect 91753 142327 91761 142361
rect 91795 142327 91803 142361
rect 91753 142303 91803 142327
rect 92089 142361 92139 142385
rect 92089 142327 92097 142361
rect 92131 142327 92139 142361
rect 92089 142303 92139 142327
rect 92425 142361 92475 142385
rect 92425 142327 92433 142361
rect 92467 142327 92475 142361
rect 92425 142303 92475 142327
rect 92761 142361 92811 142385
rect 92761 142327 92769 142361
rect 92803 142327 92811 142361
rect 92761 142303 92811 142327
rect 93097 142361 93147 142385
rect 93097 142327 93105 142361
rect 93139 142327 93147 142361
rect 93097 142303 93147 142327
rect 93433 142361 93483 142385
rect 93433 142327 93441 142361
rect 93475 142327 93483 142361
rect 93433 142303 93483 142327
rect 93769 142361 93819 142385
rect 93769 142327 93777 142361
rect 93811 142327 93819 142361
rect 93769 142303 93819 142327
rect 94105 142361 94155 142385
rect 94105 142327 94113 142361
rect 94147 142327 94155 142361
rect 94105 142303 94155 142327
rect 94441 142361 94491 142385
rect 94441 142327 94449 142361
rect 94483 142327 94491 142361
rect 94441 142303 94491 142327
rect 94777 142361 94827 142385
rect 94777 142327 94785 142361
rect 94819 142327 94827 142361
rect 94777 142303 94827 142327
rect 95113 142361 95163 142385
rect 95113 142327 95121 142361
rect 95155 142327 95163 142361
rect 95113 142303 95163 142327
rect 95449 142361 95499 142385
rect 95449 142327 95457 142361
rect 95491 142327 95499 142361
rect 95449 142303 95499 142327
rect 95785 142361 95835 142385
rect 95785 142327 95793 142361
rect 95827 142327 95835 142361
rect 95785 142303 95835 142327
rect 96121 142361 96171 142385
rect 96121 142327 96129 142361
rect 96163 142327 96171 142361
rect 96121 142303 96171 142327
rect 96457 142361 96507 142385
rect 96457 142327 96465 142361
rect 96499 142327 96507 142361
rect 96457 142303 96507 142327
rect 96793 142361 96843 142385
rect 96793 142327 96801 142361
rect 96835 142327 96843 142361
rect 96793 142303 96843 142327
rect 97129 142361 97179 142385
rect 97129 142327 97137 142361
rect 97171 142327 97179 142361
rect 97129 142303 97179 142327
rect 97465 142361 97515 142385
rect 97465 142327 97473 142361
rect 97507 142327 97515 142361
rect 97465 142303 97515 142327
rect 97801 142361 97851 142385
rect 97801 142327 97809 142361
rect 97843 142327 97851 142361
rect 97801 142303 97851 142327
rect 98137 142361 98187 142385
rect 98137 142327 98145 142361
rect 98179 142327 98187 142361
rect 98137 142303 98187 142327
rect 98473 142361 98523 142385
rect 98473 142327 98481 142361
rect 98515 142327 98523 142361
rect 98473 142303 98523 142327
rect 98809 142361 98859 142385
rect 98809 142327 98817 142361
rect 98851 142327 98859 142361
rect 98809 142303 98859 142327
rect 99145 142361 99195 142385
rect 99145 142327 99153 142361
rect 99187 142327 99195 142361
rect 99145 142303 99195 142327
rect 99481 142361 99531 142385
rect 99481 142327 99489 142361
rect 99523 142327 99531 142361
rect 99481 142303 99531 142327
rect 99817 142361 99867 142385
rect 99817 142327 99825 142361
rect 99859 142327 99867 142361
rect 99817 142303 99867 142327
rect 100153 142361 100203 142385
rect 100153 142327 100161 142361
rect 100195 142327 100203 142361
rect 100153 142303 100203 142327
rect 100489 142361 100539 142385
rect 100489 142327 100497 142361
rect 100531 142327 100539 142361
rect 100489 142303 100539 142327
rect 100825 142361 100875 142385
rect 100825 142327 100833 142361
rect 100867 142327 100875 142361
rect 100825 142303 100875 142327
rect 101161 142361 101211 142385
rect 101161 142327 101169 142361
rect 101203 142327 101211 142361
rect 101161 142303 101211 142327
rect 101497 142361 101547 142385
rect 101497 142327 101505 142361
rect 101539 142327 101547 142361
rect 101497 142303 101547 142327
rect 101833 142361 101883 142385
rect 101833 142327 101841 142361
rect 101875 142327 101883 142361
rect 101833 142303 101883 142327
rect 102169 142361 102219 142385
rect 102169 142327 102177 142361
rect 102211 142327 102219 142361
rect 102169 142303 102219 142327
rect 102505 142361 102555 142385
rect 102505 142327 102513 142361
rect 102547 142327 102555 142361
rect 102505 142303 102555 142327
rect 102841 142361 102891 142385
rect 102841 142327 102849 142361
rect 102883 142327 102891 142361
rect 102841 142303 102891 142327
rect 103177 142361 103227 142385
rect 103177 142327 103185 142361
rect 103219 142327 103227 142361
rect 103177 142303 103227 142327
rect 103513 142361 103563 142385
rect 103513 142327 103521 142361
rect 103555 142327 103563 142361
rect 103513 142303 103563 142327
rect 103849 142361 103899 142385
rect 103849 142327 103857 142361
rect 103891 142327 103899 142361
rect 103849 142303 103899 142327
rect 104185 142361 104235 142385
rect 104185 142327 104193 142361
rect 104227 142327 104235 142361
rect 104185 142303 104235 142327
rect 104521 142361 104571 142385
rect 104521 142327 104529 142361
rect 104563 142327 104571 142361
rect 104521 142303 104571 142327
rect 104857 142361 104907 142385
rect 104857 142327 104865 142361
rect 104899 142327 104907 142361
rect 104857 142303 104907 142327
rect 105193 142361 105243 142385
rect 105193 142327 105201 142361
rect 105235 142327 105243 142361
rect 105193 142303 105243 142327
rect 105529 142361 105579 142385
rect 105529 142327 105537 142361
rect 105571 142327 105579 142361
rect 105529 142303 105579 142327
rect 105865 142361 105915 142385
rect 105865 142327 105873 142361
rect 105907 142327 105915 142361
rect 105865 142303 105915 142327
rect 106201 142361 106251 142385
rect 106201 142327 106209 142361
rect 106243 142327 106251 142361
rect 106201 142303 106251 142327
rect 106537 142361 106587 142385
rect 106537 142327 106545 142361
rect 106579 142327 106587 142361
rect 106537 142303 106587 142327
rect 106873 142361 106923 142385
rect 106873 142327 106881 142361
rect 106915 142327 106923 142361
rect 106873 142303 106923 142327
rect 107209 142361 107259 142385
rect 107209 142327 107217 142361
rect 107251 142327 107259 142361
rect 107209 142303 107259 142327
rect 107545 142361 107595 142385
rect 107545 142327 107553 142361
rect 107587 142327 107595 142361
rect 107545 142303 107595 142327
rect 107881 142361 107931 142385
rect 107881 142327 107889 142361
rect 107923 142327 107931 142361
rect 107881 142303 107931 142327
rect 108217 142361 108267 142385
rect 108217 142327 108225 142361
rect 108259 142327 108267 142361
rect 108217 142303 108267 142327
rect 108553 142361 108603 142385
rect 108553 142327 108561 142361
rect 108595 142327 108603 142361
rect 108553 142303 108603 142327
rect 108889 142361 108939 142385
rect 108889 142327 108897 142361
rect 108931 142327 108939 142361
rect 108889 142303 108939 142327
rect 109225 142361 109275 142385
rect 109225 142327 109233 142361
rect 109267 142327 109275 142361
rect 109225 142303 109275 142327
rect 109561 142361 109611 142385
rect 109561 142327 109569 142361
rect 109603 142327 109611 142361
rect 109561 142303 109611 142327
rect 109897 142361 109947 142385
rect 109897 142327 109905 142361
rect 109939 142327 109947 142361
rect 109897 142303 109947 142327
rect 110233 142361 110283 142385
rect 110233 142327 110241 142361
rect 110275 142327 110283 142361
rect 110233 142303 110283 142327
rect 110569 142361 110619 142385
rect 110569 142327 110577 142361
rect 110611 142327 110619 142361
rect 110569 142303 110619 142327
rect 110905 142361 110955 142385
rect 110905 142327 110913 142361
rect 110947 142327 110955 142361
rect 110905 142303 110955 142327
rect 111241 142361 111291 142385
rect 111241 142327 111249 142361
rect 111283 142327 111291 142361
rect 111241 142303 111291 142327
rect 111577 142361 111627 142385
rect 111577 142327 111585 142361
rect 111619 142327 111627 142361
rect 111577 142303 111627 142327
rect 111913 142361 111963 142385
rect 111913 142327 111921 142361
rect 111955 142327 111963 142361
rect 111913 142303 111963 142327
rect 112249 142361 112299 142385
rect 112249 142327 112257 142361
rect 112291 142327 112299 142361
rect 112249 142303 112299 142327
rect 112585 142361 112635 142385
rect 112585 142327 112593 142361
rect 112627 142327 112635 142361
rect 112585 142303 112635 142327
rect 112921 142361 112971 142385
rect 112921 142327 112929 142361
rect 112963 142327 112971 142361
rect 112921 142303 112971 142327
rect 113257 142361 113307 142385
rect 113257 142327 113265 142361
rect 113299 142327 113307 142361
rect 113257 142303 113307 142327
rect 113593 142361 113643 142385
rect 113593 142327 113601 142361
rect 113635 142327 113643 142361
rect 113593 142303 113643 142327
rect 113929 142361 113979 142385
rect 113929 142327 113937 142361
rect 113971 142327 113979 142361
rect 113929 142303 113979 142327
rect 114265 142361 114315 142385
rect 114265 142327 114273 142361
rect 114307 142327 114315 142361
rect 114265 142303 114315 142327
rect 114601 142361 114651 142385
rect 114601 142327 114609 142361
rect 114643 142327 114651 142361
rect 114601 142303 114651 142327
rect 114937 142361 114987 142385
rect 114937 142327 114945 142361
rect 114979 142327 114987 142361
rect 114937 142303 114987 142327
rect 115273 142361 115323 142385
rect 115273 142327 115281 142361
rect 115315 142327 115323 142361
rect 115273 142303 115323 142327
rect 115609 142361 115659 142385
rect 115609 142327 115617 142361
rect 115651 142327 115659 142361
rect 115609 142303 115659 142327
rect 115945 142361 115995 142385
rect 115945 142327 115953 142361
rect 115987 142327 115995 142361
rect 115945 142303 115995 142327
rect 116281 142361 116331 142385
rect 116281 142327 116289 142361
rect 116323 142327 116331 142361
rect 116281 142303 116331 142327
rect 116617 142361 116667 142385
rect 116617 142327 116625 142361
rect 116659 142327 116667 142361
rect 116617 142303 116667 142327
rect 116953 142361 117003 142385
rect 116953 142327 116961 142361
rect 116995 142327 117003 142361
rect 116953 142303 117003 142327
rect 117289 142361 117339 142385
rect 117289 142327 117297 142361
rect 117331 142327 117339 142361
rect 117289 142303 117339 142327
rect 117625 142361 117675 142385
rect 117625 142327 117633 142361
rect 117667 142327 117675 142361
rect 117625 142303 117675 142327
rect 117961 142361 118011 142385
rect 117961 142327 117969 142361
rect 118003 142327 118011 142361
rect 117961 142303 118011 142327
rect 118297 142361 118347 142385
rect 118297 142327 118305 142361
rect 118339 142327 118347 142361
rect 118297 142303 118347 142327
rect 118633 142361 118683 142385
rect 118633 142327 118641 142361
rect 118675 142327 118683 142361
rect 118633 142303 118683 142327
rect 118969 142361 119019 142385
rect 118969 142327 118977 142361
rect 119011 142327 119019 142361
rect 118969 142303 119019 142327
rect 119305 142361 119355 142385
rect 119305 142327 119313 142361
rect 119347 142327 119355 142361
rect 119305 142303 119355 142327
rect 119641 142361 119691 142385
rect 119641 142327 119649 142361
rect 119683 142327 119691 142361
rect 119641 142303 119691 142327
rect 119977 142361 120027 142385
rect 119977 142327 119985 142361
rect 120019 142327 120027 142361
rect 119977 142303 120027 142327
rect 120313 142361 120363 142385
rect 120313 142327 120321 142361
rect 120355 142327 120363 142361
rect 120313 142303 120363 142327
rect 120649 142361 120699 142385
rect 120649 142327 120657 142361
rect 120691 142327 120699 142361
rect 120649 142303 120699 142327
rect 120985 142361 121035 142385
rect 120985 142327 120993 142361
rect 121027 142327 121035 142361
rect 120985 142303 121035 142327
rect 121321 142361 121371 142385
rect 121321 142327 121329 142361
rect 121363 142327 121371 142361
rect 121321 142303 121371 142327
rect 121657 142361 121707 142385
rect 121657 142327 121665 142361
rect 121699 142327 121707 142361
rect 121657 142303 121707 142327
rect 121993 142361 122043 142385
rect 121993 142327 122001 142361
rect 122035 142327 122043 142361
rect 121993 142303 122043 142327
rect 122329 142361 122379 142385
rect 122329 142327 122337 142361
rect 122371 142327 122379 142361
rect 122329 142303 122379 142327
rect 122665 142361 122715 142385
rect 122665 142327 122673 142361
rect 122707 142327 122715 142361
rect 122665 142303 122715 142327
rect 123001 142361 123051 142385
rect 123001 142327 123009 142361
rect 123043 142327 123051 142361
rect 123001 142303 123051 142327
rect 123337 142361 123387 142385
rect 123337 142327 123345 142361
rect 123379 142327 123387 142361
rect 123337 142303 123387 142327
rect 123673 142361 123723 142385
rect 123673 142327 123681 142361
rect 123715 142327 123723 142361
rect 123673 142303 123723 142327
rect 124009 142361 124059 142385
rect 124009 142327 124017 142361
rect 124051 142327 124059 142361
rect 124009 142303 124059 142327
rect 124345 142361 124395 142385
rect 124345 142327 124353 142361
rect 124387 142327 124395 142361
rect 124345 142303 124395 142327
rect 124681 142361 124731 142385
rect 124681 142327 124689 142361
rect 124723 142327 124731 142361
rect 124681 142303 124731 142327
rect 125017 142361 125067 142385
rect 125017 142327 125025 142361
rect 125059 142327 125067 142361
rect 125017 142303 125067 142327
rect 125353 142361 125403 142385
rect 125353 142327 125361 142361
rect 125395 142327 125403 142361
rect 125353 142303 125403 142327
rect 125689 142361 125739 142385
rect 125689 142327 125697 142361
rect 125731 142327 125739 142361
rect 125689 142303 125739 142327
rect 126025 142361 126075 142385
rect 126025 142327 126033 142361
rect 126067 142327 126075 142361
rect 126025 142303 126075 142327
rect 126361 142361 126411 142385
rect 126361 142327 126369 142361
rect 126403 142327 126411 142361
rect 126361 142303 126411 142327
rect 126697 142361 126747 142385
rect 126697 142327 126705 142361
rect 126739 142327 126747 142361
rect 126697 142303 126747 142327
rect 127033 142361 127083 142385
rect 127033 142327 127041 142361
rect 127075 142327 127083 142361
rect 127033 142303 127083 142327
rect 127369 142361 127419 142385
rect 127369 142327 127377 142361
rect 127411 142327 127419 142361
rect 127369 142303 127419 142327
rect 127705 142361 127755 142385
rect 127705 142327 127713 142361
rect 127747 142327 127755 142361
rect 127705 142303 127755 142327
rect 128041 142361 128091 142385
rect 128041 142327 128049 142361
rect 128083 142327 128091 142361
rect 128041 142303 128091 142327
rect 128377 142361 128427 142385
rect 128377 142327 128385 142361
rect 128419 142327 128427 142361
rect 128377 142303 128427 142327
rect 128713 142361 128763 142385
rect 128713 142327 128721 142361
rect 128755 142327 128763 142361
rect 128713 142303 128763 142327
rect 129049 142361 129099 142385
rect 129049 142327 129057 142361
rect 129091 142327 129099 142361
rect 129049 142303 129099 142327
rect 129385 142361 129435 142385
rect 129385 142327 129393 142361
rect 129427 142327 129435 142361
rect 129385 142303 129435 142327
rect 129721 142361 129771 142385
rect 129721 142327 129729 142361
rect 129763 142327 129771 142361
rect 129721 142303 129771 142327
rect 130057 142361 130107 142385
rect 130057 142327 130065 142361
rect 130099 142327 130107 142361
rect 130057 142303 130107 142327
rect 130393 142361 130443 142385
rect 130393 142327 130401 142361
rect 130435 142327 130443 142361
rect 130393 142303 130443 142327
rect 130729 142361 130779 142385
rect 130729 142327 130737 142361
rect 130771 142327 130779 142361
rect 130729 142303 130779 142327
rect 131065 142361 131115 142385
rect 131065 142327 131073 142361
rect 131107 142327 131115 142361
rect 131065 142303 131115 142327
rect 131401 142361 131451 142385
rect 131401 142327 131409 142361
rect 131443 142327 131451 142361
rect 131401 142303 131451 142327
rect 131737 142361 131787 142385
rect 131737 142327 131745 142361
rect 131779 142327 131787 142361
rect 131737 142303 131787 142327
rect 132073 142361 132123 142385
rect 132073 142327 132081 142361
rect 132115 142327 132123 142361
rect 132073 142303 132123 142327
rect 132409 142361 132459 142385
rect 132409 142327 132417 142361
rect 132451 142327 132459 142361
rect 132409 142303 132459 142327
rect 132745 142361 132795 142385
rect 132745 142327 132753 142361
rect 132787 142327 132795 142361
rect 132745 142303 132795 142327
rect 133081 142361 133131 142385
rect 133081 142327 133089 142361
rect 133123 142327 133131 142361
rect 133081 142303 133131 142327
rect 133417 142361 133467 142385
rect 133417 142327 133425 142361
rect 133459 142327 133467 142361
rect 133417 142303 133467 142327
rect 133753 142361 133803 142385
rect 133753 142327 133761 142361
rect 133795 142327 133803 142361
rect 133753 142303 133803 142327
rect 134089 142361 134139 142385
rect 134089 142327 134097 142361
rect 134131 142327 134139 142361
rect 134089 142303 134139 142327
rect 134425 142361 134475 142385
rect 134425 142327 134433 142361
rect 134467 142327 134475 142361
rect 134425 142303 134475 142327
rect 134761 142361 134811 142385
rect 134761 142327 134769 142361
rect 134803 142327 134811 142361
rect 134761 142303 134811 142327
rect 135097 142361 135147 142385
rect 135097 142327 135105 142361
rect 135139 142327 135147 142361
rect 135097 142303 135147 142327
rect 135433 142361 135483 142385
rect 135433 142327 135441 142361
rect 135475 142327 135483 142361
rect 135433 142303 135483 142327
rect 135769 142361 135819 142385
rect 135769 142327 135777 142361
rect 135811 142327 135819 142361
rect 135769 142303 135819 142327
rect 136105 142361 136155 142385
rect 136105 142327 136113 142361
rect 136147 142327 136155 142361
rect 136105 142303 136155 142327
rect 136441 142361 136491 142385
rect 136441 142327 136449 142361
rect 136483 142327 136491 142361
rect 136441 142303 136491 142327
rect 136777 142361 136827 142385
rect 136777 142327 136785 142361
rect 136819 142327 136827 142361
rect 136777 142303 136827 142327
rect 137113 142361 137163 142385
rect 137113 142327 137121 142361
rect 137155 142327 137163 142361
rect 137113 142303 137163 142327
rect 137449 142361 137499 142385
rect 137449 142327 137457 142361
rect 137491 142327 137499 142361
rect 137449 142303 137499 142327
rect 137785 142361 137835 142385
rect 137785 142327 137793 142361
rect 137827 142327 137835 142361
rect 137785 142303 137835 142327
rect 138121 142361 138171 142385
rect 138121 142327 138129 142361
rect 138163 142327 138171 142361
rect 138121 142303 138171 142327
rect 138457 142361 138507 142385
rect 138457 142327 138465 142361
rect 138499 142327 138507 142361
rect 138457 142303 138507 142327
rect 138793 142361 138843 142385
rect 138793 142327 138801 142361
rect 138835 142327 138843 142361
rect 138793 142303 138843 142327
rect 139129 142361 139179 142385
rect 139129 142327 139137 142361
rect 139171 142327 139179 142361
rect 139129 142303 139179 142327
rect 139465 142361 139515 142385
rect 139465 142327 139473 142361
rect 139507 142327 139515 142361
rect 139465 142303 139515 142327
rect 139801 142361 139851 142385
rect 139801 142327 139809 142361
rect 139843 142327 139851 142361
rect 139801 142303 139851 142327
rect 140137 142361 140187 142385
rect 140137 142327 140145 142361
rect 140179 142327 140187 142361
rect 140137 142303 140187 142327
rect 140473 142361 140523 142385
rect 140473 142327 140481 142361
rect 140515 142327 140523 142361
rect 140473 142303 140523 142327
rect 140809 142361 140859 142385
rect 140809 142327 140817 142361
rect 140851 142327 140859 142361
rect 140809 142303 140859 142327
rect 141145 142361 141195 142385
rect 141145 142327 141153 142361
rect 141187 142327 141195 142361
rect 141145 142303 141195 142327
rect 141481 142361 141531 142385
rect 141481 142327 141489 142361
rect 141523 142327 141531 142361
rect 141481 142303 141531 142327
rect 141817 142361 141867 142385
rect 141817 142327 141825 142361
rect 141859 142327 141867 142361
rect 141817 142303 141867 142327
rect 142153 142361 142203 142385
rect 142153 142327 142161 142361
rect 142195 142327 142203 142361
rect 142153 142303 142203 142327
rect 142489 142361 142539 142385
rect 142489 142327 142497 142361
rect 142531 142327 142539 142361
rect 142489 142303 142539 142327
rect 142825 142361 142875 142385
rect 142825 142327 142833 142361
rect 142867 142327 142875 142361
rect 142825 142303 142875 142327
rect 143161 142361 143211 142385
rect 143161 142327 143169 142361
rect 143203 142327 143211 142361
rect 143161 142303 143211 142327
rect 143497 142361 143547 142385
rect 143497 142327 143505 142361
rect 143539 142327 143547 142361
rect 143497 142303 143547 142327
rect 143833 142361 143883 142385
rect 143833 142327 143841 142361
rect 143875 142327 143883 142361
rect 143833 142303 143883 142327
rect 144169 142361 144219 142385
rect 144169 142327 144177 142361
rect 144211 142327 144219 142361
rect 144169 142303 144219 142327
rect 144505 142361 144555 142385
rect 144505 142327 144513 142361
rect 144547 142327 144555 142361
rect 144505 142303 144555 142327
rect 144841 142361 144891 142385
rect 144841 142327 144849 142361
rect 144883 142327 144891 142361
rect 144841 142303 144891 142327
rect 145177 142361 145227 142385
rect 145177 142327 145185 142361
rect 145219 142327 145227 142361
rect 145177 142303 145227 142327
rect 145513 142361 145563 142385
rect 145513 142327 145521 142361
rect 145555 142327 145563 142361
rect 145513 142303 145563 142327
rect 145849 142361 145899 142385
rect 145849 142327 145857 142361
rect 145891 142327 145899 142361
rect 145849 142303 145899 142327
rect 146185 142361 146235 142385
rect 146185 142327 146193 142361
rect 146227 142327 146235 142361
rect 146185 142303 146235 142327
rect 146521 142361 146571 142385
rect 146521 142327 146529 142361
rect 146563 142327 146571 142361
rect 146521 142303 146571 142327
rect 146857 142361 146907 142385
rect 146857 142327 146865 142361
rect 146899 142327 146907 142361
rect 146857 142303 146907 142327
rect 147193 142361 147243 142385
rect 147193 142327 147201 142361
rect 147235 142327 147243 142361
rect 147193 142303 147243 142327
rect 147529 142361 147579 142385
rect 147529 142327 147537 142361
rect 147571 142327 147579 142361
rect 147529 142303 147579 142327
rect 147865 142361 147915 142385
rect 147865 142327 147873 142361
rect 147907 142327 147915 142361
rect 147865 142303 147915 142327
rect 148201 142361 148251 142385
rect 148201 142327 148209 142361
rect 148243 142327 148251 142361
rect 148201 142303 148251 142327
rect 148537 142361 148587 142385
rect 148537 142327 148545 142361
rect 148579 142327 148587 142361
rect 148537 142303 148587 142327
rect 148873 142361 148923 142385
rect 148873 142327 148881 142361
rect 148915 142327 148923 142361
rect 148873 142303 148923 142327
rect 149209 142361 149259 142385
rect 149209 142327 149217 142361
rect 149251 142327 149259 142361
rect 149209 142303 149259 142327
rect 149545 142361 149595 142385
rect 149545 142327 149553 142361
rect 149587 142327 149595 142361
rect 149545 142303 149595 142327
rect 149881 142361 149931 142385
rect 149881 142327 149889 142361
rect 149923 142327 149931 142361
rect 149881 142303 149931 142327
rect 150217 142361 150267 142385
rect 150217 142327 150225 142361
rect 150259 142327 150267 142361
rect 150217 142303 150267 142327
rect 150553 142361 150603 142385
rect 150553 142327 150561 142361
rect 150595 142327 150603 142361
rect 150553 142303 150603 142327
rect 150889 142361 150939 142385
rect 150889 142327 150897 142361
rect 150931 142327 150939 142361
rect 150889 142303 150939 142327
rect 151225 142361 151275 142385
rect 151225 142327 151233 142361
rect 151267 142327 151275 142361
rect 151225 142303 151275 142327
rect 151561 142361 151611 142385
rect 151561 142327 151569 142361
rect 151603 142327 151611 142361
rect 151561 142303 151611 142327
rect 151897 142361 151947 142385
rect 151897 142327 151905 142361
rect 151939 142327 151947 142361
rect 151897 142303 151947 142327
rect 152233 142361 152283 142385
rect 152233 142327 152241 142361
rect 152275 142327 152283 142361
rect 152233 142303 152283 142327
rect 152569 142361 152619 142385
rect 152569 142327 152577 142361
rect 152611 142327 152619 142361
rect 152569 142303 152619 142327
rect 152905 142361 152955 142385
rect 152905 142327 152913 142361
rect 152947 142327 152955 142361
rect 152905 142303 152955 142327
rect 153241 142361 153291 142385
rect 153241 142327 153249 142361
rect 153283 142327 153291 142361
rect 153241 142303 153291 142327
rect 153577 142361 153627 142385
rect 153577 142327 153585 142361
rect 153619 142327 153627 142361
rect 153577 142303 153627 142327
rect 153913 142361 153963 142385
rect 153913 142327 153921 142361
rect 153955 142327 153963 142361
rect 153913 142303 153963 142327
rect 154249 142361 154299 142385
rect 154249 142327 154257 142361
rect 154291 142327 154299 142361
rect 154249 142303 154299 142327
rect 154585 142361 154635 142385
rect 154585 142327 154593 142361
rect 154627 142327 154635 142361
rect 154585 142303 154635 142327
rect 154921 142361 154971 142385
rect 154921 142327 154929 142361
rect 154963 142327 154971 142361
rect 154921 142303 154971 142327
rect 155257 142361 155307 142385
rect 155257 142327 155265 142361
rect 155299 142327 155307 142361
rect 155257 142303 155307 142327
rect 155593 142361 155643 142385
rect 155593 142327 155601 142361
rect 155635 142327 155643 142361
rect 155593 142303 155643 142327
rect 155929 142361 155979 142385
rect 155929 142327 155937 142361
rect 155971 142327 155979 142361
rect 155929 142303 155979 142327
rect 156265 142361 156315 142385
rect 156265 142327 156273 142361
rect 156307 142327 156315 142361
rect 156265 142303 156315 142327
rect 156601 142361 156651 142385
rect 156601 142327 156609 142361
rect 156643 142327 156651 142361
rect 156601 142303 156651 142327
rect 156937 142361 156987 142385
rect 156937 142327 156945 142361
rect 156979 142327 156987 142361
rect 156937 142303 156987 142327
rect 157273 142361 157323 142385
rect 157273 142327 157281 142361
rect 157315 142327 157323 142361
rect 157273 142303 157323 142327
rect 157609 142361 157659 142385
rect 157609 142327 157617 142361
rect 157651 142327 157659 142361
rect 157609 142303 157659 142327
rect 157945 142361 157995 142385
rect 157945 142327 157953 142361
rect 157987 142327 157995 142361
rect 157945 142303 157995 142327
rect 158281 142361 158331 142385
rect 158281 142327 158289 142361
rect 158323 142327 158331 142361
rect 158281 142303 158331 142327
rect 158617 142361 158667 142385
rect 158617 142327 158625 142361
rect 158659 142327 158667 142361
rect 158617 142303 158667 142327
rect 158953 142361 159003 142385
rect 158953 142327 158961 142361
rect 158995 142327 159003 142361
rect 158953 142303 159003 142327
rect 159289 142361 159339 142385
rect 159289 142327 159297 142361
rect 159331 142327 159339 142361
rect 159289 142303 159339 142327
rect 159625 142361 159675 142385
rect 159625 142327 159633 142361
rect 159667 142327 159675 142361
rect 159625 142303 159675 142327
rect 159961 142361 160011 142385
rect 159961 142327 159969 142361
rect 160003 142327 160011 142361
rect 159961 142303 160011 142327
rect 160297 142361 160347 142385
rect 160297 142327 160305 142361
rect 160339 142327 160347 142361
rect 160297 142303 160347 142327
rect 160633 142361 160683 142385
rect 160633 142327 160641 142361
rect 160675 142327 160683 142361
rect 160633 142303 160683 142327
rect 160969 142361 161019 142385
rect 160969 142327 160977 142361
rect 161011 142327 161019 142361
rect 160969 142303 161019 142327
rect 161305 142361 161355 142385
rect 161305 142327 161313 142361
rect 161347 142327 161355 142361
rect 161305 142303 161355 142327
rect 161641 142361 161691 142385
rect 161641 142327 161649 142361
rect 161683 142327 161691 142361
rect 161641 142303 161691 142327
rect 161977 142361 162027 142385
rect 161977 142327 161985 142361
rect 162019 142327 162027 142361
rect 161977 142303 162027 142327
rect 162313 142361 162363 142385
rect 162313 142327 162321 142361
rect 162355 142327 162363 142361
rect 162313 142303 162363 142327
rect 162649 142361 162699 142385
rect 162649 142327 162657 142361
rect 162691 142327 162699 142361
rect 162649 142303 162699 142327
rect 162985 142361 163035 142385
rect 162985 142327 162993 142361
rect 163027 142327 163035 142361
rect 162985 142303 163035 142327
rect 163321 142361 163371 142385
rect 163321 142327 163329 142361
rect 163363 142327 163371 142361
rect 163321 142303 163371 142327
rect 163657 142361 163707 142385
rect 163657 142327 163665 142361
rect 163699 142327 163707 142361
rect 163657 142303 163707 142327
rect 163993 142361 164043 142385
rect 163993 142327 164001 142361
rect 164035 142327 164043 142361
rect 163993 142303 164043 142327
rect 164329 142361 164379 142385
rect 164329 142327 164337 142361
rect 164371 142327 164379 142361
rect 164329 142303 164379 142327
rect 164665 142361 164715 142385
rect 164665 142327 164673 142361
rect 164707 142327 164715 142361
rect 164665 142303 164715 142327
rect 165001 142361 165051 142385
rect 165001 142327 165009 142361
rect 165043 142327 165051 142361
rect 165001 142303 165051 142327
rect 165337 142361 165387 142385
rect 165337 142327 165345 142361
rect 165379 142327 165387 142361
rect 165337 142303 165387 142327
rect 165673 142361 165723 142385
rect 165673 142327 165681 142361
rect 165715 142327 165723 142361
rect 165673 142303 165723 142327
rect 166009 142361 166059 142385
rect 166009 142327 166017 142361
rect 166051 142327 166059 142361
rect 166009 142303 166059 142327
rect 166345 142361 166395 142385
rect 166345 142327 166353 142361
rect 166387 142327 166395 142361
rect 166345 142303 166395 142327
rect 166681 142361 166731 142385
rect 166681 142327 166689 142361
rect 166723 142327 166731 142361
rect 166681 142303 166731 142327
rect 167017 142361 167067 142385
rect 167017 142327 167025 142361
rect 167059 142327 167067 142361
rect 167017 142303 167067 142327
rect 167353 142361 167403 142385
rect 167353 142327 167361 142361
rect 167395 142327 167403 142361
rect 167353 142303 167403 142327
rect 167689 142361 167739 142385
rect 167689 142327 167697 142361
rect 167731 142327 167739 142361
rect 167689 142303 167739 142327
rect 168025 142361 168075 142385
rect 168025 142327 168033 142361
rect 168067 142327 168075 142361
rect 168025 142303 168075 142327
rect 168361 142361 168411 142385
rect 168361 142327 168369 142361
rect 168403 142327 168411 142361
rect 168361 142303 168411 142327
rect 168697 142361 168747 142385
rect 168697 142327 168705 142361
rect 168739 142327 168747 142361
rect 168697 142303 168747 142327
rect 169033 142361 169083 142385
rect 169033 142327 169041 142361
rect 169075 142327 169083 142361
rect 169033 142303 169083 142327
rect 169369 142361 169419 142385
rect 169369 142327 169377 142361
rect 169411 142327 169419 142361
rect 169369 142303 169419 142327
rect 169705 142361 169755 142385
rect 169705 142327 169713 142361
rect 169747 142327 169755 142361
rect 169705 142303 169755 142327
rect 170041 142361 170091 142385
rect 170041 142327 170049 142361
rect 170083 142327 170091 142361
rect 170041 142303 170091 142327
rect 170377 142361 170427 142385
rect 170377 142327 170385 142361
rect 170419 142327 170427 142361
rect 170377 142303 170427 142327
rect 170713 142361 170763 142385
rect 170713 142327 170721 142361
rect 170755 142327 170763 142361
rect 170713 142303 170763 142327
rect 171049 142361 171099 142385
rect 171049 142327 171057 142361
rect 171091 142327 171099 142361
rect 171049 142303 171099 142327
rect 171385 142361 171435 142385
rect 171385 142327 171393 142361
rect 171427 142327 171435 142361
rect 171385 142303 171435 142327
rect 171721 142361 171771 142385
rect 171721 142327 171729 142361
rect 171763 142327 171771 142361
rect 171721 142303 171771 142327
rect 172057 142361 172107 142385
rect 172057 142327 172065 142361
rect 172099 142327 172107 142361
rect 172057 142303 172107 142327
rect 172393 142361 172443 142385
rect 172393 142327 172401 142361
rect 172435 142327 172443 142361
rect 172393 142303 172443 142327
rect 172729 142361 172779 142385
rect 172729 142327 172737 142361
rect 172771 142327 172779 142361
rect 172729 142303 172779 142327
rect 173065 142361 173115 142385
rect 173065 142327 173073 142361
rect 173107 142327 173115 142361
rect 173065 142303 173115 142327
rect 173401 142361 173451 142385
rect 173401 142327 173409 142361
rect 173443 142327 173451 142361
rect 173401 142303 173451 142327
rect 173737 142361 173787 142385
rect 173737 142327 173745 142361
rect 173779 142327 173787 142361
rect 173737 142303 173787 142327
rect 174073 142361 174123 142385
rect 174073 142327 174081 142361
rect 174115 142327 174123 142361
rect 174073 142303 174123 142327
rect 174409 142361 174459 142385
rect 174409 142327 174417 142361
rect 174451 142327 174459 142361
rect 174409 142303 174459 142327
rect 174745 142361 174795 142385
rect 174745 142327 174753 142361
rect 174787 142327 174795 142361
rect 174745 142303 174795 142327
rect 175081 142361 175131 142385
rect 175081 142327 175089 142361
rect 175123 142327 175131 142361
rect 175081 142303 175131 142327
rect 175417 142361 175467 142385
rect 175417 142327 175425 142361
rect 175459 142327 175467 142361
rect 175417 142303 175467 142327
rect 175753 142361 175803 142385
rect 175753 142327 175761 142361
rect 175795 142327 175803 142361
rect 175753 142303 175803 142327
rect 176089 142361 176139 142385
rect 176089 142327 176097 142361
rect 176131 142327 176139 142361
rect 176089 142303 176139 142327
rect 176425 142361 176475 142385
rect 176425 142327 176433 142361
rect 176467 142327 176475 142361
rect 176425 142303 176475 142327
rect 176761 142361 176811 142385
rect 176761 142327 176769 142361
rect 176803 142327 176811 142361
rect 176761 142303 176811 142327
rect 177097 142361 177147 142385
rect 177097 142327 177105 142361
rect 177139 142327 177147 142361
rect 177097 142303 177147 142327
rect 177433 142361 177483 142385
rect 177433 142327 177441 142361
rect 177475 142327 177483 142361
rect 177433 142303 177483 142327
rect 177769 142361 177819 142385
rect 177769 142327 177777 142361
rect 177811 142327 177819 142361
rect 177769 142303 177819 142327
rect 178105 142361 178155 142385
rect 178105 142327 178113 142361
rect 178147 142327 178155 142361
rect 178105 142303 178155 142327
rect 178441 142361 178491 142385
rect 178441 142327 178449 142361
rect 178483 142327 178491 142361
rect 178441 142303 178491 142327
rect 178777 142361 178827 142385
rect 178777 142327 178785 142361
rect 178819 142327 178827 142361
rect 178777 142303 178827 142327
rect 179113 142361 179163 142385
rect 179113 142327 179121 142361
rect 179155 142327 179163 142361
rect 179113 142303 179163 142327
rect 179449 142361 179499 142385
rect 179449 142327 179457 142361
rect 179491 142327 179499 142361
rect 179449 142303 179499 142327
rect 179785 142361 179835 142385
rect 179785 142327 179793 142361
rect 179827 142327 179835 142361
rect 179785 142303 179835 142327
rect 180121 142361 180171 142385
rect 180121 142327 180129 142361
rect 180163 142327 180171 142361
rect 180121 142303 180171 142327
rect 180457 142361 180507 142385
rect 180457 142327 180465 142361
rect 180499 142327 180507 142361
rect 180457 142303 180507 142327
rect 180793 142361 180843 142385
rect 180793 142327 180801 142361
rect 180835 142327 180843 142361
rect 180793 142303 180843 142327
rect 181129 142361 181179 142385
rect 181129 142327 181137 142361
rect 181171 142327 181179 142361
rect 181129 142303 181179 142327
rect 181465 142361 181515 142385
rect 181465 142327 181473 142361
rect 181507 142327 181515 142361
rect 181465 142303 181515 142327
rect 181801 142361 181851 142385
rect 181801 142327 181809 142361
rect 181843 142327 181851 142361
rect 181801 142303 181851 142327
rect 182137 142361 182187 142385
rect 182137 142327 182145 142361
rect 182179 142327 182187 142361
rect 182137 142303 182187 142327
rect 182473 142361 182523 142385
rect 182473 142327 182481 142361
rect 182515 142327 182523 142361
rect 182473 142303 182523 142327
rect 182809 142361 182859 142385
rect 182809 142327 182817 142361
rect 182851 142327 182859 142361
rect 182809 142303 182859 142327
rect 183145 142361 183195 142385
rect 183145 142327 183153 142361
rect 183187 142327 183195 142361
rect 183145 142303 183195 142327
rect 183481 142361 183531 142385
rect 183481 142327 183489 142361
rect 183523 142327 183531 142361
rect 183481 142303 183531 142327
rect 183817 142361 183867 142385
rect 183817 142327 183825 142361
rect 183859 142327 183867 142361
rect 183817 142303 183867 142327
rect 184153 142361 184203 142385
rect 184153 142327 184161 142361
rect 184195 142327 184203 142361
rect 184153 142303 184203 142327
rect 184489 142361 184539 142385
rect 184489 142327 184497 142361
rect 184531 142327 184539 142361
rect 184489 142303 184539 142327
rect 184825 142361 184875 142385
rect 184825 142327 184833 142361
rect 184867 142327 184875 142361
rect 184825 142303 184875 142327
rect 185161 142361 185211 142385
rect 185161 142327 185169 142361
rect 185203 142327 185211 142361
rect 185161 142303 185211 142327
rect 185497 142361 185547 142385
rect 185497 142327 185505 142361
rect 185539 142327 185547 142361
rect 185497 142303 185547 142327
rect 185833 142361 185883 142385
rect 185833 142327 185841 142361
rect 185875 142327 185883 142361
rect 185833 142303 185883 142327
rect 186169 142361 186219 142385
rect 186169 142327 186177 142361
rect 186211 142327 186219 142361
rect 186169 142303 186219 142327
rect 186505 142361 186555 142385
rect 186505 142327 186513 142361
rect 186547 142327 186555 142361
rect 186505 142303 186555 142327
rect 186841 142361 186891 142385
rect 186841 142327 186849 142361
rect 186883 142327 186891 142361
rect 186841 142303 186891 142327
rect 187177 142361 187227 142385
rect 187177 142327 187185 142361
rect 187219 142327 187227 142361
rect 187177 142303 187227 142327
rect 187513 142361 187563 142385
rect 187513 142327 187521 142361
rect 187555 142327 187563 142361
rect 187513 142303 187563 142327
rect 187849 142361 187899 142385
rect 187849 142327 187857 142361
rect 187891 142327 187899 142361
rect 187849 142303 187899 142327
rect 188185 142361 188235 142385
rect 188185 142327 188193 142361
rect 188227 142327 188235 142361
rect 188185 142303 188235 142327
rect 188521 142361 188571 142385
rect 188521 142327 188529 142361
rect 188563 142327 188571 142361
rect 188521 142303 188571 142327
rect 188857 142361 188907 142385
rect 188857 142327 188865 142361
rect 188899 142327 188907 142361
rect 188857 142303 188907 142327
rect 189193 142361 189243 142385
rect 189193 142327 189201 142361
rect 189235 142327 189243 142361
rect 189193 142303 189243 142327
rect 189529 142361 189579 142385
rect 189529 142327 189537 142361
rect 189571 142327 189579 142361
rect 189529 142303 189579 142327
rect 189865 142361 189915 142385
rect 189865 142327 189873 142361
rect 189907 142327 189915 142361
rect 189865 142303 189915 142327
rect 190201 142361 190251 142385
rect 190201 142327 190209 142361
rect 190243 142327 190251 142361
rect 190201 142303 190251 142327
rect 190537 142361 190587 142385
rect 190537 142327 190545 142361
rect 190579 142327 190587 142361
rect 190537 142303 190587 142327
rect 190873 142361 190923 142385
rect 190873 142327 190881 142361
rect 190915 142327 190923 142361
rect 190873 142303 190923 142327
rect 191209 142361 191259 142385
rect 191209 142327 191217 142361
rect 191251 142327 191259 142361
rect 191209 142303 191259 142327
rect 191545 142361 191595 142385
rect 191545 142327 191553 142361
rect 191587 142327 191595 142361
rect 191545 142303 191595 142327
rect 191881 142361 191931 142385
rect 191881 142327 191889 142361
rect 191923 142327 191931 142361
rect 191881 142303 191931 142327
rect 192217 142361 192267 142385
rect 192217 142327 192225 142361
rect 192259 142327 192267 142361
rect 192217 142303 192267 142327
rect 192553 142361 192603 142385
rect 192553 142327 192561 142361
rect 192595 142327 192603 142361
rect 192553 142303 192603 142327
rect 192889 142361 192939 142385
rect 192889 142327 192897 142361
rect 192931 142327 192939 142361
rect 192889 142303 192939 142327
rect 193225 142361 193275 142385
rect 193225 142327 193233 142361
rect 193267 142327 193275 142361
rect 193225 142303 193275 142327
rect 193561 142361 193611 142385
rect 193561 142327 193569 142361
rect 193603 142327 193611 142361
rect 193561 142303 193611 142327
rect 193897 142361 193947 142385
rect 193897 142327 193905 142361
rect 193939 142327 193947 142361
rect 193897 142303 193947 142327
rect 194233 142361 194283 142385
rect 194233 142327 194241 142361
rect 194275 142327 194283 142361
rect 194233 142303 194283 142327
rect 194569 142361 194619 142385
rect 194569 142327 194577 142361
rect 194611 142327 194619 142361
rect 194569 142303 194619 142327
rect 194905 142361 194955 142385
rect 194905 142327 194913 142361
rect 194947 142327 194955 142361
rect 194905 142303 194955 142327
rect 195241 142361 195291 142385
rect 195241 142327 195249 142361
rect 195283 142327 195291 142361
rect 195241 142303 195291 142327
rect 195577 142361 195627 142385
rect 195577 142327 195585 142361
rect 195619 142327 195627 142361
rect 195577 142303 195627 142327
rect 195913 142361 195963 142385
rect 195913 142327 195921 142361
rect 195955 142327 195963 142361
rect 195913 142303 195963 142327
rect 196249 142361 196299 142385
rect 196249 142327 196257 142361
rect 196291 142327 196299 142361
rect 196249 142303 196299 142327
rect 196585 142361 196635 142385
rect 196585 142327 196593 142361
rect 196627 142327 196635 142361
rect 196585 142303 196635 142327
rect 196921 142361 196971 142385
rect 196921 142327 196929 142361
rect 196963 142327 196971 142361
rect 196921 142303 196971 142327
rect 197257 142361 197307 142385
rect 197257 142327 197265 142361
rect 197299 142327 197307 142361
rect 197257 142303 197307 142327
rect 197593 142361 197643 142385
rect 197593 142327 197601 142361
rect 197635 142327 197643 142361
rect 197593 142303 197643 142327
rect 197929 142361 197979 142385
rect 197929 142327 197937 142361
rect 197971 142327 197979 142361
rect 197929 142303 197979 142327
rect 198265 142361 198315 142385
rect 198265 142327 198273 142361
rect 198307 142327 198315 142361
rect 198265 142303 198315 142327
rect 198601 142361 198651 142385
rect 198601 142327 198609 142361
rect 198643 142327 198651 142361
rect 198601 142303 198651 142327
rect 198937 142361 198987 142385
rect 198937 142327 198945 142361
rect 198979 142327 198987 142361
rect 198937 142303 198987 142327
rect 199273 142361 199323 142385
rect 199273 142327 199281 142361
rect 199315 142327 199323 142361
rect 199273 142303 199323 142327
rect 199609 142361 199659 142385
rect 199609 142327 199617 142361
rect 199651 142327 199659 142361
rect 199609 142303 199659 142327
rect 199945 142361 199995 142385
rect 199945 142327 199953 142361
rect 199987 142327 199995 142361
rect 199945 142303 199995 142327
rect 200281 142361 200331 142385
rect 200281 142327 200289 142361
rect 200323 142327 200331 142361
rect 200281 142303 200331 142327
rect 200617 142361 200667 142385
rect 200617 142327 200625 142361
rect 200659 142327 200667 142361
rect 200617 142303 200667 142327
rect 200953 142361 201003 142385
rect 200953 142327 200961 142361
rect 200995 142327 201003 142361
rect 200953 142303 201003 142327
rect 201289 142361 201339 142385
rect 201289 142327 201297 142361
rect 201331 142327 201339 142361
rect 201289 142303 201339 142327
rect 201625 142361 201675 142385
rect 201625 142327 201633 142361
rect 201667 142327 201675 142361
rect 201625 142303 201675 142327
rect 201961 142361 202011 142385
rect 201961 142327 201969 142361
rect 202003 142327 202011 142361
rect 201961 142303 202011 142327
rect 202297 142361 202347 142385
rect 202297 142327 202305 142361
rect 202339 142327 202347 142361
rect 202297 142303 202347 142327
rect 202633 142361 202683 142385
rect 202633 142327 202641 142361
rect 202675 142327 202683 142361
rect 202633 142303 202683 142327
rect 202969 142361 203019 142385
rect 202969 142327 202977 142361
rect 203011 142327 203019 142361
rect 202969 142303 203019 142327
rect 203305 142361 203355 142385
rect 203305 142327 203313 142361
rect 203347 142327 203355 142361
rect 203305 142303 203355 142327
rect 203641 142361 203691 142385
rect 203641 142327 203649 142361
rect 203683 142327 203691 142361
rect 203641 142303 203691 142327
rect 203977 142361 204027 142385
rect 203977 142327 203985 142361
rect 204019 142327 204027 142361
rect 203977 142303 204027 142327
rect 204313 142361 204363 142385
rect 204313 142327 204321 142361
rect 204355 142327 204363 142361
rect 204313 142303 204363 142327
rect 204649 142361 204699 142385
rect 204649 142327 204657 142361
rect 204691 142327 204699 142361
rect 204649 142303 204699 142327
rect 204985 142361 205035 142385
rect 204985 142327 204993 142361
rect 205027 142327 205035 142361
rect 204985 142303 205035 142327
rect 205321 142361 205371 142385
rect 205321 142327 205329 142361
rect 205363 142327 205371 142361
rect 205321 142303 205371 142327
rect 205657 142361 205707 142385
rect 205657 142327 205665 142361
rect 205699 142327 205707 142361
rect 205657 142303 205707 142327
rect 205993 142361 206043 142385
rect 205993 142327 206001 142361
rect 206035 142327 206043 142361
rect 205993 142303 206043 142327
rect 206329 142361 206379 142385
rect 206329 142327 206337 142361
rect 206371 142327 206379 142361
rect 206329 142303 206379 142327
rect 206665 142361 206715 142385
rect 206665 142327 206673 142361
rect 206707 142327 206715 142361
rect 206665 142303 206715 142327
rect 207001 142361 207051 142385
rect 207001 142327 207009 142361
rect 207043 142327 207051 142361
rect 207001 142303 207051 142327
rect 207337 142361 207387 142385
rect 207337 142327 207345 142361
rect 207379 142327 207387 142361
rect 207337 142303 207387 142327
rect 207673 142361 207723 142385
rect 207673 142327 207681 142361
rect 207715 142327 207723 142361
rect 207673 142303 207723 142327
rect 208009 142361 208059 142385
rect 208009 142327 208017 142361
rect 208051 142327 208059 142361
rect 208009 142303 208059 142327
rect 208345 142361 208395 142385
rect 208345 142327 208353 142361
rect 208387 142327 208395 142361
rect 208345 142303 208395 142327
rect 208681 142361 208731 142385
rect 208681 142327 208689 142361
rect 208723 142327 208731 142361
rect 208681 142303 208731 142327
rect 209017 142361 209067 142385
rect 209017 142327 209025 142361
rect 209059 142327 209067 142361
rect 209017 142303 209067 142327
rect 209353 142361 209403 142385
rect 209353 142327 209361 142361
rect 209395 142327 209403 142361
rect 209353 142303 209403 142327
rect 209689 142361 209739 142385
rect 209689 142327 209697 142361
rect 209731 142327 209739 142361
rect 209689 142303 209739 142327
rect 210025 142361 210075 142385
rect 210025 142327 210033 142361
rect 210067 142327 210075 142361
rect 210025 142303 210075 142327
rect 210361 142361 210411 142385
rect 210361 142327 210369 142361
rect 210403 142327 210411 142361
rect 210361 142303 210411 142327
rect 210697 142361 210747 142385
rect 210697 142327 210705 142361
rect 210739 142327 210747 142361
rect 210697 142303 210747 142327
rect 211033 142361 211083 142385
rect 211033 142327 211041 142361
rect 211075 142327 211083 142361
rect 211033 142303 211083 142327
rect 211369 142361 211419 142385
rect 211369 142327 211377 142361
rect 211411 142327 211419 142361
rect 211369 142303 211419 142327
rect 211705 142361 211755 142385
rect 211705 142327 211713 142361
rect 211747 142327 211755 142361
rect 211705 142303 211755 142327
rect 212041 142361 212091 142385
rect 212041 142327 212049 142361
rect 212083 142327 212091 142361
rect 212041 142303 212091 142327
rect 212377 142361 212427 142385
rect 212377 142327 212385 142361
rect 212419 142327 212427 142361
rect 212377 142303 212427 142327
rect 212713 142361 212763 142385
rect 212713 142327 212721 142361
rect 212755 142327 212763 142361
rect 212713 142303 212763 142327
rect 213049 142361 213099 142385
rect 213049 142327 213057 142361
rect 213091 142327 213099 142361
rect 213049 142303 213099 142327
rect 213385 142361 213435 142385
rect 213385 142327 213393 142361
rect 213427 142327 213435 142361
rect 213385 142303 213435 142327
rect 213721 142361 213771 142385
rect 213721 142327 213729 142361
rect 213763 142327 213771 142361
rect 213721 142303 213771 142327
rect 214057 142361 214107 142385
rect 214057 142327 214065 142361
rect 214099 142327 214107 142361
rect 214057 142303 214107 142327
rect 214393 142361 214443 142385
rect 214393 142327 214401 142361
rect 214435 142327 214443 142361
rect 214393 142303 214443 142327
rect 214729 142361 214779 142385
rect 214729 142327 214737 142361
rect 214771 142327 214779 142361
rect 214729 142303 214779 142327
rect 215065 142361 215115 142385
rect 215065 142327 215073 142361
rect 215107 142327 215115 142361
rect 215065 142303 215115 142327
rect 215401 142361 215451 142385
rect 215401 142327 215409 142361
rect 215443 142327 215451 142361
rect 215401 142303 215451 142327
rect 215737 142361 215787 142385
rect 215737 142327 215745 142361
rect 215779 142327 215787 142361
rect 215737 142303 215787 142327
rect 216073 142361 216123 142385
rect 216073 142327 216081 142361
rect 216115 142327 216123 142361
rect 216073 142303 216123 142327
rect 216409 142361 216459 142385
rect 216409 142327 216417 142361
rect 216451 142327 216459 142361
rect 216409 142303 216459 142327
rect 1705 141977 1755 142001
rect 1705 141943 1713 141977
rect 1747 141943 1755 141977
rect 1705 141919 1755 141943
rect 216911 141977 216961 142001
rect 216911 141943 216919 141977
rect 216953 141943 216961 141977
rect 216911 141919 216961 141943
rect 1705 141641 1755 141665
rect 1705 141607 1713 141641
rect 1747 141607 1755 141641
rect 1705 141583 1755 141607
rect 216911 141641 216961 141665
rect 216911 141607 216919 141641
rect 216953 141607 216961 141641
rect 216911 141583 216961 141607
rect 1705 141305 1755 141329
rect 1705 141271 1713 141305
rect 1747 141271 1755 141305
rect 1705 141247 1755 141271
rect 216911 141305 216961 141329
rect 216911 141271 216919 141305
rect 216953 141271 216961 141305
rect 216911 141247 216961 141271
rect 1705 140969 1755 140993
rect 1705 140935 1713 140969
rect 1747 140935 1755 140969
rect 1705 140911 1755 140935
rect 216911 140969 216961 140993
rect 216911 140935 216919 140969
rect 216953 140935 216961 140969
rect 216911 140911 216961 140935
rect 1705 140633 1755 140657
rect 1705 140599 1713 140633
rect 1747 140599 1755 140633
rect 1705 140575 1755 140599
rect 216911 140633 216961 140657
rect 216911 140599 216919 140633
rect 216953 140599 216961 140633
rect 216911 140575 216961 140599
rect 1705 140297 1755 140321
rect 1705 140263 1713 140297
rect 1747 140263 1755 140297
rect 1705 140239 1755 140263
rect 216911 140297 216961 140321
rect 216911 140263 216919 140297
rect 216953 140263 216961 140297
rect 216911 140239 216961 140263
rect 1705 139961 1755 139985
rect 1705 139927 1713 139961
rect 1747 139927 1755 139961
rect 1705 139903 1755 139927
rect 216911 139961 216961 139985
rect 216911 139927 216919 139961
rect 216953 139927 216961 139961
rect 216911 139903 216961 139927
rect 1705 139625 1755 139649
rect 1705 139591 1713 139625
rect 1747 139591 1755 139625
rect 1705 139567 1755 139591
rect 216911 139625 216961 139649
rect 216911 139591 216919 139625
rect 216953 139591 216961 139625
rect 216911 139567 216961 139591
rect 1705 139289 1755 139313
rect 1705 139255 1713 139289
rect 1747 139255 1755 139289
rect 1705 139231 1755 139255
rect 216911 139289 216961 139313
rect 216911 139255 216919 139289
rect 216953 139255 216961 139289
rect 216911 139231 216961 139255
rect 1705 138953 1755 138977
rect 1705 138919 1713 138953
rect 1747 138919 1755 138953
rect 1705 138895 1755 138919
rect 216911 138953 216961 138977
rect 216911 138919 216919 138953
rect 216953 138919 216961 138953
rect 216911 138895 216961 138919
rect 1705 138617 1755 138641
rect 1705 138583 1713 138617
rect 1747 138583 1755 138617
rect 1705 138559 1755 138583
rect 216911 138617 216961 138641
rect 216911 138583 216919 138617
rect 216953 138583 216961 138617
rect 216911 138559 216961 138583
rect 1705 138281 1755 138305
rect 1705 138247 1713 138281
rect 1747 138247 1755 138281
rect 1705 138223 1755 138247
rect 216911 138281 216961 138305
rect 216911 138247 216919 138281
rect 216953 138247 216961 138281
rect 216911 138223 216961 138247
rect 1705 137945 1755 137969
rect 1705 137911 1713 137945
rect 1747 137911 1755 137945
rect 1705 137887 1755 137911
rect 216911 137945 216961 137969
rect 216911 137911 216919 137945
rect 216953 137911 216961 137945
rect 216911 137887 216961 137911
rect 1705 137609 1755 137633
rect 1705 137575 1713 137609
rect 1747 137575 1755 137609
rect 1705 137551 1755 137575
rect 216911 137609 216961 137633
rect 216911 137575 216919 137609
rect 216953 137575 216961 137609
rect 216911 137551 216961 137575
rect 1705 137273 1755 137297
rect 1705 137239 1713 137273
rect 1747 137239 1755 137273
rect 1705 137215 1755 137239
rect 216911 137273 216961 137297
rect 216911 137239 216919 137273
rect 216953 137239 216961 137273
rect 216911 137215 216961 137239
rect 1705 136937 1755 136961
rect 1705 136903 1713 136937
rect 1747 136903 1755 136937
rect 1705 136879 1755 136903
rect 216911 136937 216961 136961
rect 216911 136903 216919 136937
rect 216953 136903 216961 136937
rect 216911 136879 216961 136903
rect 1705 136601 1755 136625
rect 1705 136567 1713 136601
rect 1747 136567 1755 136601
rect 1705 136543 1755 136567
rect 216911 136601 216961 136625
rect 216911 136567 216919 136601
rect 216953 136567 216961 136601
rect 216911 136543 216961 136567
rect 1705 136265 1755 136289
rect 1705 136231 1713 136265
rect 1747 136231 1755 136265
rect 1705 136207 1755 136231
rect 216911 136265 216961 136289
rect 216911 136231 216919 136265
rect 216953 136231 216961 136265
rect 216911 136207 216961 136231
rect 1705 135929 1755 135953
rect 1705 135895 1713 135929
rect 1747 135895 1755 135929
rect 1705 135871 1755 135895
rect 216911 135929 216961 135953
rect 216911 135895 216919 135929
rect 216953 135895 216961 135929
rect 216911 135871 216961 135895
rect 1705 135593 1755 135617
rect 1705 135559 1713 135593
rect 1747 135559 1755 135593
rect 1705 135535 1755 135559
rect 216911 135593 216961 135617
rect 216911 135559 216919 135593
rect 216953 135559 216961 135593
rect 216911 135535 216961 135559
rect 1705 135257 1755 135281
rect 1705 135223 1713 135257
rect 1747 135223 1755 135257
rect 1705 135199 1755 135223
rect 216911 135257 216961 135281
rect 216911 135223 216919 135257
rect 216953 135223 216961 135257
rect 216911 135199 216961 135223
rect 1705 134921 1755 134945
rect 1705 134887 1713 134921
rect 1747 134887 1755 134921
rect 1705 134863 1755 134887
rect 216911 134921 216961 134945
rect 216911 134887 216919 134921
rect 216953 134887 216961 134921
rect 216911 134863 216961 134887
rect 1705 134585 1755 134609
rect 1705 134551 1713 134585
rect 1747 134551 1755 134585
rect 1705 134527 1755 134551
rect 216911 134585 216961 134609
rect 216911 134551 216919 134585
rect 216953 134551 216961 134585
rect 216911 134527 216961 134551
rect 1705 134249 1755 134273
rect 1705 134215 1713 134249
rect 1747 134215 1755 134249
rect 1705 134191 1755 134215
rect 216911 134249 216961 134273
rect 216911 134215 216919 134249
rect 216953 134215 216961 134249
rect 216911 134191 216961 134215
rect 1705 133913 1755 133937
rect 1705 133879 1713 133913
rect 1747 133879 1755 133913
rect 1705 133855 1755 133879
rect 216911 133913 216961 133937
rect 216911 133879 216919 133913
rect 216953 133879 216961 133913
rect 216911 133855 216961 133879
rect 1705 133577 1755 133601
rect 1705 133543 1713 133577
rect 1747 133543 1755 133577
rect 1705 133519 1755 133543
rect 216911 133577 216961 133601
rect 216911 133543 216919 133577
rect 216953 133543 216961 133577
rect 216911 133519 216961 133543
rect 1705 133241 1755 133265
rect 1705 133207 1713 133241
rect 1747 133207 1755 133241
rect 1705 133183 1755 133207
rect 216911 133241 216961 133265
rect 216911 133207 216919 133241
rect 216953 133207 216961 133241
rect 216911 133183 216961 133207
rect 1705 132905 1755 132929
rect 1705 132871 1713 132905
rect 1747 132871 1755 132905
rect 1705 132847 1755 132871
rect 216911 132905 216961 132929
rect 216911 132871 216919 132905
rect 216953 132871 216961 132905
rect 216911 132847 216961 132871
rect 1705 132569 1755 132593
rect 1705 132535 1713 132569
rect 1747 132535 1755 132569
rect 1705 132511 1755 132535
rect 216911 132569 216961 132593
rect 216911 132535 216919 132569
rect 216953 132535 216961 132569
rect 216911 132511 216961 132535
rect 1705 132233 1755 132257
rect 1705 132199 1713 132233
rect 1747 132199 1755 132233
rect 1705 132175 1755 132199
rect 216911 132233 216961 132257
rect 216911 132199 216919 132233
rect 216953 132199 216961 132233
rect 216911 132175 216961 132199
rect 1705 131897 1755 131921
rect 1705 131863 1713 131897
rect 1747 131863 1755 131897
rect 1705 131839 1755 131863
rect 216911 131897 216961 131921
rect 216911 131863 216919 131897
rect 216953 131863 216961 131897
rect 216911 131839 216961 131863
rect 1705 131561 1755 131585
rect 1705 131527 1713 131561
rect 1747 131527 1755 131561
rect 1705 131503 1755 131527
rect 216911 131561 216961 131585
rect 216911 131527 216919 131561
rect 216953 131527 216961 131561
rect 216911 131503 216961 131527
rect 1705 131225 1755 131249
rect 1705 131191 1713 131225
rect 1747 131191 1755 131225
rect 1705 131167 1755 131191
rect 216911 131225 216961 131249
rect 216911 131191 216919 131225
rect 216953 131191 216961 131225
rect 216911 131167 216961 131191
rect 1705 130889 1755 130913
rect 1705 130855 1713 130889
rect 1747 130855 1755 130889
rect 1705 130831 1755 130855
rect 216911 130889 216961 130913
rect 216911 130855 216919 130889
rect 216953 130855 216961 130889
rect 216911 130831 216961 130855
rect 1705 130553 1755 130577
rect 1705 130519 1713 130553
rect 1747 130519 1755 130553
rect 1705 130495 1755 130519
rect 216911 130553 216961 130577
rect 216911 130519 216919 130553
rect 216953 130519 216961 130553
rect 216911 130495 216961 130519
rect 1705 130217 1755 130241
rect 1705 130183 1713 130217
rect 1747 130183 1755 130217
rect 1705 130159 1755 130183
rect 216911 130217 216961 130241
rect 216911 130183 216919 130217
rect 216953 130183 216961 130217
rect 216911 130159 216961 130183
rect 1705 129881 1755 129905
rect 1705 129847 1713 129881
rect 1747 129847 1755 129881
rect 1705 129823 1755 129847
rect 216911 129881 216961 129905
rect 216911 129847 216919 129881
rect 216953 129847 216961 129881
rect 216911 129823 216961 129847
rect 1705 129545 1755 129569
rect 1705 129511 1713 129545
rect 1747 129511 1755 129545
rect 1705 129487 1755 129511
rect 216911 129545 216961 129569
rect 216911 129511 216919 129545
rect 216953 129511 216961 129545
rect 216911 129487 216961 129511
rect 1705 129209 1755 129233
rect 1705 129175 1713 129209
rect 1747 129175 1755 129209
rect 1705 129151 1755 129175
rect 216911 129209 216961 129233
rect 216911 129175 216919 129209
rect 216953 129175 216961 129209
rect 216911 129151 216961 129175
rect 1705 128873 1755 128897
rect 1705 128839 1713 128873
rect 1747 128839 1755 128873
rect 1705 128815 1755 128839
rect 216911 128873 216961 128897
rect 216911 128839 216919 128873
rect 216953 128839 216961 128873
rect 216911 128815 216961 128839
rect 1705 128537 1755 128561
rect 1705 128503 1713 128537
rect 1747 128503 1755 128537
rect 1705 128479 1755 128503
rect 216911 128537 216961 128561
rect 216911 128503 216919 128537
rect 216953 128503 216961 128537
rect 216911 128479 216961 128503
rect 1705 128201 1755 128225
rect 1705 128167 1713 128201
rect 1747 128167 1755 128201
rect 1705 128143 1755 128167
rect 216911 128201 216961 128225
rect 216911 128167 216919 128201
rect 216953 128167 216961 128201
rect 216911 128143 216961 128167
rect 1705 127865 1755 127889
rect 1705 127831 1713 127865
rect 1747 127831 1755 127865
rect 1705 127807 1755 127831
rect 216911 127865 216961 127889
rect 216911 127831 216919 127865
rect 216953 127831 216961 127865
rect 216911 127807 216961 127831
rect 1705 127529 1755 127553
rect 1705 127495 1713 127529
rect 1747 127495 1755 127529
rect 1705 127471 1755 127495
rect 216911 127529 216961 127553
rect 216911 127495 216919 127529
rect 216953 127495 216961 127529
rect 216911 127471 216961 127495
rect 1705 127193 1755 127217
rect 1705 127159 1713 127193
rect 1747 127159 1755 127193
rect 1705 127135 1755 127159
rect 216911 127193 216961 127217
rect 216911 127159 216919 127193
rect 216953 127159 216961 127193
rect 216911 127135 216961 127159
rect 1705 126857 1755 126881
rect 1705 126823 1713 126857
rect 1747 126823 1755 126857
rect 1705 126799 1755 126823
rect 216911 126857 216961 126881
rect 216911 126823 216919 126857
rect 216953 126823 216961 126857
rect 216911 126799 216961 126823
rect 1705 126521 1755 126545
rect 1705 126487 1713 126521
rect 1747 126487 1755 126521
rect 1705 126463 1755 126487
rect 216911 126521 216961 126545
rect 216911 126487 216919 126521
rect 216953 126487 216961 126521
rect 216911 126463 216961 126487
rect 1705 126185 1755 126209
rect 1705 126151 1713 126185
rect 1747 126151 1755 126185
rect 1705 126127 1755 126151
rect 216911 126185 216961 126209
rect 216911 126151 216919 126185
rect 216953 126151 216961 126185
rect 216911 126127 216961 126151
rect 1705 125849 1755 125873
rect 1705 125815 1713 125849
rect 1747 125815 1755 125849
rect 1705 125791 1755 125815
rect 216911 125849 216961 125873
rect 216911 125815 216919 125849
rect 216953 125815 216961 125849
rect 216911 125791 216961 125815
rect 1705 125513 1755 125537
rect 1705 125479 1713 125513
rect 1747 125479 1755 125513
rect 1705 125455 1755 125479
rect 216911 125513 216961 125537
rect 216911 125479 216919 125513
rect 216953 125479 216961 125513
rect 216911 125455 216961 125479
rect 1705 125177 1755 125201
rect 1705 125143 1713 125177
rect 1747 125143 1755 125177
rect 1705 125119 1755 125143
rect 216911 125177 216961 125201
rect 216911 125143 216919 125177
rect 216953 125143 216961 125177
rect 216911 125119 216961 125143
rect 1705 124841 1755 124865
rect 1705 124807 1713 124841
rect 1747 124807 1755 124841
rect 1705 124783 1755 124807
rect 216911 124841 216961 124865
rect 216911 124807 216919 124841
rect 216953 124807 216961 124841
rect 216911 124783 216961 124807
rect 1705 124505 1755 124529
rect 1705 124471 1713 124505
rect 1747 124471 1755 124505
rect 1705 124447 1755 124471
rect 216911 124505 216961 124529
rect 216911 124471 216919 124505
rect 216953 124471 216961 124505
rect 216911 124447 216961 124471
rect 1705 124169 1755 124193
rect 1705 124135 1713 124169
rect 1747 124135 1755 124169
rect 1705 124111 1755 124135
rect 216911 124169 216961 124193
rect 216911 124135 216919 124169
rect 216953 124135 216961 124169
rect 216911 124111 216961 124135
rect 1705 123833 1755 123857
rect 1705 123799 1713 123833
rect 1747 123799 1755 123833
rect 1705 123775 1755 123799
rect 216911 123833 216961 123857
rect 216911 123799 216919 123833
rect 216953 123799 216961 123833
rect 216911 123775 216961 123799
rect 1705 123497 1755 123521
rect 1705 123463 1713 123497
rect 1747 123463 1755 123497
rect 1705 123439 1755 123463
rect 216911 123497 216961 123521
rect 216911 123463 216919 123497
rect 216953 123463 216961 123497
rect 216911 123439 216961 123463
rect 1705 123161 1755 123185
rect 1705 123127 1713 123161
rect 1747 123127 1755 123161
rect 1705 123103 1755 123127
rect 216911 123161 216961 123185
rect 216911 123127 216919 123161
rect 216953 123127 216961 123161
rect 216911 123103 216961 123127
rect 1705 122825 1755 122849
rect 1705 122791 1713 122825
rect 1747 122791 1755 122825
rect 1705 122767 1755 122791
rect 216911 122825 216961 122849
rect 216911 122791 216919 122825
rect 216953 122791 216961 122825
rect 216911 122767 216961 122791
rect 1705 122489 1755 122513
rect 1705 122455 1713 122489
rect 1747 122455 1755 122489
rect 1705 122431 1755 122455
rect 216911 122489 216961 122513
rect 216911 122455 216919 122489
rect 216953 122455 216961 122489
rect 216911 122431 216961 122455
rect 1705 122153 1755 122177
rect 1705 122119 1713 122153
rect 1747 122119 1755 122153
rect 1705 122095 1755 122119
rect 216911 122153 216961 122177
rect 216911 122119 216919 122153
rect 216953 122119 216961 122153
rect 216911 122095 216961 122119
rect 1705 121817 1755 121841
rect 1705 121783 1713 121817
rect 1747 121783 1755 121817
rect 1705 121759 1755 121783
rect 216911 121817 216961 121841
rect 216911 121783 216919 121817
rect 216953 121783 216961 121817
rect 216911 121759 216961 121783
rect 1705 121481 1755 121505
rect 1705 121447 1713 121481
rect 1747 121447 1755 121481
rect 1705 121423 1755 121447
rect 216911 121481 216961 121505
rect 216911 121447 216919 121481
rect 216953 121447 216961 121481
rect 216911 121423 216961 121447
rect 1705 121145 1755 121169
rect 1705 121111 1713 121145
rect 1747 121111 1755 121145
rect 1705 121087 1755 121111
rect 216911 121145 216961 121169
rect 216911 121111 216919 121145
rect 216953 121111 216961 121145
rect 216911 121087 216961 121111
rect 1705 120809 1755 120833
rect 1705 120775 1713 120809
rect 1747 120775 1755 120809
rect 1705 120751 1755 120775
rect 216911 120809 216961 120833
rect 216911 120775 216919 120809
rect 216953 120775 216961 120809
rect 216911 120751 216961 120775
rect 1705 120473 1755 120497
rect 1705 120439 1713 120473
rect 1747 120439 1755 120473
rect 1705 120415 1755 120439
rect 216911 120473 216961 120497
rect 216911 120439 216919 120473
rect 216953 120439 216961 120473
rect 216911 120415 216961 120439
rect 1705 120137 1755 120161
rect 1705 120103 1713 120137
rect 1747 120103 1755 120137
rect 1705 120079 1755 120103
rect 216911 120137 216961 120161
rect 216911 120103 216919 120137
rect 216953 120103 216961 120137
rect 216911 120079 216961 120103
rect 1705 119801 1755 119825
rect 1705 119767 1713 119801
rect 1747 119767 1755 119801
rect 1705 119743 1755 119767
rect 216911 119801 216961 119825
rect 216911 119767 216919 119801
rect 216953 119767 216961 119801
rect 216911 119743 216961 119767
rect 1705 119465 1755 119489
rect 1705 119431 1713 119465
rect 1747 119431 1755 119465
rect 1705 119407 1755 119431
rect 216911 119465 216961 119489
rect 216911 119431 216919 119465
rect 216953 119431 216961 119465
rect 216911 119407 216961 119431
rect 1705 119129 1755 119153
rect 1705 119095 1713 119129
rect 1747 119095 1755 119129
rect 1705 119071 1755 119095
rect 216911 119129 216961 119153
rect 216911 119095 216919 119129
rect 216953 119095 216961 119129
rect 216911 119071 216961 119095
rect 1705 118793 1755 118817
rect 1705 118759 1713 118793
rect 1747 118759 1755 118793
rect 1705 118735 1755 118759
rect 216911 118793 216961 118817
rect 216911 118759 216919 118793
rect 216953 118759 216961 118793
rect 216911 118735 216961 118759
rect 1705 118457 1755 118481
rect 1705 118423 1713 118457
rect 1747 118423 1755 118457
rect 1705 118399 1755 118423
rect 216911 118457 216961 118481
rect 216911 118423 216919 118457
rect 216953 118423 216961 118457
rect 216911 118399 216961 118423
rect 1705 118121 1755 118145
rect 1705 118087 1713 118121
rect 1747 118087 1755 118121
rect 1705 118063 1755 118087
rect 216911 118121 216961 118145
rect 216911 118087 216919 118121
rect 216953 118087 216961 118121
rect 216911 118063 216961 118087
rect 1705 117785 1755 117809
rect 1705 117751 1713 117785
rect 1747 117751 1755 117785
rect 1705 117727 1755 117751
rect 216911 117785 216961 117809
rect 216911 117751 216919 117785
rect 216953 117751 216961 117785
rect 216911 117727 216961 117751
rect 1705 117449 1755 117473
rect 1705 117415 1713 117449
rect 1747 117415 1755 117449
rect 1705 117391 1755 117415
rect 216911 117449 216961 117473
rect 216911 117415 216919 117449
rect 216953 117415 216961 117449
rect 216911 117391 216961 117415
rect 1705 117113 1755 117137
rect 1705 117079 1713 117113
rect 1747 117079 1755 117113
rect 1705 117055 1755 117079
rect 216911 117113 216961 117137
rect 216911 117079 216919 117113
rect 216953 117079 216961 117113
rect 216911 117055 216961 117079
rect 1705 116777 1755 116801
rect 1705 116743 1713 116777
rect 1747 116743 1755 116777
rect 1705 116719 1755 116743
rect 216911 116777 216961 116801
rect 216911 116743 216919 116777
rect 216953 116743 216961 116777
rect 216911 116719 216961 116743
rect 1705 116441 1755 116465
rect 1705 116407 1713 116441
rect 1747 116407 1755 116441
rect 1705 116383 1755 116407
rect 216911 116441 216961 116465
rect 216911 116407 216919 116441
rect 216953 116407 216961 116441
rect 216911 116383 216961 116407
rect 1705 116105 1755 116129
rect 1705 116071 1713 116105
rect 1747 116071 1755 116105
rect 1705 116047 1755 116071
rect 216911 116105 216961 116129
rect 216911 116071 216919 116105
rect 216953 116071 216961 116105
rect 216911 116047 216961 116071
rect 1705 115769 1755 115793
rect 1705 115735 1713 115769
rect 1747 115735 1755 115769
rect 1705 115711 1755 115735
rect 216911 115769 216961 115793
rect 216911 115735 216919 115769
rect 216953 115735 216961 115769
rect 216911 115711 216961 115735
rect 1705 115433 1755 115457
rect 1705 115399 1713 115433
rect 1747 115399 1755 115433
rect 1705 115375 1755 115399
rect 216911 115433 216961 115457
rect 216911 115399 216919 115433
rect 216953 115399 216961 115433
rect 216911 115375 216961 115399
rect 1705 115097 1755 115121
rect 1705 115063 1713 115097
rect 1747 115063 1755 115097
rect 1705 115039 1755 115063
rect 216911 115097 216961 115121
rect 216911 115063 216919 115097
rect 216953 115063 216961 115097
rect 216911 115039 216961 115063
rect 1705 114761 1755 114785
rect 1705 114727 1713 114761
rect 1747 114727 1755 114761
rect 1705 114703 1755 114727
rect 216911 114761 216961 114785
rect 216911 114727 216919 114761
rect 216953 114727 216961 114761
rect 216911 114703 216961 114727
rect 1705 114425 1755 114449
rect 1705 114391 1713 114425
rect 1747 114391 1755 114425
rect 1705 114367 1755 114391
rect 216911 114425 216961 114449
rect 216911 114391 216919 114425
rect 216953 114391 216961 114425
rect 216911 114367 216961 114391
rect 1705 114089 1755 114113
rect 1705 114055 1713 114089
rect 1747 114055 1755 114089
rect 1705 114031 1755 114055
rect 216911 114089 216961 114113
rect 216911 114055 216919 114089
rect 216953 114055 216961 114089
rect 216911 114031 216961 114055
rect 1705 113753 1755 113777
rect 1705 113719 1713 113753
rect 1747 113719 1755 113753
rect 1705 113695 1755 113719
rect 216911 113753 216961 113777
rect 216911 113719 216919 113753
rect 216953 113719 216961 113753
rect 216911 113695 216961 113719
rect 1705 113417 1755 113441
rect 1705 113383 1713 113417
rect 1747 113383 1755 113417
rect 1705 113359 1755 113383
rect 216911 113417 216961 113441
rect 216911 113383 216919 113417
rect 216953 113383 216961 113417
rect 216911 113359 216961 113383
rect 1705 113081 1755 113105
rect 1705 113047 1713 113081
rect 1747 113047 1755 113081
rect 1705 113023 1755 113047
rect 216911 113081 216961 113105
rect 216911 113047 216919 113081
rect 216953 113047 216961 113081
rect 216911 113023 216961 113047
rect 1705 112745 1755 112769
rect 1705 112711 1713 112745
rect 1747 112711 1755 112745
rect 1705 112687 1755 112711
rect 216911 112745 216961 112769
rect 216911 112711 216919 112745
rect 216953 112711 216961 112745
rect 216911 112687 216961 112711
rect 1705 112409 1755 112433
rect 1705 112375 1713 112409
rect 1747 112375 1755 112409
rect 1705 112351 1755 112375
rect 216911 112409 216961 112433
rect 216911 112375 216919 112409
rect 216953 112375 216961 112409
rect 216911 112351 216961 112375
rect 1705 112073 1755 112097
rect 1705 112039 1713 112073
rect 1747 112039 1755 112073
rect 1705 112015 1755 112039
rect 216911 112073 216961 112097
rect 216911 112039 216919 112073
rect 216953 112039 216961 112073
rect 216911 112015 216961 112039
rect 1705 111737 1755 111761
rect 1705 111703 1713 111737
rect 1747 111703 1755 111737
rect 1705 111679 1755 111703
rect 216911 111737 216961 111761
rect 216911 111703 216919 111737
rect 216953 111703 216961 111737
rect 216911 111679 216961 111703
rect 1705 111401 1755 111425
rect 1705 111367 1713 111401
rect 1747 111367 1755 111401
rect 1705 111343 1755 111367
rect 216911 111401 216961 111425
rect 216911 111367 216919 111401
rect 216953 111367 216961 111401
rect 216911 111343 216961 111367
rect 1705 111065 1755 111089
rect 1705 111031 1713 111065
rect 1747 111031 1755 111065
rect 1705 111007 1755 111031
rect 216911 111065 216961 111089
rect 216911 111031 216919 111065
rect 216953 111031 216961 111065
rect 216911 111007 216961 111031
rect 1705 110729 1755 110753
rect 1705 110695 1713 110729
rect 1747 110695 1755 110729
rect 1705 110671 1755 110695
rect 216911 110729 216961 110753
rect 216911 110695 216919 110729
rect 216953 110695 216961 110729
rect 216911 110671 216961 110695
rect 1705 110393 1755 110417
rect 1705 110359 1713 110393
rect 1747 110359 1755 110393
rect 1705 110335 1755 110359
rect 216911 110393 216961 110417
rect 216911 110359 216919 110393
rect 216953 110359 216961 110393
rect 216911 110335 216961 110359
rect 1705 110057 1755 110081
rect 1705 110023 1713 110057
rect 1747 110023 1755 110057
rect 1705 109999 1755 110023
rect 216911 110057 216961 110081
rect 216911 110023 216919 110057
rect 216953 110023 216961 110057
rect 216911 109999 216961 110023
rect 1705 109721 1755 109745
rect 1705 109687 1713 109721
rect 1747 109687 1755 109721
rect 1705 109663 1755 109687
rect 216911 109721 216961 109745
rect 216911 109687 216919 109721
rect 216953 109687 216961 109721
rect 216911 109663 216961 109687
rect 1705 109385 1755 109409
rect 1705 109351 1713 109385
rect 1747 109351 1755 109385
rect 1705 109327 1755 109351
rect 216911 109385 216961 109409
rect 216911 109351 216919 109385
rect 216953 109351 216961 109385
rect 216911 109327 216961 109351
rect 1705 109049 1755 109073
rect 1705 109015 1713 109049
rect 1747 109015 1755 109049
rect 1705 108991 1755 109015
rect 216911 109049 216961 109073
rect 216911 109015 216919 109049
rect 216953 109015 216961 109049
rect 216911 108991 216961 109015
rect 1705 108713 1755 108737
rect 1705 108679 1713 108713
rect 1747 108679 1755 108713
rect 1705 108655 1755 108679
rect 216911 108713 216961 108737
rect 216911 108679 216919 108713
rect 216953 108679 216961 108713
rect 216911 108655 216961 108679
rect 1705 108377 1755 108401
rect 1705 108343 1713 108377
rect 1747 108343 1755 108377
rect 1705 108319 1755 108343
rect 216911 108377 216961 108401
rect 216911 108343 216919 108377
rect 216953 108343 216961 108377
rect 216911 108319 216961 108343
rect 1705 108041 1755 108065
rect 1705 108007 1713 108041
rect 1747 108007 1755 108041
rect 1705 107983 1755 108007
rect 216911 108041 216961 108065
rect 216911 108007 216919 108041
rect 216953 108007 216961 108041
rect 216911 107983 216961 108007
rect 1705 107705 1755 107729
rect 1705 107671 1713 107705
rect 1747 107671 1755 107705
rect 1705 107647 1755 107671
rect 216911 107705 216961 107729
rect 216911 107671 216919 107705
rect 216953 107671 216961 107705
rect 216911 107647 216961 107671
rect 1705 107369 1755 107393
rect 1705 107335 1713 107369
rect 1747 107335 1755 107369
rect 1705 107311 1755 107335
rect 216911 107369 216961 107393
rect 216911 107335 216919 107369
rect 216953 107335 216961 107369
rect 216911 107311 216961 107335
rect 1705 107033 1755 107057
rect 1705 106999 1713 107033
rect 1747 106999 1755 107033
rect 1705 106975 1755 106999
rect 216911 107033 216961 107057
rect 216911 106999 216919 107033
rect 216953 106999 216961 107033
rect 216911 106975 216961 106999
rect 1705 106697 1755 106721
rect 1705 106663 1713 106697
rect 1747 106663 1755 106697
rect 1705 106639 1755 106663
rect 216911 106697 216961 106721
rect 216911 106663 216919 106697
rect 216953 106663 216961 106697
rect 216911 106639 216961 106663
rect 1705 106361 1755 106385
rect 1705 106327 1713 106361
rect 1747 106327 1755 106361
rect 1705 106303 1755 106327
rect 216911 106361 216961 106385
rect 216911 106327 216919 106361
rect 216953 106327 216961 106361
rect 216911 106303 216961 106327
rect 1705 106025 1755 106049
rect 1705 105991 1713 106025
rect 1747 105991 1755 106025
rect 1705 105967 1755 105991
rect 216911 106025 216961 106049
rect 216911 105991 216919 106025
rect 216953 105991 216961 106025
rect 216911 105967 216961 105991
rect 1705 105689 1755 105713
rect 1705 105655 1713 105689
rect 1747 105655 1755 105689
rect 1705 105631 1755 105655
rect 216911 105689 216961 105713
rect 216911 105655 216919 105689
rect 216953 105655 216961 105689
rect 216911 105631 216961 105655
rect 1705 105353 1755 105377
rect 1705 105319 1713 105353
rect 1747 105319 1755 105353
rect 1705 105295 1755 105319
rect 216911 105353 216961 105377
rect 216911 105319 216919 105353
rect 216953 105319 216961 105353
rect 216911 105295 216961 105319
rect 1705 105017 1755 105041
rect 1705 104983 1713 105017
rect 1747 104983 1755 105017
rect 1705 104959 1755 104983
rect 216911 105017 216961 105041
rect 216911 104983 216919 105017
rect 216953 104983 216961 105017
rect 216911 104959 216961 104983
rect 1705 104681 1755 104705
rect 1705 104647 1713 104681
rect 1747 104647 1755 104681
rect 1705 104623 1755 104647
rect 216911 104681 216961 104705
rect 216911 104647 216919 104681
rect 216953 104647 216961 104681
rect 216911 104623 216961 104647
rect 1705 104345 1755 104369
rect 1705 104311 1713 104345
rect 1747 104311 1755 104345
rect 1705 104287 1755 104311
rect 216911 104345 216961 104369
rect 216911 104311 216919 104345
rect 216953 104311 216961 104345
rect 216911 104287 216961 104311
rect 1705 104009 1755 104033
rect 1705 103975 1713 104009
rect 1747 103975 1755 104009
rect 1705 103951 1755 103975
rect 216911 104009 216961 104033
rect 216911 103975 216919 104009
rect 216953 103975 216961 104009
rect 216911 103951 216961 103975
rect 1705 103673 1755 103697
rect 1705 103639 1713 103673
rect 1747 103639 1755 103673
rect 1705 103615 1755 103639
rect 216911 103673 216961 103697
rect 216911 103639 216919 103673
rect 216953 103639 216961 103673
rect 216911 103615 216961 103639
rect 1705 103337 1755 103361
rect 1705 103303 1713 103337
rect 1747 103303 1755 103337
rect 1705 103279 1755 103303
rect 216911 103337 216961 103361
rect 216911 103303 216919 103337
rect 216953 103303 216961 103337
rect 216911 103279 216961 103303
rect 1705 103001 1755 103025
rect 1705 102967 1713 103001
rect 1747 102967 1755 103001
rect 1705 102943 1755 102967
rect 216911 103001 216961 103025
rect 216911 102967 216919 103001
rect 216953 102967 216961 103001
rect 216911 102943 216961 102967
rect 1705 102665 1755 102689
rect 1705 102631 1713 102665
rect 1747 102631 1755 102665
rect 1705 102607 1755 102631
rect 216911 102665 216961 102689
rect 216911 102631 216919 102665
rect 216953 102631 216961 102665
rect 216911 102607 216961 102631
rect 1705 102329 1755 102353
rect 1705 102295 1713 102329
rect 1747 102295 1755 102329
rect 1705 102271 1755 102295
rect 216911 102329 216961 102353
rect 216911 102295 216919 102329
rect 216953 102295 216961 102329
rect 216911 102271 216961 102295
rect 1705 101993 1755 102017
rect 1705 101959 1713 101993
rect 1747 101959 1755 101993
rect 1705 101935 1755 101959
rect 216911 101993 216961 102017
rect 216911 101959 216919 101993
rect 216953 101959 216961 101993
rect 216911 101935 216961 101959
rect 1705 101657 1755 101681
rect 1705 101623 1713 101657
rect 1747 101623 1755 101657
rect 1705 101599 1755 101623
rect 216911 101657 216961 101681
rect 216911 101623 216919 101657
rect 216953 101623 216961 101657
rect 216911 101599 216961 101623
rect 1705 101321 1755 101345
rect 1705 101287 1713 101321
rect 1747 101287 1755 101321
rect 1705 101263 1755 101287
rect 216911 101321 216961 101345
rect 216911 101287 216919 101321
rect 216953 101287 216961 101321
rect 216911 101263 216961 101287
rect 1705 100985 1755 101009
rect 1705 100951 1713 100985
rect 1747 100951 1755 100985
rect 1705 100927 1755 100951
rect 216911 100985 216961 101009
rect 216911 100951 216919 100985
rect 216953 100951 216961 100985
rect 216911 100927 216961 100951
rect 1705 100649 1755 100673
rect 1705 100615 1713 100649
rect 1747 100615 1755 100649
rect 1705 100591 1755 100615
rect 216911 100649 216961 100673
rect 216911 100615 216919 100649
rect 216953 100615 216961 100649
rect 216911 100591 216961 100615
rect 1705 100313 1755 100337
rect 1705 100279 1713 100313
rect 1747 100279 1755 100313
rect 1705 100255 1755 100279
rect 216911 100313 216961 100337
rect 216911 100279 216919 100313
rect 216953 100279 216961 100313
rect 216911 100255 216961 100279
rect 1705 99977 1755 100001
rect 1705 99943 1713 99977
rect 1747 99943 1755 99977
rect 1705 99919 1755 99943
rect 216911 99977 216961 100001
rect 216911 99943 216919 99977
rect 216953 99943 216961 99977
rect 216911 99919 216961 99943
rect 1705 99641 1755 99665
rect 1705 99607 1713 99641
rect 1747 99607 1755 99641
rect 1705 99583 1755 99607
rect 216911 99641 216961 99665
rect 216911 99607 216919 99641
rect 216953 99607 216961 99641
rect 216911 99583 216961 99607
rect 1705 99305 1755 99329
rect 1705 99271 1713 99305
rect 1747 99271 1755 99305
rect 1705 99247 1755 99271
rect 216911 99305 216961 99329
rect 216911 99271 216919 99305
rect 216953 99271 216961 99305
rect 216911 99247 216961 99271
rect 1705 98969 1755 98993
rect 1705 98935 1713 98969
rect 1747 98935 1755 98969
rect 1705 98911 1755 98935
rect 216911 98969 216961 98993
rect 216911 98935 216919 98969
rect 216953 98935 216961 98969
rect 216911 98911 216961 98935
rect 1705 98633 1755 98657
rect 1705 98599 1713 98633
rect 1747 98599 1755 98633
rect 1705 98575 1755 98599
rect 216911 98633 216961 98657
rect 216911 98599 216919 98633
rect 216953 98599 216961 98633
rect 216911 98575 216961 98599
rect 1705 98297 1755 98321
rect 1705 98263 1713 98297
rect 1747 98263 1755 98297
rect 1705 98239 1755 98263
rect 216911 98297 216961 98321
rect 216911 98263 216919 98297
rect 216953 98263 216961 98297
rect 216911 98239 216961 98263
rect 1705 97961 1755 97985
rect 1705 97927 1713 97961
rect 1747 97927 1755 97961
rect 1705 97903 1755 97927
rect 216911 97961 216961 97985
rect 216911 97927 216919 97961
rect 216953 97927 216961 97961
rect 216911 97903 216961 97927
rect 1705 97625 1755 97649
rect 1705 97591 1713 97625
rect 1747 97591 1755 97625
rect 1705 97567 1755 97591
rect 216911 97625 216961 97649
rect 216911 97591 216919 97625
rect 216953 97591 216961 97625
rect 216911 97567 216961 97591
rect 1705 97289 1755 97313
rect 1705 97255 1713 97289
rect 1747 97255 1755 97289
rect 1705 97231 1755 97255
rect 216911 97289 216961 97313
rect 216911 97255 216919 97289
rect 216953 97255 216961 97289
rect 216911 97231 216961 97255
rect 1705 96953 1755 96977
rect 1705 96919 1713 96953
rect 1747 96919 1755 96953
rect 1705 96895 1755 96919
rect 216911 96953 216961 96977
rect 216911 96919 216919 96953
rect 216953 96919 216961 96953
rect 216911 96895 216961 96919
rect 1705 96617 1755 96641
rect 1705 96583 1713 96617
rect 1747 96583 1755 96617
rect 1705 96559 1755 96583
rect 216911 96617 216961 96641
rect 216911 96583 216919 96617
rect 216953 96583 216961 96617
rect 216911 96559 216961 96583
rect 1705 96281 1755 96305
rect 1705 96247 1713 96281
rect 1747 96247 1755 96281
rect 1705 96223 1755 96247
rect 216911 96281 216961 96305
rect 216911 96247 216919 96281
rect 216953 96247 216961 96281
rect 216911 96223 216961 96247
rect 1705 95945 1755 95969
rect 1705 95911 1713 95945
rect 1747 95911 1755 95945
rect 1705 95887 1755 95911
rect 216911 95945 216961 95969
rect 216911 95911 216919 95945
rect 216953 95911 216961 95945
rect 216911 95887 216961 95911
rect 1705 95609 1755 95633
rect 1705 95575 1713 95609
rect 1747 95575 1755 95609
rect 1705 95551 1755 95575
rect 216911 95609 216961 95633
rect 216911 95575 216919 95609
rect 216953 95575 216961 95609
rect 216911 95551 216961 95575
rect 1705 95273 1755 95297
rect 1705 95239 1713 95273
rect 1747 95239 1755 95273
rect 1705 95215 1755 95239
rect 216911 95273 216961 95297
rect 216911 95239 216919 95273
rect 216953 95239 216961 95273
rect 216911 95215 216961 95239
rect 1705 94937 1755 94961
rect 1705 94903 1713 94937
rect 1747 94903 1755 94937
rect 1705 94879 1755 94903
rect 216911 94937 216961 94961
rect 216911 94903 216919 94937
rect 216953 94903 216961 94937
rect 216911 94879 216961 94903
rect 1705 94601 1755 94625
rect 1705 94567 1713 94601
rect 1747 94567 1755 94601
rect 1705 94543 1755 94567
rect 216911 94601 216961 94625
rect 216911 94567 216919 94601
rect 216953 94567 216961 94601
rect 216911 94543 216961 94567
rect 1705 94265 1755 94289
rect 1705 94231 1713 94265
rect 1747 94231 1755 94265
rect 1705 94207 1755 94231
rect 216911 94265 216961 94289
rect 216911 94231 216919 94265
rect 216953 94231 216961 94265
rect 216911 94207 216961 94231
rect 1705 93929 1755 93953
rect 1705 93895 1713 93929
rect 1747 93895 1755 93929
rect 1705 93871 1755 93895
rect 216911 93929 216961 93953
rect 216911 93895 216919 93929
rect 216953 93895 216961 93929
rect 216911 93871 216961 93895
rect 1705 93593 1755 93617
rect 1705 93559 1713 93593
rect 1747 93559 1755 93593
rect 1705 93535 1755 93559
rect 216911 93593 216961 93617
rect 216911 93559 216919 93593
rect 216953 93559 216961 93593
rect 216911 93535 216961 93559
rect 1705 93257 1755 93281
rect 1705 93223 1713 93257
rect 1747 93223 1755 93257
rect 1705 93199 1755 93223
rect 216911 93257 216961 93281
rect 216911 93223 216919 93257
rect 216953 93223 216961 93257
rect 216911 93199 216961 93223
rect 1705 92921 1755 92945
rect 1705 92887 1713 92921
rect 1747 92887 1755 92921
rect 1705 92863 1755 92887
rect 216911 92921 216961 92945
rect 216911 92887 216919 92921
rect 216953 92887 216961 92921
rect 216911 92863 216961 92887
rect 1705 92585 1755 92609
rect 1705 92551 1713 92585
rect 1747 92551 1755 92585
rect 1705 92527 1755 92551
rect 216911 92585 216961 92609
rect 216911 92551 216919 92585
rect 216953 92551 216961 92585
rect 216911 92527 216961 92551
rect 1705 92249 1755 92273
rect 1705 92215 1713 92249
rect 1747 92215 1755 92249
rect 1705 92191 1755 92215
rect 216911 92249 216961 92273
rect 216911 92215 216919 92249
rect 216953 92215 216961 92249
rect 216911 92191 216961 92215
rect 1705 91913 1755 91937
rect 1705 91879 1713 91913
rect 1747 91879 1755 91913
rect 1705 91855 1755 91879
rect 216911 91913 216961 91937
rect 216911 91879 216919 91913
rect 216953 91879 216961 91913
rect 216911 91855 216961 91879
rect 1705 91577 1755 91601
rect 1705 91543 1713 91577
rect 1747 91543 1755 91577
rect 1705 91519 1755 91543
rect 216911 91577 216961 91601
rect 216911 91543 216919 91577
rect 216953 91543 216961 91577
rect 216911 91519 216961 91543
rect 1705 91241 1755 91265
rect 1705 91207 1713 91241
rect 1747 91207 1755 91241
rect 1705 91183 1755 91207
rect 216911 91241 216961 91265
rect 216911 91207 216919 91241
rect 216953 91207 216961 91241
rect 216911 91183 216961 91207
rect 1705 90905 1755 90929
rect 1705 90871 1713 90905
rect 1747 90871 1755 90905
rect 1705 90847 1755 90871
rect 216911 90905 216961 90929
rect 216911 90871 216919 90905
rect 216953 90871 216961 90905
rect 216911 90847 216961 90871
rect 1705 90569 1755 90593
rect 1705 90535 1713 90569
rect 1747 90535 1755 90569
rect 1705 90511 1755 90535
rect 216911 90569 216961 90593
rect 216911 90535 216919 90569
rect 216953 90535 216961 90569
rect 216911 90511 216961 90535
rect 1705 90233 1755 90257
rect 1705 90199 1713 90233
rect 1747 90199 1755 90233
rect 1705 90175 1755 90199
rect 216911 90233 216961 90257
rect 216911 90199 216919 90233
rect 216953 90199 216961 90233
rect 216911 90175 216961 90199
rect 1705 89897 1755 89921
rect 1705 89863 1713 89897
rect 1747 89863 1755 89897
rect 1705 89839 1755 89863
rect 216911 89897 216961 89921
rect 216911 89863 216919 89897
rect 216953 89863 216961 89897
rect 216911 89839 216961 89863
rect 1705 89561 1755 89585
rect 1705 89527 1713 89561
rect 1747 89527 1755 89561
rect 1705 89503 1755 89527
rect 216911 89561 216961 89585
rect 216911 89527 216919 89561
rect 216953 89527 216961 89561
rect 216911 89503 216961 89527
rect 1705 89225 1755 89249
rect 1705 89191 1713 89225
rect 1747 89191 1755 89225
rect 1705 89167 1755 89191
rect 216911 89225 216961 89249
rect 216911 89191 216919 89225
rect 216953 89191 216961 89225
rect 216911 89167 216961 89191
rect 1705 88889 1755 88913
rect 1705 88855 1713 88889
rect 1747 88855 1755 88889
rect 1705 88831 1755 88855
rect 216911 88889 216961 88913
rect 216911 88855 216919 88889
rect 216953 88855 216961 88889
rect 216911 88831 216961 88855
rect 1705 88553 1755 88577
rect 1705 88519 1713 88553
rect 1747 88519 1755 88553
rect 1705 88495 1755 88519
rect 216911 88553 216961 88577
rect 216911 88519 216919 88553
rect 216953 88519 216961 88553
rect 216911 88495 216961 88519
rect 1705 88217 1755 88241
rect 1705 88183 1713 88217
rect 1747 88183 1755 88217
rect 1705 88159 1755 88183
rect 216911 88217 216961 88241
rect 216911 88183 216919 88217
rect 216953 88183 216961 88217
rect 216911 88159 216961 88183
rect 1705 87881 1755 87905
rect 1705 87847 1713 87881
rect 1747 87847 1755 87881
rect 1705 87823 1755 87847
rect 216911 87881 216961 87905
rect 216911 87847 216919 87881
rect 216953 87847 216961 87881
rect 216911 87823 216961 87847
rect 1705 87545 1755 87569
rect 1705 87511 1713 87545
rect 1747 87511 1755 87545
rect 1705 87487 1755 87511
rect 216911 87545 216961 87569
rect 216911 87511 216919 87545
rect 216953 87511 216961 87545
rect 216911 87487 216961 87511
rect 1705 87209 1755 87233
rect 1705 87175 1713 87209
rect 1747 87175 1755 87209
rect 1705 87151 1755 87175
rect 216911 87209 216961 87233
rect 216911 87175 216919 87209
rect 216953 87175 216961 87209
rect 216911 87151 216961 87175
rect 1705 86873 1755 86897
rect 1705 86839 1713 86873
rect 1747 86839 1755 86873
rect 1705 86815 1755 86839
rect 216911 86873 216961 86897
rect 216911 86839 216919 86873
rect 216953 86839 216961 86873
rect 216911 86815 216961 86839
rect 1705 86537 1755 86561
rect 1705 86503 1713 86537
rect 1747 86503 1755 86537
rect 1705 86479 1755 86503
rect 216911 86537 216961 86561
rect 216911 86503 216919 86537
rect 216953 86503 216961 86537
rect 216911 86479 216961 86503
rect 1705 86201 1755 86225
rect 1705 86167 1713 86201
rect 1747 86167 1755 86201
rect 1705 86143 1755 86167
rect 216911 86201 216961 86225
rect 216911 86167 216919 86201
rect 216953 86167 216961 86201
rect 216911 86143 216961 86167
rect 1705 85865 1755 85889
rect 1705 85831 1713 85865
rect 1747 85831 1755 85865
rect 1705 85807 1755 85831
rect 216911 85865 216961 85889
rect 216911 85831 216919 85865
rect 216953 85831 216961 85865
rect 216911 85807 216961 85831
rect 1705 85529 1755 85553
rect 1705 85495 1713 85529
rect 1747 85495 1755 85529
rect 1705 85471 1755 85495
rect 216911 85529 216961 85553
rect 216911 85495 216919 85529
rect 216953 85495 216961 85529
rect 216911 85471 216961 85495
rect 1705 85193 1755 85217
rect 1705 85159 1713 85193
rect 1747 85159 1755 85193
rect 1705 85135 1755 85159
rect 216911 85193 216961 85217
rect 216911 85159 216919 85193
rect 216953 85159 216961 85193
rect 216911 85135 216961 85159
rect 1705 84857 1755 84881
rect 1705 84823 1713 84857
rect 1747 84823 1755 84857
rect 1705 84799 1755 84823
rect 216911 84857 216961 84881
rect 216911 84823 216919 84857
rect 216953 84823 216961 84857
rect 216911 84799 216961 84823
rect 1705 84521 1755 84545
rect 1705 84487 1713 84521
rect 1747 84487 1755 84521
rect 1705 84463 1755 84487
rect 216911 84521 216961 84545
rect 216911 84487 216919 84521
rect 216953 84487 216961 84521
rect 216911 84463 216961 84487
rect 1705 84185 1755 84209
rect 1705 84151 1713 84185
rect 1747 84151 1755 84185
rect 1705 84127 1755 84151
rect 216911 84185 216961 84209
rect 216911 84151 216919 84185
rect 216953 84151 216961 84185
rect 216911 84127 216961 84151
rect 1705 83849 1755 83873
rect 1705 83815 1713 83849
rect 1747 83815 1755 83849
rect 1705 83791 1755 83815
rect 216911 83849 216961 83873
rect 216911 83815 216919 83849
rect 216953 83815 216961 83849
rect 216911 83791 216961 83815
rect 1705 83513 1755 83537
rect 1705 83479 1713 83513
rect 1747 83479 1755 83513
rect 1705 83455 1755 83479
rect 216911 83513 216961 83537
rect 216911 83479 216919 83513
rect 216953 83479 216961 83513
rect 216911 83455 216961 83479
rect 1705 83177 1755 83201
rect 1705 83143 1713 83177
rect 1747 83143 1755 83177
rect 1705 83119 1755 83143
rect 216911 83177 216961 83201
rect 216911 83143 216919 83177
rect 216953 83143 216961 83177
rect 216911 83119 216961 83143
rect 1705 82841 1755 82865
rect 1705 82807 1713 82841
rect 1747 82807 1755 82841
rect 1705 82783 1755 82807
rect 216911 82841 216961 82865
rect 216911 82807 216919 82841
rect 216953 82807 216961 82841
rect 216911 82783 216961 82807
rect 1705 82505 1755 82529
rect 1705 82471 1713 82505
rect 1747 82471 1755 82505
rect 1705 82447 1755 82471
rect 216911 82505 216961 82529
rect 216911 82471 216919 82505
rect 216953 82471 216961 82505
rect 216911 82447 216961 82471
rect 1705 82169 1755 82193
rect 1705 82135 1713 82169
rect 1747 82135 1755 82169
rect 1705 82111 1755 82135
rect 216911 82169 216961 82193
rect 216911 82135 216919 82169
rect 216953 82135 216961 82169
rect 216911 82111 216961 82135
rect 1705 81833 1755 81857
rect 1705 81799 1713 81833
rect 1747 81799 1755 81833
rect 1705 81775 1755 81799
rect 216911 81833 216961 81857
rect 216911 81799 216919 81833
rect 216953 81799 216961 81833
rect 216911 81775 216961 81799
rect 1705 81497 1755 81521
rect 1705 81463 1713 81497
rect 1747 81463 1755 81497
rect 1705 81439 1755 81463
rect 216911 81497 216961 81521
rect 216911 81463 216919 81497
rect 216953 81463 216961 81497
rect 216911 81439 216961 81463
rect 1705 81161 1755 81185
rect 1705 81127 1713 81161
rect 1747 81127 1755 81161
rect 1705 81103 1755 81127
rect 216911 81161 216961 81185
rect 216911 81127 216919 81161
rect 216953 81127 216961 81161
rect 216911 81103 216961 81127
rect 1705 80825 1755 80849
rect 1705 80791 1713 80825
rect 1747 80791 1755 80825
rect 1705 80767 1755 80791
rect 216911 80825 216961 80849
rect 216911 80791 216919 80825
rect 216953 80791 216961 80825
rect 216911 80767 216961 80791
rect 1705 80489 1755 80513
rect 1705 80455 1713 80489
rect 1747 80455 1755 80489
rect 1705 80431 1755 80455
rect 216911 80489 216961 80513
rect 216911 80455 216919 80489
rect 216953 80455 216961 80489
rect 216911 80431 216961 80455
rect 1705 80153 1755 80177
rect 1705 80119 1713 80153
rect 1747 80119 1755 80153
rect 1705 80095 1755 80119
rect 216911 80153 216961 80177
rect 216911 80119 216919 80153
rect 216953 80119 216961 80153
rect 216911 80095 216961 80119
rect 1705 79817 1755 79841
rect 1705 79783 1713 79817
rect 1747 79783 1755 79817
rect 1705 79759 1755 79783
rect 216911 79817 216961 79841
rect 216911 79783 216919 79817
rect 216953 79783 216961 79817
rect 216911 79759 216961 79783
rect 1705 79481 1755 79505
rect 1705 79447 1713 79481
rect 1747 79447 1755 79481
rect 1705 79423 1755 79447
rect 216911 79481 216961 79505
rect 216911 79447 216919 79481
rect 216953 79447 216961 79481
rect 216911 79423 216961 79447
rect 1705 79145 1755 79169
rect 1705 79111 1713 79145
rect 1747 79111 1755 79145
rect 1705 79087 1755 79111
rect 216911 79145 216961 79169
rect 216911 79111 216919 79145
rect 216953 79111 216961 79145
rect 216911 79087 216961 79111
rect 1705 78809 1755 78833
rect 1705 78775 1713 78809
rect 1747 78775 1755 78809
rect 1705 78751 1755 78775
rect 216911 78809 216961 78833
rect 216911 78775 216919 78809
rect 216953 78775 216961 78809
rect 216911 78751 216961 78775
rect 1705 78473 1755 78497
rect 1705 78439 1713 78473
rect 1747 78439 1755 78473
rect 1705 78415 1755 78439
rect 216911 78473 216961 78497
rect 216911 78439 216919 78473
rect 216953 78439 216961 78473
rect 216911 78415 216961 78439
rect 1705 78137 1755 78161
rect 1705 78103 1713 78137
rect 1747 78103 1755 78137
rect 1705 78079 1755 78103
rect 216911 78137 216961 78161
rect 216911 78103 216919 78137
rect 216953 78103 216961 78137
rect 216911 78079 216961 78103
rect 1705 77801 1755 77825
rect 1705 77767 1713 77801
rect 1747 77767 1755 77801
rect 1705 77743 1755 77767
rect 216911 77801 216961 77825
rect 216911 77767 216919 77801
rect 216953 77767 216961 77801
rect 216911 77743 216961 77767
rect 1705 77465 1755 77489
rect 1705 77431 1713 77465
rect 1747 77431 1755 77465
rect 1705 77407 1755 77431
rect 216911 77465 216961 77489
rect 216911 77431 216919 77465
rect 216953 77431 216961 77465
rect 216911 77407 216961 77431
rect 1705 77129 1755 77153
rect 1705 77095 1713 77129
rect 1747 77095 1755 77129
rect 1705 77071 1755 77095
rect 216911 77129 216961 77153
rect 216911 77095 216919 77129
rect 216953 77095 216961 77129
rect 216911 77071 216961 77095
rect 1705 76793 1755 76817
rect 1705 76759 1713 76793
rect 1747 76759 1755 76793
rect 1705 76735 1755 76759
rect 216911 76793 216961 76817
rect 216911 76759 216919 76793
rect 216953 76759 216961 76793
rect 216911 76735 216961 76759
rect 1705 76457 1755 76481
rect 1705 76423 1713 76457
rect 1747 76423 1755 76457
rect 1705 76399 1755 76423
rect 216911 76457 216961 76481
rect 216911 76423 216919 76457
rect 216953 76423 216961 76457
rect 216911 76399 216961 76423
rect 1705 76121 1755 76145
rect 1705 76087 1713 76121
rect 1747 76087 1755 76121
rect 1705 76063 1755 76087
rect 216911 76121 216961 76145
rect 216911 76087 216919 76121
rect 216953 76087 216961 76121
rect 216911 76063 216961 76087
rect 1705 75785 1755 75809
rect 1705 75751 1713 75785
rect 1747 75751 1755 75785
rect 1705 75727 1755 75751
rect 216911 75785 216961 75809
rect 216911 75751 216919 75785
rect 216953 75751 216961 75785
rect 216911 75727 216961 75751
rect 1705 75449 1755 75473
rect 1705 75415 1713 75449
rect 1747 75415 1755 75449
rect 1705 75391 1755 75415
rect 216911 75449 216961 75473
rect 216911 75415 216919 75449
rect 216953 75415 216961 75449
rect 216911 75391 216961 75415
rect 1705 75113 1755 75137
rect 1705 75079 1713 75113
rect 1747 75079 1755 75113
rect 1705 75055 1755 75079
rect 216911 75113 216961 75137
rect 216911 75079 216919 75113
rect 216953 75079 216961 75113
rect 216911 75055 216961 75079
rect 1705 74777 1755 74801
rect 1705 74743 1713 74777
rect 1747 74743 1755 74777
rect 1705 74719 1755 74743
rect 216911 74777 216961 74801
rect 216911 74743 216919 74777
rect 216953 74743 216961 74777
rect 216911 74719 216961 74743
rect 1705 74441 1755 74465
rect 1705 74407 1713 74441
rect 1747 74407 1755 74441
rect 1705 74383 1755 74407
rect 216911 74441 216961 74465
rect 216911 74407 216919 74441
rect 216953 74407 216961 74441
rect 216911 74383 216961 74407
rect 1705 74105 1755 74129
rect 1705 74071 1713 74105
rect 1747 74071 1755 74105
rect 1705 74047 1755 74071
rect 216911 74105 216961 74129
rect 216911 74071 216919 74105
rect 216953 74071 216961 74105
rect 216911 74047 216961 74071
rect 1705 73769 1755 73793
rect 1705 73735 1713 73769
rect 1747 73735 1755 73769
rect 1705 73711 1755 73735
rect 216911 73769 216961 73793
rect 216911 73735 216919 73769
rect 216953 73735 216961 73769
rect 216911 73711 216961 73735
rect 1705 73433 1755 73457
rect 1705 73399 1713 73433
rect 1747 73399 1755 73433
rect 1705 73375 1755 73399
rect 216911 73433 216961 73457
rect 216911 73399 216919 73433
rect 216953 73399 216961 73433
rect 216911 73375 216961 73399
rect 1705 73097 1755 73121
rect 1705 73063 1713 73097
rect 1747 73063 1755 73097
rect 1705 73039 1755 73063
rect 216911 73097 216961 73121
rect 216911 73063 216919 73097
rect 216953 73063 216961 73097
rect 216911 73039 216961 73063
rect 1705 72761 1755 72785
rect 1705 72727 1713 72761
rect 1747 72727 1755 72761
rect 1705 72703 1755 72727
rect 216911 72761 216961 72785
rect 216911 72727 216919 72761
rect 216953 72727 216961 72761
rect 216911 72703 216961 72727
rect 1705 72425 1755 72449
rect 1705 72391 1713 72425
rect 1747 72391 1755 72425
rect 1705 72367 1755 72391
rect 216911 72425 216961 72449
rect 216911 72391 216919 72425
rect 216953 72391 216961 72425
rect 216911 72367 216961 72391
rect 1705 72089 1755 72113
rect 1705 72055 1713 72089
rect 1747 72055 1755 72089
rect 1705 72031 1755 72055
rect 216911 72089 216961 72113
rect 216911 72055 216919 72089
rect 216953 72055 216961 72089
rect 216911 72031 216961 72055
rect 1705 71753 1755 71777
rect 1705 71719 1713 71753
rect 1747 71719 1755 71753
rect 1705 71695 1755 71719
rect 216911 71753 216961 71777
rect 216911 71719 216919 71753
rect 216953 71719 216961 71753
rect 216911 71695 216961 71719
rect 1705 71417 1755 71441
rect 1705 71383 1713 71417
rect 1747 71383 1755 71417
rect 1705 71359 1755 71383
rect 216911 71417 216961 71441
rect 216911 71383 216919 71417
rect 216953 71383 216961 71417
rect 216911 71359 216961 71383
rect 1705 71081 1755 71105
rect 1705 71047 1713 71081
rect 1747 71047 1755 71081
rect 1705 71023 1755 71047
rect 216911 71081 216961 71105
rect 216911 71047 216919 71081
rect 216953 71047 216961 71081
rect 216911 71023 216961 71047
rect 1705 70745 1755 70769
rect 1705 70711 1713 70745
rect 1747 70711 1755 70745
rect 1705 70687 1755 70711
rect 216911 70745 216961 70769
rect 216911 70711 216919 70745
rect 216953 70711 216961 70745
rect 216911 70687 216961 70711
rect 1705 70409 1755 70433
rect 1705 70375 1713 70409
rect 1747 70375 1755 70409
rect 1705 70351 1755 70375
rect 216911 70409 216961 70433
rect 216911 70375 216919 70409
rect 216953 70375 216961 70409
rect 216911 70351 216961 70375
rect 1705 70073 1755 70097
rect 1705 70039 1713 70073
rect 1747 70039 1755 70073
rect 1705 70015 1755 70039
rect 216911 70073 216961 70097
rect 216911 70039 216919 70073
rect 216953 70039 216961 70073
rect 216911 70015 216961 70039
rect 1705 69737 1755 69761
rect 1705 69703 1713 69737
rect 1747 69703 1755 69737
rect 1705 69679 1755 69703
rect 216911 69737 216961 69761
rect 216911 69703 216919 69737
rect 216953 69703 216961 69737
rect 216911 69679 216961 69703
rect 1705 69401 1755 69425
rect 1705 69367 1713 69401
rect 1747 69367 1755 69401
rect 1705 69343 1755 69367
rect 216911 69401 216961 69425
rect 216911 69367 216919 69401
rect 216953 69367 216961 69401
rect 216911 69343 216961 69367
rect 1705 69065 1755 69089
rect 1705 69031 1713 69065
rect 1747 69031 1755 69065
rect 1705 69007 1755 69031
rect 216911 69065 216961 69089
rect 216911 69031 216919 69065
rect 216953 69031 216961 69065
rect 216911 69007 216961 69031
rect 1705 68729 1755 68753
rect 1705 68695 1713 68729
rect 1747 68695 1755 68729
rect 1705 68671 1755 68695
rect 216911 68729 216961 68753
rect 216911 68695 216919 68729
rect 216953 68695 216961 68729
rect 216911 68671 216961 68695
rect 1705 68393 1755 68417
rect 1705 68359 1713 68393
rect 1747 68359 1755 68393
rect 1705 68335 1755 68359
rect 216911 68393 216961 68417
rect 216911 68359 216919 68393
rect 216953 68359 216961 68393
rect 216911 68335 216961 68359
rect 1705 68057 1755 68081
rect 1705 68023 1713 68057
rect 1747 68023 1755 68057
rect 1705 67999 1755 68023
rect 216911 68057 216961 68081
rect 216911 68023 216919 68057
rect 216953 68023 216961 68057
rect 216911 67999 216961 68023
rect 1705 67721 1755 67745
rect 1705 67687 1713 67721
rect 1747 67687 1755 67721
rect 1705 67663 1755 67687
rect 216911 67721 216961 67745
rect 216911 67687 216919 67721
rect 216953 67687 216961 67721
rect 216911 67663 216961 67687
rect 1705 67385 1755 67409
rect 1705 67351 1713 67385
rect 1747 67351 1755 67385
rect 1705 67327 1755 67351
rect 216911 67385 216961 67409
rect 216911 67351 216919 67385
rect 216953 67351 216961 67385
rect 216911 67327 216961 67351
rect 1705 67049 1755 67073
rect 1705 67015 1713 67049
rect 1747 67015 1755 67049
rect 1705 66991 1755 67015
rect 216911 67049 216961 67073
rect 216911 67015 216919 67049
rect 216953 67015 216961 67049
rect 216911 66991 216961 67015
rect 1705 66713 1755 66737
rect 1705 66679 1713 66713
rect 1747 66679 1755 66713
rect 1705 66655 1755 66679
rect 216911 66713 216961 66737
rect 216911 66679 216919 66713
rect 216953 66679 216961 66713
rect 216911 66655 216961 66679
rect 1705 66377 1755 66401
rect 1705 66343 1713 66377
rect 1747 66343 1755 66377
rect 1705 66319 1755 66343
rect 216911 66377 216961 66401
rect 216911 66343 216919 66377
rect 216953 66343 216961 66377
rect 216911 66319 216961 66343
rect 1705 66041 1755 66065
rect 1705 66007 1713 66041
rect 1747 66007 1755 66041
rect 1705 65983 1755 66007
rect 216911 66041 216961 66065
rect 216911 66007 216919 66041
rect 216953 66007 216961 66041
rect 216911 65983 216961 66007
rect 1705 65705 1755 65729
rect 1705 65671 1713 65705
rect 1747 65671 1755 65705
rect 1705 65647 1755 65671
rect 216911 65705 216961 65729
rect 216911 65671 216919 65705
rect 216953 65671 216961 65705
rect 216911 65647 216961 65671
rect 1705 65369 1755 65393
rect 1705 65335 1713 65369
rect 1747 65335 1755 65369
rect 1705 65311 1755 65335
rect 216911 65369 216961 65393
rect 216911 65335 216919 65369
rect 216953 65335 216961 65369
rect 216911 65311 216961 65335
rect 1705 65033 1755 65057
rect 1705 64999 1713 65033
rect 1747 64999 1755 65033
rect 1705 64975 1755 64999
rect 216911 65033 216961 65057
rect 216911 64999 216919 65033
rect 216953 64999 216961 65033
rect 216911 64975 216961 64999
rect 1705 64697 1755 64721
rect 1705 64663 1713 64697
rect 1747 64663 1755 64697
rect 1705 64639 1755 64663
rect 216911 64697 216961 64721
rect 216911 64663 216919 64697
rect 216953 64663 216961 64697
rect 216911 64639 216961 64663
rect 1705 64361 1755 64385
rect 1705 64327 1713 64361
rect 1747 64327 1755 64361
rect 1705 64303 1755 64327
rect 216911 64361 216961 64385
rect 216911 64327 216919 64361
rect 216953 64327 216961 64361
rect 216911 64303 216961 64327
rect 1705 64025 1755 64049
rect 1705 63991 1713 64025
rect 1747 63991 1755 64025
rect 1705 63967 1755 63991
rect 216911 64025 216961 64049
rect 216911 63991 216919 64025
rect 216953 63991 216961 64025
rect 216911 63967 216961 63991
rect 1705 63689 1755 63713
rect 1705 63655 1713 63689
rect 1747 63655 1755 63689
rect 1705 63631 1755 63655
rect 216911 63689 216961 63713
rect 216911 63655 216919 63689
rect 216953 63655 216961 63689
rect 216911 63631 216961 63655
rect 1705 63353 1755 63377
rect 1705 63319 1713 63353
rect 1747 63319 1755 63353
rect 1705 63295 1755 63319
rect 216911 63353 216961 63377
rect 216911 63319 216919 63353
rect 216953 63319 216961 63353
rect 216911 63295 216961 63319
rect 1705 63017 1755 63041
rect 1705 62983 1713 63017
rect 1747 62983 1755 63017
rect 1705 62959 1755 62983
rect 216911 63017 216961 63041
rect 216911 62983 216919 63017
rect 216953 62983 216961 63017
rect 216911 62959 216961 62983
rect 1705 62681 1755 62705
rect 1705 62647 1713 62681
rect 1747 62647 1755 62681
rect 1705 62623 1755 62647
rect 216911 62681 216961 62705
rect 216911 62647 216919 62681
rect 216953 62647 216961 62681
rect 216911 62623 216961 62647
rect 1705 62345 1755 62369
rect 1705 62311 1713 62345
rect 1747 62311 1755 62345
rect 1705 62287 1755 62311
rect 216911 62345 216961 62369
rect 216911 62311 216919 62345
rect 216953 62311 216961 62345
rect 216911 62287 216961 62311
rect 1705 62009 1755 62033
rect 1705 61975 1713 62009
rect 1747 61975 1755 62009
rect 1705 61951 1755 61975
rect 216911 62009 216961 62033
rect 216911 61975 216919 62009
rect 216953 61975 216961 62009
rect 216911 61951 216961 61975
rect 1705 61673 1755 61697
rect 1705 61639 1713 61673
rect 1747 61639 1755 61673
rect 1705 61615 1755 61639
rect 216911 61673 216961 61697
rect 216911 61639 216919 61673
rect 216953 61639 216961 61673
rect 216911 61615 216961 61639
rect 1705 61337 1755 61361
rect 1705 61303 1713 61337
rect 1747 61303 1755 61337
rect 1705 61279 1755 61303
rect 216911 61337 216961 61361
rect 216911 61303 216919 61337
rect 216953 61303 216961 61337
rect 216911 61279 216961 61303
rect 1705 61001 1755 61025
rect 1705 60967 1713 61001
rect 1747 60967 1755 61001
rect 1705 60943 1755 60967
rect 216911 61001 216961 61025
rect 216911 60967 216919 61001
rect 216953 60967 216961 61001
rect 216911 60943 216961 60967
rect 1705 60665 1755 60689
rect 1705 60631 1713 60665
rect 1747 60631 1755 60665
rect 1705 60607 1755 60631
rect 216911 60665 216961 60689
rect 216911 60631 216919 60665
rect 216953 60631 216961 60665
rect 216911 60607 216961 60631
rect 1705 60329 1755 60353
rect 1705 60295 1713 60329
rect 1747 60295 1755 60329
rect 1705 60271 1755 60295
rect 216911 60329 216961 60353
rect 216911 60295 216919 60329
rect 216953 60295 216961 60329
rect 216911 60271 216961 60295
rect 1705 59993 1755 60017
rect 1705 59959 1713 59993
rect 1747 59959 1755 59993
rect 1705 59935 1755 59959
rect 216911 59993 216961 60017
rect 216911 59959 216919 59993
rect 216953 59959 216961 59993
rect 216911 59935 216961 59959
rect 1705 59657 1755 59681
rect 1705 59623 1713 59657
rect 1747 59623 1755 59657
rect 1705 59599 1755 59623
rect 216911 59657 216961 59681
rect 216911 59623 216919 59657
rect 216953 59623 216961 59657
rect 216911 59599 216961 59623
rect 1705 59321 1755 59345
rect 1705 59287 1713 59321
rect 1747 59287 1755 59321
rect 1705 59263 1755 59287
rect 216911 59321 216961 59345
rect 216911 59287 216919 59321
rect 216953 59287 216961 59321
rect 216911 59263 216961 59287
rect 1705 58985 1755 59009
rect 1705 58951 1713 58985
rect 1747 58951 1755 58985
rect 1705 58927 1755 58951
rect 216911 58985 216961 59009
rect 216911 58951 216919 58985
rect 216953 58951 216961 58985
rect 216911 58927 216961 58951
rect 1705 58649 1755 58673
rect 1705 58615 1713 58649
rect 1747 58615 1755 58649
rect 1705 58591 1755 58615
rect 216911 58649 216961 58673
rect 216911 58615 216919 58649
rect 216953 58615 216961 58649
rect 216911 58591 216961 58615
rect 1705 58313 1755 58337
rect 1705 58279 1713 58313
rect 1747 58279 1755 58313
rect 1705 58255 1755 58279
rect 216911 58313 216961 58337
rect 216911 58279 216919 58313
rect 216953 58279 216961 58313
rect 216911 58255 216961 58279
rect 1705 57977 1755 58001
rect 1705 57943 1713 57977
rect 1747 57943 1755 57977
rect 1705 57919 1755 57943
rect 216911 57977 216961 58001
rect 216911 57943 216919 57977
rect 216953 57943 216961 57977
rect 216911 57919 216961 57943
rect 1705 57641 1755 57665
rect 1705 57607 1713 57641
rect 1747 57607 1755 57641
rect 1705 57583 1755 57607
rect 216911 57641 216961 57665
rect 216911 57607 216919 57641
rect 216953 57607 216961 57641
rect 216911 57583 216961 57607
rect 1705 57305 1755 57329
rect 1705 57271 1713 57305
rect 1747 57271 1755 57305
rect 1705 57247 1755 57271
rect 216911 57305 216961 57329
rect 216911 57271 216919 57305
rect 216953 57271 216961 57305
rect 216911 57247 216961 57271
rect 1705 56969 1755 56993
rect 1705 56935 1713 56969
rect 1747 56935 1755 56969
rect 1705 56911 1755 56935
rect 216911 56969 216961 56993
rect 216911 56935 216919 56969
rect 216953 56935 216961 56969
rect 216911 56911 216961 56935
rect 1705 56633 1755 56657
rect 1705 56599 1713 56633
rect 1747 56599 1755 56633
rect 1705 56575 1755 56599
rect 216911 56633 216961 56657
rect 216911 56599 216919 56633
rect 216953 56599 216961 56633
rect 216911 56575 216961 56599
rect 1705 56297 1755 56321
rect 1705 56263 1713 56297
rect 1747 56263 1755 56297
rect 1705 56239 1755 56263
rect 216911 56297 216961 56321
rect 216911 56263 216919 56297
rect 216953 56263 216961 56297
rect 216911 56239 216961 56263
rect 1705 55961 1755 55985
rect 1705 55927 1713 55961
rect 1747 55927 1755 55961
rect 1705 55903 1755 55927
rect 216911 55961 216961 55985
rect 216911 55927 216919 55961
rect 216953 55927 216961 55961
rect 216911 55903 216961 55927
rect 1705 55625 1755 55649
rect 1705 55591 1713 55625
rect 1747 55591 1755 55625
rect 1705 55567 1755 55591
rect 216911 55625 216961 55649
rect 216911 55591 216919 55625
rect 216953 55591 216961 55625
rect 216911 55567 216961 55591
rect 1705 55289 1755 55313
rect 1705 55255 1713 55289
rect 1747 55255 1755 55289
rect 1705 55231 1755 55255
rect 216911 55289 216961 55313
rect 216911 55255 216919 55289
rect 216953 55255 216961 55289
rect 216911 55231 216961 55255
rect 1705 54953 1755 54977
rect 1705 54919 1713 54953
rect 1747 54919 1755 54953
rect 1705 54895 1755 54919
rect 216911 54953 216961 54977
rect 216911 54919 216919 54953
rect 216953 54919 216961 54953
rect 216911 54895 216961 54919
rect 1705 54617 1755 54641
rect 1705 54583 1713 54617
rect 1747 54583 1755 54617
rect 1705 54559 1755 54583
rect 216911 54617 216961 54641
rect 216911 54583 216919 54617
rect 216953 54583 216961 54617
rect 216911 54559 216961 54583
rect 1705 54281 1755 54305
rect 1705 54247 1713 54281
rect 1747 54247 1755 54281
rect 1705 54223 1755 54247
rect 216911 54281 216961 54305
rect 216911 54247 216919 54281
rect 216953 54247 216961 54281
rect 216911 54223 216961 54247
rect 1705 53945 1755 53969
rect 1705 53911 1713 53945
rect 1747 53911 1755 53945
rect 1705 53887 1755 53911
rect 216911 53945 216961 53969
rect 216911 53911 216919 53945
rect 216953 53911 216961 53945
rect 216911 53887 216961 53911
rect 1705 53609 1755 53633
rect 1705 53575 1713 53609
rect 1747 53575 1755 53609
rect 1705 53551 1755 53575
rect 216911 53609 216961 53633
rect 216911 53575 216919 53609
rect 216953 53575 216961 53609
rect 216911 53551 216961 53575
rect 1705 53273 1755 53297
rect 1705 53239 1713 53273
rect 1747 53239 1755 53273
rect 1705 53215 1755 53239
rect 216911 53273 216961 53297
rect 216911 53239 216919 53273
rect 216953 53239 216961 53273
rect 216911 53215 216961 53239
rect 1705 52937 1755 52961
rect 1705 52903 1713 52937
rect 1747 52903 1755 52937
rect 1705 52879 1755 52903
rect 216911 52937 216961 52961
rect 216911 52903 216919 52937
rect 216953 52903 216961 52937
rect 216911 52879 216961 52903
rect 1705 52601 1755 52625
rect 1705 52567 1713 52601
rect 1747 52567 1755 52601
rect 1705 52543 1755 52567
rect 216911 52601 216961 52625
rect 216911 52567 216919 52601
rect 216953 52567 216961 52601
rect 216911 52543 216961 52567
rect 1705 52265 1755 52289
rect 1705 52231 1713 52265
rect 1747 52231 1755 52265
rect 1705 52207 1755 52231
rect 216911 52265 216961 52289
rect 216911 52231 216919 52265
rect 216953 52231 216961 52265
rect 216911 52207 216961 52231
rect 1705 51929 1755 51953
rect 1705 51895 1713 51929
rect 1747 51895 1755 51929
rect 1705 51871 1755 51895
rect 216911 51929 216961 51953
rect 216911 51895 216919 51929
rect 216953 51895 216961 51929
rect 216911 51871 216961 51895
rect 1705 51593 1755 51617
rect 1705 51559 1713 51593
rect 1747 51559 1755 51593
rect 1705 51535 1755 51559
rect 216911 51593 216961 51617
rect 216911 51559 216919 51593
rect 216953 51559 216961 51593
rect 216911 51535 216961 51559
rect 1705 51257 1755 51281
rect 1705 51223 1713 51257
rect 1747 51223 1755 51257
rect 1705 51199 1755 51223
rect 216911 51257 216961 51281
rect 216911 51223 216919 51257
rect 216953 51223 216961 51257
rect 216911 51199 216961 51223
rect 1705 50921 1755 50945
rect 1705 50887 1713 50921
rect 1747 50887 1755 50921
rect 1705 50863 1755 50887
rect 216911 50921 216961 50945
rect 216911 50887 216919 50921
rect 216953 50887 216961 50921
rect 216911 50863 216961 50887
rect 1705 50585 1755 50609
rect 1705 50551 1713 50585
rect 1747 50551 1755 50585
rect 1705 50527 1755 50551
rect 216911 50585 216961 50609
rect 216911 50551 216919 50585
rect 216953 50551 216961 50585
rect 216911 50527 216961 50551
rect 1705 50249 1755 50273
rect 1705 50215 1713 50249
rect 1747 50215 1755 50249
rect 1705 50191 1755 50215
rect 216911 50249 216961 50273
rect 216911 50215 216919 50249
rect 216953 50215 216961 50249
rect 216911 50191 216961 50215
rect 1705 49913 1755 49937
rect 1705 49879 1713 49913
rect 1747 49879 1755 49913
rect 1705 49855 1755 49879
rect 216911 49913 216961 49937
rect 216911 49879 216919 49913
rect 216953 49879 216961 49913
rect 216911 49855 216961 49879
rect 1705 49577 1755 49601
rect 1705 49543 1713 49577
rect 1747 49543 1755 49577
rect 1705 49519 1755 49543
rect 216911 49577 216961 49601
rect 216911 49543 216919 49577
rect 216953 49543 216961 49577
rect 216911 49519 216961 49543
rect 1705 49241 1755 49265
rect 1705 49207 1713 49241
rect 1747 49207 1755 49241
rect 1705 49183 1755 49207
rect 216911 49241 216961 49265
rect 216911 49207 216919 49241
rect 216953 49207 216961 49241
rect 216911 49183 216961 49207
rect 1705 48905 1755 48929
rect 1705 48871 1713 48905
rect 1747 48871 1755 48905
rect 1705 48847 1755 48871
rect 216911 48905 216961 48929
rect 216911 48871 216919 48905
rect 216953 48871 216961 48905
rect 216911 48847 216961 48871
rect 1705 48569 1755 48593
rect 1705 48535 1713 48569
rect 1747 48535 1755 48569
rect 1705 48511 1755 48535
rect 216911 48569 216961 48593
rect 216911 48535 216919 48569
rect 216953 48535 216961 48569
rect 216911 48511 216961 48535
rect 1705 48233 1755 48257
rect 1705 48199 1713 48233
rect 1747 48199 1755 48233
rect 1705 48175 1755 48199
rect 216911 48233 216961 48257
rect 216911 48199 216919 48233
rect 216953 48199 216961 48233
rect 216911 48175 216961 48199
rect 1705 47897 1755 47921
rect 1705 47863 1713 47897
rect 1747 47863 1755 47897
rect 1705 47839 1755 47863
rect 216911 47897 216961 47921
rect 216911 47863 216919 47897
rect 216953 47863 216961 47897
rect 216911 47839 216961 47863
rect 1705 47561 1755 47585
rect 1705 47527 1713 47561
rect 1747 47527 1755 47561
rect 1705 47503 1755 47527
rect 216911 47561 216961 47585
rect 216911 47527 216919 47561
rect 216953 47527 216961 47561
rect 216911 47503 216961 47527
rect 1705 47225 1755 47249
rect 1705 47191 1713 47225
rect 1747 47191 1755 47225
rect 1705 47167 1755 47191
rect 216911 47225 216961 47249
rect 216911 47191 216919 47225
rect 216953 47191 216961 47225
rect 216911 47167 216961 47191
rect 1705 46889 1755 46913
rect 1705 46855 1713 46889
rect 1747 46855 1755 46889
rect 1705 46831 1755 46855
rect 216911 46889 216961 46913
rect 216911 46855 216919 46889
rect 216953 46855 216961 46889
rect 216911 46831 216961 46855
rect 1705 46553 1755 46577
rect 1705 46519 1713 46553
rect 1747 46519 1755 46553
rect 1705 46495 1755 46519
rect 216911 46553 216961 46577
rect 216911 46519 216919 46553
rect 216953 46519 216961 46553
rect 216911 46495 216961 46519
rect 1705 46217 1755 46241
rect 1705 46183 1713 46217
rect 1747 46183 1755 46217
rect 1705 46159 1755 46183
rect 216911 46217 216961 46241
rect 216911 46183 216919 46217
rect 216953 46183 216961 46217
rect 216911 46159 216961 46183
rect 1705 45881 1755 45905
rect 1705 45847 1713 45881
rect 1747 45847 1755 45881
rect 1705 45823 1755 45847
rect 216911 45881 216961 45905
rect 216911 45847 216919 45881
rect 216953 45847 216961 45881
rect 216911 45823 216961 45847
rect 1705 45545 1755 45569
rect 1705 45511 1713 45545
rect 1747 45511 1755 45545
rect 1705 45487 1755 45511
rect 216911 45545 216961 45569
rect 216911 45511 216919 45545
rect 216953 45511 216961 45545
rect 216911 45487 216961 45511
rect 1705 45209 1755 45233
rect 1705 45175 1713 45209
rect 1747 45175 1755 45209
rect 1705 45151 1755 45175
rect 216911 45209 216961 45233
rect 216911 45175 216919 45209
rect 216953 45175 216961 45209
rect 216911 45151 216961 45175
rect 1705 44873 1755 44897
rect 1705 44839 1713 44873
rect 1747 44839 1755 44873
rect 1705 44815 1755 44839
rect 216911 44873 216961 44897
rect 216911 44839 216919 44873
rect 216953 44839 216961 44873
rect 216911 44815 216961 44839
rect 1705 44537 1755 44561
rect 1705 44503 1713 44537
rect 1747 44503 1755 44537
rect 1705 44479 1755 44503
rect 216911 44537 216961 44561
rect 216911 44503 216919 44537
rect 216953 44503 216961 44537
rect 216911 44479 216961 44503
rect 1705 44201 1755 44225
rect 1705 44167 1713 44201
rect 1747 44167 1755 44201
rect 1705 44143 1755 44167
rect 216911 44201 216961 44225
rect 216911 44167 216919 44201
rect 216953 44167 216961 44201
rect 216911 44143 216961 44167
rect 1705 43865 1755 43889
rect 1705 43831 1713 43865
rect 1747 43831 1755 43865
rect 1705 43807 1755 43831
rect 216911 43865 216961 43889
rect 216911 43831 216919 43865
rect 216953 43831 216961 43865
rect 216911 43807 216961 43831
rect 1705 43529 1755 43553
rect 1705 43495 1713 43529
rect 1747 43495 1755 43529
rect 1705 43471 1755 43495
rect 216911 43529 216961 43553
rect 216911 43495 216919 43529
rect 216953 43495 216961 43529
rect 216911 43471 216961 43495
rect 1705 43193 1755 43217
rect 1705 43159 1713 43193
rect 1747 43159 1755 43193
rect 1705 43135 1755 43159
rect 216911 43193 216961 43217
rect 216911 43159 216919 43193
rect 216953 43159 216961 43193
rect 216911 43135 216961 43159
rect 1705 42857 1755 42881
rect 1705 42823 1713 42857
rect 1747 42823 1755 42857
rect 1705 42799 1755 42823
rect 216911 42857 216961 42881
rect 216911 42823 216919 42857
rect 216953 42823 216961 42857
rect 216911 42799 216961 42823
rect 1705 42521 1755 42545
rect 1705 42487 1713 42521
rect 1747 42487 1755 42521
rect 1705 42463 1755 42487
rect 216911 42521 216961 42545
rect 216911 42487 216919 42521
rect 216953 42487 216961 42521
rect 216911 42463 216961 42487
rect 1705 42185 1755 42209
rect 1705 42151 1713 42185
rect 1747 42151 1755 42185
rect 1705 42127 1755 42151
rect 216911 42185 216961 42209
rect 216911 42151 216919 42185
rect 216953 42151 216961 42185
rect 216911 42127 216961 42151
rect 1705 41849 1755 41873
rect 1705 41815 1713 41849
rect 1747 41815 1755 41849
rect 1705 41791 1755 41815
rect 216911 41849 216961 41873
rect 216911 41815 216919 41849
rect 216953 41815 216961 41849
rect 216911 41791 216961 41815
rect 1705 41513 1755 41537
rect 1705 41479 1713 41513
rect 1747 41479 1755 41513
rect 1705 41455 1755 41479
rect 216911 41513 216961 41537
rect 216911 41479 216919 41513
rect 216953 41479 216961 41513
rect 216911 41455 216961 41479
rect 1705 41177 1755 41201
rect 1705 41143 1713 41177
rect 1747 41143 1755 41177
rect 1705 41119 1755 41143
rect 216911 41177 216961 41201
rect 216911 41143 216919 41177
rect 216953 41143 216961 41177
rect 216911 41119 216961 41143
rect 1705 40841 1755 40865
rect 1705 40807 1713 40841
rect 1747 40807 1755 40841
rect 1705 40783 1755 40807
rect 216911 40841 216961 40865
rect 216911 40807 216919 40841
rect 216953 40807 216961 40841
rect 216911 40783 216961 40807
rect 1705 40505 1755 40529
rect 1705 40471 1713 40505
rect 1747 40471 1755 40505
rect 1705 40447 1755 40471
rect 216911 40505 216961 40529
rect 216911 40471 216919 40505
rect 216953 40471 216961 40505
rect 216911 40447 216961 40471
rect 1705 40169 1755 40193
rect 1705 40135 1713 40169
rect 1747 40135 1755 40169
rect 1705 40111 1755 40135
rect 216911 40169 216961 40193
rect 216911 40135 216919 40169
rect 216953 40135 216961 40169
rect 216911 40111 216961 40135
rect 1705 39833 1755 39857
rect 1705 39799 1713 39833
rect 1747 39799 1755 39833
rect 1705 39775 1755 39799
rect 216911 39833 216961 39857
rect 216911 39799 216919 39833
rect 216953 39799 216961 39833
rect 216911 39775 216961 39799
rect 1705 39497 1755 39521
rect 1705 39463 1713 39497
rect 1747 39463 1755 39497
rect 1705 39439 1755 39463
rect 216911 39497 216961 39521
rect 216911 39463 216919 39497
rect 216953 39463 216961 39497
rect 216911 39439 216961 39463
rect 1705 39161 1755 39185
rect 1705 39127 1713 39161
rect 1747 39127 1755 39161
rect 1705 39103 1755 39127
rect 216911 39161 216961 39185
rect 216911 39127 216919 39161
rect 216953 39127 216961 39161
rect 216911 39103 216961 39127
rect 1705 38825 1755 38849
rect 1705 38791 1713 38825
rect 1747 38791 1755 38825
rect 1705 38767 1755 38791
rect 216911 38825 216961 38849
rect 216911 38791 216919 38825
rect 216953 38791 216961 38825
rect 216911 38767 216961 38791
rect 1705 38489 1755 38513
rect 1705 38455 1713 38489
rect 1747 38455 1755 38489
rect 1705 38431 1755 38455
rect 216911 38489 216961 38513
rect 216911 38455 216919 38489
rect 216953 38455 216961 38489
rect 216911 38431 216961 38455
rect 1705 38153 1755 38177
rect 1705 38119 1713 38153
rect 1747 38119 1755 38153
rect 1705 38095 1755 38119
rect 216911 38153 216961 38177
rect 216911 38119 216919 38153
rect 216953 38119 216961 38153
rect 216911 38095 216961 38119
rect 1705 37817 1755 37841
rect 1705 37783 1713 37817
rect 1747 37783 1755 37817
rect 1705 37759 1755 37783
rect 216911 37817 216961 37841
rect 216911 37783 216919 37817
rect 216953 37783 216961 37817
rect 216911 37759 216961 37783
rect 1705 37481 1755 37505
rect 1705 37447 1713 37481
rect 1747 37447 1755 37481
rect 1705 37423 1755 37447
rect 216911 37481 216961 37505
rect 216911 37447 216919 37481
rect 216953 37447 216961 37481
rect 216911 37423 216961 37447
rect 1705 37145 1755 37169
rect 1705 37111 1713 37145
rect 1747 37111 1755 37145
rect 1705 37087 1755 37111
rect 216911 37145 216961 37169
rect 216911 37111 216919 37145
rect 216953 37111 216961 37145
rect 216911 37087 216961 37111
rect 1705 36809 1755 36833
rect 1705 36775 1713 36809
rect 1747 36775 1755 36809
rect 1705 36751 1755 36775
rect 216911 36809 216961 36833
rect 216911 36775 216919 36809
rect 216953 36775 216961 36809
rect 216911 36751 216961 36775
rect 1705 36473 1755 36497
rect 1705 36439 1713 36473
rect 1747 36439 1755 36473
rect 1705 36415 1755 36439
rect 216911 36473 216961 36497
rect 216911 36439 216919 36473
rect 216953 36439 216961 36473
rect 216911 36415 216961 36439
rect 1705 36137 1755 36161
rect 1705 36103 1713 36137
rect 1747 36103 1755 36137
rect 1705 36079 1755 36103
rect 216911 36137 216961 36161
rect 216911 36103 216919 36137
rect 216953 36103 216961 36137
rect 216911 36079 216961 36103
rect 1705 35801 1755 35825
rect 1705 35767 1713 35801
rect 1747 35767 1755 35801
rect 1705 35743 1755 35767
rect 216911 35801 216961 35825
rect 216911 35767 216919 35801
rect 216953 35767 216961 35801
rect 216911 35743 216961 35767
rect 1705 35465 1755 35489
rect 1705 35431 1713 35465
rect 1747 35431 1755 35465
rect 1705 35407 1755 35431
rect 216911 35465 216961 35489
rect 216911 35431 216919 35465
rect 216953 35431 216961 35465
rect 216911 35407 216961 35431
rect 1705 35129 1755 35153
rect 1705 35095 1713 35129
rect 1747 35095 1755 35129
rect 1705 35071 1755 35095
rect 216911 35129 216961 35153
rect 216911 35095 216919 35129
rect 216953 35095 216961 35129
rect 216911 35071 216961 35095
rect 1705 34793 1755 34817
rect 1705 34759 1713 34793
rect 1747 34759 1755 34793
rect 1705 34735 1755 34759
rect 216911 34793 216961 34817
rect 216911 34759 216919 34793
rect 216953 34759 216961 34793
rect 216911 34735 216961 34759
rect 1705 34457 1755 34481
rect 1705 34423 1713 34457
rect 1747 34423 1755 34457
rect 1705 34399 1755 34423
rect 216911 34457 216961 34481
rect 216911 34423 216919 34457
rect 216953 34423 216961 34457
rect 216911 34399 216961 34423
rect 1705 34121 1755 34145
rect 1705 34087 1713 34121
rect 1747 34087 1755 34121
rect 1705 34063 1755 34087
rect 216911 34121 216961 34145
rect 216911 34087 216919 34121
rect 216953 34087 216961 34121
rect 216911 34063 216961 34087
rect 1705 33785 1755 33809
rect 1705 33751 1713 33785
rect 1747 33751 1755 33785
rect 1705 33727 1755 33751
rect 216911 33785 216961 33809
rect 216911 33751 216919 33785
rect 216953 33751 216961 33785
rect 216911 33727 216961 33751
rect 1705 33449 1755 33473
rect 1705 33415 1713 33449
rect 1747 33415 1755 33449
rect 1705 33391 1755 33415
rect 216911 33449 216961 33473
rect 216911 33415 216919 33449
rect 216953 33415 216961 33449
rect 216911 33391 216961 33415
rect 1705 33113 1755 33137
rect 1705 33079 1713 33113
rect 1747 33079 1755 33113
rect 1705 33055 1755 33079
rect 216911 33113 216961 33137
rect 216911 33079 216919 33113
rect 216953 33079 216961 33113
rect 216911 33055 216961 33079
rect 1705 32777 1755 32801
rect 1705 32743 1713 32777
rect 1747 32743 1755 32777
rect 1705 32719 1755 32743
rect 216911 32777 216961 32801
rect 216911 32743 216919 32777
rect 216953 32743 216961 32777
rect 216911 32719 216961 32743
rect 1705 32441 1755 32465
rect 1705 32407 1713 32441
rect 1747 32407 1755 32441
rect 1705 32383 1755 32407
rect 216911 32441 216961 32465
rect 216911 32407 216919 32441
rect 216953 32407 216961 32441
rect 216911 32383 216961 32407
rect 1705 32105 1755 32129
rect 1705 32071 1713 32105
rect 1747 32071 1755 32105
rect 1705 32047 1755 32071
rect 216911 32105 216961 32129
rect 216911 32071 216919 32105
rect 216953 32071 216961 32105
rect 216911 32047 216961 32071
rect 1705 31769 1755 31793
rect 1705 31735 1713 31769
rect 1747 31735 1755 31769
rect 1705 31711 1755 31735
rect 216911 31769 216961 31793
rect 216911 31735 216919 31769
rect 216953 31735 216961 31769
rect 216911 31711 216961 31735
rect 1705 31433 1755 31457
rect 1705 31399 1713 31433
rect 1747 31399 1755 31433
rect 1705 31375 1755 31399
rect 216911 31433 216961 31457
rect 216911 31399 216919 31433
rect 216953 31399 216961 31433
rect 216911 31375 216961 31399
rect 1705 31097 1755 31121
rect 1705 31063 1713 31097
rect 1747 31063 1755 31097
rect 1705 31039 1755 31063
rect 216911 31097 216961 31121
rect 216911 31063 216919 31097
rect 216953 31063 216961 31097
rect 216911 31039 216961 31063
rect 1705 30761 1755 30785
rect 1705 30727 1713 30761
rect 1747 30727 1755 30761
rect 1705 30703 1755 30727
rect 216911 30761 216961 30785
rect 216911 30727 216919 30761
rect 216953 30727 216961 30761
rect 216911 30703 216961 30727
rect 1705 30425 1755 30449
rect 1705 30391 1713 30425
rect 1747 30391 1755 30425
rect 1705 30367 1755 30391
rect 216911 30425 216961 30449
rect 216911 30391 216919 30425
rect 216953 30391 216961 30425
rect 216911 30367 216961 30391
rect 1705 30089 1755 30113
rect 1705 30055 1713 30089
rect 1747 30055 1755 30089
rect 1705 30031 1755 30055
rect 216911 30089 216961 30113
rect 216911 30055 216919 30089
rect 216953 30055 216961 30089
rect 216911 30031 216961 30055
rect 1705 29753 1755 29777
rect 1705 29719 1713 29753
rect 1747 29719 1755 29753
rect 1705 29695 1755 29719
rect 216911 29753 216961 29777
rect 216911 29719 216919 29753
rect 216953 29719 216961 29753
rect 216911 29695 216961 29719
rect 1705 29417 1755 29441
rect 1705 29383 1713 29417
rect 1747 29383 1755 29417
rect 1705 29359 1755 29383
rect 216911 29417 216961 29441
rect 216911 29383 216919 29417
rect 216953 29383 216961 29417
rect 216911 29359 216961 29383
rect 1705 29081 1755 29105
rect 1705 29047 1713 29081
rect 1747 29047 1755 29081
rect 1705 29023 1755 29047
rect 216911 29081 216961 29105
rect 216911 29047 216919 29081
rect 216953 29047 216961 29081
rect 216911 29023 216961 29047
rect 1705 28745 1755 28769
rect 1705 28711 1713 28745
rect 1747 28711 1755 28745
rect 1705 28687 1755 28711
rect 216911 28745 216961 28769
rect 216911 28711 216919 28745
rect 216953 28711 216961 28745
rect 216911 28687 216961 28711
rect 1705 28409 1755 28433
rect 1705 28375 1713 28409
rect 1747 28375 1755 28409
rect 1705 28351 1755 28375
rect 216911 28409 216961 28433
rect 216911 28375 216919 28409
rect 216953 28375 216961 28409
rect 216911 28351 216961 28375
rect 1705 28073 1755 28097
rect 1705 28039 1713 28073
rect 1747 28039 1755 28073
rect 1705 28015 1755 28039
rect 216911 28073 216961 28097
rect 216911 28039 216919 28073
rect 216953 28039 216961 28073
rect 216911 28015 216961 28039
rect 1705 27737 1755 27761
rect 1705 27703 1713 27737
rect 1747 27703 1755 27737
rect 1705 27679 1755 27703
rect 216911 27737 216961 27761
rect 216911 27703 216919 27737
rect 216953 27703 216961 27737
rect 216911 27679 216961 27703
rect 1705 27401 1755 27425
rect 1705 27367 1713 27401
rect 1747 27367 1755 27401
rect 1705 27343 1755 27367
rect 216911 27401 216961 27425
rect 216911 27367 216919 27401
rect 216953 27367 216961 27401
rect 216911 27343 216961 27367
rect 1705 27065 1755 27089
rect 1705 27031 1713 27065
rect 1747 27031 1755 27065
rect 1705 27007 1755 27031
rect 216911 27065 216961 27089
rect 216911 27031 216919 27065
rect 216953 27031 216961 27065
rect 216911 27007 216961 27031
rect 1705 26729 1755 26753
rect 1705 26695 1713 26729
rect 1747 26695 1755 26729
rect 1705 26671 1755 26695
rect 216911 26729 216961 26753
rect 216911 26695 216919 26729
rect 216953 26695 216961 26729
rect 216911 26671 216961 26695
rect 1705 26393 1755 26417
rect 1705 26359 1713 26393
rect 1747 26359 1755 26393
rect 1705 26335 1755 26359
rect 216911 26393 216961 26417
rect 216911 26359 216919 26393
rect 216953 26359 216961 26393
rect 216911 26335 216961 26359
rect 1705 26057 1755 26081
rect 1705 26023 1713 26057
rect 1747 26023 1755 26057
rect 1705 25999 1755 26023
rect 216911 26057 216961 26081
rect 216911 26023 216919 26057
rect 216953 26023 216961 26057
rect 216911 25999 216961 26023
rect 1705 25721 1755 25745
rect 1705 25687 1713 25721
rect 1747 25687 1755 25721
rect 1705 25663 1755 25687
rect 216911 25721 216961 25745
rect 216911 25687 216919 25721
rect 216953 25687 216961 25721
rect 216911 25663 216961 25687
rect 1705 25385 1755 25409
rect 1705 25351 1713 25385
rect 1747 25351 1755 25385
rect 1705 25327 1755 25351
rect 216911 25385 216961 25409
rect 216911 25351 216919 25385
rect 216953 25351 216961 25385
rect 216911 25327 216961 25351
rect 1705 25049 1755 25073
rect 1705 25015 1713 25049
rect 1747 25015 1755 25049
rect 1705 24991 1755 25015
rect 216911 25049 216961 25073
rect 216911 25015 216919 25049
rect 216953 25015 216961 25049
rect 216911 24991 216961 25015
rect 1705 24713 1755 24737
rect 1705 24679 1713 24713
rect 1747 24679 1755 24713
rect 1705 24655 1755 24679
rect 216911 24713 216961 24737
rect 216911 24679 216919 24713
rect 216953 24679 216961 24713
rect 216911 24655 216961 24679
rect 1705 24377 1755 24401
rect 1705 24343 1713 24377
rect 1747 24343 1755 24377
rect 1705 24319 1755 24343
rect 216911 24377 216961 24401
rect 216911 24343 216919 24377
rect 216953 24343 216961 24377
rect 216911 24319 216961 24343
rect 1705 24041 1755 24065
rect 1705 24007 1713 24041
rect 1747 24007 1755 24041
rect 1705 23983 1755 24007
rect 216911 24041 216961 24065
rect 216911 24007 216919 24041
rect 216953 24007 216961 24041
rect 216911 23983 216961 24007
rect 1705 23705 1755 23729
rect 1705 23671 1713 23705
rect 1747 23671 1755 23705
rect 1705 23647 1755 23671
rect 216911 23705 216961 23729
rect 216911 23671 216919 23705
rect 216953 23671 216961 23705
rect 216911 23647 216961 23671
rect 1705 23369 1755 23393
rect 1705 23335 1713 23369
rect 1747 23335 1755 23369
rect 1705 23311 1755 23335
rect 216911 23369 216961 23393
rect 216911 23335 216919 23369
rect 216953 23335 216961 23369
rect 216911 23311 216961 23335
rect 1705 23033 1755 23057
rect 1705 22999 1713 23033
rect 1747 22999 1755 23033
rect 1705 22975 1755 22999
rect 216911 23033 216961 23057
rect 216911 22999 216919 23033
rect 216953 22999 216961 23033
rect 216911 22975 216961 22999
rect 1705 22697 1755 22721
rect 1705 22663 1713 22697
rect 1747 22663 1755 22697
rect 1705 22639 1755 22663
rect 216911 22697 216961 22721
rect 216911 22663 216919 22697
rect 216953 22663 216961 22697
rect 216911 22639 216961 22663
rect 1705 22361 1755 22385
rect 1705 22327 1713 22361
rect 1747 22327 1755 22361
rect 1705 22303 1755 22327
rect 216911 22361 216961 22385
rect 216911 22327 216919 22361
rect 216953 22327 216961 22361
rect 216911 22303 216961 22327
rect 1705 22025 1755 22049
rect 1705 21991 1713 22025
rect 1747 21991 1755 22025
rect 1705 21967 1755 21991
rect 216911 22025 216961 22049
rect 216911 21991 216919 22025
rect 216953 21991 216961 22025
rect 216911 21967 216961 21991
rect 1705 21689 1755 21713
rect 1705 21655 1713 21689
rect 1747 21655 1755 21689
rect 1705 21631 1755 21655
rect 216911 21689 216961 21713
rect 216911 21655 216919 21689
rect 216953 21655 216961 21689
rect 216911 21631 216961 21655
rect 1705 21353 1755 21377
rect 1705 21319 1713 21353
rect 1747 21319 1755 21353
rect 1705 21295 1755 21319
rect 216911 21353 216961 21377
rect 216911 21319 216919 21353
rect 216953 21319 216961 21353
rect 216911 21295 216961 21319
rect 1705 21017 1755 21041
rect 1705 20983 1713 21017
rect 1747 20983 1755 21017
rect 1705 20959 1755 20983
rect 216911 21017 216961 21041
rect 216911 20983 216919 21017
rect 216953 20983 216961 21017
rect 216911 20959 216961 20983
rect 1705 20681 1755 20705
rect 1705 20647 1713 20681
rect 1747 20647 1755 20681
rect 1705 20623 1755 20647
rect 216911 20681 216961 20705
rect 216911 20647 216919 20681
rect 216953 20647 216961 20681
rect 216911 20623 216961 20647
rect 1705 20345 1755 20369
rect 1705 20311 1713 20345
rect 1747 20311 1755 20345
rect 1705 20287 1755 20311
rect 216911 20345 216961 20369
rect 216911 20311 216919 20345
rect 216953 20311 216961 20345
rect 216911 20287 216961 20311
rect 1705 20009 1755 20033
rect 1705 19975 1713 20009
rect 1747 19975 1755 20009
rect 1705 19951 1755 19975
rect 216911 20009 216961 20033
rect 216911 19975 216919 20009
rect 216953 19975 216961 20009
rect 216911 19951 216961 19975
rect 1705 19673 1755 19697
rect 1705 19639 1713 19673
rect 1747 19639 1755 19673
rect 1705 19615 1755 19639
rect 216911 19673 216961 19697
rect 216911 19639 216919 19673
rect 216953 19639 216961 19673
rect 216911 19615 216961 19639
rect 1705 19337 1755 19361
rect 1705 19303 1713 19337
rect 1747 19303 1755 19337
rect 1705 19279 1755 19303
rect 216911 19337 216961 19361
rect 216911 19303 216919 19337
rect 216953 19303 216961 19337
rect 216911 19279 216961 19303
rect 1705 19001 1755 19025
rect 1705 18967 1713 19001
rect 1747 18967 1755 19001
rect 1705 18943 1755 18967
rect 216911 19001 216961 19025
rect 216911 18967 216919 19001
rect 216953 18967 216961 19001
rect 216911 18943 216961 18967
rect 1705 18665 1755 18689
rect 1705 18631 1713 18665
rect 1747 18631 1755 18665
rect 1705 18607 1755 18631
rect 216911 18665 216961 18689
rect 216911 18631 216919 18665
rect 216953 18631 216961 18665
rect 216911 18607 216961 18631
rect 1705 18329 1755 18353
rect 1705 18295 1713 18329
rect 1747 18295 1755 18329
rect 1705 18271 1755 18295
rect 216911 18329 216961 18353
rect 216911 18295 216919 18329
rect 216953 18295 216961 18329
rect 216911 18271 216961 18295
rect 1705 17993 1755 18017
rect 1705 17959 1713 17993
rect 1747 17959 1755 17993
rect 1705 17935 1755 17959
rect 216911 17993 216961 18017
rect 216911 17959 216919 17993
rect 216953 17959 216961 17993
rect 216911 17935 216961 17959
rect 1705 17657 1755 17681
rect 1705 17623 1713 17657
rect 1747 17623 1755 17657
rect 1705 17599 1755 17623
rect 216911 17657 216961 17681
rect 216911 17623 216919 17657
rect 216953 17623 216961 17657
rect 216911 17599 216961 17623
rect 1705 17321 1755 17345
rect 1705 17287 1713 17321
rect 1747 17287 1755 17321
rect 1705 17263 1755 17287
rect 216911 17321 216961 17345
rect 216911 17287 216919 17321
rect 216953 17287 216961 17321
rect 216911 17263 216961 17287
rect 1705 16985 1755 17009
rect 1705 16951 1713 16985
rect 1747 16951 1755 16985
rect 1705 16927 1755 16951
rect 216911 16985 216961 17009
rect 216911 16951 216919 16985
rect 216953 16951 216961 16985
rect 216911 16927 216961 16951
rect 1705 16649 1755 16673
rect 1705 16615 1713 16649
rect 1747 16615 1755 16649
rect 1705 16591 1755 16615
rect 216911 16649 216961 16673
rect 216911 16615 216919 16649
rect 216953 16615 216961 16649
rect 216911 16591 216961 16615
rect 1705 16313 1755 16337
rect 1705 16279 1713 16313
rect 1747 16279 1755 16313
rect 1705 16255 1755 16279
rect 216911 16313 216961 16337
rect 216911 16279 216919 16313
rect 216953 16279 216961 16313
rect 216911 16255 216961 16279
rect 1705 15977 1755 16001
rect 1705 15943 1713 15977
rect 1747 15943 1755 15977
rect 1705 15919 1755 15943
rect 216911 15977 216961 16001
rect 216911 15943 216919 15977
rect 216953 15943 216961 15977
rect 216911 15919 216961 15943
rect 1705 15641 1755 15665
rect 1705 15607 1713 15641
rect 1747 15607 1755 15641
rect 1705 15583 1755 15607
rect 216911 15641 216961 15665
rect 216911 15607 216919 15641
rect 216953 15607 216961 15641
rect 216911 15583 216961 15607
rect 1705 15305 1755 15329
rect 1705 15271 1713 15305
rect 1747 15271 1755 15305
rect 1705 15247 1755 15271
rect 216911 15305 216961 15329
rect 216911 15271 216919 15305
rect 216953 15271 216961 15305
rect 216911 15247 216961 15271
rect 1705 14969 1755 14993
rect 1705 14935 1713 14969
rect 1747 14935 1755 14969
rect 1705 14911 1755 14935
rect 216911 14969 216961 14993
rect 216911 14935 216919 14969
rect 216953 14935 216961 14969
rect 216911 14911 216961 14935
rect 1705 14633 1755 14657
rect 1705 14599 1713 14633
rect 1747 14599 1755 14633
rect 1705 14575 1755 14599
rect 216911 14633 216961 14657
rect 216911 14599 216919 14633
rect 216953 14599 216961 14633
rect 216911 14575 216961 14599
rect 1705 14297 1755 14321
rect 1705 14263 1713 14297
rect 1747 14263 1755 14297
rect 1705 14239 1755 14263
rect 216911 14297 216961 14321
rect 216911 14263 216919 14297
rect 216953 14263 216961 14297
rect 216911 14239 216961 14263
rect 1705 13961 1755 13985
rect 1705 13927 1713 13961
rect 1747 13927 1755 13961
rect 1705 13903 1755 13927
rect 216911 13961 216961 13985
rect 216911 13927 216919 13961
rect 216953 13927 216961 13961
rect 216911 13903 216961 13927
rect 1705 13625 1755 13649
rect 1705 13591 1713 13625
rect 1747 13591 1755 13625
rect 1705 13567 1755 13591
rect 216911 13625 216961 13649
rect 216911 13591 216919 13625
rect 216953 13591 216961 13625
rect 216911 13567 216961 13591
rect 1705 13289 1755 13313
rect 1705 13255 1713 13289
rect 1747 13255 1755 13289
rect 1705 13231 1755 13255
rect 216911 13289 216961 13313
rect 216911 13255 216919 13289
rect 216953 13255 216961 13289
rect 216911 13231 216961 13255
rect 1705 12953 1755 12977
rect 1705 12919 1713 12953
rect 1747 12919 1755 12953
rect 1705 12895 1755 12919
rect 216911 12953 216961 12977
rect 216911 12919 216919 12953
rect 216953 12919 216961 12953
rect 216911 12895 216961 12919
rect 1705 12617 1755 12641
rect 1705 12583 1713 12617
rect 1747 12583 1755 12617
rect 1705 12559 1755 12583
rect 216911 12617 216961 12641
rect 216911 12583 216919 12617
rect 216953 12583 216961 12617
rect 216911 12559 216961 12583
rect 1705 12281 1755 12305
rect 1705 12247 1713 12281
rect 1747 12247 1755 12281
rect 1705 12223 1755 12247
rect 216911 12281 216961 12305
rect 216911 12247 216919 12281
rect 216953 12247 216961 12281
rect 216911 12223 216961 12247
rect 1705 11945 1755 11969
rect 1705 11911 1713 11945
rect 1747 11911 1755 11945
rect 1705 11887 1755 11911
rect 216911 11945 216961 11969
rect 216911 11911 216919 11945
rect 216953 11911 216961 11945
rect 216911 11887 216961 11911
rect 1705 11609 1755 11633
rect 1705 11575 1713 11609
rect 1747 11575 1755 11609
rect 1705 11551 1755 11575
rect 216911 11609 216961 11633
rect 216911 11575 216919 11609
rect 216953 11575 216961 11609
rect 216911 11551 216961 11575
rect 1705 11273 1755 11297
rect 1705 11239 1713 11273
rect 1747 11239 1755 11273
rect 1705 11215 1755 11239
rect 216911 11273 216961 11297
rect 216911 11239 216919 11273
rect 216953 11239 216961 11273
rect 216911 11215 216961 11239
rect 1705 10937 1755 10961
rect 1705 10903 1713 10937
rect 1747 10903 1755 10937
rect 1705 10879 1755 10903
rect 216911 10937 216961 10961
rect 216911 10903 216919 10937
rect 216953 10903 216961 10937
rect 216911 10879 216961 10903
rect 1705 10601 1755 10625
rect 1705 10567 1713 10601
rect 1747 10567 1755 10601
rect 1705 10543 1755 10567
rect 216911 10601 216961 10625
rect 216911 10567 216919 10601
rect 216953 10567 216961 10601
rect 216911 10543 216961 10567
rect 1705 10265 1755 10289
rect 1705 10231 1713 10265
rect 1747 10231 1755 10265
rect 1705 10207 1755 10231
rect 216911 10265 216961 10289
rect 216911 10231 216919 10265
rect 216953 10231 216961 10265
rect 216911 10207 216961 10231
rect 1705 9929 1755 9953
rect 1705 9895 1713 9929
rect 1747 9895 1755 9929
rect 1705 9871 1755 9895
rect 216911 9929 216961 9953
rect 216911 9895 216919 9929
rect 216953 9895 216961 9929
rect 216911 9871 216961 9895
rect 1705 9593 1755 9617
rect 1705 9559 1713 9593
rect 1747 9559 1755 9593
rect 1705 9535 1755 9559
rect 216911 9593 216961 9617
rect 216911 9559 216919 9593
rect 216953 9559 216961 9593
rect 216911 9535 216961 9559
rect 1705 9257 1755 9281
rect 1705 9223 1713 9257
rect 1747 9223 1755 9257
rect 1705 9199 1755 9223
rect 216911 9257 216961 9281
rect 216911 9223 216919 9257
rect 216953 9223 216961 9257
rect 216911 9199 216961 9223
rect 1705 8921 1755 8945
rect 1705 8887 1713 8921
rect 1747 8887 1755 8921
rect 1705 8863 1755 8887
rect 216911 8921 216961 8945
rect 216911 8887 216919 8921
rect 216953 8887 216961 8921
rect 216911 8863 216961 8887
rect 1705 8585 1755 8609
rect 1705 8551 1713 8585
rect 1747 8551 1755 8585
rect 1705 8527 1755 8551
rect 216911 8585 216961 8609
rect 216911 8551 216919 8585
rect 216953 8551 216961 8585
rect 216911 8527 216961 8551
rect 1705 8249 1755 8273
rect 1705 8215 1713 8249
rect 1747 8215 1755 8249
rect 1705 8191 1755 8215
rect 216911 8249 216961 8273
rect 216911 8215 216919 8249
rect 216953 8215 216961 8249
rect 216911 8191 216961 8215
rect 1705 7913 1755 7937
rect 1705 7879 1713 7913
rect 1747 7879 1755 7913
rect 1705 7855 1755 7879
rect 216911 7913 216961 7937
rect 216911 7879 216919 7913
rect 216953 7879 216961 7913
rect 216911 7855 216961 7879
rect 1705 7577 1755 7601
rect 1705 7543 1713 7577
rect 1747 7543 1755 7577
rect 1705 7519 1755 7543
rect 216911 7577 216961 7601
rect 216911 7543 216919 7577
rect 216953 7543 216961 7577
rect 216911 7519 216961 7543
rect 1705 7241 1755 7265
rect 1705 7207 1713 7241
rect 1747 7207 1755 7241
rect 1705 7183 1755 7207
rect 216911 7241 216961 7265
rect 216911 7207 216919 7241
rect 216953 7207 216961 7241
rect 216911 7183 216961 7207
rect 1705 6905 1755 6929
rect 1705 6871 1713 6905
rect 1747 6871 1755 6905
rect 1705 6847 1755 6871
rect 216911 6905 216961 6929
rect 216911 6871 216919 6905
rect 216953 6871 216961 6905
rect 216911 6847 216961 6871
rect 1705 6569 1755 6593
rect 1705 6535 1713 6569
rect 1747 6535 1755 6569
rect 1705 6511 1755 6535
rect 216911 6569 216961 6593
rect 216911 6535 216919 6569
rect 216953 6535 216961 6569
rect 216911 6511 216961 6535
rect 1705 6233 1755 6257
rect 1705 6199 1713 6233
rect 1747 6199 1755 6233
rect 1705 6175 1755 6199
rect 216911 6233 216961 6257
rect 216911 6199 216919 6233
rect 216953 6199 216961 6233
rect 216911 6175 216961 6199
rect 1705 5897 1755 5921
rect 1705 5863 1713 5897
rect 1747 5863 1755 5897
rect 1705 5839 1755 5863
rect 216911 5897 216961 5921
rect 216911 5863 216919 5897
rect 216953 5863 216961 5897
rect 216911 5839 216961 5863
rect 1705 5561 1755 5585
rect 1705 5527 1713 5561
rect 1747 5527 1755 5561
rect 1705 5503 1755 5527
rect 216911 5561 216961 5585
rect 216911 5527 216919 5561
rect 216953 5527 216961 5561
rect 216911 5503 216961 5527
rect 1705 5225 1755 5249
rect 1705 5191 1713 5225
rect 1747 5191 1755 5225
rect 1705 5167 1755 5191
rect 216911 5225 216961 5249
rect 216911 5191 216919 5225
rect 216953 5191 216961 5225
rect 216911 5167 216961 5191
rect 1705 4889 1755 4913
rect 1705 4855 1713 4889
rect 1747 4855 1755 4889
rect 1705 4831 1755 4855
rect 216911 4889 216961 4913
rect 216911 4855 216919 4889
rect 216953 4855 216961 4889
rect 216911 4831 216961 4855
rect 1705 4553 1755 4577
rect 1705 4519 1713 4553
rect 1747 4519 1755 4553
rect 1705 4495 1755 4519
rect 216911 4553 216961 4577
rect 216911 4519 216919 4553
rect 216953 4519 216961 4553
rect 216911 4495 216961 4519
rect 1705 4217 1755 4241
rect 1705 4183 1713 4217
rect 1747 4183 1755 4217
rect 1705 4159 1755 4183
rect 216911 4217 216961 4241
rect 216911 4183 216919 4217
rect 216953 4183 216961 4217
rect 216911 4159 216961 4183
rect 1705 3881 1755 3905
rect 1705 3847 1713 3881
rect 1747 3847 1755 3881
rect 1705 3823 1755 3847
rect 216911 3881 216961 3905
rect 216911 3847 216919 3881
rect 216953 3847 216961 3881
rect 216911 3823 216961 3847
rect 1705 3545 1755 3569
rect 1705 3511 1713 3545
rect 1747 3511 1755 3545
rect 1705 3487 1755 3511
rect 216911 3545 216961 3569
rect 216911 3511 216919 3545
rect 216953 3511 216961 3545
rect 216911 3487 216961 3511
rect 1705 3209 1755 3233
rect 1705 3175 1713 3209
rect 1747 3175 1755 3209
rect 1705 3151 1755 3175
rect 216911 3209 216961 3233
rect 216911 3175 216919 3209
rect 216953 3175 216961 3209
rect 216911 3151 216961 3175
rect 1705 2873 1755 2897
rect 1705 2839 1713 2873
rect 1747 2839 1755 2873
rect 1705 2815 1755 2839
rect 216911 2873 216961 2897
rect 216911 2839 216919 2873
rect 216953 2839 216961 2873
rect 216911 2815 216961 2839
rect 1705 2537 1755 2561
rect 1705 2503 1713 2537
rect 1747 2503 1755 2537
rect 1705 2479 1755 2503
rect 216911 2537 216961 2561
rect 216911 2503 216919 2537
rect 216953 2503 216961 2537
rect 216911 2479 216961 2503
rect 1705 2201 1755 2225
rect 1705 2167 1713 2201
rect 1747 2167 1755 2201
rect 1705 2143 1755 2167
rect 216911 2201 216961 2225
rect 216911 2167 216919 2201
rect 216953 2167 216961 2201
rect 216911 2143 216961 2167
rect 2041 1865 2091 1889
rect 2041 1831 2049 1865
rect 2083 1831 2091 1865
rect 2041 1807 2091 1831
rect 2377 1865 2427 1889
rect 2377 1831 2385 1865
rect 2419 1831 2427 1865
rect 2377 1807 2427 1831
rect 2713 1865 2763 1889
rect 2713 1831 2721 1865
rect 2755 1831 2763 1865
rect 2713 1807 2763 1831
rect 3049 1865 3099 1889
rect 3049 1831 3057 1865
rect 3091 1831 3099 1865
rect 3049 1807 3099 1831
rect 3385 1865 3435 1889
rect 3385 1831 3393 1865
rect 3427 1831 3435 1865
rect 3385 1807 3435 1831
rect 3721 1865 3771 1889
rect 3721 1831 3729 1865
rect 3763 1831 3771 1865
rect 3721 1807 3771 1831
rect 4057 1865 4107 1889
rect 4057 1831 4065 1865
rect 4099 1831 4107 1865
rect 4057 1807 4107 1831
rect 4393 1865 4443 1889
rect 4393 1831 4401 1865
rect 4435 1831 4443 1865
rect 4393 1807 4443 1831
rect 4729 1865 4779 1889
rect 4729 1831 4737 1865
rect 4771 1831 4779 1865
rect 4729 1807 4779 1831
rect 5065 1865 5115 1889
rect 5065 1831 5073 1865
rect 5107 1831 5115 1865
rect 5065 1807 5115 1831
rect 5401 1865 5451 1889
rect 5401 1831 5409 1865
rect 5443 1831 5451 1865
rect 5401 1807 5451 1831
rect 5737 1865 5787 1889
rect 5737 1831 5745 1865
rect 5779 1831 5787 1865
rect 5737 1807 5787 1831
rect 6073 1865 6123 1889
rect 6073 1831 6081 1865
rect 6115 1831 6123 1865
rect 6073 1807 6123 1831
rect 6409 1865 6459 1889
rect 6409 1831 6417 1865
rect 6451 1831 6459 1865
rect 6409 1807 6459 1831
rect 6745 1865 6795 1889
rect 6745 1831 6753 1865
rect 6787 1831 6795 1865
rect 6745 1807 6795 1831
rect 7081 1865 7131 1889
rect 7081 1831 7089 1865
rect 7123 1831 7131 1865
rect 7081 1807 7131 1831
rect 7417 1865 7467 1889
rect 7417 1831 7425 1865
rect 7459 1831 7467 1865
rect 7417 1807 7467 1831
rect 7753 1865 7803 1889
rect 7753 1831 7761 1865
rect 7795 1831 7803 1865
rect 7753 1807 7803 1831
rect 8089 1865 8139 1889
rect 8089 1831 8097 1865
rect 8131 1831 8139 1865
rect 8089 1807 8139 1831
rect 8425 1865 8475 1889
rect 8425 1831 8433 1865
rect 8467 1831 8475 1865
rect 8425 1807 8475 1831
rect 8761 1865 8811 1889
rect 8761 1831 8769 1865
rect 8803 1831 8811 1865
rect 8761 1807 8811 1831
rect 9097 1865 9147 1889
rect 9097 1831 9105 1865
rect 9139 1831 9147 1865
rect 9097 1807 9147 1831
rect 9433 1865 9483 1889
rect 9433 1831 9441 1865
rect 9475 1831 9483 1865
rect 9433 1807 9483 1831
rect 9769 1865 9819 1889
rect 9769 1831 9777 1865
rect 9811 1831 9819 1865
rect 9769 1807 9819 1831
rect 10105 1865 10155 1889
rect 10105 1831 10113 1865
rect 10147 1831 10155 1865
rect 10105 1807 10155 1831
rect 10441 1865 10491 1889
rect 10441 1831 10449 1865
rect 10483 1831 10491 1865
rect 10441 1807 10491 1831
rect 10777 1865 10827 1889
rect 10777 1831 10785 1865
rect 10819 1831 10827 1865
rect 10777 1807 10827 1831
rect 11113 1865 11163 1889
rect 11113 1831 11121 1865
rect 11155 1831 11163 1865
rect 11113 1807 11163 1831
rect 11449 1865 11499 1889
rect 11449 1831 11457 1865
rect 11491 1831 11499 1865
rect 11449 1807 11499 1831
rect 11785 1865 11835 1889
rect 11785 1831 11793 1865
rect 11827 1831 11835 1865
rect 11785 1807 11835 1831
rect 12121 1865 12171 1889
rect 12121 1831 12129 1865
rect 12163 1831 12171 1865
rect 12121 1807 12171 1831
rect 12457 1865 12507 1889
rect 12457 1831 12465 1865
rect 12499 1831 12507 1865
rect 12457 1807 12507 1831
rect 12793 1865 12843 1889
rect 12793 1831 12801 1865
rect 12835 1831 12843 1865
rect 12793 1807 12843 1831
rect 13129 1865 13179 1889
rect 13129 1831 13137 1865
rect 13171 1831 13179 1865
rect 13129 1807 13179 1831
rect 13465 1865 13515 1889
rect 13465 1831 13473 1865
rect 13507 1831 13515 1865
rect 13465 1807 13515 1831
rect 13801 1865 13851 1889
rect 13801 1831 13809 1865
rect 13843 1831 13851 1865
rect 13801 1807 13851 1831
rect 14137 1865 14187 1889
rect 14137 1831 14145 1865
rect 14179 1831 14187 1865
rect 14137 1807 14187 1831
rect 14473 1865 14523 1889
rect 14473 1831 14481 1865
rect 14515 1831 14523 1865
rect 14473 1807 14523 1831
rect 14809 1865 14859 1889
rect 14809 1831 14817 1865
rect 14851 1831 14859 1865
rect 14809 1807 14859 1831
rect 15145 1865 15195 1889
rect 15145 1831 15153 1865
rect 15187 1831 15195 1865
rect 15145 1807 15195 1831
rect 15481 1865 15531 1889
rect 15481 1831 15489 1865
rect 15523 1831 15531 1865
rect 15481 1807 15531 1831
rect 15817 1865 15867 1889
rect 15817 1831 15825 1865
rect 15859 1831 15867 1865
rect 15817 1807 15867 1831
rect 16153 1865 16203 1889
rect 16153 1831 16161 1865
rect 16195 1831 16203 1865
rect 16153 1807 16203 1831
rect 16489 1865 16539 1889
rect 16489 1831 16497 1865
rect 16531 1831 16539 1865
rect 16489 1807 16539 1831
rect 16825 1865 16875 1889
rect 16825 1831 16833 1865
rect 16867 1831 16875 1865
rect 16825 1807 16875 1831
rect 17161 1865 17211 1889
rect 17161 1831 17169 1865
rect 17203 1831 17211 1865
rect 17161 1807 17211 1831
rect 17497 1865 17547 1889
rect 17497 1831 17505 1865
rect 17539 1831 17547 1865
rect 17497 1807 17547 1831
rect 17833 1865 17883 1889
rect 17833 1831 17841 1865
rect 17875 1831 17883 1865
rect 17833 1807 17883 1831
rect 18169 1865 18219 1889
rect 18169 1831 18177 1865
rect 18211 1831 18219 1865
rect 18169 1807 18219 1831
rect 18505 1865 18555 1889
rect 18505 1831 18513 1865
rect 18547 1831 18555 1865
rect 18505 1807 18555 1831
rect 18841 1865 18891 1889
rect 18841 1831 18849 1865
rect 18883 1831 18891 1865
rect 18841 1807 18891 1831
rect 19177 1865 19227 1889
rect 19177 1831 19185 1865
rect 19219 1831 19227 1865
rect 19177 1807 19227 1831
rect 19513 1865 19563 1889
rect 19513 1831 19521 1865
rect 19555 1831 19563 1865
rect 19513 1807 19563 1831
rect 19849 1865 19899 1889
rect 19849 1831 19857 1865
rect 19891 1831 19899 1865
rect 19849 1807 19899 1831
rect 20185 1865 20235 1889
rect 20185 1831 20193 1865
rect 20227 1831 20235 1865
rect 20185 1807 20235 1831
rect 20521 1865 20571 1889
rect 20521 1831 20529 1865
rect 20563 1831 20571 1865
rect 20521 1807 20571 1831
rect 20857 1865 20907 1889
rect 20857 1831 20865 1865
rect 20899 1831 20907 1865
rect 20857 1807 20907 1831
rect 21193 1865 21243 1889
rect 21193 1831 21201 1865
rect 21235 1831 21243 1865
rect 21193 1807 21243 1831
rect 21529 1865 21579 1889
rect 21529 1831 21537 1865
rect 21571 1831 21579 1865
rect 21529 1807 21579 1831
rect 21865 1865 21915 1889
rect 21865 1831 21873 1865
rect 21907 1831 21915 1865
rect 21865 1807 21915 1831
rect 22201 1865 22251 1889
rect 22201 1831 22209 1865
rect 22243 1831 22251 1865
rect 22201 1807 22251 1831
rect 22537 1865 22587 1889
rect 22537 1831 22545 1865
rect 22579 1831 22587 1865
rect 22537 1807 22587 1831
rect 22873 1865 22923 1889
rect 22873 1831 22881 1865
rect 22915 1831 22923 1865
rect 22873 1807 22923 1831
rect 23209 1865 23259 1889
rect 23209 1831 23217 1865
rect 23251 1831 23259 1865
rect 23209 1807 23259 1831
rect 23545 1865 23595 1889
rect 23545 1831 23553 1865
rect 23587 1831 23595 1865
rect 23545 1807 23595 1831
rect 23881 1865 23931 1889
rect 23881 1831 23889 1865
rect 23923 1831 23931 1865
rect 23881 1807 23931 1831
rect 24217 1865 24267 1889
rect 24217 1831 24225 1865
rect 24259 1831 24267 1865
rect 24217 1807 24267 1831
rect 24553 1865 24603 1889
rect 24553 1831 24561 1865
rect 24595 1831 24603 1865
rect 24553 1807 24603 1831
rect 24889 1865 24939 1889
rect 24889 1831 24897 1865
rect 24931 1831 24939 1865
rect 24889 1807 24939 1831
rect 25225 1865 25275 1889
rect 25225 1831 25233 1865
rect 25267 1831 25275 1865
rect 25225 1807 25275 1831
rect 25561 1865 25611 1889
rect 25561 1831 25569 1865
rect 25603 1831 25611 1865
rect 25561 1807 25611 1831
rect 25897 1865 25947 1889
rect 25897 1831 25905 1865
rect 25939 1831 25947 1865
rect 25897 1807 25947 1831
rect 26233 1865 26283 1889
rect 26233 1831 26241 1865
rect 26275 1831 26283 1865
rect 26233 1807 26283 1831
rect 26569 1865 26619 1889
rect 26569 1831 26577 1865
rect 26611 1831 26619 1865
rect 26569 1807 26619 1831
rect 26905 1865 26955 1889
rect 26905 1831 26913 1865
rect 26947 1831 26955 1865
rect 26905 1807 26955 1831
rect 27241 1865 27291 1889
rect 27241 1831 27249 1865
rect 27283 1831 27291 1865
rect 27241 1807 27291 1831
rect 27577 1865 27627 1889
rect 27577 1831 27585 1865
rect 27619 1831 27627 1865
rect 27577 1807 27627 1831
rect 27913 1865 27963 1889
rect 27913 1831 27921 1865
rect 27955 1831 27963 1865
rect 27913 1807 27963 1831
rect 28249 1865 28299 1889
rect 28249 1831 28257 1865
rect 28291 1831 28299 1865
rect 28249 1807 28299 1831
rect 28585 1865 28635 1889
rect 28585 1831 28593 1865
rect 28627 1831 28635 1865
rect 28585 1807 28635 1831
rect 28921 1865 28971 1889
rect 28921 1831 28929 1865
rect 28963 1831 28971 1865
rect 28921 1807 28971 1831
rect 29257 1865 29307 1889
rect 29257 1831 29265 1865
rect 29299 1831 29307 1865
rect 29257 1807 29307 1831
rect 29593 1865 29643 1889
rect 29593 1831 29601 1865
rect 29635 1831 29643 1865
rect 29593 1807 29643 1831
rect 29929 1865 29979 1889
rect 29929 1831 29937 1865
rect 29971 1831 29979 1865
rect 29929 1807 29979 1831
rect 30265 1865 30315 1889
rect 30265 1831 30273 1865
rect 30307 1831 30315 1865
rect 30265 1807 30315 1831
rect 30601 1865 30651 1889
rect 30601 1831 30609 1865
rect 30643 1831 30651 1865
rect 30601 1807 30651 1831
rect 30937 1865 30987 1889
rect 30937 1831 30945 1865
rect 30979 1831 30987 1865
rect 30937 1807 30987 1831
rect 31273 1865 31323 1889
rect 31273 1831 31281 1865
rect 31315 1831 31323 1865
rect 31273 1807 31323 1831
rect 31609 1865 31659 1889
rect 31609 1831 31617 1865
rect 31651 1831 31659 1865
rect 31609 1807 31659 1831
rect 31945 1865 31995 1889
rect 31945 1831 31953 1865
rect 31987 1831 31995 1865
rect 31945 1807 31995 1831
rect 32281 1865 32331 1889
rect 32281 1831 32289 1865
rect 32323 1831 32331 1865
rect 32281 1807 32331 1831
rect 32617 1865 32667 1889
rect 32617 1831 32625 1865
rect 32659 1831 32667 1865
rect 32617 1807 32667 1831
rect 32953 1865 33003 1889
rect 32953 1831 32961 1865
rect 32995 1831 33003 1865
rect 32953 1807 33003 1831
rect 33289 1865 33339 1889
rect 33289 1831 33297 1865
rect 33331 1831 33339 1865
rect 33289 1807 33339 1831
rect 33625 1865 33675 1889
rect 33625 1831 33633 1865
rect 33667 1831 33675 1865
rect 33625 1807 33675 1831
rect 33961 1865 34011 1889
rect 33961 1831 33969 1865
rect 34003 1831 34011 1865
rect 33961 1807 34011 1831
rect 34297 1865 34347 1889
rect 34297 1831 34305 1865
rect 34339 1831 34347 1865
rect 34297 1807 34347 1831
rect 34633 1865 34683 1889
rect 34633 1831 34641 1865
rect 34675 1831 34683 1865
rect 34633 1807 34683 1831
rect 34969 1865 35019 1889
rect 34969 1831 34977 1865
rect 35011 1831 35019 1865
rect 34969 1807 35019 1831
rect 35305 1865 35355 1889
rect 35305 1831 35313 1865
rect 35347 1831 35355 1865
rect 35305 1807 35355 1831
rect 35641 1865 35691 1889
rect 35641 1831 35649 1865
rect 35683 1831 35691 1865
rect 35641 1807 35691 1831
rect 35977 1865 36027 1889
rect 35977 1831 35985 1865
rect 36019 1831 36027 1865
rect 35977 1807 36027 1831
rect 36313 1865 36363 1889
rect 36313 1831 36321 1865
rect 36355 1831 36363 1865
rect 36313 1807 36363 1831
rect 36649 1865 36699 1889
rect 36649 1831 36657 1865
rect 36691 1831 36699 1865
rect 36649 1807 36699 1831
rect 36985 1865 37035 1889
rect 36985 1831 36993 1865
rect 37027 1831 37035 1865
rect 36985 1807 37035 1831
rect 37321 1865 37371 1889
rect 37321 1831 37329 1865
rect 37363 1831 37371 1865
rect 37321 1807 37371 1831
rect 37657 1865 37707 1889
rect 37657 1831 37665 1865
rect 37699 1831 37707 1865
rect 37657 1807 37707 1831
rect 37993 1865 38043 1889
rect 37993 1831 38001 1865
rect 38035 1831 38043 1865
rect 37993 1807 38043 1831
rect 38329 1865 38379 1889
rect 38329 1831 38337 1865
rect 38371 1831 38379 1865
rect 38329 1807 38379 1831
rect 38665 1865 38715 1889
rect 38665 1831 38673 1865
rect 38707 1831 38715 1865
rect 38665 1807 38715 1831
rect 39001 1865 39051 1889
rect 39001 1831 39009 1865
rect 39043 1831 39051 1865
rect 39001 1807 39051 1831
rect 39337 1865 39387 1889
rect 39337 1831 39345 1865
rect 39379 1831 39387 1865
rect 39337 1807 39387 1831
rect 39673 1865 39723 1889
rect 39673 1831 39681 1865
rect 39715 1831 39723 1865
rect 39673 1807 39723 1831
rect 40009 1865 40059 1889
rect 40009 1831 40017 1865
rect 40051 1831 40059 1865
rect 40009 1807 40059 1831
rect 40345 1865 40395 1889
rect 40345 1831 40353 1865
rect 40387 1831 40395 1865
rect 40345 1807 40395 1831
rect 40681 1865 40731 1889
rect 40681 1831 40689 1865
rect 40723 1831 40731 1865
rect 40681 1807 40731 1831
rect 41017 1865 41067 1889
rect 41017 1831 41025 1865
rect 41059 1831 41067 1865
rect 41017 1807 41067 1831
rect 41353 1865 41403 1889
rect 41353 1831 41361 1865
rect 41395 1831 41403 1865
rect 41353 1807 41403 1831
rect 41689 1865 41739 1889
rect 41689 1831 41697 1865
rect 41731 1831 41739 1865
rect 41689 1807 41739 1831
rect 42025 1865 42075 1889
rect 42025 1831 42033 1865
rect 42067 1831 42075 1865
rect 42025 1807 42075 1831
rect 42361 1865 42411 1889
rect 42361 1831 42369 1865
rect 42403 1831 42411 1865
rect 42361 1807 42411 1831
rect 42697 1865 42747 1889
rect 42697 1831 42705 1865
rect 42739 1831 42747 1865
rect 42697 1807 42747 1831
rect 43033 1865 43083 1889
rect 43033 1831 43041 1865
rect 43075 1831 43083 1865
rect 43033 1807 43083 1831
rect 43369 1865 43419 1889
rect 43369 1831 43377 1865
rect 43411 1831 43419 1865
rect 43369 1807 43419 1831
rect 43705 1865 43755 1889
rect 43705 1831 43713 1865
rect 43747 1831 43755 1865
rect 43705 1807 43755 1831
rect 44041 1865 44091 1889
rect 44041 1831 44049 1865
rect 44083 1831 44091 1865
rect 44041 1807 44091 1831
rect 44377 1865 44427 1889
rect 44377 1831 44385 1865
rect 44419 1831 44427 1865
rect 44377 1807 44427 1831
rect 44713 1865 44763 1889
rect 44713 1831 44721 1865
rect 44755 1831 44763 1865
rect 44713 1807 44763 1831
rect 45049 1865 45099 1889
rect 45049 1831 45057 1865
rect 45091 1831 45099 1865
rect 45049 1807 45099 1831
rect 45385 1865 45435 1889
rect 45385 1831 45393 1865
rect 45427 1831 45435 1865
rect 45385 1807 45435 1831
rect 45721 1865 45771 1889
rect 45721 1831 45729 1865
rect 45763 1831 45771 1865
rect 45721 1807 45771 1831
rect 46057 1865 46107 1889
rect 46057 1831 46065 1865
rect 46099 1831 46107 1865
rect 46057 1807 46107 1831
rect 46393 1865 46443 1889
rect 46393 1831 46401 1865
rect 46435 1831 46443 1865
rect 46393 1807 46443 1831
rect 46729 1865 46779 1889
rect 46729 1831 46737 1865
rect 46771 1831 46779 1865
rect 46729 1807 46779 1831
rect 47065 1865 47115 1889
rect 47065 1831 47073 1865
rect 47107 1831 47115 1865
rect 47065 1807 47115 1831
rect 47401 1865 47451 1889
rect 47401 1831 47409 1865
rect 47443 1831 47451 1865
rect 47401 1807 47451 1831
rect 47737 1865 47787 1889
rect 47737 1831 47745 1865
rect 47779 1831 47787 1865
rect 47737 1807 47787 1831
rect 48073 1865 48123 1889
rect 48073 1831 48081 1865
rect 48115 1831 48123 1865
rect 48073 1807 48123 1831
rect 48409 1865 48459 1889
rect 48409 1831 48417 1865
rect 48451 1831 48459 1865
rect 48409 1807 48459 1831
rect 48745 1865 48795 1889
rect 48745 1831 48753 1865
rect 48787 1831 48795 1865
rect 48745 1807 48795 1831
rect 49081 1865 49131 1889
rect 49081 1831 49089 1865
rect 49123 1831 49131 1865
rect 49081 1807 49131 1831
rect 49417 1865 49467 1889
rect 49417 1831 49425 1865
rect 49459 1831 49467 1865
rect 49417 1807 49467 1831
rect 49753 1865 49803 1889
rect 49753 1831 49761 1865
rect 49795 1831 49803 1865
rect 49753 1807 49803 1831
rect 50089 1865 50139 1889
rect 50089 1831 50097 1865
rect 50131 1831 50139 1865
rect 50089 1807 50139 1831
rect 50425 1865 50475 1889
rect 50425 1831 50433 1865
rect 50467 1831 50475 1865
rect 50425 1807 50475 1831
rect 50761 1865 50811 1889
rect 50761 1831 50769 1865
rect 50803 1831 50811 1865
rect 50761 1807 50811 1831
rect 51097 1865 51147 1889
rect 51097 1831 51105 1865
rect 51139 1831 51147 1865
rect 51097 1807 51147 1831
rect 51433 1865 51483 1889
rect 51433 1831 51441 1865
rect 51475 1831 51483 1865
rect 51433 1807 51483 1831
rect 51769 1865 51819 1889
rect 51769 1831 51777 1865
rect 51811 1831 51819 1865
rect 51769 1807 51819 1831
rect 52105 1865 52155 1889
rect 52105 1831 52113 1865
rect 52147 1831 52155 1865
rect 52105 1807 52155 1831
rect 52441 1865 52491 1889
rect 52441 1831 52449 1865
rect 52483 1831 52491 1865
rect 52441 1807 52491 1831
rect 52777 1865 52827 1889
rect 52777 1831 52785 1865
rect 52819 1831 52827 1865
rect 52777 1807 52827 1831
rect 53113 1865 53163 1889
rect 53113 1831 53121 1865
rect 53155 1831 53163 1865
rect 53113 1807 53163 1831
rect 53449 1865 53499 1889
rect 53449 1831 53457 1865
rect 53491 1831 53499 1865
rect 53449 1807 53499 1831
rect 53785 1865 53835 1889
rect 53785 1831 53793 1865
rect 53827 1831 53835 1865
rect 53785 1807 53835 1831
rect 54121 1865 54171 1889
rect 54121 1831 54129 1865
rect 54163 1831 54171 1865
rect 54121 1807 54171 1831
rect 54457 1865 54507 1889
rect 54457 1831 54465 1865
rect 54499 1831 54507 1865
rect 54457 1807 54507 1831
rect 54793 1865 54843 1889
rect 54793 1831 54801 1865
rect 54835 1831 54843 1865
rect 54793 1807 54843 1831
rect 55129 1865 55179 1889
rect 55129 1831 55137 1865
rect 55171 1831 55179 1865
rect 55129 1807 55179 1831
rect 55465 1865 55515 1889
rect 55465 1831 55473 1865
rect 55507 1831 55515 1865
rect 55465 1807 55515 1831
rect 55801 1865 55851 1889
rect 55801 1831 55809 1865
rect 55843 1831 55851 1865
rect 55801 1807 55851 1831
rect 56137 1865 56187 1889
rect 56137 1831 56145 1865
rect 56179 1831 56187 1865
rect 56137 1807 56187 1831
rect 56473 1865 56523 1889
rect 56473 1831 56481 1865
rect 56515 1831 56523 1865
rect 56473 1807 56523 1831
rect 56809 1865 56859 1889
rect 56809 1831 56817 1865
rect 56851 1831 56859 1865
rect 56809 1807 56859 1831
rect 57145 1865 57195 1889
rect 57145 1831 57153 1865
rect 57187 1831 57195 1865
rect 57145 1807 57195 1831
rect 57481 1865 57531 1889
rect 57481 1831 57489 1865
rect 57523 1831 57531 1865
rect 57481 1807 57531 1831
rect 57817 1865 57867 1889
rect 57817 1831 57825 1865
rect 57859 1831 57867 1865
rect 57817 1807 57867 1831
rect 58153 1865 58203 1889
rect 58153 1831 58161 1865
rect 58195 1831 58203 1865
rect 58153 1807 58203 1831
rect 58489 1865 58539 1889
rect 58489 1831 58497 1865
rect 58531 1831 58539 1865
rect 58489 1807 58539 1831
rect 58825 1865 58875 1889
rect 58825 1831 58833 1865
rect 58867 1831 58875 1865
rect 58825 1807 58875 1831
rect 59161 1865 59211 1889
rect 59161 1831 59169 1865
rect 59203 1831 59211 1865
rect 59161 1807 59211 1831
rect 59497 1865 59547 1889
rect 59497 1831 59505 1865
rect 59539 1831 59547 1865
rect 59497 1807 59547 1831
rect 59833 1865 59883 1889
rect 59833 1831 59841 1865
rect 59875 1831 59883 1865
rect 59833 1807 59883 1831
rect 60169 1865 60219 1889
rect 60169 1831 60177 1865
rect 60211 1831 60219 1865
rect 60169 1807 60219 1831
rect 60505 1865 60555 1889
rect 60505 1831 60513 1865
rect 60547 1831 60555 1865
rect 60505 1807 60555 1831
rect 60841 1865 60891 1889
rect 60841 1831 60849 1865
rect 60883 1831 60891 1865
rect 60841 1807 60891 1831
rect 61177 1865 61227 1889
rect 61177 1831 61185 1865
rect 61219 1831 61227 1865
rect 61177 1807 61227 1831
rect 61513 1865 61563 1889
rect 61513 1831 61521 1865
rect 61555 1831 61563 1865
rect 61513 1807 61563 1831
rect 61849 1865 61899 1889
rect 61849 1831 61857 1865
rect 61891 1831 61899 1865
rect 61849 1807 61899 1831
rect 62185 1865 62235 1889
rect 62185 1831 62193 1865
rect 62227 1831 62235 1865
rect 62185 1807 62235 1831
rect 62521 1865 62571 1889
rect 62521 1831 62529 1865
rect 62563 1831 62571 1865
rect 62521 1807 62571 1831
rect 62857 1865 62907 1889
rect 62857 1831 62865 1865
rect 62899 1831 62907 1865
rect 62857 1807 62907 1831
rect 63193 1865 63243 1889
rect 63193 1831 63201 1865
rect 63235 1831 63243 1865
rect 63193 1807 63243 1831
rect 63529 1865 63579 1889
rect 63529 1831 63537 1865
rect 63571 1831 63579 1865
rect 63529 1807 63579 1831
rect 63865 1865 63915 1889
rect 63865 1831 63873 1865
rect 63907 1831 63915 1865
rect 63865 1807 63915 1831
rect 64201 1865 64251 1889
rect 64201 1831 64209 1865
rect 64243 1831 64251 1865
rect 64201 1807 64251 1831
rect 64537 1865 64587 1889
rect 64537 1831 64545 1865
rect 64579 1831 64587 1865
rect 64537 1807 64587 1831
rect 64873 1865 64923 1889
rect 64873 1831 64881 1865
rect 64915 1831 64923 1865
rect 64873 1807 64923 1831
rect 65209 1865 65259 1889
rect 65209 1831 65217 1865
rect 65251 1831 65259 1865
rect 65209 1807 65259 1831
rect 65545 1865 65595 1889
rect 65545 1831 65553 1865
rect 65587 1831 65595 1865
rect 65545 1807 65595 1831
rect 65881 1865 65931 1889
rect 65881 1831 65889 1865
rect 65923 1831 65931 1865
rect 65881 1807 65931 1831
rect 66217 1865 66267 1889
rect 66217 1831 66225 1865
rect 66259 1831 66267 1865
rect 66217 1807 66267 1831
rect 66553 1865 66603 1889
rect 66553 1831 66561 1865
rect 66595 1831 66603 1865
rect 66553 1807 66603 1831
rect 66889 1865 66939 1889
rect 66889 1831 66897 1865
rect 66931 1831 66939 1865
rect 66889 1807 66939 1831
rect 67225 1865 67275 1889
rect 67225 1831 67233 1865
rect 67267 1831 67275 1865
rect 67225 1807 67275 1831
rect 67561 1865 67611 1889
rect 67561 1831 67569 1865
rect 67603 1831 67611 1865
rect 67561 1807 67611 1831
rect 67897 1865 67947 1889
rect 67897 1831 67905 1865
rect 67939 1831 67947 1865
rect 67897 1807 67947 1831
rect 68233 1865 68283 1889
rect 68233 1831 68241 1865
rect 68275 1831 68283 1865
rect 68233 1807 68283 1831
rect 68569 1865 68619 1889
rect 68569 1831 68577 1865
rect 68611 1831 68619 1865
rect 68569 1807 68619 1831
rect 68905 1865 68955 1889
rect 68905 1831 68913 1865
rect 68947 1831 68955 1865
rect 68905 1807 68955 1831
rect 69241 1865 69291 1889
rect 69241 1831 69249 1865
rect 69283 1831 69291 1865
rect 69241 1807 69291 1831
rect 69577 1865 69627 1889
rect 69577 1831 69585 1865
rect 69619 1831 69627 1865
rect 69577 1807 69627 1831
rect 69913 1865 69963 1889
rect 69913 1831 69921 1865
rect 69955 1831 69963 1865
rect 69913 1807 69963 1831
rect 70249 1865 70299 1889
rect 70249 1831 70257 1865
rect 70291 1831 70299 1865
rect 70249 1807 70299 1831
rect 70585 1865 70635 1889
rect 70585 1831 70593 1865
rect 70627 1831 70635 1865
rect 70585 1807 70635 1831
rect 70921 1865 70971 1889
rect 70921 1831 70929 1865
rect 70963 1831 70971 1865
rect 70921 1807 70971 1831
rect 71257 1865 71307 1889
rect 71257 1831 71265 1865
rect 71299 1831 71307 1865
rect 71257 1807 71307 1831
rect 71593 1865 71643 1889
rect 71593 1831 71601 1865
rect 71635 1831 71643 1865
rect 71593 1807 71643 1831
rect 71929 1865 71979 1889
rect 71929 1831 71937 1865
rect 71971 1831 71979 1865
rect 71929 1807 71979 1831
rect 72265 1865 72315 1889
rect 72265 1831 72273 1865
rect 72307 1831 72315 1865
rect 72265 1807 72315 1831
rect 72601 1865 72651 1889
rect 72601 1831 72609 1865
rect 72643 1831 72651 1865
rect 72601 1807 72651 1831
rect 72937 1865 72987 1889
rect 72937 1831 72945 1865
rect 72979 1831 72987 1865
rect 72937 1807 72987 1831
rect 73273 1865 73323 1889
rect 73273 1831 73281 1865
rect 73315 1831 73323 1865
rect 73273 1807 73323 1831
rect 73609 1865 73659 1889
rect 73609 1831 73617 1865
rect 73651 1831 73659 1865
rect 73609 1807 73659 1831
rect 73945 1865 73995 1889
rect 73945 1831 73953 1865
rect 73987 1831 73995 1865
rect 73945 1807 73995 1831
rect 74281 1865 74331 1889
rect 74281 1831 74289 1865
rect 74323 1831 74331 1865
rect 74281 1807 74331 1831
rect 74617 1865 74667 1889
rect 74617 1831 74625 1865
rect 74659 1831 74667 1865
rect 74617 1807 74667 1831
rect 74953 1865 75003 1889
rect 74953 1831 74961 1865
rect 74995 1831 75003 1865
rect 74953 1807 75003 1831
rect 75289 1865 75339 1889
rect 75289 1831 75297 1865
rect 75331 1831 75339 1865
rect 75289 1807 75339 1831
rect 75625 1865 75675 1889
rect 75625 1831 75633 1865
rect 75667 1831 75675 1865
rect 75625 1807 75675 1831
rect 75961 1865 76011 1889
rect 75961 1831 75969 1865
rect 76003 1831 76011 1865
rect 75961 1807 76011 1831
rect 76297 1865 76347 1889
rect 76297 1831 76305 1865
rect 76339 1831 76347 1865
rect 76297 1807 76347 1831
rect 76633 1865 76683 1889
rect 76633 1831 76641 1865
rect 76675 1831 76683 1865
rect 76633 1807 76683 1831
rect 76969 1865 77019 1889
rect 76969 1831 76977 1865
rect 77011 1831 77019 1865
rect 76969 1807 77019 1831
rect 77305 1865 77355 1889
rect 77305 1831 77313 1865
rect 77347 1831 77355 1865
rect 77305 1807 77355 1831
rect 77641 1865 77691 1889
rect 77641 1831 77649 1865
rect 77683 1831 77691 1865
rect 77641 1807 77691 1831
rect 77977 1865 78027 1889
rect 77977 1831 77985 1865
rect 78019 1831 78027 1865
rect 77977 1807 78027 1831
rect 78313 1865 78363 1889
rect 78313 1831 78321 1865
rect 78355 1831 78363 1865
rect 78313 1807 78363 1831
rect 78649 1865 78699 1889
rect 78649 1831 78657 1865
rect 78691 1831 78699 1865
rect 78649 1807 78699 1831
rect 78985 1865 79035 1889
rect 78985 1831 78993 1865
rect 79027 1831 79035 1865
rect 78985 1807 79035 1831
rect 79321 1865 79371 1889
rect 79321 1831 79329 1865
rect 79363 1831 79371 1865
rect 79321 1807 79371 1831
rect 79657 1865 79707 1889
rect 79657 1831 79665 1865
rect 79699 1831 79707 1865
rect 79657 1807 79707 1831
rect 79993 1865 80043 1889
rect 79993 1831 80001 1865
rect 80035 1831 80043 1865
rect 79993 1807 80043 1831
rect 80329 1865 80379 1889
rect 80329 1831 80337 1865
rect 80371 1831 80379 1865
rect 80329 1807 80379 1831
rect 80665 1865 80715 1889
rect 80665 1831 80673 1865
rect 80707 1831 80715 1865
rect 80665 1807 80715 1831
rect 81001 1865 81051 1889
rect 81001 1831 81009 1865
rect 81043 1831 81051 1865
rect 81001 1807 81051 1831
rect 81337 1865 81387 1889
rect 81337 1831 81345 1865
rect 81379 1831 81387 1865
rect 81337 1807 81387 1831
rect 81673 1865 81723 1889
rect 81673 1831 81681 1865
rect 81715 1831 81723 1865
rect 81673 1807 81723 1831
rect 82009 1865 82059 1889
rect 82009 1831 82017 1865
rect 82051 1831 82059 1865
rect 82009 1807 82059 1831
rect 82345 1865 82395 1889
rect 82345 1831 82353 1865
rect 82387 1831 82395 1865
rect 82345 1807 82395 1831
rect 82681 1865 82731 1889
rect 82681 1831 82689 1865
rect 82723 1831 82731 1865
rect 82681 1807 82731 1831
rect 83017 1865 83067 1889
rect 83017 1831 83025 1865
rect 83059 1831 83067 1865
rect 83017 1807 83067 1831
rect 83353 1865 83403 1889
rect 83353 1831 83361 1865
rect 83395 1831 83403 1865
rect 83353 1807 83403 1831
rect 83689 1865 83739 1889
rect 83689 1831 83697 1865
rect 83731 1831 83739 1865
rect 83689 1807 83739 1831
rect 84025 1865 84075 1889
rect 84025 1831 84033 1865
rect 84067 1831 84075 1865
rect 84025 1807 84075 1831
rect 84361 1865 84411 1889
rect 84361 1831 84369 1865
rect 84403 1831 84411 1865
rect 84361 1807 84411 1831
rect 84697 1865 84747 1889
rect 84697 1831 84705 1865
rect 84739 1831 84747 1865
rect 84697 1807 84747 1831
rect 85033 1865 85083 1889
rect 85033 1831 85041 1865
rect 85075 1831 85083 1865
rect 85033 1807 85083 1831
rect 85369 1865 85419 1889
rect 85369 1831 85377 1865
rect 85411 1831 85419 1865
rect 85369 1807 85419 1831
rect 85705 1865 85755 1889
rect 85705 1831 85713 1865
rect 85747 1831 85755 1865
rect 85705 1807 85755 1831
rect 86041 1865 86091 1889
rect 86041 1831 86049 1865
rect 86083 1831 86091 1865
rect 86041 1807 86091 1831
rect 86377 1865 86427 1889
rect 86377 1831 86385 1865
rect 86419 1831 86427 1865
rect 86377 1807 86427 1831
rect 86713 1865 86763 1889
rect 86713 1831 86721 1865
rect 86755 1831 86763 1865
rect 86713 1807 86763 1831
rect 87049 1865 87099 1889
rect 87049 1831 87057 1865
rect 87091 1831 87099 1865
rect 87049 1807 87099 1831
rect 87385 1865 87435 1889
rect 87385 1831 87393 1865
rect 87427 1831 87435 1865
rect 87385 1807 87435 1831
rect 87721 1865 87771 1889
rect 87721 1831 87729 1865
rect 87763 1831 87771 1865
rect 87721 1807 87771 1831
rect 88057 1865 88107 1889
rect 88057 1831 88065 1865
rect 88099 1831 88107 1865
rect 88057 1807 88107 1831
rect 88393 1865 88443 1889
rect 88393 1831 88401 1865
rect 88435 1831 88443 1865
rect 88393 1807 88443 1831
rect 88729 1865 88779 1889
rect 88729 1831 88737 1865
rect 88771 1831 88779 1865
rect 88729 1807 88779 1831
rect 89065 1865 89115 1889
rect 89065 1831 89073 1865
rect 89107 1831 89115 1865
rect 89065 1807 89115 1831
rect 89401 1865 89451 1889
rect 89401 1831 89409 1865
rect 89443 1831 89451 1865
rect 89401 1807 89451 1831
rect 89737 1865 89787 1889
rect 89737 1831 89745 1865
rect 89779 1831 89787 1865
rect 89737 1807 89787 1831
rect 90073 1865 90123 1889
rect 90073 1831 90081 1865
rect 90115 1831 90123 1865
rect 90073 1807 90123 1831
rect 90409 1865 90459 1889
rect 90409 1831 90417 1865
rect 90451 1831 90459 1865
rect 90409 1807 90459 1831
rect 90745 1865 90795 1889
rect 90745 1831 90753 1865
rect 90787 1831 90795 1865
rect 90745 1807 90795 1831
rect 91081 1865 91131 1889
rect 91081 1831 91089 1865
rect 91123 1831 91131 1865
rect 91081 1807 91131 1831
rect 91417 1865 91467 1889
rect 91417 1831 91425 1865
rect 91459 1831 91467 1865
rect 91417 1807 91467 1831
rect 91753 1865 91803 1889
rect 91753 1831 91761 1865
rect 91795 1831 91803 1865
rect 91753 1807 91803 1831
rect 92089 1865 92139 1889
rect 92089 1831 92097 1865
rect 92131 1831 92139 1865
rect 92089 1807 92139 1831
rect 92425 1865 92475 1889
rect 92425 1831 92433 1865
rect 92467 1831 92475 1865
rect 92425 1807 92475 1831
rect 92761 1865 92811 1889
rect 92761 1831 92769 1865
rect 92803 1831 92811 1865
rect 92761 1807 92811 1831
rect 93097 1865 93147 1889
rect 93097 1831 93105 1865
rect 93139 1831 93147 1865
rect 93097 1807 93147 1831
rect 93433 1865 93483 1889
rect 93433 1831 93441 1865
rect 93475 1831 93483 1865
rect 93433 1807 93483 1831
rect 93769 1865 93819 1889
rect 93769 1831 93777 1865
rect 93811 1831 93819 1865
rect 93769 1807 93819 1831
rect 94105 1865 94155 1889
rect 94105 1831 94113 1865
rect 94147 1831 94155 1865
rect 94105 1807 94155 1831
rect 94441 1865 94491 1889
rect 94441 1831 94449 1865
rect 94483 1831 94491 1865
rect 94441 1807 94491 1831
rect 94777 1865 94827 1889
rect 94777 1831 94785 1865
rect 94819 1831 94827 1865
rect 94777 1807 94827 1831
rect 95113 1865 95163 1889
rect 95113 1831 95121 1865
rect 95155 1831 95163 1865
rect 95113 1807 95163 1831
rect 95449 1865 95499 1889
rect 95449 1831 95457 1865
rect 95491 1831 95499 1865
rect 95449 1807 95499 1831
rect 95785 1865 95835 1889
rect 95785 1831 95793 1865
rect 95827 1831 95835 1865
rect 95785 1807 95835 1831
rect 96121 1865 96171 1889
rect 96121 1831 96129 1865
rect 96163 1831 96171 1865
rect 96121 1807 96171 1831
rect 96457 1865 96507 1889
rect 96457 1831 96465 1865
rect 96499 1831 96507 1865
rect 96457 1807 96507 1831
rect 96793 1865 96843 1889
rect 96793 1831 96801 1865
rect 96835 1831 96843 1865
rect 96793 1807 96843 1831
rect 97129 1865 97179 1889
rect 97129 1831 97137 1865
rect 97171 1831 97179 1865
rect 97129 1807 97179 1831
rect 97465 1865 97515 1889
rect 97465 1831 97473 1865
rect 97507 1831 97515 1865
rect 97465 1807 97515 1831
rect 97801 1865 97851 1889
rect 97801 1831 97809 1865
rect 97843 1831 97851 1865
rect 97801 1807 97851 1831
rect 98137 1865 98187 1889
rect 98137 1831 98145 1865
rect 98179 1831 98187 1865
rect 98137 1807 98187 1831
rect 98473 1865 98523 1889
rect 98473 1831 98481 1865
rect 98515 1831 98523 1865
rect 98473 1807 98523 1831
rect 98809 1865 98859 1889
rect 98809 1831 98817 1865
rect 98851 1831 98859 1865
rect 98809 1807 98859 1831
rect 99145 1865 99195 1889
rect 99145 1831 99153 1865
rect 99187 1831 99195 1865
rect 99145 1807 99195 1831
rect 99481 1865 99531 1889
rect 99481 1831 99489 1865
rect 99523 1831 99531 1865
rect 99481 1807 99531 1831
rect 99817 1865 99867 1889
rect 99817 1831 99825 1865
rect 99859 1831 99867 1865
rect 99817 1807 99867 1831
rect 100153 1865 100203 1889
rect 100153 1831 100161 1865
rect 100195 1831 100203 1865
rect 100153 1807 100203 1831
rect 100489 1865 100539 1889
rect 100489 1831 100497 1865
rect 100531 1831 100539 1865
rect 100489 1807 100539 1831
rect 100825 1865 100875 1889
rect 100825 1831 100833 1865
rect 100867 1831 100875 1865
rect 100825 1807 100875 1831
rect 101161 1865 101211 1889
rect 101161 1831 101169 1865
rect 101203 1831 101211 1865
rect 101161 1807 101211 1831
rect 101497 1865 101547 1889
rect 101497 1831 101505 1865
rect 101539 1831 101547 1865
rect 101497 1807 101547 1831
rect 101833 1865 101883 1889
rect 101833 1831 101841 1865
rect 101875 1831 101883 1865
rect 101833 1807 101883 1831
rect 102169 1865 102219 1889
rect 102169 1831 102177 1865
rect 102211 1831 102219 1865
rect 102169 1807 102219 1831
rect 102505 1865 102555 1889
rect 102505 1831 102513 1865
rect 102547 1831 102555 1865
rect 102505 1807 102555 1831
rect 102841 1865 102891 1889
rect 102841 1831 102849 1865
rect 102883 1831 102891 1865
rect 102841 1807 102891 1831
rect 103177 1865 103227 1889
rect 103177 1831 103185 1865
rect 103219 1831 103227 1865
rect 103177 1807 103227 1831
rect 103513 1865 103563 1889
rect 103513 1831 103521 1865
rect 103555 1831 103563 1865
rect 103513 1807 103563 1831
rect 103849 1865 103899 1889
rect 103849 1831 103857 1865
rect 103891 1831 103899 1865
rect 103849 1807 103899 1831
rect 104185 1865 104235 1889
rect 104185 1831 104193 1865
rect 104227 1831 104235 1865
rect 104185 1807 104235 1831
rect 104521 1865 104571 1889
rect 104521 1831 104529 1865
rect 104563 1831 104571 1865
rect 104521 1807 104571 1831
rect 104857 1865 104907 1889
rect 104857 1831 104865 1865
rect 104899 1831 104907 1865
rect 104857 1807 104907 1831
rect 105193 1865 105243 1889
rect 105193 1831 105201 1865
rect 105235 1831 105243 1865
rect 105193 1807 105243 1831
rect 105529 1865 105579 1889
rect 105529 1831 105537 1865
rect 105571 1831 105579 1865
rect 105529 1807 105579 1831
rect 105865 1865 105915 1889
rect 105865 1831 105873 1865
rect 105907 1831 105915 1865
rect 105865 1807 105915 1831
rect 106201 1865 106251 1889
rect 106201 1831 106209 1865
rect 106243 1831 106251 1865
rect 106201 1807 106251 1831
rect 106537 1865 106587 1889
rect 106537 1831 106545 1865
rect 106579 1831 106587 1865
rect 106537 1807 106587 1831
rect 106873 1865 106923 1889
rect 106873 1831 106881 1865
rect 106915 1831 106923 1865
rect 106873 1807 106923 1831
rect 107209 1865 107259 1889
rect 107209 1831 107217 1865
rect 107251 1831 107259 1865
rect 107209 1807 107259 1831
rect 107545 1865 107595 1889
rect 107545 1831 107553 1865
rect 107587 1831 107595 1865
rect 107545 1807 107595 1831
rect 107881 1865 107931 1889
rect 107881 1831 107889 1865
rect 107923 1831 107931 1865
rect 107881 1807 107931 1831
rect 108217 1865 108267 1889
rect 108217 1831 108225 1865
rect 108259 1831 108267 1865
rect 108217 1807 108267 1831
rect 108553 1865 108603 1889
rect 108553 1831 108561 1865
rect 108595 1831 108603 1865
rect 108553 1807 108603 1831
rect 108889 1865 108939 1889
rect 108889 1831 108897 1865
rect 108931 1831 108939 1865
rect 108889 1807 108939 1831
rect 109225 1865 109275 1889
rect 109225 1831 109233 1865
rect 109267 1831 109275 1865
rect 109225 1807 109275 1831
rect 109561 1865 109611 1889
rect 109561 1831 109569 1865
rect 109603 1831 109611 1865
rect 109561 1807 109611 1831
rect 109897 1865 109947 1889
rect 109897 1831 109905 1865
rect 109939 1831 109947 1865
rect 109897 1807 109947 1831
rect 110233 1865 110283 1889
rect 110233 1831 110241 1865
rect 110275 1831 110283 1865
rect 110233 1807 110283 1831
rect 110569 1865 110619 1889
rect 110569 1831 110577 1865
rect 110611 1831 110619 1865
rect 110569 1807 110619 1831
rect 110905 1865 110955 1889
rect 110905 1831 110913 1865
rect 110947 1831 110955 1865
rect 110905 1807 110955 1831
rect 111241 1865 111291 1889
rect 111241 1831 111249 1865
rect 111283 1831 111291 1865
rect 111241 1807 111291 1831
rect 111577 1865 111627 1889
rect 111577 1831 111585 1865
rect 111619 1831 111627 1865
rect 111577 1807 111627 1831
rect 111913 1865 111963 1889
rect 111913 1831 111921 1865
rect 111955 1831 111963 1865
rect 111913 1807 111963 1831
rect 112249 1865 112299 1889
rect 112249 1831 112257 1865
rect 112291 1831 112299 1865
rect 112249 1807 112299 1831
rect 112585 1865 112635 1889
rect 112585 1831 112593 1865
rect 112627 1831 112635 1865
rect 112585 1807 112635 1831
rect 112921 1865 112971 1889
rect 112921 1831 112929 1865
rect 112963 1831 112971 1865
rect 112921 1807 112971 1831
rect 113257 1865 113307 1889
rect 113257 1831 113265 1865
rect 113299 1831 113307 1865
rect 113257 1807 113307 1831
rect 113593 1865 113643 1889
rect 113593 1831 113601 1865
rect 113635 1831 113643 1865
rect 113593 1807 113643 1831
rect 113929 1865 113979 1889
rect 113929 1831 113937 1865
rect 113971 1831 113979 1865
rect 113929 1807 113979 1831
rect 114265 1865 114315 1889
rect 114265 1831 114273 1865
rect 114307 1831 114315 1865
rect 114265 1807 114315 1831
rect 114601 1865 114651 1889
rect 114601 1831 114609 1865
rect 114643 1831 114651 1865
rect 114601 1807 114651 1831
rect 114937 1865 114987 1889
rect 114937 1831 114945 1865
rect 114979 1831 114987 1865
rect 114937 1807 114987 1831
rect 115273 1865 115323 1889
rect 115273 1831 115281 1865
rect 115315 1831 115323 1865
rect 115273 1807 115323 1831
rect 115609 1865 115659 1889
rect 115609 1831 115617 1865
rect 115651 1831 115659 1865
rect 115609 1807 115659 1831
rect 115945 1865 115995 1889
rect 115945 1831 115953 1865
rect 115987 1831 115995 1865
rect 115945 1807 115995 1831
rect 116281 1865 116331 1889
rect 116281 1831 116289 1865
rect 116323 1831 116331 1865
rect 116281 1807 116331 1831
rect 116617 1865 116667 1889
rect 116617 1831 116625 1865
rect 116659 1831 116667 1865
rect 116617 1807 116667 1831
rect 116953 1865 117003 1889
rect 116953 1831 116961 1865
rect 116995 1831 117003 1865
rect 116953 1807 117003 1831
rect 117289 1865 117339 1889
rect 117289 1831 117297 1865
rect 117331 1831 117339 1865
rect 117289 1807 117339 1831
rect 117625 1865 117675 1889
rect 117625 1831 117633 1865
rect 117667 1831 117675 1865
rect 117625 1807 117675 1831
rect 117961 1865 118011 1889
rect 117961 1831 117969 1865
rect 118003 1831 118011 1865
rect 117961 1807 118011 1831
rect 118297 1865 118347 1889
rect 118297 1831 118305 1865
rect 118339 1831 118347 1865
rect 118297 1807 118347 1831
rect 118633 1865 118683 1889
rect 118633 1831 118641 1865
rect 118675 1831 118683 1865
rect 118633 1807 118683 1831
rect 118969 1865 119019 1889
rect 118969 1831 118977 1865
rect 119011 1831 119019 1865
rect 118969 1807 119019 1831
rect 119305 1865 119355 1889
rect 119305 1831 119313 1865
rect 119347 1831 119355 1865
rect 119305 1807 119355 1831
rect 119641 1865 119691 1889
rect 119641 1831 119649 1865
rect 119683 1831 119691 1865
rect 119641 1807 119691 1831
rect 119977 1865 120027 1889
rect 119977 1831 119985 1865
rect 120019 1831 120027 1865
rect 119977 1807 120027 1831
rect 120313 1865 120363 1889
rect 120313 1831 120321 1865
rect 120355 1831 120363 1865
rect 120313 1807 120363 1831
rect 120649 1865 120699 1889
rect 120649 1831 120657 1865
rect 120691 1831 120699 1865
rect 120649 1807 120699 1831
rect 120985 1865 121035 1889
rect 120985 1831 120993 1865
rect 121027 1831 121035 1865
rect 120985 1807 121035 1831
rect 121321 1865 121371 1889
rect 121321 1831 121329 1865
rect 121363 1831 121371 1865
rect 121321 1807 121371 1831
rect 121657 1865 121707 1889
rect 121657 1831 121665 1865
rect 121699 1831 121707 1865
rect 121657 1807 121707 1831
rect 121993 1865 122043 1889
rect 121993 1831 122001 1865
rect 122035 1831 122043 1865
rect 121993 1807 122043 1831
rect 122329 1865 122379 1889
rect 122329 1831 122337 1865
rect 122371 1831 122379 1865
rect 122329 1807 122379 1831
rect 122665 1865 122715 1889
rect 122665 1831 122673 1865
rect 122707 1831 122715 1865
rect 122665 1807 122715 1831
rect 123001 1865 123051 1889
rect 123001 1831 123009 1865
rect 123043 1831 123051 1865
rect 123001 1807 123051 1831
rect 123337 1865 123387 1889
rect 123337 1831 123345 1865
rect 123379 1831 123387 1865
rect 123337 1807 123387 1831
rect 123673 1865 123723 1889
rect 123673 1831 123681 1865
rect 123715 1831 123723 1865
rect 123673 1807 123723 1831
rect 124009 1865 124059 1889
rect 124009 1831 124017 1865
rect 124051 1831 124059 1865
rect 124009 1807 124059 1831
rect 124345 1865 124395 1889
rect 124345 1831 124353 1865
rect 124387 1831 124395 1865
rect 124345 1807 124395 1831
rect 124681 1865 124731 1889
rect 124681 1831 124689 1865
rect 124723 1831 124731 1865
rect 124681 1807 124731 1831
rect 125017 1865 125067 1889
rect 125017 1831 125025 1865
rect 125059 1831 125067 1865
rect 125017 1807 125067 1831
rect 125353 1865 125403 1889
rect 125353 1831 125361 1865
rect 125395 1831 125403 1865
rect 125353 1807 125403 1831
rect 125689 1865 125739 1889
rect 125689 1831 125697 1865
rect 125731 1831 125739 1865
rect 125689 1807 125739 1831
rect 126025 1865 126075 1889
rect 126025 1831 126033 1865
rect 126067 1831 126075 1865
rect 126025 1807 126075 1831
rect 126361 1865 126411 1889
rect 126361 1831 126369 1865
rect 126403 1831 126411 1865
rect 126361 1807 126411 1831
rect 126697 1865 126747 1889
rect 126697 1831 126705 1865
rect 126739 1831 126747 1865
rect 126697 1807 126747 1831
rect 127033 1865 127083 1889
rect 127033 1831 127041 1865
rect 127075 1831 127083 1865
rect 127033 1807 127083 1831
rect 127369 1865 127419 1889
rect 127369 1831 127377 1865
rect 127411 1831 127419 1865
rect 127369 1807 127419 1831
rect 127705 1865 127755 1889
rect 127705 1831 127713 1865
rect 127747 1831 127755 1865
rect 127705 1807 127755 1831
rect 128041 1865 128091 1889
rect 128041 1831 128049 1865
rect 128083 1831 128091 1865
rect 128041 1807 128091 1831
rect 128377 1865 128427 1889
rect 128377 1831 128385 1865
rect 128419 1831 128427 1865
rect 128377 1807 128427 1831
rect 128713 1865 128763 1889
rect 128713 1831 128721 1865
rect 128755 1831 128763 1865
rect 128713 1807 128763 1831
rect 129049 1865 129099 1889
rect 129049 1831 129057 1865
rect 129091 1831 129099 1865
rect 129049 1807 129099 1831
rect 129385 1865 129435 1889
rect 129385 1831 129393 1865
rect 129427 1831 129435 1865
rect 129385 1807 129435 1831
rect 129721 1865 129771 1889
rect 129721 1831 129729 1865
rect 129763 1831 129771 1865
rect 129721 1807 129771 1831
rect 130057 1865 130107 1889
rect 130057 1831 130065 1865
rect 130099 1831 130107 1865
rect 130057 1807 130107 1831
rect 130393 1865 130443 1889
rect 130393 1831 130401 1865
rect 130435 1831 130443 1865
rect 130393 1807 130443 1831
rect 130729 1865 130779 1889
rect 130729 1831 130737 1865
rect 130771 1831 130779 1865
rect 130729 1807 130779 1831
rect 131065 1865 131115 1889
rect 131065 1831 131073 1865
rect 131107 1831 131115 1865
rect 131065 1807 131115 1831
rect 131401 1865 131451 1889
rect 131401 1831 131409 1865
rect 131443 1831 131451 1865
rect 131401 1807 131451 1831
rect 131737 1865 131787 1889
rect 131737 1831 131745 1865
rect 131779 1831 131787 1865
rect 131737 1807 131787 1831
rect 132073 1865 132123 1889
rect 132073 1831 132081 1865
rect 132115 1831 132123 1865
rect 132073 1807 132123 1831
rect 132409 1865 132459 1889
rect 132409 1831 132417 1865
rect 132451 1831 132459 1865
rect 132409 1807 132459 1831
rect 132745 1865 132795 1889
rect 132745 1831 132753 1865
rect 132787 1831 132795 1865
rect 132745 1807 132795 1831
rect 133081 1865 133131 1889
rect 133081 1831 133089 1865
rect 133123 1831 133131 1865
rect 133081 1807 133131 1831
rect 133417 1865 133467 1889
rect 133417 1831 133425 1865
rect 133459 1831 133467 1865
rect 133417 1807 133467 1831
rect 133753 1865 133803 1889
rect 133753 1831 133761 1865
rect 133795 1831 133803 1865
rect 133753 1807 133803 1831
rect 134089 1865 134139 1889
rect 134089 1831 134097 1865
rect 134131 1831 134139 1865
rect 134089 1807 134139 1831
rect 134425 1865 134475 1889
rect 134425 1831 134433 1865
rect 134467 1831 134475 1865
rect 134425 1807 134475 1831
rect 134761 1865 134811 1889
rect 134761 1831 134769 1865
rect 134803 1831 134811 1865
rect 134761 1807 134811 1831
rect 135097 1865 135147 1889
rect 135097 1831 135105 1865
rect 135139 1831 135147 1865
rect 135097 1807 135147 1831
rect 135433 1865 135483 1889
rect 135433 1831 135441 1865
rect 135475 1831 135483 1865
rect 135433 1807 135483 1831
rect 135769 1865 135819 1889
rect 135769 1831 135777 1865
rect 135811 1831 135819 1865
rect 135769 1807 135819 1831
rect 136105 1865 136155 1889
rect 136105 1831 136113 1865
rect 136147 1831 136155 1865
rect 136105 1807 136155 1831
rect 136441 1865 136491 1889
rect 136441 1831 136449 1865
rect 136483 1831 136491 1865
rect 136441 1807 136491 1831
rect 136777 1865 136827 1889
rect 136777 1831 136785 1865
rect 136819 1831 136827 1865
rect 136777 1807 136827 1831
rect 137113 1865 137163 1889
rect 137113 1831 137121 1865
rect 137155 1831 137163 1865
rect 137113 1807 137163 1831
rect 137449 1865 137499 1889
rect 137449 1831 137457 1865
rect 137491 1831 137499 1865
rect 137449 1807 137499 1831
rect 137785 1865 137835 1889
rect 137785 1831 137793 1865
rect 137827 1831 137835 1865
rect 137785 1807 137835 1831
rect 138121 1865 138171 1889
rect 138121 1831 138129 1865
rect 138163 1831 138171 1865
rect 138121 1807 138171 1831
rect 138457 1865 138507 1889
rect 138457 1831 138465 1865
rect 138499 1831 138507 1865
rect 138457 1807 138507 1831
rect 138793 1865 138843 1889
rect 138793 1831 138801 1865
rect 138835 1831 138843 1865
rect 138793 1807 138843 1831
rect 139129 1865 139179 1889
rect 139129 1831 139137 1865
rect 139171 1831 139179 1865
rect 139129 1807 139179 1831
rect 139465 1865 139515 1889
rect 139465 1831 139473 1865
rect 139507 1831 139515 1865
rect 139465 1807 139515 1831
rect 139801 1865 139851 1889
rect 139801 1831 139809 1865
rect 139843 1831 139851 1865
rect 139801 1807 139851 1831
rect 140137 1865 140187 1889
rect 140137 1831 140145 1865
rect 140179 1831 140187 1865
rect 140137 1807 140187 1831
rect 140473 1865 140523 1889
rect 140473 1831 140481 1865
rect 140515 1831 140523 1865
rect 140473 1807 140523 1831
rect 140809 1865 140859 1889
rect 140809 1831 140817 1865
rect 140851 1831 140859 1865
rect 140809 1807 140859 1831
rect 141145 1865 141195 1889
rect 141145 1831 141153 1865
rect 141187 1831 141195 1865
rect 141145 1807 141195 1831
rect 141481 1865 141531 1889
rect 141481 1831 141489 1865
rect 141523 1831 141531 1865
rect 141481 1807 141531 1831
rect 141817 1865 141867 1889
rect 141817 1831 141825 1865
rect 141859 1831 141867 1865
rect 141817 1807 141867 1831
rect 142153 1865 142203 1889
rect 142153 1831 142161 1865
rect 142195 1831 142203 1865
rect 142153 1807 142203 1831
rect 142489 1865 142539 1889
rect 142489 1831 142497 1865
rect 142531 1831 142539 1865
rect 142489 1807 142539 1831
rect 142825 1865 142875 1889
rect 142825 1831 142833 1865
rect 142867 1831 142875 1865
rect 142825 1807 142875 1831
rect 143161 1865 143211 1889
rect 143161 1831 143169 1865
rect 143203 1831 143211 1865
rect 143161 1807 143211 1831
rect 143497 1865 143547 1889
rect 143497 1831 143505 1865
rect 143539 1831 143547 1865
rect 143497 1807 143547 1831
rect 143833 1865 143883 1889
rect 143833 1831 143841 1865
rect 143875 1831 143883 1865
rect 143833 1807 143883 1831
rect 144169 1865 144219 1889
rect 144169 1831 144177 1865
rect 144211 1831 144219 1865
rect 144169 1807 144219 1831
rect 144505 1865 144555 1889
rect 144505 1831 144513 1865
rect 144547 1831 144555 1865
rect 144505 1807 144555 1831
rect 144841 1865 144891 1889
rect 144841 1831 144849 1865
rect 144883 1831 144891 1865
rect 144841 1807 144891 1831
rect 145177 1865 145227 1889
rect 145177 1831 145185 1865
rect 145219 1831 145227 1865
rect 145177 1807 145227 1831
rect 145513 1865 145563 1889
rect 145513 1831 145521 1865
rect 145555 1831 145563 1865
rect 145513 1807 145563 1831
rect 145849 1865 145899 1889
rect 145849 1831 145857 1865
rect 145891 1831 145899 1865
rect 145849 1807 145899 1831
rect 146185 1865 146235 1889
rect 146185 1831 146193 1865
rect 146227 1831 146235 1865
rect 146185 1807 146235 1831
rect 146521 1865 146571 1889
rect 146521 1831 146529 1865
rect 146563 1831 146571 1865
rect 146521 1807 146571 1831
rect 146857 1865 146907 1889
rect 146857 1831 146865 1865
rect 146899 1831 146907 1865
rect 146857 1807 146907 1831
rect 147193 1865 147243 1889
rect 147193 1831 147201 1865
rect 147235 1831 147243 1865
rect 147193 1807 147243 1831
rect 147529 1865 147579 1889
rect 147529 1831 147537 1865
rect 147571 1831 147579 1865
rect 147529 1807 147579 1831
rect 147865 1865 147915 1889
rect 147865 1831 147873 1865
rect 147907 1831 147915 1865
rect 147865 1807 147915 1831
rect 148201 1865 148251 1889
rect 148201 1831 148209 1865
rect 148243 1831 148251 1865
rect 148201 1807 148251 1831
rect 148537 1865 148587 1889
rect 148537 1831 148545 1865
rect 148579 1831 148587 1865
rect 148537 1807 148587 1831
rect 148873 1865 148923 1889
rect 148873 1831 148881 1865
rect 148915 1831 148923 1865
rect 148873 1807 148923 1831
rect 149209 1865 149259 1889
rect 149209 1831 149217 1865
rect 149251 1831 149259 1865
rect 149209 1807 149259 1831
rect 149545 1865 149595 1889
rect 149545 1831 149553 1865
rect 149587 1831 149595 1865
rect 149545 1807 149595 1831
rect 149881 1865 149931 1889
rect 149881 1831 149889 1865
rect 149923 1831 149931 1865
rect 149881 1807 149931 1831
rect 150217 1865 150267 1889
rect 150217 1831 150225 1865
rect 150259 1831 150267 1865
rect 150217 1807 150267 1831
rect 150553 1865 150603 1889
rect 150553 1831 150561 1865
rect 150595 1831 150603 1865
rect 150553 1807 150603 1831
rect 150889 1865 150939 1889
rect 150889 1831 150897 1865
rect 150931 1831 150939 1865
rect 150889 1807 150939 1831
rect 151225 1865 151275 1889
rect 151225 1831 151233 1865
rect 151267 1831 151275 1865
rect 151225 1807 151275 1831
rect 151561 1865 151611 1889
rect 151561 1831 151569 1865
rect 151603 1831 151611 1865
rect 151561 1807 151611 1831
rect 151897 1865 151947 1889
rect 151897 1831 151905 1865
rect 151939 1831 151947 1865
rect 151897 1807 151947 1831
rect 152233 1865 152283 1889
rect 152233 1831 152241 1865
rect 152275 1831 152283 1865
rect 152233 1807 152283 1831
rect 152569 1865 152619 1889
rect 152569 1831 152577 1865
rect 152611 1831 152619 1865
rect 152569 1807 152619 1831
rect 152905 1865 152955 1889
rect 152905 1831 152913 1865
rect 152947 1831 152955 1865
rect 152905 1807 152955 1831
rect 153241 1865 153291 1889
rect 153241 1831 153249 1865
rect 153283 1831 153291 1865
rect 153241 1807 153291 1831
rect 153577 1865 153627 1889
rect 153577 1831 153585 1865
rect 153619 1831 153627 1865
rect 153577 1807 153627 1831
rect 153913 1865 153963 1889
rect 153913 1831 153921 1865
rect 153955 1831 153963 1865
rect 153913 1807 153963 1831
rect 154249 1865 154299 1889
rect 154249 1831 154257 1865
rect 154291 1831 154299 1865
rect 154249 1807 154299 1831
rect 154585 1865 154635 1889
rect 154585 1831 154593 1865
rect 154627 1831 154635 1865
rect 154585 1807 154635 1831
rect 154921 1865 154971 1889
rect 154921 1831 154929 1865
rect 154963 1831 154971 1865
rect 154921 1807 154971 1831
rect 155257 1865 155307 1889
rect 155257 1831 155265 1865
rect 155299 1831 155307 1865
rect 155257 1807 155307 1831
rect 155593 1865 155643 1889
rect 155593 1831 155601 1865
rect 155635 1831 155643 1865
rect 155593 1807 155643 1831
rect 155929 1865 155979 1889
rect 155929 1831 155937 1865
rect 155971 1831 155979 1865
rect 155929 1807 155979 1831
rect 156265 1865 156315 1889
rect 156265 1831 156273 1865
rect 156307 1831 156315 1865
rect 156265 1807 156315 1831
rect 156601 1865 156651 1889
rect 156601 1831 156609 1865
rect 156643 1831 156651 1865
rect 156601 1807 156651 1831
rect 156937 1865 156987 1889
rect 156937 1831 156945 1865
rect 156979 1831 156987 1865
rect 156937 1807 156987 1831
rect 157273 1865 157323 1889
rect 157273 1831 157281 1865
rect 157315 1831 157323 1865
rect 157273 1807 157323 1831
rect 157609 1865 157659 1889
rect 157609 1831 157617 1865
rect 157651 1831 157659 1865
rect 157609 1807 157659 1831
rect 157945 1865 157995 1889
rect 157945 1831 157953 1865
rect 157987 1831 157995 1865
rect 157945 1807 157995 1831
rect 158281 1865 158331 1889
rect 158281 1831 158289 1865
rect 158323 1831 158331 1865
rect 158281 1807 158331 1831
rect 158617 1865 158667 1889
rect 158617 1831 158625 1865
rect 158659 1831 158667 1865
rect 158617 1807 158667 1831
rect 158953 1865 159003 1889
rect 158953 1831 158961 1865
rect 158995 1831 159003 1865
rect 158953 1807 159003 1831
rect 159289 1865 159339 1889
rect 159289 1831 159297 1865
rect 159331 1831 159339 1865
rect 159289 1807 159339 1831
rect 159625 1865 159675 1889
rect 159625 1831 159633 1865
rect 159667 1831 159675 1865
rect 159625 1807 159675 1831
rect 159961 1865 160011 1889
rect 159961 1831 159969 1865
rect 160003 1831 160011 1865
rect 159961 1807 160011 1831
rect 160297 1865 160347 1889
rect 160297 1831 160305 1865
rect 160339 1831 160347 1865
rect 160297 1807 160347 1831
rect 160633 1865 160683 1889
rect 160633 1831 160641 1865
rect 160675 1831 160683 1865
rect 160633 1807 160683 1831
rect 160969 1865 161019 1889
rect 160969 1831 160977 1865
rect 161011 1831 161019 1865
rect 160969 1807 161019 1831
rect 161305 1865 161355 1889
rect 161305 1831 161313 1865
rect 161347 1831 161355 1865
rect 161305 1807 161355 1831
rect 161641 1865 161691 1889
rect 161641 1831 161649 1865
rect 161683 1831 161691 1865
rect 161641 1807 161691 1831
rect 161977 1865 162027 1889
rect 161977 1831 161985 1865
rect 162019 1831 162027 1865
rect 161977 1807 162027 1831
rect 162313 1865 162363 1889
rect 162313 1831 162321 1865
rect 162355 1831 162363 1865
rect 162313 1807 162363 1831
rect 162649 1865 162699 1889
rect 162649 1831 162657 1865
rect 162691 1831 162699 1865
rect 162649 1807 162699 1831
rect 162985 1865 163035 1889
rect 162985 1831 162993 1865
rect 163027 1831 163035 1865
rect 162985 1807 163035 1831
rect 163321 1865 163371 1889
rect 163321 1831 163329 1865
rect 163363 1831 163371 1865
rect 163321 1807 163371 1831
rect 163657 1865 163707 1889
rect 163657 1831 163665 1865
rect 163699 1831 163707 1865
rect 163657 1807 163707 1831
rect 163993 1865 164043 1889
rect 163993 1831 164001 1865
rect 164035 1831 164043 1865
rect 163993 1807 164043 1831
rect 164329 1865 164379 1889
rect 164329 1831 164337 1865
rect 164371 1831 164379 1865
rect 164329 1807 164379 1831
rect 164665 1865 164715 1889
rect 164665 1831 164673 1865
rect 164707 1831 164715 1865
rect 164665 1807 164715 1831
rect 165001 1865 165051 1889
rect 165001 1831 165009 1865
rect 165043 1831 165051 1865
rect 165001 1807 165051 1831
rect 165337 1865 165387 1889
rect 165337 1831 165345 1865
rect 165379 1831 165387 1865
rect 165337 1807 165387 1831
rect 165673 1865 165723 1889
rect 165673 1831 165681 1865
rect 165715 1831 165723 1865
rect 165673 1807 165723 1831
rect 166009 1865 166059 1889
rect 166009 1831 166017 1865
rect 166051 1831 166059 1865
rect 166009 1807 166059 1831
rect 166345 1865 166395 1889
rect 166345 1831 166353 1865
rect 166387 1831 166395 1865
rect 166345 1807 166395 1831
rect 166681 1865 166731 1889
rect 166681 1831 166689 1865
rect 166723 1831 166731 1865
rect 166681 1807 166731 1831
rect 167017 1865 167067 1889
rect 167017 1831 167025 1865
rect 167059 1831 167067 1865
rect 167017 1807 167067 1831
rect 167353 1865 167403 1889
rect 167353 1831 167361 1865
rect 167395 1831 167403 1865
rect 167353 1807 167403 1831
rect 167689 1865 167739 1889
rect 167689 1831 167697 1865
rect 167731 1831 167739 1865
rect 167689 1807 167739 1831
rect 168025 1865 168075 1889
rect 168025 1831 168033 1865
rect 168067 1831 168075 1865
rect 168025 1807 168075 1831
rect 168361 1865 168411 1889
rect 168361 1831 168369 1865
rect 168403 1831 168411 1865
rect 168361 1807 168411 1831
rect 168697 1865 168747 1889
rect 168697 1831 168705 1865
rect 168739 1831 168747 1865
rect 168697 1807 168747 1831
rect 169033 1865 169083 1889
rect 169033 1831 169041 1865
rect 169075 1831 169083 1865
rect 169033 1807 169083 1831
rect 169369 1865 169419 1889
rect 169369 1831 169377 1865
rect 169411 1831 169419 1865
rect 169369 1807 169419 1831
rect 169705 1865 169755 1889
rect 169705 1831 169713 1865
rect 169747 1831 169755 1865
rect 169705 1807 169755 1831
rect 170041 1865 170091 1889
rect 170041 1831 170049 1865
rect 170083 1831 170091 1865
rect 170041 1807 170091 1831
rect 170377 1865 170427 1889
rect 170377 1831 170385 1865
rect 170419 1831 170427 1865
rect 170377 1807 170427 1831
rect 170713 1865 170763 1889
rect 170713 1831 170721 1865
rect 170755 1831 170763 1865
rect 170713 1807 170763 1831
rect 171049 1865 171099 1889
rect 171049 1831 171057 1865
rect 171091 1831 171099 1865
rect 171049 1807 171099 1831
rect 171385 1865 171435 1889
rect 171385 1831 171393 1865
rect 171427 1831 171435 1865
rect 171385 1807 171435 1831
rect 171721 1865 171771 1889
rect 171721 1831 171729 1865
rect 171763 1831 171771 1865
rect 171721 1807 171771 1831
rect 172057 1865 172107 1889
rect 172057 1831 172065 1865
rect 172099 1831 172107 1865
rect 172057 1807 172107 1831
rect 172393 1865 172443 1889
rect 172393 1831 172401 1865
rect 172435 1831 172443 1865
rect 172393 1807 172443 1831
rect 172729 1865 172779 1889
rect 172729 1831 172737 1865
rect 172771 1831 172779 1865
rect 172729 1807 172779 1831
rect 173065 1865 173115 1889
rect 173065 1831 173073 1865
rect 173107 1831 173115 1865
rect 173065 1807 173115 1831
rect 173401 1865 173451 1889
rect 173401 1831 173409 1865
rect 173443 1831 173451 1865
rect 173401 1807 173451 1831
rect 173737 1865 173787 1889
rect 173737 1831 173745 1865
rect 173779 1831 173787 1865
rect 173737 1807 173787 1831
rect 174073 1865 174123 1889
rect 174073 1831 174081 1865
rect 174115 1831 174123 1865
rect 174073 1807 174123 1831
rect 174409 1865 174459 1889
rect 174409 1831 174417 1865
rect 174451 1831 174459 1865
rect 174409 1807 174459 1831
rect 174745 1865 174795 1889
rect 174745 1831 174753 1865
rect 174787 1831 174795 1865
rect 174745 1807 174795 1831
rect 175081 1865 175131 1889
rect 175081 1831 175089 1865
rect 175123 1831 175131 1865
rect 175081 1807 175131 1831
rect 175417 1865 175467 1889
rect 175417 1831 175425 1865
rect 175459 1831 175467 1865
rect 175417 1807 175467 1831
rect 175753 1865 175803 1889
rect 175753 1831 175761 1865
rect 175795 1831 175803 1865
rect 175753 1807 175803 1831
rect 176089 1865 176139 1889
rect 176089 1831 176097 1865
rect 176131 1831 176139 1865
rect 176089 1807 176139 1831
rect 176425 1865 176475 1889
rect 176425 1831 176433 1865
rect 176467 1831 176475 1865
rect 176425 1807 176475 1831
rect 176761 1865 176811 1889
rect 176761 1831 176769 1865
rect 176803 1831 176811 1865
rect 176761 1807 176811 1831
rect 177097 1865 177147 1889
rect 177097 1831 177105 1865
rect 177139 1831 177147 1865
rect 177097 1807 177147 1831
rect 177433 1865 177483 1889
rect 177433 1831 177441 1865
rect 177475 1831 177483 1865
rect 177433 1807 177483 1831
rect 177769 1865 177819 1889
rect 177769 1831 177777 1865
rect 177811 1831 177819 1865
rect 177769 1807 177819 1831
rect 178105 1865 178155 1889
rect 178105 1831 178113 1865
rect 178147 1831 178155 1865
rect 178105 1807 178155 1831
rect 178441 1865 178491 1889
rect 178441 1831 178449 1865
rect 178483 1831 178491 1865
rect 178441 1807 178491 1831
rect 178777 1865 178827 1889
rect 178777 1831 178785 1865
rect 178819 1831 178827 1865
rect 178777 1807 178827 1831
rect 179113 1865 179163 1889
rect 179113 1831 179121 1865
rect 179155 1831 179163 1865
rect 179113 1807 179163 1831
rect 179449 1865 179499 1889
rect 179449 1831 179457 1865
rect 179491 1831 179499 1865
rect 179449 1807 179499 1831
rect 179785 1865 179835 1889
rect 179785 1831 179793 1865
rect 179827 1831 179835 1865
rect 179785 1807 179835 1831
rect 180121 1865 180171 1889
rect 180121 1831 180129 1865
rect 180163 1831 180171 1865
rect 180121 1807 180171 1831
rect 180457 1865 180507 1889
rect 180457 1831 180465 1865
rect 180499 1831 180507 1865
rect 180457 1807 180507 1831
rect 180793 1865 180843 1889
rect 180793 1831 180801 1865
rect 180835 1831 180843 1865
rect 180793 1807 180843 1831
rect 181129 1865 181179 1889
rect 181129 1831 181137 1865
rect 181171 1831 181179 1865
rect 181129 1807 181179 1831
rect 181465 1865 181515 1889
rect 181465 1831 181473 1865
rect 181507 1831 181515 1865
rect 181465 1807 181515 1831
rect 181801 1865 181851 1889
rect 181801 1831 181809 1865
rect 181843 1831 181851 1865
rect 181801 1807 181851 1831
rect 182137 1865 182187 1889
rect 182137 1831 182145 1865
rect 182179 1831 182187 1865
rect 182137 1807 182187 1831
rect 182473 1865 182523 1889
rect 182473 1831 182481 1865
rect 182515 1831 182523 1865
rect 182473 1807 182523 1831
rect 182809 1865 182859 1889
rect 182809 1831 182817 1865
rect 182851 1831 182859 1865
rect 182809 1807 182859 1831
rect 183145 1865 183195 1889
rect 183145 1831 183153 1865
rect 183187 1831 183195 1865
rect 183145 1807 183195 1831
rect 183481 1865 183531 1889
rect 183481 1831 183489 1865
rect 183523 1831 183531 1865
rect 183481 1807 183531 1831
rect 183817 1865 183867 1889
rect 183817 1831 183825 1865
rect 183859 1831 183867 1865
rect 183817 1807 183867 1831
rect 184153 1865 184203 1889
rect 184153 1831 184161 1865
rect 184195 1831 184203 1865
rect 184153 1807 184203 1831
rect 184489 1865 184539 1889
rect 184489 1831 184497 1865
rect 184531 1831 184539 1865
rect 184489 1807 184539 1831
rect 184825 1865 184875 1889
rect 184825 1831 184833 1865
rect 184867 1831 184875 1865
rect 184825 1807 184875 1831
rect 185161 1865 185211 1889
rect 185161 1831 185169 1865
rect 185203 1831 185211 1865
rect 185161 1807 185211 1831
rect 185497 1865 185547 1889
rect 185497 1831 185505 1865
rect 185539 1831 185547 1865
rect 185497 1807 185547 1831
rect 185833 1865 185883 1889
rect 185833 1831 185841 1865
rect 185875 1831 185883 1865
rect 185833 1807 185883 1831
rect 186169 1865 186219 1889
rect 186169 1831 186177 1865
rect 186211 1831 186219 1865
rect 186169 1807 186219 1831
rect 186505 1865 186555 1889
rect 186505 1831 186513 1865
rect 186547 1831 186555 1865
rect 186505 1807 186555 1831
rect 186841 1865 186891 1889
rect 186841 1831 186849 1865
rect 186883 1831 186891 1865
rect 186841 1807 186891 1831
rect 187177 1865 187227 1889
rect 187177 1831 187185 1865
rect 187219 1831 187227 1865
rect 187177 1807 187227 1831
rect 187513 1865 187563 1889
rect 187513 1831 187521 1865
rect 187555 1831 187563 1865
rect 187513 1807 187563 1831
rect 187849 1865 187899 1889
rect 187849 1831 187857 1865
rect 187891 1831 187899 1865
rect 187849 1807 187899 1831
rect 188185 1865 188235 1889
rect 188185 1831 188193 1865
rect 188227 1831 188235 1865
rect 188185 1807 188235 1831
rect 188521 1865 188571 1889
rect 188521 1831 188529 1865
rect 188563 1831 188571 1865
rect 188521 1807 188571 1831
rect 188857 1865 188907 1889
rect 188857 1831 188865 1865
rect 188899 1831 188907 1865
rect 188857 1807 188907 1831
rect 189193 1865 189243 1889
rect 189193 1831 189201 1865
rect 189235 1831 189243 1865
rect 189193 1807 189243 1831
rect 189529 1865 189579 1889
rect 189529 1831 189537 1865
rect 189571 1831 189579 1865
rect 189529 1807 189579 1831
rect 189865 1865 189915 1889
rect 189865 1831 189873 1865
rect 189907 1831 189915 1865
rect 189865 1807 189915 1831
rect 190201 1865 190251 1889
rect 190201 1831 190209 1865
rect 190243 1831 190251 1865
rect 190201 1807 190251 1831
rect 190537 1865 190587 1889
rect 190537 1831 190545 1865
rect 190579 1831 190587 1865
rect 190537 1807 190587 1831
rect 190873 1865 190923 1889
rect 190873 1831 190881 1865
rect 190915 1831 190923 1865
rect 190873 1807 190923 1831
rect 191209 1865 191259 1889
rect 191209 1831 191217 1865
rect 191251 1831 191259 1865
rect 191209 1807 191259 1831
rect 191545 1865 191595 1889
rect 191545 1831 191553 1865
rect 191587 1831 191595 1865
rect 191545 1807 191595 1831
rect 191881 1865 191931 1889
rect 191881 1831 191889 1865
rect 191923 1831 191931 1865
rect 191881 1807 191931 1831
rect 192217 1865 192267 1889
rect 192217 1831 192225 1865
rect 192259 1831 192267 1865
rect 192217 1807 192267 1831
rect 192553 1865 192603 1889
rect 192553 1831 192561 1865
rect 192595 1831 192603 1865
rect 192553 1807 192603 1831
rect 192889 1865 192939 1889
rect 192889 1831 192897 1865
rect 192931 1831 192939 1865
rect 192889 1807 192939 1831
rect 193225 1865 193275 1889
rect 193225 1831 193233 1865
rect 193267 1831 193275 1865
rect 193225 1807 193275 1831
rect 193561 1865 193611 1889
rect 193561 1831 193569 1865
rect 193603 1831 193611 1865
rect 193561 1807 193611 1831
rect 193897 1865 193947 1889
rect 193897 1831 193905 1865
rect 193939 1831 193947 1865
rect 193897 1807 193947 1831
rect 194233 1865 194283 1889
rect 194233 1831 194241 1865
rect 194275 1831 194283 1865
rect 194233 1807 194283 1831
rect 194569 1865 194619 1889
rect 194569 1831 194577 1865
rect 194611 1831 194619 1865
rect 194569 1807 194619 1831
rect 194905 1865 194955 1889
rect 194905 1831 194913 1865
rect 194947 1831 194955 1865
rect 194905 1807 194955 1831
rect 195241 1865 195291 1889
rect 195241 1831 195249 1865
rect 195283 1831 195291 1865
rect 195241 1807 195291 1831
rect 195577 1865 195627 1889
rect 195577 1831 195585 1865
rect 195619 1831 195627 1865
rect 195577 1807 195627 1831
rect 195913 1865 195963 1889
rect 195913 1831 195921 1865
rect 195955 1831 195963 1865
rect 195913 1807 195963 1831
rect 196249 1865 196299 1889
rect 196249 1831 196257 1865
rect 196291 1831 196299 1865
rect 196249 1807 196299 1831
rect 196585 1865 196635 1889
rect 196585 1831 196593 1865
rect 196627 1831 196635 1865
rect 196585 1807 196635 1831
rect 196921 1865 196971 1889
rect 196921 1831 196929 1865
rect 196963 1831 196971 1865
rect 196921 1807 196971 1831
rect 197257 1865 197307 1889
rect 197257 1831 197265 1865
rect 197299 1831 197307 1865
rect 197257 1807 197307 1831
rect 197593 1865 197643 1889
rect 197593 1831 197601 1865
rect 197635 1831 197643 1865
rect 197593 1807 197643 1831
rect 197929 1865 197979 1889
rect 197929 1831 197937 1865
rect 197971 1831 197979 1865
rect 197929 1807 197979 1831
rect 198265 1865 198315 1889
rect 198265 1831 198273 1865
rect 198307 1831 198315 1865
rect 198265 1807 198315 1831
rect 198601 1865 198651 1889
rect 198601 1831 198609 1865
rect 198643 1831 198651 1865
rect 198601 1807 198651 1831
rect 198937 1865 198987 1889
rect 198937 1831 198945 1865
rect 198979 1831 198987 1865
rect 198937 1807 198987 1831
rect 199273 1865 199323 1889
rect 199273 1831 199281 1865
rect 199315 1831 199323 1865
rect 199273 1807 199323 1831
rect 199609 1865 199659 1889
rect 199609 1831 199617 1865
rect 199651 1831 199659 1865
rect 199609 1807 199659 1831
rect 199945 1865 199995 1889
rect 199945 1831 199953 1865
rect 199987 1831 199995 1865
rect 199945 1807 199995 1831
rect 200281 1865 200331 1889
rect 200281 1831 200289 1865
rect 200323 1831 200331 1865
rect 200281 1807 200331 1831
rect 200617 1865 200667 1889
rect 200617 1831 200625 1865
rect 200659 1831 200667 1865
rect 200617 1807 200667 1831
rect 200953 1865 201003 1889
rect 200953 1831 200961 1865
rect 200995 1831 201003 1865
rect 200953 1807 201003 1831
rect 201289 1865 201339 1889
rect 201289 1831 201297 1865
rect 201331 1831 201339 1865
rect 201289 1807 201339 1831
rect 201625 1865 201675 1889
rect 201625 1831 201633 1865
rect 201667 1831 201675 1865
rect 201625 1807 201675 1831
rect 201961 1865 202011 1889
rect 201961 1831 201969 1865
rect 202003 1831 202011 1865
rect 201961 1807 202011 1831
rect 202297 1865 202347 1889
rect 202297 1831 202305 1865
rect 202339 1831 202347 1865
rect 202297 1807 202347 1831
rect 202633 1865 202683 1889
rect 202633 1831 202641 1865
rect 202675 1831 202683 1865
rect 202633 1807 202683 1831
rect 202969 1865 203019 1889
rect 202969 1831 202977 1865
rect 203011 1831 203019 1865
rect 202969 1807 203019 1831
rect 203305 1865 203355 1889
rect 203305 1831 203313 1865
rect 203347 1831 203355 1865
rect 203305 1807 203355 1831
rect 203641 1865 203691 1889
rect 203641 1831 203649 1865
rect 203683 1831 203691 1865
rect 203641 1807 203691 1831
rect 203977 1865 204027 1889
rect 203977 1831 203985 1865
rect 204019 1831 204027 1865
rect 203977 1807 204027 1831
rect 204313 1865 204363 1889
rect 204313 1831 204321 1865
rect 204355 1831 204363 1865
rect 204313 1807 204363 1831
rect 204649 1865 204699 1889
rect 204649 1831 204657 1865
rect 204691 1831 204699 1865
rect 204649 1807 204699 1831
rect 204985 1865 205035 1889
rect 204985 1831 204993 1865
rect 205027 1831 205035 1865
rect 204985 1807 205035 1831
rect 205321 1865 205371 1889
rect 205321 1831 205329 1865
rect 205363 1831 205371 1865
rect 205321 1807 205371 1831
rect 205657 1865 205707 1889
rect 205657 1831 205665 1865
rect 205699 1831 205707 1865
rect 205657 1807 205707 1831
rect 205993 1865 206043 1889
rect 205993 1831 206001 1865
rect 206035 1831 206043 1865
rect 205993 1807 206043 1831
rect 206329 1865 206379 1889
rect 206329 1831 206337 1865
rect 206371 1831 206379 1865
rect 206329 1807 206379 1831
rect 206665 1865 206715 1889
rect 206665 1831 206673 1865
rect 206707 1831 206715 1865
rect 206665 1807 206715 1831
rect 207001 1865 207051 1889
rect 207001 1831 207009 1865
rect 207043 1831 207051 1865
rect 207001 1807 207051 1831
rect 207337 1865 207387 1889
rect 207337 1831 207345 1865
rect 207379 1831 207387 1865
rect 207337 1807 207387 1831
rect 207673 1865 207723 1889
rect 207673 1831 207681 1865
rect 207715 1831 207723 1865
rect 207673 1807 207723 1831
rect 208009 1865 208059 1889
rect 208009 1831 208017 1865
rect 208051 1831 208059 1865
rect 208009 1807 208059 1831
rect 208345 1865 208395 1889
rect 208345 1831 208353 1865
rect 208387 1831 208395 1865
rect 208345 1807 208395 1831
rect 208681 1865 208731 1889
rect 208681 1831 208689 1865
rect 208723 1831 208731 1865
rect 208681 1807 208731 1831
rect 209017 1865 209067 1889
rect 209017 1831 209025 1865
rect 209059 1831 209067 1865
rect 209017 1807 209067 1831
rect 209353 1865 209403 1889
rect 209353 1831 209361 1865
rect 209395 1831 209403 1865
rect 209353 1807 209403 1831
rect 209689 1865 209739 1889
rect 209689 1831 209697 1865
rect 209731 1831 209739 1865
rect 209689 1807 209739 1831
rect 210025 1865 210075 1889
rect 210025 1831 210033 1865
rect 210067 1831 210075 1865
rect 210025 1807 210075 1831
rect 210361 1865 210411 1889
rect 210361 1831 210369 1865
rect 210403 1831 210411 1865
rect 210361 1807 210411 1831
rect 210697 1865 210747 1889
rect 210697 1831 210705 1865
rect 210739 1831 210747 1865
rect 210697 1807 210747 1831
rect 211033 1865 211083 1889
rect 211033 1831 211041 1865
rect 211075 1831 211083 1865
rect 211033 1807 211083 1831
rect 211369 1865 211419 1889
rect 211369 1831 211377 1865
rect 211411 1831 211419 1865
rect 211369 1807 211419 1831
rect 211705 1865 211755 1889
rect 211705 1831 211713 1865
rect 211747 1831 211755 1865
rect 211705 1807 211755 1831
rect 212041 1865 212091 1889
rect 212041 1831 212049 1865
rect 212083 1831 212091 1865
rect 212041 1807 212091 1831
rect 212377 1865 212427 1889
rect 212377 1831 212385 1865
rect 212419 1831 212427 1865
rect 212377 1807 212427 1831
rect 212713 1865 212763 1889
rect 212713 1831 212721 1865
rect 212755 1831 212763 1865
rect 212713 1807 212763 1831
rect 213049 1865 213099 1889
rect 213049 1831 213057 1865
rect 213091 1831 213099 1865
rect 213049 1807 213099 1831
rect 213385 1865 213435 1889
rect 213385 1831 213393 1865
rect 213427 1831 213435 1865
rect 213385 1807 213435 1831
rect 213721 1865 213771 1889
rect 213721 1831 213729 1865
rect 213763 1831 213771 1865
rect 213721 1807 213771 1831
rect 214057 1865 214107 1889
rect 214057 1831 214065 1865
rect 214099 1831 214107 1865
rect 214057 1807 214107 1831
rect 214393 1865 214443 1889
rect 214393 1831 214401 1865
rect 214435 1831 214443 1865
rect 214393 1807 214443 1831
rect 214729 1865 214779 1889
rect 214729 1831 214737 1865
rect 214771 1831 214779 1865
rect 214729 1807 214779 1831
rect 215065 1865 215115 1889
rect 215065 1831 215073 1865
rect 215107 1831 215115 1865
rect 215065 1807 215115 1831
rect 215401 1865 215451 1889
rect 215401 1831 215409 1865
rect 215443 1831 215451 1865
rect 215401 1807 215451 1831
rect 215737 1865 215787 1889
rect 215737 1831 215745 1865
rect 215779 1831 215787 1865
rect 215737 1807 215787 1831
rect 216073 1865 216123 1889
rect 216073 1831 216081 1865
rect 216115 1831 216123 1865
rect 216073 1807 216123 1831
rect 216409 1865 216459 1889
rect 216409 1831 216417 1865
rect 216451 1831 216459 1865
rect 216409 1807 216459 1831
<< nsubdiffcont >>
rect 2049 142327 2083 142361
rect 2385 142327 2419 142361
rect 2721 142327 2755 142361
rect 3057 142327 3091 142361
rect 3393 142327 3427 142361
rect 3729 142327 3763 142361
rect 4065 142327 4099 142361
rect 4401 142327 4435 142361
rect 4737 142327 4771 142361
rect 5073 142327 5107 142361
rect 5409 142327 5443 142361
rect 5745 142327 5779 142361
rect 6081 142327 6115 142361
rect 6417 142327 6451 142361
rect 6753 142327 6787 142361
rect 7089 142327 7123 142361
rect 7425 142327 7459 142361
rect 7761 142327 7795 142361
rect 8097 142327 8131 142361
rect 8433 142327 8467 142361
rect 8769 142327 8803 142361
rect 9105 142327 9139 142361
rect 9441 142327 9475 142361
rect 9777 142327 9811 142361
rect 10113 142327 10147 142361
rect 10449 142327 10483 142361
rect 10785 142327 10819 142361
rect 11121 142327 11155 142361
rect 11457 142327 11491 142361
rect 11793 142327 11827 142361
rect 12129 142327 12163 142361
rect 12465 142327 12499 142361
rect 12801 142327 12835 142361
rect 13137 142327 13171 142361
rect 13473 142327 13507 142361
rect 13809 142327 13843 142361
rect 14145 142327 14179 142361
rect 14481 142327 14515 142361
rect 14817 142327 14851 142361
rect 15153 142327 15187 142361
rect 15489 142327 15523 142361
rect 15825 142327 15859 142361
rect 16161 142327 16195 142361
rect 16497 142327 16531 142361
rect 16833 142327 16867 142361
rect 17169 142327 17203 142361
rect 17505 142327 17539 142361
rect 17841 142327 17875 142361
rect 18177 142327 18211 142361
rect 18513 142327 18547 142361
rect 18849 142327 18883 142361
rect 19185 142327 19219 142361
rect 19521 142327 19555 142361
rect 19857 142327 19891 142361
rect 20193 142327 20227 142361
rect 20529 142327 20563 142361
rect 20865 142327 20899 142361
rect 21201 142327 21235 142361
rect 21537 142327 21571 142361
rect 21873 142327 21907 142361
rect 22209 142327 22243 142361
rect 22545 142327 22579 142361
rect 22881 142327 22915 142361
rect 23217 142327 23251 142361
rect 23553 142327 23587 142361
rect 23889 142327 23923 142361
rect 24225 142327 24259 142361
rect 24561 142327 24595 142361
rect 24897 142327 24931 142361
rect 25233 142327 25267 142361
rect 25569 142327 25603 142361
rect 25905 142327 25939 142361
rect 26241 142327 26275 142361
rect 26577 142327 26611 142361
rect 26913 142327 26947 142361
rect 27249 142327 27283 142361
rect 27585 142327 27619 142361
rect 27921 142327 27955 142361
rect 28257 142327 28291 142361
rect 28593 142327 28627 142361
rect 28929 142327 28963 142361
rect 29265 142327 29299 142361
rect 29601 142327 29635 142361
rect 29937 142327 29971 142361
rect 30273 142327 30307 142361
rect 30609 142327 30643 142361
rect 30945 142327 30979 142361
rect 31281 142327 31315 142361
rect 31617 142327 31651 142361
rect 31953 142327 31987 142361
rect 32289 142327 32323 142361
rect 32625 142327 32659 142361
rect 32961 142327 32995 142361
rect 33297 142327 33331 142361
rect 33633 142327 33667 142361
rect 33969 142327 34003 142361
rect 34305 142327 34339 142361
rect 34641 142327 34675 142361
rect 34977 142327 35011 142361
rect 35313 142327 35347 142361
rect 35649 142327 35683 142361
rect 35985 142327 36019 142361
rect 36321 142327 36355 142361
rect 36657 142327 36691 142361
rect 36993 142327 37027 142361
rect 37329 142327 37363 142361
rect 37665 142327 37699 142361
rect 38001 142327 38035 142361
rect 38337 142327 38371 142361
rect 38673 142327 38707 142361
rect 39009 142327 39043 142361
rect 39345 142327 39379 142361
rect 39681 142327 39715 142361
rect 40017 142327 40051 142361
rect 40353 142327 40387 142361
rect 40689 142327 40723 142361
rect 41025 142327 41059 142361
rect 41361 142327 41395 142361
rect 41697 142327 41731 142361
rect 42033 142327 42067 142361
rect 42369 142327 42403 142361
rect 42705 142327 42739 142361
rect 43041 142327 43075 142361
rect 43377 142327 43411 142361
rect 43713 142327 43747 142361
rect 44049 142327 44083 142361
rect 44385 142327 44419 142361
rect 44721 142327 44755 142361
rect 45057 142327 45091 142361
rect 45393 142327 45427 142361
rect 45729 142327 45763 142361
rect 46065 142327 46099 142361
rect 46401 142327 46435 142361
rect 46737 142327 46771 142361
rect 47073 142327 47107 142361
rect 47409 142327 47443 142361
rect 47745 142327 47779 142361
rect 48081 142327 48115 142361
rect 48417 142327 48451 142361
rect 48753 142327 48787 142361
rect 49089 142327 49123 142361
rect 49425 142327 49459 142361
rect 49761 142327 49795 142361
rect 50097 142327 50131 142361
rect 50433 142327 50467 142361
rect 50769 142327 50803 142361
rect 51105 142327 51139 142361
rect 51441 142327 51475 142361
rect 51777 142327 51811 142361
rect 52113 142327 52147 142361
rect 52449 142327 52483 142361
rect 52785 142327 52819 142361
rect 53121 142327 53155 142361
rect 53457 142327 53491 142361
rect 53793 142327 53827 142361
rect 54129 142327 54163 142361
rect 54465 142327 54499 142361
rect 54801 142327 54835 142361
rect 55137 142327 55171 142361
rect 55473 142327 55507 142361
rect 55809 142327 55843 142361
rect 56145 142327 56179 142361
rect 56481 142327 56515 142361
rect 56817 142327 56851 142361
rect 57153 142327 57187 142361
rect 57489 142327 57523 142361
rect 57825 142327 57859 142361
rect 58161 142327 58195 142361
rect 58497 142327 58531 142361
rect 58833 142327 58867 142361
rect 59169 142327 59203 142361
rect 59505 142327 59539 142361
rect 59841 142327 59875 142361
rect 60177 142327 60211 142361
rect 60513 142327 60547 142361
rect 60849 142327 60883 142361
rect 61185 142327 61219 142361
rect 61521 142327 61555 142361
rect 61857 142327 61891 142361
rect 62193 142327 62227 142361
rect 62529 142327 62563 142361
rect 62865 142327 62899 142361
rect 63201 142327 63235 142361
rect 63537 142327 63571 142361
rect 63873 142327 63907 142361
rect 64209 142327 64243 142361
rect 64545 142327 64579 142361
rect 64881 142327 64915 142361
rect 65217 142327 65251 142361
rect 65553 142327 65587 142361
rect 65889 142327 65923 142361
rect 66225 142327 66259 142361
rect 66561 142327 66595 142361
rect 66897 142327 66931 142361
rect 67233 142327 67267 142361
rect 67569 142327 67603 142361
rect 67905 142327 67939 142361
rect 68241 142327 68275 142361
rect 68577 142327 68611 142361
rect 68913 142327 68947 142361
rect 69249 142327 69283 142361
rect 69585 142327 69619 142361
rect 69921 142327 69955 142361
rect 70257 142327 70291 142361
rect 70593 142327 70627 142361
rect 70929 142327 70963 142361
rect 71265 142327 71299 142361
rect 71601 142327 71635 142361
rect 71937 142327 71971 142361
rect 72273 142327 72307 142361
rect 72609 142327 72643 142361
rect 72945 142327 72979 142361
rect 73281 142327 73315 142361
rect 73617 142327 73651 142361
rect 73953 142327 73987 142361
rect 74289 142327 74323 142361
rect 74625 142327 74659 142361
rect 74961 142327 74995 142361
rect 75297 142327 75331 142361
rect 75633 142327 75667 142361
rect 75969 142327 76003 142361
rect 76305 142327 76339 142361
rect 76641 142327 76675 142361
rect 76977 142327 77011 142361
rect 77313 142327 77347 142361
rect 77649 142327 77683 142361
rect 77985 142327 78019 142361
rect 78321 142327 78355 142361
rect 78657 142327 78691 142361
rect 78993 142327 79027 142361
rect 79329 142327 79363 142361
rect 79665 142327 79699 142361
rect 80001 142327 80035 142361
rect 80337 142327 80371 142361
rect 80673 142327 80707 142361
rect 81009 142327 81043 142361
rect 81345 142327 81379 142361
rect 81681 142327 81715 142361
rect 82017 142327 82051 142361
rect 82353 142327 82387 142361
rect 82689 142327 82723 142361
rect 83025 142327 83059 142361
rect 83361 142327 83395 142361
rect 83697 142327 83731 142361
rect 84033 142327 84067 142361
rect 84369 142327 84403 142361
rect 84705 142327 84739 142361
rect 85041 142327 85075 142361
rect 85377 142327 85411 142361
rect 85713 142327 85747 142361
rect 86049 142327 86083 142361
rect 86385 142327 86419 142361
rect 86721 142327 86755 142361
rect 87057 142327 87091 142361
rect 87393 142327 87427 142361
rect 87729 142327 87763 142361
rect 88065 142327 88099 142361
rect 88401 142327 88435 142361
rect 88737 142327 88771 142361
rect 89073 142327 89107 142361
rect 89409 142327 89443 142361
rect 89745 142327 89779 142361
rect 90081 142327 90115 142361
rect 90417 142327 90451 142361
rect 90753 142327 90787 142361
rect 91089 142327 91123 142361
rect 91425 142327 91459 142361
rect 91761 142327 91795 142361
rect 92097 142327 92131 142361
rect 92433 142327 92467 142361
rect 92769 142327 92803 142361
rect 93105 142327 93139 142361
rect 93441 142327 93475 142361
rect 93777 142327 93811 142361
rect 94113 142327 94147 142361
rect 94449 142327 94483 142361
rect 94785 142327 94819 142361
rect 95121 142327 95155 142361
rect 95457 142327 95491 142361
rect 95793 142327 95827 142361
rect 96129 142327 96163 142361
rect 96465 142327 96499 142361
rect 96801 142327 96835 142361
rect 97137 142327 97171 142361
rect 97473 142327 97507 142361
rect 97809 142327 97843 142361
rect 98145 142327 98179 142361
rect 98481 142327 98515 142361
rect 98817 142327 98851 142361
rect 99153 142327 99187 142361
rect 99489 142327 99523 142361
rect 99825 142327 99859 142361
rect 100161 142327 100195 142361
rect 100497 142327 100531 142361
rect 100833 142327 100867 142361
rect 101169 142327 101203 142361
rect 101505 142327 101539 142361
rect 101841 142327 101875 142361
rect 102177 142327 102211 142361
rect 102513 142327 102547 142361
rect 102849 142327 102883 142361
rect 103185 142327 103219 142361
rect 103521 142327 103555 142361
rect 103857 142327 103891 142361
rect 104193 142327 104227 142361
rect 104529 142327 104563 142361
rect 104865 142327 104899 142361
rect 105201 142327 105235 142361
rect 105537 142327 105571 142361
rect 105873 142327 105907 142361
rect 106209 142327 106243 142361
rect 106545 142327 106579 142361
rect 106881 142327 106915 142361
rect 107217 142327 107251 142361
rect 107553 142327 107587 142361
rect 107889 142327 107923 142361
rect 108225 142327 108259 142361
rect 108561 142327 108595 142361
rect 108897 142327 108931 142361
rect 109233 142327 109267 142361
rect 109569 142327 109603 142361
rect 109905 142327 109939 142361
rect 110241 142327 110275 142361
rect 110577 142327 110611 142361
rect 110913 142327 110947 142361
rect 111249 142327 111283 142361
rect 111585 142327 111619 142361
rect 111921 142327 111955 142361
rect 112257 142327 112291 142361
rect 112593 142327 112627 142361
rect 112929 142327 112963 142361
rect 113265 142327 113299 142361
rect 113601 142327 113635 142361
rect 113937 142327 113971 142361
rect 114273 142327 114307 142361
rect 114609 142327 114643 142361
rect 114945 142327 114979 142361
rect 115281 142327 115315 142361
rect 115617 142327 115651 142361
rect 115953 142327 115987 142361
rect 116289 142327 116323 142361
rect 116625 142327 116659 142361
rect 116961 142327 116995 142361
rect 117297 142327 117331 142361
rect 117633 142327 117667 142361
rect 117969 142327 118003 142361
rect 118305 142327 118339 142361
rect 118641 142327 118675 142361
rect 118977 142327 119011 142361
rect 119313 142327 119347 142361
rect 119649 142327 119683 142361
rect 119985 142327 120019 142361
rect 120321 142327 120355 142361
rect 120657 142327 120691 142361
rect 120993 142327 121027 142361
rect 121329 142327 121363 142361
rect 121665 142327 121699 142361
rect 122001 142327 122035 142361
rect 122337 142327 122371 142361
rect 122673 142327 122707 142361
rect 123009 142327 123043 142361
rect 123345 142327 123379 142361
rect 123681 142327 123715 142361
rect 124017 142327 124051 142361
rect 124353 142327 124387 142361
rect 124689 142327 124723 142361
rect 125025 142327 125059 142361
rect 125361 142327 125395 142361
rect 125697 142327 125731 142361
rect 126033 142327 126067 142361
rect 126369 142327 126403 142361
rect 126705 142327 126739 142361
rect 127041 142327 127075 142361
rect 127377 142327 127411 142361
rect 127713 142327 127747 142361
rect 128049 142327 128083 142361
rect 128385 142327 128419 142361
rect 128721 142327 128755 142361
rect 129057 142327 129091 142361
rect 129393 142327 129427 142361
rect 129729 142327 129763 142361
rect 130065 142327 130099 142361
rect 130401 142327 130435 142361
rect 130737 142327 130771 142361
rect 131073 142327 131107 142361
rect 131409 142327 131443 142361
rect 131745 142327 131779 142361
rect 132081 142327 132115 142361
rect 132417 142327 132451 142361
rect 132753 142327 132787 142361
rect 133089 142327 133123 142361
rect 133425 142327 133459 142361
rect 133761 142327 133795 142361
rect 134097 142327 134131 142361
rect 134433 142327 134467 142361
rect 134769 142327 134803 142361
rect 135105 142327 135139 142361
rect 135441 142327 135475 142361
rect 135777 142327 135811 142361
rect 136113 142327 136147 142361
rect 136449 142327 136483 142361
rect 136785 142327 136819 142361
rect 137121 142327 137155 142361
rect 137457 142327 137491 142361
rect 137793 142327 137827 142361
rect 138129 142327 138163 142361
rect 138465 142327 138499 142361
rect 138801 142327 138835 142361
rect 139137 142327 139171 142361
rect 139473 142327 139507 142361
rect 139809 142327 139843 142361
rect 140145 142327 140179 142361
rect 140481 142327 140515 142361
rect 140817 142327 140851 142361
rect 141153 142327 141187 142361
rect 141489 142327 141523 142361
rect 141825 142327 141859 142361
rect 142161 142327 142195 142361
rect 142497 142327 142531 142361
rect 142833 142327 142867 142361
rect 143169 142327 143203 142361
rect 143505 142327 143539 142361
rect 143841 142327 143875 142361
rect 144177 142327 144211 142361
rect 144513 142327 144547 142361
rect 144849 142327 144883 142361
rect 145185 142327 145219 142361
rect 145521 142327 145555 142361
rect 145857 142327 145891 142361
rect 146193 142327 146227 142361
rect 146529 142327 146563 142361
rect 146865 142327 146899 142361
rect 147201 142327 147235 142361
rect 147537 142327 147571 142361
rect 147873 142327 147907 142361
rect 148209 142327 148243 142361
rect 148545 142327 148579 142361
rect 148881 142327 148915 142361
rect 149217 142327 149251 142361
rect 149553 142327 149587 142361
rect 149889 142327 149923 142361
rect 150225 142327 150259 142361
rect 150561 142327 150595 142361
rect 150897 142327 150931 142361
rect 151233 142327 151267 142361
rect 151569 142327 151603 142361
rect 151905 142327 151939 142361
rect 152241 142327 152275 142361
rect 152577 142327 152611 142361
rect 152913 142327 152947 142361
rect 153249 142327 153283 142361
rect 153585 142327 153619 142361
rect 153921 142327 153955 142361
rect 154257 142327 154291 142361
rect 154593 142327 154627 142361
rect 154929 142327 154963 142361
rect 155265 142327 155299 142361
rect 155601 142327 155635 142361
rect 155937 142327 155971 142361
rect 156273 142327 156307 142361
rect 156609 142327 156643 142361
rect 156945 142327 156979 142361
rect 157281 142327 157315 142361
rect 157617 142327 157651 142361
rect 157953 142327 157987 142361
rect 158289 142327 158323 142361
rect 158625 142327 158659 142361
rect 158961 142327 158995 142361
rect 159297 142327 159331 142361
rect 159633 142327 159667 142361
rect 159969 142327 160003 142361
rect 160305 142327 160339 142361
rect 160641 142327 160675 142361
rect 160977 142327 161011 142361
rect 161313 142327 161347 142361
rect 161649 142327 161683 142361
rect 161985 142327 162019 142361
rect 162321 142327 162355 142361
rect 162657 142327 162691 142361
rect 162993 142327 163027 142361
rect 163329 142327 163363 142361
rect 163665 142327 163699 142361
rect 164001 142327 164035 142361
rect 164337 142327 164371 142361
rect 164673 142327 164707 142361
rect 165009 142327 165043 142361
rect 165345 142327 165379 142361
rect 165681 142327 165715 142361
rect 166017 142327 166051 142361
rect 166353 142327 166387 142361
rect 166689 142327 166723 142361
rect 167025 142327 167059 142361
rect 167361 142327 167395 142361
rect 167697 142327 167731 142361
rect 168033 142327 168067 142361
rect 168369 142327 168403 142361
rect 168705 142327 168739 142361
rect 169041 142327 169075 142361
rect 169377 142327 169411 142361
rect 169713 142327 169747 142361
rect 170049 142327 170083 142361
rect 170385 142327 170419 142361
rect 170721 142327 170755 142361
rect 171057 142327 171091 142361
rect 171393 142327 171427 142361
rect 171729 142327 171763 142361
rect 172065 142327 172099 142361
rect 172401 142327 172435 142361
rect 172737 142327 172771 142361
rect 173073 142327 173107 142361
rect 173409 142327 173443 142361
rect 173745 142327 173779 142361
rect 174081 142327 174115 142361
rect 174417 142327 174451 142361
rect 174753 142327 174787 142361
rect 175089 142327 175123 142361
rect 175425 142327 175459 142361
rect 175761 142327 175795 142361
rect 176097 142327 176131 142361
rect 176433 142327 176467 142361
rect 176769 142327 176803 142361
rect 177105 142327 177139 142361
rect 177441 142327 177475 142361
rect 177777 142327 177811 142361
rect 178113 142327 178147 142361
rect 178449 142327 178483 142361
rect 178785 142327 178819 142361
rect 179121 142327 179155 142361
rect 179457 142327 179491 142361
rect 179793 142327 179827 142361
rect 180129 142327 180163 142361
rect 180465 142327 180499 142361
rect 180801 142327 180835 142361
rect 181137 142327 181171 142361
rect 181473 142327 181507 142361
rect 181809 142327 181843 142361
rect 182145 142327 182179 142361
rect 182481 142327 182515 142361
rect 182817 142327 182851 142361
rect 183153 142327 183187 142361
rect 183489 142327 183523 142361
rect 183825 142327 183859 142361
rect 184161 142327 184195 142361
rect 184497 142327 184531 142361
rect 184833 142327 184867 142361
rect 185169 142327 185203 142361
rect 185505 142327 185539 142361
rect 185841 142327 185875 142361
rect 186177 142327 186211 142361
rect 186513 142327 186547 142361
rect 186849 142327 186883 142361
rect 187185 142327 187219 142361
rect 187521 142327 187555 142361
rect 187857 142327 187891 142361
rect 188193 142327 188227 142361
rect 188529 142327 188563 142361
rect 188865 142327 188899 142361
rect 189201 142327 189235 142361
rect 189537 142327 189571 142361
rect 189873 142327 189907 142361
rect 190209 142327 190243 142361
rect 190545 142327 190579 142361
rect 190881 142327 190915 142361
rect 191217 142327 191251 142361
rect 191553 142327 191587 142361
rect 191889 142327 191923 142361
rect 192225 142327 192259 142361
rect 192561 142327 192595 142361
rect 192897 142327 192931 142361
rect 193233 142327 193267 142361
rect 193569 142327 193603 142361
rect 193905 142327 193939 142361
rect 194241 142327 194275 142361
rect 194577 142327 194611 142361
rect 194913 142327 194947 142361
rect 195249 142327 195283 142361
rect 195585 142327 195619 142361
rect 195921 142327 195955 142361
rect 196257 142327 196291 142361
rect 196593 142327 196627 142361
rect 196929 142327 196963 142361
rect 197265 142327 197299 142361
rect 197601 142327 197635 142361
rect 197937 142327 197971 142361
rect 198273 142327 198307 142361
rect 198609 142327 198643 142361
rect 198945 142327 198979 142361
rect 199281 142327 199315 142361
rect 199617 142327 199651 142361
rect 199953 142327 199987 142361
rect 200289 142327 200323 142361
rect 200625 142327 200659 142361
rect 200961 142327 200995 142361
rect 201297 142327 201331 142361
rect 201633 142327 201667 142361
rect 201969 142327 202003 142361
rect 202305 142327 202339 142361
rect 202641 142327 202675 142361
rect 202977 142327 203011 142361
rect 203313 142327 203347 142361
rect 203649 142327 203683 142361
rect 203985 142327 204019 142361
rect 204321 142327 204355 142361
rect 204657 142327 204691 142361
rect 204993 142327 205027 142361
rect 205329 142327 205363 142361
rect 205665 142327 205699 142361
rect 206001 142327 206035 142361
rect 206337 142327 206371 142361
rect 206673 142327 206707 142361
rect 207009 142327 207043 142361
rect 207345 142327 207379 142361
rect 207681 142327 207715 142361
rect 208017 142327 208051 142361
rect 208353 142327 208387 142361
rect 208689 142327 208723 142361
rect 209025 142327 209059 142361
rect 209361 142327 209395 142361
rect 209697 142327 209731 142361
rect 210033 142327 210067 142361
rect 210369 142327 210403 142361
rect 210705 142327 210739 142361
rect 211041 142327 211075 142361
rect 211377 142327 211411 142361
rect 211713 142327 211747 142361
rect 212049 142327 212083 142361
rect 212385 142327 212419 142361
rect 212721 142327 212755 142361
rect 213057 142327 213091 142361
rect 213393 142327 213427 142361
rect 213729 142327 213763 142361
rect 214065 142327 214099 142361
rect 214401 142327 214435 142361
rect 214737 142327 214771 142361
rect 215073 142327 215107 142361
rect 215409 142327 215443 142361
rect 215745 142327 215779 142361
rect 216081 142327 216115 142361
rect 216417 142327 216451 142361
rect 1713 141943 1747 141977
rect 216919 141943 216953 141977
rect 1713 141607 1747 141641
rect 216919 141607 216953 141641
rect 1713 141271 1747 141305
rect 216919 141271 216953 141305
rect 1713 140935 1747 140969
rect 216919 140935 216953 140969
rect 1713 140599 1747 140633
rect 216919 140599 216953 140633
rect 1713 140263 1747 140297
rect 216919 140263 216953 140297
rect 1713 139927 1747 139961
rect 216919 139927 216953 139961
rect 1713 139591 1747 139625
rect 216919 139591 216953 139625
rect 1713 139255 1747 139289
rect 216919 139255 216953 139289
rect 1713 138919 1747 138953
rect 216919 138919 216953 138953
rect 1713 138583 1747 138617
rect 216919 138583 216953 138617
rect 1713 138247 1747 138281
rect 216919 138247 216953 138281
rect 1713 137911 1747 137945
rect 216919 137911 216953 137945
rect 1713 137575 1747 137609
rect 216919 137575 216953 137609
rect 1713 137239 1747 137273
rect 216919 137239 216953 137273
rect 1713 136903 1747 136937
rect 216919 136903 216953 136937
rect 1713 136567 1747 136601
rect 216919 136567 216953 136601
rect 1713 136231 1747 136265
rect 216919 136231 216953 136265
rect 1713 135895 1747 135929
rect 216919 135895 216953 135929
rect 1713 135559 1747 135593
rect 216919 135559 216953 135593
rect 1713 135223 1747 135257
rect 216919 135223 216953 135257
rect 1713 134887 1747 134921
rect 216919 134887 216953 134921
rect 1713 134551 1747 134585
rect 216919 134551 216953 134585
rect 1713 134215 1747 134249
rect 216919 134215 216953 134249
rect 1713 133879 1747 133913
rect 216919 133879 216953 133913
rect 1713 133543 1747 133577
rect 216919 133543 216953 133577
rect 1713 133207 1747 133241
rect 216919 133207 216953 133241
rect 1713 132871 1747 132905
rect 216919 132871 216953 132905
rect 1713 132535 1747 132569
rect 216919 132535 216953 132569
rect 1713 132199 1747 132233
rect 216919 132199 216953 132233
rect 1713 131863 1747 131897
rect 216919 131863 216953 131897
rect 1713 131527 1747 131561
rect 216919 131527 216953 131561
rect 1713 131191 1747 131225
rect 216919 131191 216953 131225
rect 1713 130855 1747 130889
rect 216919 130855 216953 130889
rect 1713 130519 1747 130553
rect 216919 130519 216953 130553
rect 1713 130183 1747 130217
rect 216919 130183 216953 130217
rect 1713 129847 1747 129881
rect 216919 129847 216953 129881
rect 1713 129511 1747 129545
rect 216919 129511 216953 129545
rect 1713 129175 1747 129209
rect 216919 129175 216953 129209
rect 1713 128839 1747 128873
rect 216919 128839 216953 128873
rect 1713 128503 1747 128537
rect 216919 128503 216953 128537
rect 1713 128167 1747 128201
rect 216919 128167 216953 128201
rect 1713 127831 1747 127865
rect 216919 127831 216953 127865
rect 1713 127495 1747 127529
rect 216919 127495 216953 127529
rect 1713 127159 1747 127193
rect 216919 127159 216953 127193
rect 1713 126823 1747 126857
rect 216919 126823 216953 126857
rect 1713 126487 1747 126521
rect 216919 126487 216953 126521
rect 1713 126151 1747 126185
rect 216919 126151 216953 126185
rect 1713 125815 1747 125849
rect 216919 125815 216953 125849
rect 1713 125479 1747 125513
rect 216919 125479 216953 125513
rect 1713 125143 1747 125177
rect 216919 125143 216953 125177
rect 1713 124807 1747 124841
rect 216919 124807 216953 124841
rect 1713 124471 1747 124505
rect 216919 124471 216953 124505
rect 1713 124135 1747 124169
rect 216919 124135 216953 124169
rect 1713 123799 1747 123833
rect 216919 123799 216953 123833
rect 1713 123463 1747 123497
rect 216919 123463 216953 123497
rect 1713 123127 1747 123161
rect 216919 123127 216953 123161
rect 1713 122791 1747 122825
rect 216919 122791 216953 122825
rect 1713 122455 1747 122489
rect 216919 122455 216953 122489
rect 1713 122119 1747 122153
rect 216919 122119 216953 122153
rect 1713 121783 1747 121817
rect 216919 121783 216953 121817
rect 1713 121447 1747 121481
rect 216919 121447 216953 121481
rect 1713 121111 1747 121145
rect 216919 121111 216953 121145
rect 1713 120775 1747 120809
rect 216919 120775 216953 120809
rect 1713 120439 1747 120473
rect 216919 120439 216953 120473
rect 1713 120103 1747 120137
rect 216919 120103 216953 120137
rect 1713 119767 1747 119801
rect 216919 119767 216953 119801
rect 1713 119431 1747 119465
rect 216919 119431 216953 119465
rect 1713 119095 1747 119129
rect 216919 119095 216953 119129
rect 1713 118759 1747 118793
rect 216919 118759 216953 118793
rect 1713 118423 1747 118457
rect 216919 118423 216953 118457
rect 1713 118087 1747 118121
rect 216919 118087 216953 118121
rect 1713 117751 1747 117785
rect 216919 117751 216953 117785
rect 1713 117415 1747 117449
rect 216919 117415 216953 117449
rect 1713 117079 1747 117113
rect 216919 117079 216953 117113
rect 1713 116743 1747 116777
rect 216919 116743 216953 116777
rect 1713 116407 1747 116441
rect 216919 116407 216953 116441
rect 1713 116071 1747 116105
rect 216919 116071 216953 116105
rect 1713 115735 1747 115769
rect 216919 115735 216953 115769
rect 1713 115399 1747 115433
rect 216919 115399 216953 115433
rect 1713 115063 1747 115097
rect 216919 115063 216953 115097
rect 1713 114727 1747 114761
rect 216919 114727 216953 114761
rect 1713 114391 1747 114425
rect 216919 114391 216953 114425
rect 1713 114055 1747 114089
rect 216919 114055 216953 114089
rect 1713 113719 1747 113753
rect 216919 113719 216953 113753
rect 1713 113383 1747 113417
rect 216919 113383 216953 113417
rect 1713 113047 1747 113081
rect 216919 113047 216953 113081
rect 1713 112711 1747 112745
rect 216919 112711 216953 112745
rect 1713 112375 1747 112409
rect 216919 112375 216953 112409
rect 1713 112039 1747 112073
rect 216919 112039 216953 112073
rect 1713 111703 1747 111737
rect 216919 111703 216953 111737
rect 1713 111367 1747 111401
rect 216919 111367 216953 111401
rect 1713 111031 1747 111065
rect 216919 111031 216953 111065
rect 1713 110695 1747 110729
rect 216919 110695 216953 110729
rect 1713 110359 1747 110393
rect 216919 110359 216953 110393
rect 1713 110023 1747 110057
rect 216919 110023 216953 110057
rect 1713 109687 1747 109721
rect 216919 109687 216953 109721
rect 1713 109351 1747 109385
rect 216919 109351 216953 109385
rect 1713 109015 1747 109049
rect 216919 109015 216953 109049
rect 1713 108679 1747 108713
rect 216919 108679 216953 108713
rect 1713 108343 1747 108377
rect 216919 108343 216953 108377
rect 1713 108007 1747 108041
rect 216919 108007 216953 108041
rect 1713 107671 1747 107705
rect 216919 107671 216953 107705
rect 1713 107335 1747 107369
rect 216919 107335 216953 107369
rect 1713 106999 1747 107033
rect 216919 106999 216953 107033
rect 1713 106663 1747 106697
rect 216919 106663 216953 106697
rect 1713 106327 1747 106361
rect 216919 106327 216953 106361
rect 1713 105991 1747 106025
rect 216919 105991 216953 106025
rect 1713 105655 1747 105689
rect 216919 105655 216953 105689
rect 1713 105319 1747 105353
rect 216919 105319 216953 105353
rect 1713 104983 1747 105017
rect 216919 104983 216953 105017
rect 1713 104647 1747 104681
rect 216919 104647 216953 104681
rect 1713 104311 1747 104345
rect 216919 104311 216953 104345
rect 1713 103975 1747 104009
rect 216919 103975 216953 104009
rect 1713 103639 1747 103673
rect 216919 103639 216953 103673
rect 1713 103303 1747 103337
rect 216919 103303 216953 103337
rect 1713 102967 1747 103001
rect 216919 102967 216953 103001
rect 1713 102631 1747 102665
rect 216919 102631 216953 102665
rect 1713 102295 1747 102329
rect 216919 102295 216953 102329
rect 1713 101959 1747 101993
rect 216919 101959 216953 101993
rect 1713 101623 1747 101657
rect 216919 101623 216953 101657
rect 1713 101287 1747 101321
rect 216919 101287 216953 101321
rect 1713 100951 1747 100985
rect 216919 100951 216953 100985
rect 1713 100615 1747 100649
rect 216919 100615 216953 100649
rect 1713 100279 1747 100313
rect 216919 100279 216953 100313
rect 1713 99943 1747 99977
rect 216919 99943 216953 99977
rect 1713 99607 1747 99641
rect 216919 99607 216953 99641
rect 1713 99271 1747 99305
rect 216919 99271 216953 99305
rect 1713 98935 1747 98969
rect 216919 98935 216953 98969
rect 1713 98599 1747 98633
rect 216919 98599 216953 98633
rect 1713 98263 1747 98297
rect 216919 98263 216953 98297
rect 1713 97927 1747 97961
rect 216919 97927 216953 97961
rect 1713 97591 1747 97625
rect 216919 97591 216953 97625
rect 1713 97255 1747 97289
rect 216919 97255 216953 97289
rect 1713 96919 1747 96953
rect 216919 96919 216953 96953
rect 1713 96583 1747 96617
rect 216919 96583 216953 96617
rect 1713 96247 1747 96281
rect 216919 96247 216953 96281
rect 1713 95911 1747 95945
rect 216919 95911 216953 95945
rect 1713 95575 1747 95609
rect 216919 95575 216953 95609
rect 1713 95239 1747 95273
rect 216919 95239 216953 95273
rect 1713 94903 1747 94937
rect 216919 94903 216953 94937
rect 1713 94567 1747 94601
rect 216919 94567 216953 94601
rect 1713 94231 1747 94265
rect 216919 94231 216953 94265
rect 1713 93895 1747 93929
rect 216919 93895 216953 93929
rect 1713 93559 1747 93593
rect 216919 93559 216953 93593
rect 1713 93223 1747 93257
rect 216919 93223 216953 93257
rect 1713 92887 1747 92921
rect 216919 92887 216953 92921
rect 1713 92551 1747 92585
rect 216919 92551 216953 92585
rect 1713 92215 1747 92249
rect 216919 92215 216953 92249
rect 1713 91879 1747 91913
rect 216919 91879 216953 91913
rect 1713 91543 1747 91577
rect 216919 91543 216953 91577
rect 1713 91207 1747 91241
rect 216919 91207 216953 91241
rect 1713 90871 1747 90905
rect 216919 90871 216953 90905
rect 1713 90535 1747 90569
rect 216919 90535 216953 90569
rect 1713 90199 1747 90233
rect 216919 90199 216953 90233
rect 1713 89863 1747 89897
rect 216919 89863 216953 89897
rect 1713 89527 1747 89561
rect 216919 89527 216953 89561
rect 1713 89191 1747 89225
rect 216919 89191 216953 89225
rect 1713 88855 1747 88889
rect 216919 88855 216953 88889
rect 1713 88519 1747 88553
rect 216919 88519 216953 88553
rect 1713 88183 1747 88217
rect 216919 88183 216953 88217
rect 1713 87847 1747 87881
rect 216919 87847 216953 87881
rect 1713 87511 1747 87545
rect 216919 87511 216953 87545
rect 1713 87175 1747 87209
rect 216919 87175 216953 87209
rect 1713 86839 1747 86873
rect 216919 86839 216953 86873
rect 1713 86503 1747 86537
rect 216919 86503 216953 86537
rect 1713 86167 1747 86201
rect 216919 86167 216953 86201
rect 1713 85831 1747 85865
rect 216919 85831 216953 85865
rect 1713 85495 1747 85529
rect 216919 85495 216953 85529
rect 1713 85159 1747 85193
rect 216919 85159 216953 85193
rect 1713 84823 1747 84857
rect 216919 84823 216953 84857
rect 1713 84487 1747 84521
rect 216919 84487 216953 84521
rect 1713 84151 1747 84185
rect 216919 84151 216953 84185
rect 1713 83815 1747 83849
rect 216919 83815 216953 83849
rect 1713 83479 1747 83513
rect 216919 83479 216953 83513
rect 1713 83143 1747 83177
rect 216919 83143 216953 83177
rect 1713 82807 1747 82841
rect 216919 82807 216953 82841
rect 1713 82471 1747 82505
rect 216919 82471 216953 82505
rect 1713 82135 1747 82169
rect 216919 82135 216953 82169
rect 1713 81799 1747 81833
rect 216919 81799 216953 81833
rect 1713 81463 1747 81497
rect 216919 81463 216953 81497
rect 1713 81127 1747 81161
rect 216919 81127 216953 81161
rect 1713 80791 1747 80825
rect 216919 80791 216953 80825
rect 1713 80455 1747 80489
rect 216919 80455 216953 80489
rect 1713 80119 1747 80153
rect 216919 80119 216953 80153
rect 1713 79783 1747 79817
rect 216919 79783 216953 79817
rect 1713 79447 1747 79481
rect 216919 79447 216953 79481
rect 1713 79111 1747 79145
rect 216919 79111 216953 79145
rect 1713 78775 1747 78809
rect 216919 78775 216953 78809
rect 1713 78439 1747 78473
rect 216919 78439 216953 78473
rect 1713 78103 1747 78137
rect 216919 78103 216953 78137
rect 1713 77767 1747 77801
rect 216919 77767 216953 77801
rect 1713 77431 1747 77465
rect 216919 77431 216953 77465
rect 1713 77095 1747 77129
rect 216919 77095 216953 77129
rect 1713 76759 1747 76793
rect 216919 76759 216953 76793
rect 1713 76423 1747 76457
rect 216919 76423 216953 76457
rect 1713 76087 1747 76121
rect 216919 76087 216953 76121
rect 1713 75751 1747 75785
rect 216919 75751 216953 75785
rect 1713 75415 1747 75449
rect 216919 75415 216953 75449
rect 1713 75079 1747 75113
rect 216919 75079 216953 75113
rect 1713 74743 1747 74777
rect 216919 74743 216953 74777
rect 1713 74407 1747 74441
rect 216919 74407 216953 74441
rect 1713 74071 1747 74105
rect 216919 74071 216953 74105
rect 1713 73735 1747 73769
rect 216919 73735 216953 73769
rect 1713 73399 1747 73433
rect 216919 73399 216953 73433
rect 1713 73063 1747 73097
rect 216919 73063 216953 73097
rect 1713 72727 1747 72761
rect 216919 72727 216953 72761
rect 1713 72391 1747 72425
rect 216919 72391 216953 72425
rect 1713 72055 1747 72089
rect 216919 72055 216953 72089
rect 1713 71719 1747 71753
rect 216919 71719 216953 71753
rect 1713 71383 1747 71417
rect 216919 71383 216953 71417
rect 1713 71047 1747 71081
rect 216919 71047 216953 71081
rect 1713 70711 1747 70745
rect 216919 70711 216953 70745
rect 1713 70375 1747 70409
rect 216919 70375 216953 70409
rect 1713 70039 1747 70073
rect 216919 70039 216953 70073
rect 1713 69703 1747 69737
rect 216919 69703 216953 69737
rect 1713 69367 1747 69401
rect 216919 69367 216953 69401
rect 1713 69031 1747 69065
rect 216919 69031 216953 69065
rect 1713 68695 1747 68729
rect 216919 68695 216953 68729
rect 1713 68359 1747 68393
rect 216919 68359 216953 68393
rect 1713 68023 1747 68057
rect 216919 68023 216953 68057
rect 1713 67687 1747 67721
rect 216919 67687 216953 67721
rect 1713 67351 1747 67385
rect 216919 67351 216953 67385
rect 1713 67015 1747 67049
rect 216919 67015 216953 67049
rect 1713 66679 1747 66713
rect 216919 66679 216953 66713
rect 1713 66343 1747 66377
rect 216919 66343 216953 66377
rect 1713 66007 1747 66041
rect 216919 66007 216953 66041
rect 1713 65671 1747 65705
rect 216919 65671 216953 65705
rect 1713 65335 1747 65369
rect 216919 65335 216953 65369
rect 1713 64999 1747 65033
rect 216919 64999 216953 65033
rect 1713 64663 1747 64697
rect 216919 64663 216953 64697
rect 1713 64327 1747 64361
rect 216919 64327 216953 64361
rect 1713 63991 1747 64025
rect 216919 63991 216953 64025
rect 1713 63655 1747 63689
rect 216919 63655 216953 63689
rect 1713 63319 1747 63353
rect 216919 63319 216953 63353
rect 1713 62983 1747 63017
rect 216919 62983 216953 63017
rect 1713 62647 1747 62681
rect 216919 62647 216953 62681
rect 1713 62311 1747 62345
rect 216919 62311 216953 62345
rect 1713 61975 1747 62009
rect 216919 61975 216953 62009
rect 1713 61639 1747 61673
rect 216919 61639 216953 61673
rect 1713 61303 1747 61337
rect 216919 61303 216953 61337
rect 1713 60967 1747 61001
rect 216919 60967 216953 61001
rect 1713 60631 1747 60665
rect 216919 60631 216953 60665
rect 1713 60295 1747 60329
rect 216919 60295 216953 60329
rect 1713 59959 1747 59993
rect 216919 59959 216953 59993
rect 1713 59623 1747 59657
rect 216919 59623 216953 59657
rect 1713 59287 1747 59321
rect 216919 59287 216953 59321
rect 1713 58951 1747 58985
rect 216919 58951 216953 58985
rect 1713 58615 1747 58649
rect 216919 58615 216953 58649
rect 1713 58279 1747 58313
rect 216919 58279 216953 58313
rect 1713 57943 1747 57977
rect 216919 57943 216953 57977
rect 1713 57607 1747 57641
rect 216919 57607 216953 57641
rect 1713 57271 1747 57305
rect 216919 57271 216953 57305
rect 1713 56935 1747 56969
rect 216919 56935 216953 56969
rect 1713 56599 1747 56633
rect 216919 56599 216953 56633
rect 1713 56263 1747 56297
rect 216919 56263 216953 56297
rect 1713 55927 1747 55961
rect 216919 55927 216953 55961
rect 1713 55591 1747 55625
rect 216919 55591 216953 55625
rect 1713 55255 1747 55289
rect 216919 55255 216953 55289
rect 1713 54919 1747 54953
rect 216919 54919 216953 54953
rect 1713 54583 1747 54617
rect 216919 54583 216953 54617
rect 1713 54247 1747 54281
rect 216919 54247 216953 54281
rect 1713 53911 1747 53945
rect 216919 53911 216953 53945
rect 1713 53575 1747 53609
rect 216919 53575 216953 53609
rect 1713 53239 1747 53273
rect 216919 53239 216953 53273
rect 1713 52903 1747 52937
rect 216919 52903 216953 52937
rect 1713 52567 1747 52601
rect 216919 52567 216953 52601
rect 1713 52231 1747 52265
rect 216919 52231 216953 52265
rect 1713 51895 1747 51929
rect 216919 51895 216953 51929
rect 1713 51559 1747 51593
rect 216919 51559 216953 51593
rect 1713 51223 1747 51257
rect 216919 51223 216953 51257
rect 1713 50887 1747 50921
rect 216919 50887 216953 50921
rect 1713 50551 1747 50585
rect 216919 50551 216953 50585
rect 1713 50215 1747 50249
rect 216919 50215 216953 50249
rect 1713 49879 1747 49913
rect 216919 49879 216953 49913
rect 1713 49543 1747 49577
rect 216919 49543 216953 49577
rect 1713 49207 1747 49241
rect 216919 49207 216953 49241
rect 1713 48871 1747 48905
rect 216919 48871 216953 48905
rect 1713 48535 1747 48569
rect 216919 48535 216953 48569
rect 1713 48199 1747 48233
rect 216919 48199 216953 48233
rect 1713 47863 1747 47897
rect 216919 47863 216953 47897
rect 1713 47527 1747 47561
rect 216919 47527 216953 47561
rect 1713 47191 1747 47225
rect 216919 47191 216953 47225
rect 1713 46855 1747 46889
rect 216919 46855 216953 46889
rect 1713 46519 1747 46553
rect 216919 46519 216953 46553
rect 1713 46183 1747 46217
rect 216919 46183 216953 46217
rect 1713 45847 1747 45881
rect 216919 45847 216953 45881
rect 1713 45511 1747 45545
rect 216919 45511 216953 45545
rect 1713 45175 1747 45209
rect 216919 45175 216953 45209
rect 1713 44839 1747 44873
rect 216919 44839 216953 44873
rect 1713 44503 1747 44537
rect 216919 44503 216953 44537
rect 1713 44167 1747 44201
rect 216919 44167 216953 44201
rect 1713 43831 1747 43865
rect 216919 43831 216953 43865
rect 1713 43495 1747 43529
rect 216919 43495 216953 43529
rect 1713 43159 1747 43193
rect 216919 43159 216953 43193
rect 1713 42823 1747 42857
rect 216919 42823 216953 42857
rect 1713 42487 1747 42521
rect 216919 42487 216953 42521
rect 1713 42151 1747 42185
rect 216919 42151 216953 42185
rect 1713 41815 1747 41849
rect 216919 41815 216953 41849
rect 1713 41479 1747 41513
rect 216919 41479 216953 41513
rect 1713 41143 1747 41177
rect 216919 41143 216953 41177
rect 1713 40807 1747 40841
rect 216919 40807 216953 40841
rect 1713 40471 1747 40505
rect 216919 40471 216953 40505
rect 1713 40135 1747 40169
rect 216919 40135 216953 40169
rect 1713 39799 1747 39833
rect 216919 39799 216953 39833
rect 1713 39463 1747 39497
rect 216919 39463 216953 39497
rect 1713 39127 1747 39161
rect 216919 39127 216953 39161
rect 1713 38791 1747 38825
rect 216919 38791 216953 38825
rect 1713 38455 1747 38489
rect 216919 38455 216953 38489
rect 1713 38119 1747 38153
rect 216919 38119 216953 38153
rect 1713 37783 1747 37817
rect 216919 37783 216953 37817
rect 1713 37447 1747 37481
rect 216919 37447 216953 37481
rect 1713 37111 1747 37145
rect 216919 37111 216953 37145
rect 1713 36775 1747 36809
rect 216919 36775 216953 36809
rect 1713 36439 1747 36473
rect 216919 36439 216953 36473
rect 1713 36103 1747 36137
rect 216919 36103 216953 36137
rect 1713 35767 1747 35801
rect 216919 35767 216953 35801
rect 1713 35431 1747 35465
rect 216919 35431 216953 35465
rect 1713 35095 1747 35129
rect 216919 35095 216953 35129
rect 1713 34759 1747 34793
rect 216919 34759 216953 34793
rect 1713 34423 1747 34457
rect 216919 34423 216953 34457
rect 1713 34087 1747 34121
rect 216919 34087 216953 34121
rect 1713 33751 1747 33785
rect 216919 33751 216953 33785
rect 1713 33415 1747 33449
rect 216919 33415 216953 33449
rect 1713 33079 1747 33113
rect 216919 33079 216953 33113
rect 1713 32743 1747 32777
rect 216919 32743 216953 32777
rect 1713 32407 1747 32441
rect 216919 32407 216953 32441
rect 1713 32071 1747 32105
rect 216919 32071 216953 32105
rect 1713 31735 1747 31769
rect 216919 31735 216953 31769
rect 1713 31399 1747 31433
rect 216919 31399 216953 31433
rect 1713 31063 1747 31097
rect 216919 31063 216953 31097
rect 1713 30727 1747 30761
rect 216919 30727 216953 30761
rect 1713 30391 1747 30425
rect 216919 30391 216953 30425
rect 1713 30055 1747 30089
rect 216919 30055 216953 30089
rect 1713 29719 1747 29753
rect 216919 29719 216953 29753
rect 1713 29383 1747 29417
rect 216919 29383 216953 29417
rect 1713 29047 1747 29081
rect 216919 29047 216953 29081
rect 1713 28711 1747 28745
rect 216919 28711 216953 28745
rect 1713 28375 1747 28409
rect 216919 28375 216953 28409
rect 1713 28039 1747 28073
rect 216919 28039 216953 28073
rect 1713 27703 1747 27737
rect 216919 27703 216953 27737
rect 1713 27367 1747 27401
rect 216919 27367 216953 27401
rect 1713 27031 1747 27065
rect 216919 27031 216953 27065
rect 1713 26695 1747 26729
rect 216919 26695 216953 26729
rect 1713 26359 1747 26393
rect 216919 26359 216953 26393
rect 1713 26023 1747 26057
rect 216919 26023 216953 26057
rect 1713 25687 1747 25721
rect 216919 25687 216953 25721
rect 1713 25351 1747 25385
rect 216919 25351 216953 25385
rect 1713 25015 1747 25049
rect 216919 25015 216953 25049
rect 1713 24679 1747 24713
rect 216919 24679 216953 24713
rect 1713 24343 1747 24377
rect 216919 24343 216953 24377
rect 1713 24007 1747 24041
rect 216919 24007 216953 24041
rect 1713 23671 1747 23705
rect 216919 23671 216953 23705
rect 1713 23335 1747 23369
rect 216919 23335 216953 23369
rect 1713 22999 1747 23033
rect 216919 22999 216953 23033
rect 1713 22663 1747 22697
rect 216919 22663 216953 22697
rect 1713 22327 1747 22361
rect 216919 22327 216953 22361
rect 1713 21991 1747 22025
rect 216919 21991 216953 22025
rect 1713 21655 1747 21689
rect 216919 21655 216953 21689
rect 1713 21319 1747 21353
rect 216919 21319 216953 21353
rect 1713 20983 1747 21017
rect 216919 20983 216953 21017
rect 1713 20647 1747 20681
rect 216919 20647 216953 20681
rect 1713 20311 1747 20345
rect 216919 20311 216953 20345
rect 1713 19975 1747 20009
rect 216919 19975 216953 20009
rect 1713 19639 1747 19673
rect 216919 19639 216953 19673
rect 1713 19303 1747 19337
rect 216919 19303 216953 19337
rect 1713 18967 1747 19001
rect 216919 18967 216953 19001
rect 1713 18631 1747 18665
rect 216919 18631 216953 18665
rect 1713 18295 1747 18329
rect 216919 18295 216953 18329
rect 1713 17959 1747 17993
rect 216919 17959 216953 17993
rect 1713 17623 1747 17657
rect 216919 17623 216953 17657
rect 1713 17287 1747 17321
rect 216919 17287 216953 17321
rect 1713 16951 1747 16985
rect 216919 16951 216953 16985
rect 1713 16615 1747 16649
rect 216919 16615 216953 16649
rect 1713 16279 1747 16313
rect 216919 16279 216953 16313
rect 1713 15943 1747 15977
rect 216919 15943 216953 15977
rect 1713 15607 1747 15641
rect 216919 15607 216953 15641
rect 1713 15271 1747 15305
rect 216919 15271 216953 15305
rect 1713 14935 1747 14969
rect 216919 14935 216953 14969
rect 1713 14599 1747 14633
rect 216919 14599 216953 14633
rect 1713 14263 1747 14297
rect 216919 14263 216953 14297
rect 1713 13927 1747 13961
rect 216919 13927 216953 13961
rect 1713 13591 1747 13625
rect 216919 13591 216953 13625
rect 1713 13255 1747 13289
rect 216919 13255 216953 13289
rect 1713 12919 1747 12953
rect 216919 12919 216953 12953
rect 1713 12583 1747 12617
rect 216919 12583 216953 12617
rect 1713 12247 1747 12281
rect 216919 12247 216953 12281
rect 1713 11911 1747 11945
rect 216919 11911 216953 11945
rect 1713 11575 1747 11609
rect 216919 11575 216953 11609
rect 1713 11239 1747 11273
rect 216919 11239 216953 11273
rect 1713 10903 1747 10937
rect 216919 10903 216953 10937
rect 1713 10567 1747 10601
rect 216919 10567 216953 10601
rect 1713 10231 1747 10265
rect 216919 10231 216953 10265
rect 1713 9895 1747 9929
rect 216919 9895 216953 9929
rect 1713 9559 1747 9593
rect 216919 9559 216953 9593
rect 1713 9223 1747 9257
rect 216919 9223 216953 9257
rect 1713 8887 1747 8921
rect 216919 8887 216953 8921
rect 1713 8551 1747 8585
rect 216919 8551 216953 8585
rect 1713 8215 1747 8249
rect 216919 8215 216953 8249
rect 1713 7879 1747 7913
rect 216919 7879 216953 7913
rect 1713 7543 1747 7577
rect 216919 7543 216953 7577
rect 1713 7207 1747 7241
rect 216919 7207 216953 7241
rect 1713 6871 1747 6905
rect 216919 6871 216953 6905
rect 1713 6535 1747 6569
rect 216919 6535 216953 6569
rect 1713 6199 1747 6233
rect 216919 6199 216953 6233
rect 1713 5863 1747 5897
rect 216919 5863 216953 5897
rect 1713 5527 1747 5561
rect 216919 5527 216953 5561
rect 1713 5191 1747 5225
rect 216919 5191 216953 5225
rect 1713 4855 1747 4889
rect 216919 4855 216953 4889
rect 1713 4519 1747 4553
rect 216919 4519 216953 4553
rect 1713 4183 1747 4217
rect 216919 4183 216953 4217
rect 1713 3847 1747 3881
rect 216919 3847 216953 3881
rect 1713 3511 1747 3545
rect 216919 3511 216953 3545
rect 1713 3175 1747 3209
rect 216919 3175 216953 3209
rect 1713 2839 1747 2873
rect 216919 2839 216953 2873
rect 1713 2503 1747 2537
rect 216919 2503 216953 2537
rect 1713 2167 1747 2201
rect 216919 2167 216953 2201
rect 2049 1831 2083 1865
rect 2385 1831 2419 1865
rect 2721 1831 2755 1865
rect 3057 1831 3091 1865
rect 3393 1831 3427 1865
rect 3729 1831 3763 1865
rect 4065 1831 4099 1865
rect 4401 1831 4435 1865
rect 4737 1831 4771 1865
rect 5073 1831 5107 1865
rect 5409 1831 5443 1865
rect 5745 1831 5779 1865
rect 6081 1831 6115 1865
rect 6417 1831 6451 1865
rect 6753 1831 6787 1865
rect 7089 1831 7123 1865
rect 7425 1831 7459 1865
rect 7761 1831 7795 1865
rect 8097 1831 8131 1865
rect 8433 1831 8467 1865
rect 8769 1831 8803 1865
rect 9105 1831 9139 1865
rect 9441 1831 9475 1865
rect 9777 1831 9811 1865
rect 10113 1831 10147 1865
rect 10449 1831 10483 1865
rect 10785 1831 10819 1865
rect 11121 1831 11155 1865
rect 11457 1831 11491 1865
rect 11793 1831 11827 1865
rect 12129 1831 12163 1865
rect 12465 1831 12499 1865
rect 12801 1831 12835 1865
rect 13137 1831 13171 1865
rect 13473 1831 13507 1865
rect 13809 1831 13843 1865
rect 14145 1831 14179 1865
rect 14481 1831 14515 1865
rect 14817 1831 14851 1865
rect 15153 1831 15187 1865
rect 15489 1831 15523 1865
rect 15825 1831 15859 1865
rect 16161 1831 16195 1865
rect 16497 1831 16531 1865
rect 16833 1831 16867 1865
rect 17169 1831 17203 1865
rect 17505 1831 17539 1865
rect 17841 1831 17875 1865
rect 18177 1831 18211 1865
rect 18513 1831 18547 1865
rect 18849 1831 18883 1865
rect 19185 1831 19219 1865
rect 19521 1831 19555 1865
rect 19857 1831 19891 1865
rect 20193 1831 20227 1865
rect 20529 1831 20563 1865
rect 20865 1831 20899 1865
rect 21201 1831 21235 1865
rect 21537 1831 21571 1865
rect 21873 1831 21907 1865
rect 22209 1831 22243 1865
rect 22545 1831 22579 1865
rect 22881 1831 22915 1865
rect 23217 1831 23251 1865
rect 23553 1831 23587 1865
rect 23889 1831 23923 1865
rect 24225 1831 24259 1865
rect 24561 1831 24595 1865
rect 24897 1831 24931 1865
rect 25233 1831 25267 1865
rect 25569 1831 25603 1865
rect 25905 1831 25939 1865
rect 26241 1831 26275 1865
rect 26577 1831 26611 1865
rect 26913 1831 26947 1865
rect 27249 1831 27283 1865
rect 27585 1831 27619 1865
rect 27921 1831 27955 1865
rect 28257 1831 28291 1865
rect 28593 1831 28627 1865
rect 28929 1831 28963 1865
rect 29265 1831 29299 1865
rect 29601 1831 29635 1865
rect 29937 1831 29971 1865
rect 30273 1831 30307 1865
rect 30609 1831 30643 1865
rect 30945 1831 30979 1865
rect 31281 1831 31315 1865
rect 31617 1831 31651 1865
rect 31953 1831 31987 1865
rect 32289 1831 32323 1865
rect 32625 1831 32659 1865
rect 32961 1831 32995 1865
rect 33297 1831 33331 1865
rect 33633 1831 33667 1865
rect 33969 1831 34003 1865
rect 34305 1831 34339 1865
rect 34641 1831 34675 1865
rect 34977 1831 35011 1865
rect 35313 1831 35347 1865
rect 35649 1831 35683 1865
rect 35985 1831 36019 1865
rect 36321 1831 36355 1865
rect 36657 1831 36691 1865
rect 36993 1831 37027 1865
rect 37329 1831 37363 1865
rect 37665 1831 37699 1865
rect 38001 1831 38035 1865
rect 38337 1831 38371 1865
rect 38673 1831 38707 1865
rect 39009 1831 39043 1865
rect 39345 1831 39379 1865
rect 39681 1831 39715 1865
rect 40017 1831 40051 1865
rect 40353 1831 40387 1865
rect 40689 1831 40723 1865
rect 41025 1831 41059 1865
rect 41361 1831 41395 1865
rect 41697 1831 41731 1865
rect 42033 1831 42067 1865
rect 42369 1831 42403 1865
rect 42705 1831 42739 1865
rect 43041 1831 43075 1865
rect 43377 1831 43411 1865
rect 43713 1831 43747 1865
rect 44049 1831 44083 1865
rect 44385 1831 44419 1865
rect 44721 1831 44755 1865
rect 45057 1831 45091 1865
rect 45393 1831 45427 1865
rect 45729 1831 45763 1865
rect 46065 1831 46099 1865
rect 46401 1831 46435 1865
rect 46737 1831 46771 1865
rect 47073 1831 47107 1865
rect 47409 1831 47443 1865
rect 47745 1831 47779 1865
rect 48081 1831 48115 1865
rect 48417 1831 48451 1865
rect 48753 1831 48787 1865
rect 49089 1831 49123 1865
rect 49425 1831 49459 1865
rect 49761 1831 49795 1865
rect 50097 1831 50131 1865
rect 50433 1831 50467 1865
rect 50769 1831 50803 1865
rect 51105 1831 51139 1865
rect 51441 1831 51475 1865
rect 51777 1831 51811 1865
rect 52113 1831 52147 1865
rect 52449 1831 52483 1865
rect 52785 1831 52819 1865
rect 53121 1831 53155 1865
rect 53457 1831 53491 1865
rect 53793 1831 53827 1865
rect 54129 1831 54163 1865
rect 54465 1831 54499 1865
rect 54801 1831 54835 1865
rect 55137 1831 55171 1865
rect 55473 1831 55507 1865
rect 55809 1831 55843 1865
rect 56145 1831 56179 1865
rect 56481 1831 56515 1865
rect 56817 1831 56851 1865
rect 57153 1831 57187 1865
rect 57489 1831 57523 1865
rect 57825 1831 57859 1865
rect 58161 1831 58195 1865
rect 58497 1831 58531 1865
rect 58833 1831 58867 1865
rect 59169 1831 59203 1865
rect 59505 1831 59539 1865
rect 59841 1831 59875 1865
rect 60177 1831 60211 1865
rect 60513 1831 60547 1865
rect 60849 1831 60883 1865
rect 61185 1831 61219 1865
rect 61521 1831 61555 1865
rect 61857 1831 61891 1865
rect 62193 1831 62227 1865
rect 62529 1831 62563 1865
rect 62865 1831 62899 1865
rect 63201 1831 63235 1865
rect 63537 1831 63571 1865
rect 63873 1831 63907 1865
rect 64209 1831 64243 1865
rect 64545 1831 64579 1865
rect 64881 1831 64915 1865
rect 65217 1831 65251 1865
rect 65553 1831 65587 1865
rect 65889 1831 65923 1865
rect 66225 1831 66259 1865
rect 66561 1831 66595 1865
rect 66897 1831 66931 1865
rect 67233 1831 67267 1865
rect 67569 1831 67603 1865
rect 67905 1831 67939 1865
rect 68241 1831 68275 1865
rect 68577 1831 68611 1865
rect 68913 1831 68947 1865
rect 69249 1831 69283 1865
rect 69585 1831 69619 1865
rect 69921 1831 69955 1865
rect 70257 1831 70291 1865
rect 70593 1831 70627 1865
rect 70929 1831 70963 1865
rect 71265 1831 71299 1865
rect 71601 1831 71635 1865
rect 71937 1831 71971 1865
rect 72273 1831 72307 1865
rect 72609 1831 72643 1865
rect 72945 1831 72979 1865
rect 73281 1831 73315 1865
rect 73617 1831 73651 1865
rect 73953 1831 73987 1865
rect 74289 1831 74323 1865
rect 74625 1831 74659 1865
rect 74961 1831 74995 1865
rect 75297 1831 75331 1865
rect 75633 1831 75667 1865
rect 75969 1831 76003 1865
rect 76305 1831 76339 1865
rect 76641 1831 76675 1865
rect 76977 1831 77011 1865
rect 77313 1831 77347 1865
rect 77649 1831 77683 1865
rect 77985 1831 78019 1865
rect 78321 1831 78355 1865
rect 78657 1831 78691 1865
rect 78993 1831 79027 1865
rect 79329 1831 79363 1865
rect 79665 1831 79699 1865
rect 80001 1831 80035 1865
rect 80337 1831 80371 1865
rect 80673 1831 80707 1865
rect 81009 1831 81043 1865
rect 81345 1831 81379 1865
rect 81681 1831 81715 1865
rect 82017 1831 82051 1865
rect 82353 1831 82387 1865
rect 82689 1831 82723 1865
rect 83025 1831 83059 1865
rect 83361 1831 83395 1865
rect 83697 1831 83731 1865
rect 84033 1831 84067 1865
rect 84369 1831 84403 1865
rect 84705 1831 84739 1865
rect 85041 1831 85075 1865
rect 85377 1831 85411 1865
rect 85713 1831 85747 1865
rect 86049 1831 86083 1865
rect 86385 1831 86419 1865
rect 86721 1831 86755 1865
rect 87057 1831 87091 1865
rect 87393 1831 87427 1865
rect 87729 1831 87763 1865
rect 88065 1831 88099 1865
rect 88401 1831 88435 1865
rect 88737 1831 88771 1865
rect 89073 1831 89107 1865
rect 89409 1831 89443 1865
rect 89745 1831 89779 1865
rect 90081 1831 90115 1865
rect 90417 1831 90451 1865
rect 90753 1831 90787 1865
rect 91089 1831 91123 1865
rect 91425 1831 91459 1865
rect 91761 1831 91795 1865
rect 92097 1831 92131 1865
rect 92433 1831 92467 1865
rect 92769 1831 92803 1865
rect 93105 1831 93139 1865
rect 93441 1831 93475 1865
rect 93777 1831 93811 1865
rect 94113 1831 94147 1865
rect 94449 1831 94483 1865
rect 94785 1831 94819 1865
rect 95121 1831 95155 1865
rect 95457 1831 95491 1865
rect 95793 1831 95827 1865
rect 96129 1831 96163 1865
rect 96465 1831 96499 1865
rect 96801 1831 96835 1865
rect 97137 1831 97171 1865
rect 97473 1831 97507 1865
rect 97809 1831 97843 1865
rect 98145 1831 98179 1865
rect 98481 1831 98515 1865
rect 98817 1831 98851 1865
rect 99153 1831 99187 1865
rect 99489 1831 99523 1865
rect 99825 1831 99859 1865
rect 100161 1831 100195 1865
rect 100497 1831 100531 1865
rect 100833 1831 100867 1865
rect 101169 1831 101203 1865
rect 101505 1831 101539 1865
rect 101841 1831 101875 1865
rect 102177 1831 102211 1865
rect 102513 1831 102547 1865
rect 102849 1831 102883 1865
rect 103185 1831 103219 1865
rect 103521 1831 103555 1865
rect 103857 1831 103891 1865
rect 104193 1831 104227 1865
rect 104529 1831 104563 1865
rect 104865 1831 104899 1865
rect 105201 1831 105235 1865
rect 105537 1831 105571 1865
rect 105873 1831 105907 1865
rect 106209 1831 106243 1865
rect 106545 1831 106579 1865
rect 106881 1831 106915 1865
rect 107217 1831 107251 1865
rect 107553 1831 107587 1865
rect 107889 1831 107923 1865
rect 108225 1831 108259 1865
rect 108561 1831 108595 1865
rect 108897 1831 108931 1865
rect 109233 1831 109267 1865
rect 109569 1831 109603 1865
rect 109905 1831 109939 1865
rect 110241 1831 110275 1865
rect 110577 1831 110611 1865
rect 110913 1831 110947 1865
rect 111249 1831 111283 1865
rect 111585 1831 111619 1865
rect 111921 1831 111955 1865
rect 112257 1831 112291 1865
rect 112593 1831 112627 1865
rect 112929 1831 112963 1865
rect 113265 1831 113299 1865
rect 113601 1831 113635 1865
rect 113937 1831 113971 1865
rect 114273 1831 114307 1865
rect 114609 1831 114643 1865
rect 114945 1831 114979 1865
rect 115281 1831 115315 1865
rect 115617 1831 115651 1865
rect 115953 1831 115987 1865
rect 116289 1831 116323 1865
rect 116625 1831 116659 1865
rect 116961 1831 116995 1865
rect 117297 1831 117331 1865
rect 117633 1831 117667 1865
rect 117969 1831 118003 1865
rect 118305 1831 118339 1865
rect 118641 1831 118675 1865
rect 118977 1831 119011 1865
rect 119313 1831 119347 1865
rect 119649 1831 119683 1865
rect 119985 1831 120019 1865
rect 120321 1831 120355 1865
rect 120657 1831 120691 1865
rect 120993 1831 121027 1865
rect 121329 1831 121363 1865
rect 121665 1831 121699 1865
rect 122001 1831 122035 1865
rect 122337 1831 122371 1865
rect 122673 1831 122707 1865
rect 123009 1831 123043 1865
rect 123345 1831 123379 1865
rect 123681 1831 123715 1865
rect 124017 1831 124051 1865
rect 124353 1831 124387 1865
rect 124689 1831 124723 1865
rect 125025 1831 125059 1865
rect 125361 1831 125395 1865
rect 125697 1831 125731 1865
rect 126033 1831 126067 1865
rect 126369 1831 126403 1865
rect 126705 1831 126739 1865
rect 127041 1831 127075 1865
rect 127377 1831 127411 1865
rect 127713 1831 127747 1865
rect 128049 1831 128083 1865
rect 128385 1831 128419 1865
rect 128721 1831 128755 1865
rect 129057 1831 129091 1865
rect 129393 1831 129427 1865
rect 129729 1831 129763 1865
rect 130065 1831 130099 1865
rect 130401 1831 130435 1865
rect 130737 1831 130771 1865
rect 131073 1831 131107 1865
rect 131409 1831 131443 1865
rect 131745 1831 131779 1865
rect 132081 1831 132115 1865
rect 132417 1831 132451 1865
rect 132753 1831 132787 1865
rect 133089 1831 133123 1865
rect 133425 1831 133459 1865
rect 133761 1831 133795 1865
rect 134097 1831 134131 1865
rect 134433 1831 134467 1865
rect 134769 1831 134803 1865
rect 135105 1831 135139 1865
rect 135441 1831 135475 1865
rect 135777 1831 135811 1865
rect 136113 1831 136147 1865
rect 136449 1831 136483 1865
rect 136785 1831 136819 1865
rect 137121 1831 137155 1865
rect 137457 1831 137491 1865
rect 137793 1831 137827 1865
rect 138129 1831 138163 1865
rect 138465 1831 138499 1865
rect 138801 1831 138835 1865
rect 139137 1831 139171 1865
rect 139473 1831 139507 1865
rect 139809 1831 139843 1865
rect 140145 1831 140179 1865
rect 140481 1831 140515 1865
rect 140817 1831 140851 1865
rect 141153 1831 141187 1865
rect 141489 1831 141523 1865
rect 141825 1831 141859 1865
rect 142161 1831 142195 1865
rect 142497 1831 142531 1865
rect 142833 1831 142867 1865
rect 143169 1831 143203 1865
rect 143505 1831 143539 1865
rect 143841 1831 143875 1865
rect 144177 1831 144211 1865
rect 144513 1831 144547 1865
rect 144849 1831 144883 1865
rect 145185 1831 145219 1865
rect 145521 1831 145555 1865
rect 145857 1831 145891 1865
rect 146193 1831 146227 1865
rect 146529 1831 146563 1865
rect 146865 1831 146899 1865
rect 147201 1831 147235 1865
rect 147537 1831 147571 1865
rect 147873 1831 147907 1865
rect 148209 1831 148243 1865
rect 148545 1831 148579 1865
rect 148881 1831 148915 1865
rect 149217 1831 149251 1865
rect 149553 1831 149587 1865
rect 149889 1831 149923 1865
rect 150225 1831 150259 1865
rect 150561 1831 150595 1865
rect 150897 1831 150931 1865
rect 151233 1831 151267 1865
rect 151569 1831 151603 1865
rect 151905 1831 151939 1865
rect 152241 1831 152275 1865
rect 152577 1831 152611 1865
rect 152913 1831 152947 1865
rect 153249 1831 153283 1865
rect 153585 1831 153619 1865
rect 153921 1831 153955 1865
rect 154257 1831 154291 1865
rect 154593 1831 154627 1865
rect 154929 1831 154963 1865
rect 155265 1831 155299 1865
rect 155601 1831 155635 1865
rect 155937 1831 155971 1865
rect 156273 1831 156307 1865
rect 156609 1831 156643 1865
rect 156945 1831 156979 1865
rect 157281 1831 157315 1865
rect 157617 1831 157651 1865
rect 157953 1831 157987 1865
rect 158289 1831 158323 1865
rect 158625 1831 158659 1865
rect 158961 1831 158995 1865
rect 159297 1831 159331 1865
rect 159633 1831 159667 1865
rect 159969 1831 160003 1865
rect 160305 1831 160339 1865
rect 160641 1831 160675 1865
rect 160977 1831 161011 1865
rect 161313 1831 161347 1865
rect 161649 1831 161683 1865
rect 161985 1831 162019 1865
rect 162321 1831 162355 1865
rect 162657 1831 162691 1865
rect 162993 1831 163027 1865
rect 163329 1831 163363 1865
rect 163665 1831 163699 1865
rect 164001 1831 164035 1865
rect 164337 1831 164371 1865
rect 164673 1831 164707 1865
rect 165009 1831 165043 1865
rect 165345 1831 165379 1865
rect 165681 1831 165715 1865
rect 166017 1831 166051 1865
rect 166353 1831 166387 1865
rect 166689 1831 166723 1865
rect 167025 1831 167059 1865
rect 167361 1831 167395 1865
rect 167697 1831 167731 1865
rect 168033 1831 168067 1865
rect 168369 1831 168403 1865
rect 168705 1831 168739 1865
rect 169041 1831 169075 1865
rect 169377 1831 169411 1865
rect 169713 1831 169747 1865
rect 170049 1831 170083 1865
rect 170385 1831 170419 1865
rect 170721 1831 170755 1865
rect 171057 1831 171091 1865
rect 171393 1831 171427 1865
rect 171729 1831 171763 1865
rect 172065 1831 172099 1865
rect 172401 1831 172435 1865
rect 172737 1831 172771 1865
rect 173073 1831 173107 1865
rect 173409 1831 173443 1865
rect 173745 1831 173779 1865
rect 174081 1831 174115 1865
rect 174417 1831 174451 1865
rect 174753 1831 174787 1865
rect 175089 1831 175123 1865
rect 175425 1831 175459 1865
rect 175761 1831 175795 1865
rect 176097 1831 176131 1865
rect 176433 1831 176467 1865
rect 176769 1831 176803 1865
rect 177105 1831 177139 1865
rect 177441 1831 177475 1865
rect 177777 1831 177811 1865
rect 178113 1831 178147 1865
rect 178449 1831 178483 1865
rect 178785 1831 178819 1865
rect 179121 1831 179155 1865
rect 179457 1831 179491 1865
rect 179793 1831 179827 1865
rect 180129 1831 180163 1865
rect 180465 1831 180499 1865
rect 180801 1831 180835 1865
rect 181137 1831 181171 1865
rect 181473 1831 181507 1865
rect 181809 1831 181843 1865
rect 182145 1831 182179 1865
rect 182481 1831 182515 1865
rect 182817 1831 182851 1865
rect 183153 1831 183187 1865
rect 183489 1831 183523 1865
rect 183825 1831 183859 1865
rect 184161 1831 184195 1865
rect 184497 1831 184531 1865
rect 184833 1831 184867 1865
rect 185169 1831 185203 1865
rect 185505 1831 185539 1865
rect 185841 1831 185875 1865
rect 186177 1831 186211 1865
rect 186513 1831 186547 1865
rect 186849 1831 186883 1865
rect 187185 1831 187219 1865
rect 187521 1831 187555 1865
rect 187857 1831 187891 1865
rect 188193 1831 188227 1865
rect 188529 1831 188563 1865
rect 188865 1831 188899 1865
rect 189201 1831 189235 1865
rect 189537 1831 189571 1865
rect 189873 1831 189907 1865
rect 190209 1831 190243 1865
rect 190545 1831 190579 1865
rect 190881 1831 190915 1865
rect 191217 1831 191251 1865
rect 191553 1831 191587 1865
rect 191889 1831 191923 1865
rect 192225 1831 192259 1865
rect 192561 1831 192595 1865
rect 192897 1831 192931 1865
rect 193233 1831 193267 1865
rect 193569 1831 193603 1865
rect 193905 1831 193939 1865
rect 194241 1831 194275 1865
rect 194577 1831 194611 1865
rect 194913 1831 194947 1865
rect 195249 1831 195283 1865
rect 195585 1831 195619 1865
rect 195921 1831 195955 1865
rect 196257 1831 196291 1865
rect 196593 1831 196627 1865
rect 196929 1831 196963 1865
rect 197265 1831 197299 1865
rect 197601 1831 197635 1865
rect 197937 1831 197971 1865
rect 198273 1831 198307 1865
rect 198609 1831 198643 1865
rect 198945 1831 198979 1865
rect 199281 1831 199315 1865
rect 199617 1831 199651 1865
rect 199953 1831 199987 1865
rect 200289 1831 200323 1865
rect 200625 1831 200659 1865
rect 200961 1831 200995 1865
rect 201297 1831 201331 1865
rect 201633 1831 201667 1865
rect 201969 1831 202003 1865
rect 202305 1831 202339 1865
rect 202641 1831 202675 1865
rect 202977 1831 203011 1865
rect 203313 1831 203347 1865
rect 203649 1831 203683 1865
rect 203985 1831 204019 1865
rect 204321 1831 204355 1865
rect 204657 1831 204691 1865
rect 204993 1831 205027 1865
rect 205329 1831 205363 1865
rect 205665 1831 205699 1865
rect 206001 1831 206035 1865
rect 206337 1831 206371 1865
rect 206673 1831 206707 1865
rect 207009 1831 207043 1865
rect 207345 1831 207379 1865
rect 207681 1831 207715 1865
rect 208017 1831 208051 1865
rect 208353 1831 208387 1865
rect 208689 1831 208723 1865
rect 209025 1831 209059 1865
rect 209361 1831 209395 1865
rect 209697 1831 209731 1865
rect 210033 1831 210067 1865
rect 210369 1831 210403 1865
rect 210705 1831 210739 1865
rect 211041 1831 211075 1865
rect 211377 1831 211411 1865
rect 211713 1831 211747 1865
rect 212049 1831 212083 1865
rect 212385 1831 212419 1865
rect 212721 1831 212755 1865
rect 213057 1831 213091 1865
rect 213393 1831 213427 1865
rect 213729 1831 213763 1865
rect 214065 1831 214099 1865
rect 214401 1831 214435 1865
rect 214737 1831 214771 1865
rect 215073 1831 215107 1865
rect 215409 1831 215443 1865
rect 215745 1831 215779 1865
rect 216081 1831 216115 1865
rect 216417 1831 216451 1865
<< locali >>
rect 2049 142361 2083 142377
rect 2049 142311 2083 142327
rect 2385 142361 2419 142377
rect 2385 142311 2419 142327
rect 2721 142361 2755 142377
rect 2721 142311 2755 142327
rect 3057 142361 3091 142377
rect 3057 142311 3091 142327
rect 3393 142361 3427 142377
rect 3393 142311 3427 142327
rect 3729 142361 3763 142377
rect 3729 142311 3763 142327
rect 4065 142361 4099 142377
rect 4065 142311 4099 142327
rect 4401 142361 4435 142377
rect 4401 142311 4435 142327
rect 4737 142361 4771 142377
rect 4737 142311 4771 142327
rect 5073 142361 5107 142377
rect 5073 142311 5107 142327
rect 5409 142361 5443 142377
rect 5409 142311 5443 142327
rect 5745 142361 5779 142377
rect 5745 142311 5779 142327
rect 6081 142361 6115 142377
rect 6081 142311 6115 142327
rect 6417 142361 6451 142377
rect 6417 142311 6451 142327
rect 6753 142361 6787 142377
rect 6753 142311 6787 142327
rect 7089 142361 7123 142377
rect 7089 142311 7123 142327
rect 7425 142361 7459 142377
rect 7425 142311 7459 142327
rect 7761 142361 7795 142377
rect 7761 142311 7795 142327
rect 8097 142361 8131 142377
rect 8097 142311 8131 142327
rect 8433 142361 8467 142377
rect 8433 142311 8467 142327
rect 8769 142361 8803 142377
rect 8769 142311 8803 142327
rect 9105 142361 9139 142377
rect 9105 142311 9139 142327
rect 9441 142361 9475 142377
rect 9441 142311 9475 142327
rect 9777 142361 9811 142377
rect 9777 142311 9811 142327
rect 10113 142361 10147 142377
rect 10113 142311 10147 142327
rect 10449 142361 10483 142377
rect 10449 142311 10483 142327
rect 10785 142361 10819 142377
rect 10785 142311 10819 142327
rect 11121 142361 11155 142377
rect 11121 142311 11155 142327
rect 11457 142361 11491 142377
rect 11457 142311 11491 142327
rect 11793 142361 11827 142377
rect 11793 142311 11827 142327
rect 12129 142361 12163 142377
rect 12129 142311 12163 142327
rect 12465 142361 12499 142377
rect 12465 142311 12499 142327
rect 12801 142361 12835 142377
rect 12801 142311 12835 142327
rect 13137 142361 13171 142377
rect 13137 142311 13171 142327
rect 13473 142361 13507 142377
rect 13473 142311 13507 142327
rect 13809 142361 13843 142377
rect 13809 142311 13843 142327
rect 14145 142361 14179 142377
rect 14145 142311 14179 142327
rect 14481 142361 14515 142377
rect 14481 142311 14515 142327
rect 14817 142361 14851 142377
rect 14817 142311 14851 142327
rect 15153 142361 15187 142377
rect 15153 142311 15187 142327
rect 15489 142361 15523 142377
rect 15489 142311 15523 142327
rect 15825 142361 15859 142377
rect 15825 142311 15859 142327
rect 16161 142361 16195 142377
rect 16161 142311 16195 142327
rect 16497 142361 16531 142377
rect 16497 142311 16531 142327
rect 16833 142361 16867 142377
rect 16833 142311 16867 142327
rect 17169 142361 17203 142377
rect 17169 142311 17203 142327
rect 17505 142361 17539 142377
rect 17505 142311 17539 142327
rect 17841 142361 17875 142377
rect 17841 142311 17875 142327
rect 18177 142361 18211 142377
rect 18177 142311 18211 142327
rect 18513 142361 18547 142377
rect 18513 142311 18547 142327
rect 18849 142361 18883 142377
rect 18849 142311 18883 142327
rect 19185 142361 19219 142377
rect 19185 142311 19219 142327
rect 19521 142361 19555 142377
rect 19521 142311 19555 142327
rect 19857 142361 19891 142377
rect 19857 142311 19891 142327
rect 20193 142361 20227 142377
rect 20193 142311 20227 142327
rect 20529 142361 20563 142377
rect 20529 142311 20563 142327
rect 20865 142361 20899 142377
rect 20865 142311 20899 142327
rect 21201 142361 21235 142377
rect 21201 142311 21235 142327
rect 21537 142361 21571 142377
rect 21537 142311 21571 142327
rect 21873 142361 21907 142377
rect 21873 142311 21907 142327
rect 22209 142361 22243 142377
rect 22209 142311 22243 142327
rect 22545 142361 22579 142377
rect 22545 142311 22579 142327
rect 22881 142361 22915 142377
rect 22881 142311 22915 142327
rect 23217 142361 23251 142377
rect 23217 142311 23251 142327
rect 23553 142361 23587 142377
rect 23553 142311 23587 142327
rect 23889 142361 23923 142377
rect 23889 142311 23923 142327
rect 24225 142361 24259 142377
rect 24225 142311 24259 142327
rect 24561 142361 24595 142377
rect 24561 142311 24595 142327
rect 24897 142361 24931 142377
rect 24897 142311 24931 142327
rect 25233 142361 25267 142377
rect 25233 142311 25267 142327
rect 25569 142361 25603 142377
rect 25569 142311 25603 142327
rect 25905 142361 25939 142377
rect 25905 142311 25939 142327
rect 26241 142361 26275 142377
rect 26241 142311 26275 142327
rect 26577 142361 26611 142377
rect 26577 142311 26611 142327
rect 26913 142361 26947 142377
rect 26913 142311 26947 142327
rect 27249 142361 27283 142377
rect 27249 142311 27283 142327
rect 27585 142361 27619 142377
rect 27585 142311 27619 142327
rect 27921 142361 27955 142377
rect 27921 142311 27955 142327
rect 28257 142361 28291 142377
rect 28257 142311 28291 142327
rect 28593 142361 28627 142377
rect 28593 142311 28627 142327
rect 28929 142361 28963 142377
rect 28929 142311 28963 142327
rect 29265 142361 29299 142377
rect 29265 142311 29299 142327
rect 29601 142361 29635 142377
rect 29601 142311 29635 142327
rect 29937 142361 29971 142377
rect 29937 142311 29971 142327
rect 30273 142361 30307 142377
rect 30273 142311 30307 142327
rect 30609 142361 30643 142377
rect 30609 142311 30643 142327
rect 30945 142361 30979 142377
rect 30945 142311 30979 142327
rect 31281 142361 31315 142377
rect 31281 142311 31315 142327
rect 31617 142361 31651 142377
rect 31617 142311 31651 142327
rect 31953 142361 31987 142377
rect 31953 142311 31987 142327
rect 32289 142361 32323 142377
rect 32289 142311 32323 142327
rect 32625 142361 32659 142377
rect 32625 142311 32659 142327
rect 32961 142361 32995 142377
rect 32961 142311 32995 142327
rect 33297 142361 33331 142377
rect 33297 142311 33331 142327
rect 33633 142361 33667 142377
rect 33633 142311 33667 142327
rect 33969 142361 34003 142377
rect 33969 142311 34003 142327
rect 34305 142361 34339 142377
rect 34305 142311 34339 142327
rect 34641 142361 34675 142377
rect 34641 142311 34675 142327
rect 34977 142361 35011 142377
rect 34977 142311 35011 142327
rect 35313 142361 35347 142377
rect 35313 142311 35347 142327
rect 35649 142361 35683 142377
rect 35649 142311 35683 142327
rect 35985 142361 36019 142377
rect 35985 142311 36019 142327
rect 36321 142361 36355 142377
rect 36321 142311 36355 142327
rect 36657 142361 36691 142377
rect 36657 142311 36691 142327
rect 36993 142361 37027 142377
rect 36993 142311 37027 142327
rect 37329 142361 37363 142377
rect 37329 142311 37363 142327
rect 37665 142361 37699 142377
rect 37665 142311 37699 142327
rect 38001 142361 38035 142377
rect 38001 142311 38035 142327
rect 38337 142361 38371 142377
rect 38337 142311 38371 142327
rect 38673 142361 38707 142377
rect 38673 142311 38707 142327
rect 39009 142361 39043 142377
rect 39009 142311 39043 142327
rect 39345 142361 39379 142377
rect 39345 142311 39379 142327
rect 39681 142361 39715 142377
rect 39681 142311 39715 142327
rect 40017 142361 40051 142377
rect 40017 142311 40051 142327
rect 40353 142361 40387 142377
rect 40353 142311 40387 142327
rect 40689 142361 40723 142377
rect 40689 142311 40723 142327
rect 41025 142361 41059 142377
rect 41025 142311 41059 142327
rect 41361 142361 41395 142377
rect 41361 142311 41395 142327
rect 41697 142361 41731 142377
rect 41697 142311 41731 142327
rect 42033 142361 42067 142377
rect 42033 142311 42067 142327
rect 42369 142361 42403 142377
rect 42369 142311 42403 142327
rect 42705 142361 42739 142377
rect 42705 142311 42739 142327
rect 43041 142361 43075 142377
rect 43041 142311 43075 142327
rect 43377 142361 43411 142377
rect 43377 142311 43411 142327
rect 43713 142361 43747 142377
rect 43713 142311 43747 142327
rect 44049 142361 44083 142377
rect 44049 142311 44083 142327
rect 44385 142361 44419 142377
rect 44385 142311 44419 142327
rect 44721 142361 44755 142377
rect 44721 142311 44755 142327
rect 45057 142361 45091 142377
rect 45057 142311 45091 142327
rect 45393 142361 45427 142377
rect 45393 142311 45427 142327
rect 45729 142361 45763 142377
rect 45729 142311 45763 142327
rect 46065 142361 46099 142377
rect 46065 142311 46099 142327
rect 46401 142361 46435 142377
rect 46401 142311 46435 142327
rect 46737 142361 46771 142377
rect 46737 142311 46771 142327
rect 47073 142361 47107 142377
rect 47073 142311 47107 142327
rect 47409 142361 47443 142377
rect 47409 142311 47443 142327
rect 47745 142361 47779 142377
rect 47745 142311 47779 142327
rect 48081 142361 48115 142377
rect 48081 142311 48115 142327
rect 48417 142361 48451 142377
rect 48417 142311 48451 142327
rect 48753 142361 48787 142377
rect 48753 142311 48787 142327
rect 49089 142361 49123 142377
rect 49089 142311 49123 142327
rect 49425 142361 49459 142377
rect 49425 142311 49459 142327
rect 49761 142361 49795 142377
rect 49761 142311 49795 142327
rect 50097 142361 50131 142377
rect 50097 142311 50131 142327
rect 50433 142361 50467 142377
rect 50433 142311 50467 142327
rect 50769 142361 50803 142377
rect 50769 142311 50803 142327
rect 51105 142361 51139 142377
rect 51105 142311 51139 142327
rect 51441 142361 51475 142377
rect 51441 142311 51475 142327
rect 51777 142361 51811 142377
rect 51777 142311 51811 142327
rect 52113 142361 52147 142377
rect 52113 142311 52147 142327
rect 52449 142361 52483 142377
rect 52449 142311 52483 142327
rect 52785 142361 52819 142377
rect 52785 142311 52819 142327
rect 53121 142361 53155 142377
rect 53121 142311 53155 142327
rect 53457 142361 53491 142377
rect 53457 142311 53491 142327
rect 53793 142361 53827 142377
rect 53793 142311 53827 142327
rect 54129 142361 54163 142377
rect 54129 142311 54163 142327
rect 54465 142361 54499 142377
rect 54465 142311 54499 142327
rect 54801 142361 54835 142377
rect 54801 142311 54835 142327
rect 55137 142361 55171 142377
rect 55137 142311 55171 142327
rect 55473 142361 55507 142377
rect 55473 142311 55507 142327
rect 55809 142361 55843 142377
rect 55809 142311 55843 142327
rect 56145 142361 56179 142377
rect 56145 142311 56179 142327
rect 56481 142361 56515 142377
rect 56481 142311 56515 142327
rect 56817 142361 56851 142377
rect 56817 142311 56851 142327
rect 57153 142361 57187 142377
rect 57153 142311 57187 142327
rect 57489 142361 57523 142377
rect 57489 142311 57523 142327
rect 57825 142361 57859 142377
rect 57825 142311 57859 142327
rect 58161 142361 58195 142377
rect 58161 142311 58195 142327
rect 58497 142361 58531 142377
rect 58497 142311 58531 142327
rect 58833 142361 58867 142377
rect 58833 142311 58867 142327
rect 59169 142361 59203 142377
rect 59169 142311 59203 142327
rect 59505 142361 59539 142377
rect 59505 142311 59539 142327
rect 59841 142361 59875 142377
rect 59841 142311 59875 142327
rect 60177 142361 60211 142377
rect 60177 142311 60211 142327
rect 60513 142361 60547 142377
rect 60513 142311 60547 142327
rect 60849 142361 60883 142377
rect 60849 142311 60883 142327
rect 61185 142361 61219 142377
rect 61185 142311 61219 142327
rect 61521 142361 61555 142377
rect 61521 142311 61555 142327
rect 61857 142361 61891 142377
rect 61857 142311 61891 142327
rect 62193 142361 62227 142377
rect 62193 142311 62227 142327
rect 62529 142361 62563 142377
rect 62529 142311 62563 142327
rect 62865 142361 62899 142377
rect 62865 142311 62899 142327
rect 63201 142361 63235 142377
rect 63201 142311 63235 142327
rect 63537 142361 63571 142377
rect 63537 142311 63571 142327
rect 63873 142361 63907 142377
rect 63873 142311 63907 142327
rect 64209 142361 64243 142377
rect 64209 142311 64243 142327
rect 64545 142361 64579 142377
rect 64545 142311 64579 142327
rect 64881 142361 64915 142377
rect 64881 142311 64915 142327
rect 65217 142361 65251 142377
rect 65217 142311 65251 142327
rect 65553 142361 65587 142377
rect 65553 142311 65587 142327
rect 65889 142361 65923 142377
rect 65889 142311 65923 142327
rect 66225 142361 66259 142377
rect 66225 142311 66259 142327
rect 66561 142361 66595 142377
rect 66561 142311 66595 142327
rect 66897 142361 66931 142377
rect 66897 142311 66931 142327
rect 67233 142361 67267 142377
rect 67233 142311 67267 142327
rect 67569 142361 67603 142377
rect 67569 142311 67603 142327
rect 67905 142361 67939 142377
rect 67905 142311 67939 142327
rect 68241 142361 68275 142377
rect 68241 142311 68275 142327
rect 68577 142361 68611 142377
rect 68577 142311 68611 142327
rect 68913 142361 68947 142377
rect 68913 142311 68947 142327
rect 69249 142361 69283 142377
rect 69249 142311 69283 142327
rect 69585 142361 69619 142377
rect 69585 142311 69619 142327
rect 69921 142361 69955 142377
rect 69921 142311 69955 142327
rect 70257 142361 70291 142377
rect 70257 142311 70291 142327
rect 70593 142361 70627 142377
rect 70593 142311 70627 142327
rect 70929 142361 70963 142377
rect 70929 142311 70963 142327
rect 71265 142361 71299 142377
rect 71265 142311 71299 142327
rect 71601 142361 71635 142377
rect 71601 142311 71635 142327
rect 71937 142361 71971 142377
rect 71937 142311 71971 142327
rect 72273 142361 72307 142377
rect 72273 142311 72307 142327
rect 72609 142361 72643 142377
rect 72609 142311 72643 142327
rect 72945 142361 72979 142377
rect 72945 142311 72979 142327
rect 73281 142361 73315 142377
rect 73281 142311 73315 142327
rect 73617 142361 73651 142377
rect 73617 142311 73651 142327
rect 73953 142361 73987 142377
rect 73953 142311 73987 142327
rect 74289 142361 74323 142377
rect 74289 142311 74323 142327
rect 74625 142361 74659 142377
rect 74625 142311 74659 142327
rect 74961 142361 74995 142377
rect 74961 142311 74995 142327
rect 75297 142361 75331 142377
rect 75297 142311 75331 142327
rect 75633 142361 75667 142377
rect 75633 142311 75667 142327
rect 75969 142361 76003 142377
rect 75969 142311 76003 142327
rect 76305 142361 76339 142377
rect 76305 142311 76339 142327
rect 76641 142361 76675 142377
rect 76641 142311 76675 142327
rect 76977 142361 77011 142377
rect 76977 142311 77011 142327
rect 77313 142361 77347 142377
rect 77313 142311 77347 142327
rect 77649 142361 77683 142377
rect 77649 142311 77683 142327
rect 77985 142361 78019 142377
rect 77985 142311 78019 142327
rect 78321 142361 78355 142377
rect 78321 142311 78355 142327
rect 78657 142361 78691 142377
rect 78657 142311 78691 142327
rect 78993 142361 79027 142377
rect 78993 142311 79027 142327
rect 79329 142361 79363 142377
rect 79329 142311 79363 142327
rect 79665 142361 79699 142377
rect 79665 142311 79699 142327
rect 80001 142361 80035 142377
rect 80001 142311 80035 142327
rect 80337 142361 80371 142377
rect 80337 142311 80371 142327
rect 80673 142361 80707 142377
rect 80673 142311 80707 142327
rect 81009 142361 81043 142377
rect 81009 142311 81043 142327
rect 81345 142361 81379 142377
rect 81345 142311 81379 142327
rect 81681 142361 81715 142377
rect 81681 142311 81715 142327
rect 82017 142361 82051 142377
rect 82017 142311 82051 142327
rect 82353 142361 82387 142377
rect 82353 142311 82387 142327
rect 82689 142361 82723 142377
rect 82689 142311 82723 142327
rect 83025 142361 83059 142377
rect 83025 142311 83059 142327
rect 83361 142361 83395 142377
rect 83361 142311 83395 142327
rect 83697 142361 83731 142377
rect 83697 142311 83731 142327
rect 84033 142361 84067 142377
rect 84033 142311 84067 142327
rect 84369 142361 84403 142377
rect 84369 142311 84403 142327
rect 84705 142361 84739 142377
rect 84705 142311 84739 142327
rect 85041 142361 85075 142377
rect 85041 142311 85075 142327
rect 85377 142361 85411 142377
rect 85377 142311 85411 142327
rect 85713 142361 85747 142377
rect 85713 142311 85747 142327
rect 86049 142361 86083 142377
rect 86049 142311 86083 142327
rect 86385 142361 86419 142377
rect 86385 142311 86419 142327
rect 86721 142361 86755 142377
rect 86721 142311 86755 142327
rect 87057 142361 87091 142377
rect 87057 142311 87091 142327
rect 87393 142361 87427 142377
rect 87393 142311 87427 142327
rect 87729 142361 87763 142377
rect 87729 142311 87763 142327
rect 88065 142361 88099 142377
rect 88065 142311 88099 142327
rect 88401 142361 88435 142377
rect 88401 142311 88435 142327
rect 88737 142361 88771 142377
rect 88737 142311 88771 142327
rect 89073 142361 89107 142377
rect 89073 142311 89107 142327
rect 89409 142361 89443 142377
rect 89409 142311 89443 142327
rect 89745 142361 89779 142377
rect 89745 142311 89779 142327
rect 90081 142361 90115 142377
rect 90081 142311 90115 142327
rect 90417 142361 90451 142377
rect 90417 142311 90451 142327
rect 90753 142361 90787 142377
rect 90753 142311 90787 142327
rect 91089 142361 91123 142377
rect 91089 142311 91123 142327
rect 91425 142361 91459 142377
rect 91425 142311 91459 142327
rect 91761 142361 91795 142377
rect 91761 142311 91795 142327
rect 92097 142361 92131 142377
rect 92097 142311 92131 142327
rect 92433 142361 92467 142377
rect 92433 142311 92467 142327
rect 92769 142361 92803 142377
rect 92769 142311 92803 142327
rect 93105 142361 93139 142377
rect 93105 142311 93139 142327
rect 93441 142361 93475 142377
rect 93441 142311 93475 142327
rect 93777 142361 93811 142377
rect 93777 142311 93811 142327
rect 94113 142361 94147 142377
rect 94113 142311 94147 142327
rect 94449 142361 94483 142377
rect 94449 142311 94483 142327
rect 94785 142361 94819 142377
rect 94785 142311 94819 142327
rect 95121 142361 95155 142377
rect 95121 142311 95155 142327
rect 95457 142361 95491 142377
rect 95457 142311 95491 142327
rect 95793 142361 95827 142377
rect 95793 142311 95827 142327
rect 96129 142361 96163 142377
rect 96129 142311 96163 142327
rect 96465 142361 96499 142377
rect 96465 142311 96499 142327
rect 96801 142361 96835 142377
rect 96801 142311 96835 142327
rect 97137 142361 97171 142377
rect 97137 142311 97171 142327
rect 97473 142361 97507 142377
rect 97473 142311 97507 142327
rect 97809 142361 97843 142377
rect 97809 142311 97843 142327
rect 98145 142361 98179 142377
rect 98145 142311 98179 142327
rect 98481 142361 98515 142377
rect 98481 142311 98515 142327
rect 98817 142361 98851 142377
rect 98817 142311 98851 142327
rect 99153 142361 99187 142377
rect 99153 142311 99187 142327
rect 99489 142361 99523 142377
rect 99489 142311 99523 142327
rect 99825 142361 99859 142377
rect 99825 142311 99859 142327
rect 100161 142361 100195 142377
rect 100161 142311 100195 142327
rect 100497 142361 100531 142377
rect 100497 142311 100531 142327
rect 100833 142361 100867 142377
rect 100833 142311 100867 142327
rect 101169 142361 101203 142377
rect 101169 142311 101203 142327
rect 101505 142361 101539 142377
rect 101505 142311 101539 142327
rect 101841 142361 101875 142377
rect 101841 142311 101875 142327
rect 102177 142361 102211 142377
rect 102177 142311 102211 142327
rect 102513 142361 102547 142377
rect 102513 142311 102547 142327
rect 102849 142361 102883 142377
rect 102849 142311 102883 142327
rect 103185 142361 103219 142377
rect 103185 142311 103219 142327
rect 103521 142361 103555 142377
rect 103521 142311 103555 142327
rect 103857 142361 103891 142377
rect 103857 142311 103891 142327
rect 104193 142361 104227 142377
rect 104193 142311 104227 142327
rect 104529 142361 104563 142377
rect 104529 142311 104563 142327
rect 104865 142361 104899 142377
rect 104865 142311 104899 142327
rect 105201 142361 105235 142377
rect 105201 142311 105235 142327
rect 105537 142361 105571 142377
rect 105537 142311 105571 142327
rect 105873 142361 105907 142377
rect 105873 142311 105907 142327
rect 106209 142361 106243 142377
rect 106209 142311 106243 142327
rect 106545 142361 106579 142377
rect 106545 142311 106579 142327
rect 106881 142361 106915 142377
rect 106881 142311 106915 142327
rect 107217 142361 107251 142377
rect 107217 142311 107251 142327
rect 107553 142361 107587 142377
rect 107553 142311 107587 142327
rect 107889 142361 107923 142377
rect 107889 142311 107923 142327
rect 108225 142361 108259 142377
rect 108225 142311 108259 142327
rect 108561 142361 108595 142377
rect 108561 142311 108595 142327
rect 108897 142361 108931 142377
rect 108897 142311 108931 142327
rect 109233 142361 109267 142377
rect 109233 142311 109267 142327
rect 109569 142361 109603 142377
rect 109569 142311 109603 142327
rect 109905 142361 109939 142377
rect 109905 142311 109939 142327
rect 110241 142361 110275 142377
rect 110241 142311 110275 142327
rect 110577 142361 110611 142377
rect 110577 142311 110611 142327
rect 110913 142361 110947 142377
rect 110913 142311 110947 142327
rect 111249 142361 111283 142377
rect 111249 142311 111283 142327
rect 111585 142361 111619 142377
rect 111585 142311 111619 142327
rect 111921 142361 111955 142377
rect 111921 142311 111955 142327
rect 112257 142361 112291 142377
rect 112257 142311 112291 142327
rect 112593 142361 112627 142377
rect 112593 142311 112627 142327
rect 112929 142361 112963 142377
rect 112929 142311 112963 142327
rect 113265 142361 113299 142377
rect 113265 142311 113299 142327
rect 113601 142361 113635 142377
rect 113601 142311 113635 142327
rect 113937 142361 113971 142377
rect 113937 142311 113971 142327
rect 114273 142361 114307 142377
rect 114273 142311 114307 142327
rect 114609 142361 114643 142377
rect 114609 142311 114643 142327
rect 114945 142361 114979 142377
rect 114945 142311 114979 142327
rect 115281 142361 115315 142377
rect 115281 142311 115315 142327
rect 115617 142361 115651 142377
rect 115617 142311 115651 142327
rect 115953 142361 115987 142377
rect 115953 142311 115987 142327
rect 116289 142361 116323 142377
rect 116289 142311 116323 142327
rect 116625 142361 116659 142377
rect 116625 142311 116659 142327
rect 116961 142361 116995 142377
rect 116961 142311 116995 142327
rect 117297 142361 117331 142377
rect 117297 142311 117331 142327
rect 117633 142361 117667 142377
rect 117633 142311 117667 142327
rect 117969 142361 118003 142377
rect 117969 142311 118003 142327
rect 118305 142361 118339 142377
rect 118305 142311 118339 142327
rect 118641 142361 118675 142377
rect 118641 142311 118675 142327
rect 118977 142361 119011 142377
rect 118977 142311 119011 142327
rect 119313 142361 119347 142377
rect 119313 142311 119347 142327
rect 119649 142361 119683 142377
rect 119649 142311 119683 142327
rect 119985 142361 120019 142377
rect 119985 142311 120019 142327
rect 120321 142361 120355 142377
rect 120321 142311 120355 142327
rect 120657 142361 120691 142377
rect 120657 142311 120691 142327
rect 120993 142361 121027 142377
rect 120993 142311 121027 142327
rect 121329 142361 121363 142377
rect 121329 142311 121363 142327
rect 121665 142361 121699 142377
rect 121665 142311 121699 142327
rect 122001 142361 122035 142377
rect 122001 142311 122035 142327
rect 122337 142361 122371 142377
rect 122337 142311 122371 142327
rect 122673 142361 122707 142377
rect 122673 142311 122707 142327
rect 123009 142361 123043 142377
rect 123009 142311 123043 142327
rect 123345 142361 123379 142377
rect 123345 142311 123379 142327
rect 123681 142361 123715 142377
rect 123681 142311 123715 142327
rect 124017 142361 124051 142377
rect 124017 142311 124051 142327
rect 124353 142361 124387 142377
rect 124353 142311 124387 142327
rect 124689 142361 124723 142377
rect 124689 142311 124723 142327
rect 125025 142361 125059 142377
rect 125025 142311 125059 142327
rect 125361 142361 125395 142377
rect 125361 142311 125395 142327
rect 125697 142361 125731 142377
rect 125697 142311 125731 142327
rect 126033 142361 126067 142377
rect 126033 142311 126067 142327
rect 126369 142361 126403 142377
rect 126369 142311 126403 142327
rect 126705 142361 126739 142377
rect 126705 142311 126739 142327
rect 127041 142361 127075 142377
rect 127041 142311 127075 142327
rect 127377 142361 127411 142377
rect 127377 142311 127411 142327
rect 127713 142361 127747 142377
rect 127713 142311 127747 142327
rect 128049 142361 128083 142377
rect 128049 142311 128083 142327
rect 128385 142361 128419 142377
rect 128385 142311 128419 142327
rect 128721 142361 128755 142377
rect 128721 142311 128755 142327
rect 129057 142361 129091 142377
rect 129057 142311 129091 142327
rect 129393 142361 129427 142377
rect 129393 142311 129427 142327
rect 129729 142361 129763 142377
rect 129729 142311 129763 142327
rect 130065 142361 130099 142377
rect 130065 142311 130099 142327
rect 130401 142361 130435 142377
rect 130401 142311 130435 142327
rect 130737 142361 130771 142377
rect 130737 142311 130771 142327
rect 131073 142361 131107 142377
rect 131073 142311 131107 142327
rect 131409 142361 131443 142377
rect 131409 142311 131443 142327
rect 131745 142361 131779 142377
rect 131745 142311 131779 142327
rect 132081 142361 132115 142377
rect 132081 142311 132115 142327
rect 132417 142361 132451 142377
rect 132417 142311 132451 142327
rect 132753 142361 132787 142377
rect 132753 142311 132787 142327
rect 133089 142361 133123 142377
rect 133089 142311 133123 142327
rect 133425 142361 133459 142377
rect 133425 142311 133459 142327
rect 133761 142361 133795 142377
rect 133761 142311 133795 142327
rect 134097 142361 134131 142377
rect 134097 142311 134131 142327
rect 134433 142361 134467 142377
rect 134433 142311 134467 142327
rect 134769 142361 134803 142377
rect 134769 142311 134803 142327
rect 135105 142361 135139 142377
rect 135105 142311 135139 142327
rect 135441 142361 135475 142377
rect 135441 142311 135475 142327
rect 135777 142361 135811 142377
rect 135777 142311 135811 142327
rect 136113 142361 136147 142377
rect 136113 142311 136147 142327
rect 136449 142361 136483 142377
rect 136449 142311 136483 142327
rect 136785 142361 136819 142377
rect 136785 142311 136819 142327
rect 137121 142361 137155 142377
rect 137121 142311 137155 142327
rect 137457 142361 137491 142377
rect 137457 142311 137491 142327
rect 137793 142361 137827 142377
rect 137793 142311 137827 142327
rect 138129 142361 138163 142377
rect 138129 142311 138163 142327
rect 138465 142361 138499 142377
rect 138465 142311 138499 142327
rect 138801 142361 138835 142377
rect 138801 142311 138835 142327
rect 139137 142361 139171 142377
rect 139137 142311 139171 142327
rect 139473 142361 139507 142377
rect 139473 142311 139507 142327
rect 139809 142361 139843 142377
rect 139809 142311 139843 142327
rect 140145 142361 140179 142377
rect 140145 142311 140179 142327
rect 140481 142361 140515 142377
rect 140481 142311 140515 142327
rect 140817 142361 140851 142377
rect 140817 142311 140851 142327
rect 141153 142361 141187 142377
rect 141153 142311 141187 142327
rect 141489 142361 141523 142377
rect 141489 142311 141523 142327
rect 141825 142361 141859 142377
rect 141825 142311 141859 142327
rect 142161 142361 142195 142377
rect 142161 142311 142195 142327
rect 142497 142361 142531 142377
rect 142497 142311 142531 142327
rect 142833 142361 142867 142377
rect 142833 142311 142867 142327
rect 143169 142361 143203 142377
rect 143169 142311 143203 142327
rect 143505 142361 143539 142377
rect 143505 142311 143539 142327
rect 143841 142361 143875 142377
rect 143841 142311 143875 142327
rect 144177 142361 144211 142377
rect 144177 142311 144211 142327
rect 144513 142361 144547 142377
rect 144513 142311 144547 142327
rect 144849 142361 144883 142377
rect 144849 142311 144883 142327
rect 145185 142361 145219 142377
rect 145185 142311 145219 142327
rect 145521 142361 145555 142377
rect 145521 142311 145555 142327
rect 145857 142361 145891 142377
rect 145857 142311 145891 142327
rect 146193 142361 146227 142377
rect 146193 142311 146227 142327
rect 146529 142361 146563 142377
rect 146529 142311 146563 142327
rect 146865 142361 146899 142377
rect 146865 142311 146899 142327
rect 147201 142361 147235 142377
rect 147201 142311 147235 142327
rect 147537 142361 147571 142377
rect 147537 142311 147571 142327
rect 147873 142361 147907 142377
rect 147873 142311 147907 142327
rect 148209 142361 148243 142377
rect 148209 142311 148243 142327
rect 148545 142361 148579 142377
rect 148545 142311 148579 142327
rect 148881 142361 148915 142377
rect 148881 142311 148915 142327
rect 149217 142361 149251 142377
rect 149217 142311 149251 142327
rect 149553 142361 149587 142377
rect 149553 142311 149587 142327
rect 149889 142361 149923 142377
rect 149889 142311 149923 142327
rect 150225 142361 150259 142377
rect 150225 142311 150259 142327
rect 150561 142361 150595 142377
rect 150561 142311 150595 142327
rect 150897 142361 150931 142377
rect 150897 142311 150931 142327
rect 151233 142361 151267 142377
rect 151233 142311 151267 142327
rect 151569 142361 151603 142377
rect 151569 142311 151603 142327
rect 151905 142361 151939 142377
rect 151905 142311 151939 142327
rect 152241 142361 152275 142377
rect 152241 142311 152275 142327
rect 152577 142361 152611 142377
rect 152577 142311 152611 142327
rect 152913 142361 152947 142377
rect 152913 142311 152947 142327
rect 153249 142361 153283 142377
rect 153249 142311 153283 142327
rect 153585 142361 153619 142377
rect 153585 142311 153619 142327
rect 153921 142361 153955 142377
rect 153921 142311 153955 142327
rect 154257 142361 154291 142377
rect 154257 142311 154291 142327
rect 154593 142361 154627 142377
rect 154593 142311 154627 142327
rect 154929 142361 154963 142377
rect 154929 142311 154963 142327
rect 155265 142361 155299 142377
rect 155265 142311 155299 142327
rect 155601 142361 155635 142377
rect 155601 142311 155635 142327
rect 155937 142361 155971 142377
rect 155937 142311 155971 142327
rect 156273 142361 156307 142377
rect 156273 142311 156307 142327
rect 156609 142361 156643 142377
rect 156609 142311 156643 142327
rect 156945 142361 156979 142377
rect 156945 142311 156979 142327
rect 157281 142361 157315 142377
rect 157281 142311 157315 142327
rect 157617 142361 157651 142377
rect 157617 142311 157651 142327
rect 157953 142361 157987 142377
rect 157953 142311 157987 142327
rect 158289 142361 158323 142377
rect 158289 142311 158323 142327
rect 158625 142361 158659 142377
rect 158625 142311 158659 142327
rect 158961 142361 158995 142377
rect 158961 142311 158995 142327
rect 159297 142361 159331 142377
rect 159297 142311 159331 142327
rect 159633 142361 159667 142377
rect 159633 142311 159667 142327
rect 159969 142361 160003 142377
rect 159969 142311 160003 142327
rect 160305 142361 160339 142377
rect 160305 142311 160339 142327
rect 160641 142361 160675 142377
rect 160641 142311 160675 142327
rect 160977 142361 161011 142377
rect 160977 142311 161011 142327
rect 161313 142361 161347 142377
rect 161313 142311 161347 142327
rect 161649 142361 161683 142377
rect 161649 142311 161683 142327
rect 161985 142361 162019 142377
rect 161985 142311 162019 142327
rect 162321 142361 162355 142377
rect 162321 142311 162355 142327
rect 162657 142361 162691 142377
rect 162657 142311 162691 142327
rect 162993 142361 163027 142377
rect 162993 142311 163027 142327
rect 163329 142361 163363 142377
rect 163329 142311 163363 142327
rect 163665 142361 163699 142377
rect 163665 142311 163699 142327
rect 164001 142361 164035 142377
rect 164001 142311 164035 142327
rect 164337 142361 164371 142377
rect 164337 142311 164371 142327
rect 164673 142361 164707 142377
rect 164673 142311 164707 142327
rect 165009 142361 165043 142377
rect 165009 142311 165043 142327
rect 165345 142361 165379 142377
rect 165345 142311 165379 142327
rect 165681 142361 165715 142377
rect 165681 142311 165715 142327
rect 166017 142361 166051 142377
rect 166017 142311 166051 142327
rect 166353 142361 166387 142377
rect 166353 142311 166387 142327
rect 166689 142361 166723 142377
rect 166689 142311 166723 142327
rect 167025 142361 167059 142377
rect 167025 142311 167059 142327
rect 167361 142361 167395 142377
rect 167361 142311 167395 142327
rect 167697 142361 167731 142377
rect 167697 142311 167731 142327
rect 168033 142361 168067 142377
rect 168033 142311 168067 142327
rect 168369 142361 168403 142377
rect 168369 142311 168403 142327
rect 168705 142361 168739 142377
rect 168705 142311 168739 142327
rect 169041 142361 169075 142377
rect 169041 142311 169075 142327
rect 169377 142361 169411 142377
rect 169377 142311 169411 142327
rect 169713 142361 169747 142377
rect 169713 142311 169747 142327
rect 170049 142361 170083 142377
rect 170049 142311 170083 142327
rect 170385 142361 170419 142377
rect 170385 142311 170419 142327
rect 170721 142361 170755 142377
rect 170721 142311 170755 142327
rect 171057 142361 171091 142377
rect 171057 142311 171091 142327
rect 171393 142361 171427 142377
rect 171393 142311 171427 142327
rect 171729 142361 171763 142377
rect 171729 142311 171763 142327
rect 172065 142361 172099 142377
rect 172065 142311 172099 142327
rect 172401 142361 172435 142377
rect 172401 142311 172435 142327
rect 172737 142361 172771 142377
rect 172737 142311 172771 142327
rect 173073 142361 173107 142377
rect 173073 142311 173107 142327
rect 173409 142361 173443 142377
rect 173409 142311 173443 142327
rect 173745 142361 173779 142377
rect 173745 142311 173779 142327
rect 174081 142361 174115 142377
rect 174081 142311 174115 142327
rect 174417 142361 174451 142377
rect 174417 142311 174451 142327
rect 174753 142361 174787 142377
rect 174753 142311 174787 142327
rect 175089 142361 175123 142377
rect 175089 142311 175123 142327
rect 175425 142361 175459 142377
rect 175425 142311 175459 142327
rect 175761 142361 175795 142377
rect 175761 142311 175795 142327
rect 176097 142361 176131 142377
rect 176097 142311 176131 142327
rect 176433 142361 176467 142377
rect 176433 142311 176467 142327
rect 176769 142361 176803 142377
rect 176769 142311 176803 142327
rect 177105 142361 177139 142377
rect 177105 142311 177139 142327
rect 177441 142361 177475 142377
rect 177441 142311 177475 142327
rect 177777 142361 177811 142377
rect 177777 142311 177811 142327
rect 178113 142361 178147 142377
rect 178113 142311 178147 142327
rect 178449 142361 178483 142377
rect 178449 142311 178483 142327
rect 178785 142361 178819 142377
rect 178785 142311 178819 142327
rect 179121 142361 179155 142377
rect 179121 142311 179155 142327
rect 179457 142361 179491 142377
rect 179457 142311 179491 142327
rect 179793 142361 179827 142377
rect 179793 142311 179827 142327
rect 180129 142361 180163 142377
rect 180129 142311 180163 142327
rect 180465 142361 180499 142377
rect 180465 142311 180499 142327
rect 180801 142361 180835 142377
rect 180801 142311 180835 142327
rect 181137 142361 181171 142377
rect 181137 142311 181171 142327
rect 181473 142361 181507 142377
rect 181473 142311 181507 142327
rect 181809 142361 181843 142377
rect 181809 142311 181843 142327
rect 182145 142361 182179 142377
rect 182145 142311 182179 142327
rect 182481 142361 182515 142377
rect 182481 142311 182515 142327
rect 182817 142361 182851 142377
rect 182817 142311 182851 142327
rect 183153 142361 183187 142377
rect 183153 142311 183187 142327
rect 183489 142361 183523 142377
rect 183489 142311 183523 142327
rect 183825 142361 183859 142377
rect 183825 142311 183859 142327
rect 184161 142361 184195 142377
rect 184161 142311 184195 142327
rect 184497 142361 184531 142377
rect 184497 142311 184531 142327
rect 184833 142361 184867 142377
rect 184833 142311 184867 142327
rect 185169 142361 185203 142377
rect 185169 142311 185203 142327
rect 185505 142361 185539 142377
rect 185505 142311 185539 142327
rect 185841 142361 185875 142377
rect 185841 142311 185875 142327
rect 186177 142361 186211 142377
rect 186177 142311 186211 142327
rect 186513 142361 186547 142377
rect 186513 142311 186547 142327
rect 186849 142361 186883 142377
rect 186849 142311 186883 142327
rect 187185 142361 187219 142377
rect 187185 142311 187219 142327
rect 187521 142361 187555 142377
rect 187521 142311 187555 142327
rect 187857 142361 187891 142377
rect 187857 142311 187891 142327
rect 188193 142361 188227 142377
rect 188193 142311 188227 142327
rect 188529 142361 188563 142377
rect 188529 142311 188563 142327
rect 188865 142361 188899 142377
rect 188865 142311 188899 142327
rect 189201 142361 189235 142377
rect 189201 142311 189235 142327
rect 189537 142361 189571 142377
rect 189537 142311 189571 142327
rect 189873 142361 189907 142377
rect 189873 142311 189907 142327
rect 190209 142361 190243 142377
rect 190209 142311 190243 142327
rect 190545 142361 190579 142377
rect 190545 142311 190579 142327
rect 190881 142361 190915 142377
rect 190881 142311 190915 142327
rect 191217 142361 191251 142377
rect 191217 142311 191251 142327
rect 191553 142361 191587 142377
rect 191553 142311 191587 142327
rect 191889 142361 191923 142377
rect 191889 142311 191923 142327
rect 192225 142361 192259 142377
rect 192225 142311 192259 142327
rect 192561 142361 192595 142377
rect 192561 142311 192595 142327
rect 192897 142361 192931 142377
rect 192897 142311 192931 142327
rect 193233 142361 193267 142377
rect 193233 142311 193267 142327
rect 193569 142361 193603 142377
rect 193569 142311 193603 142327
rect 193905 142361 193939 142377
rect 193905 142311 193939 142327
rect 194241 142361 194275 142377
rect 194241 142311 194275 142327
rect 194577 142361 194611 142377
rect 194577 142311 194611 142327
rect 194913 142361 194947 142377
rect 194913 142311 194947 142327
rect 195249 142361 195283 142377
rect 195249 142311 195283 142327
rect 195585 142361 195619 142377
rect 195585 142311 195619 142327
rect 195921 142361 195955 142377
rect 195921 142311 195955 142327
rect 196257 142361 196291 142377
rect 196257 142311 196291 142327
rect 196593 142361 196627 142377
rect 196593 142311 196627 142327
rect 196929 142361 196963 142377
rect 196929 142311 196963 142327
rect 197265 142361 197299 142377
rect 197265 142311 197299 142327
rect 197601 142361 197635 142377
rect 197601 142311 197635 142327
rect 197937 142361 197971 142377
rect 197937 142311 197971 142327
rect 198273 142361 198307 142377
rect 198273 142311 198307 142327
rect 198609 142361 198643 142377
rect 198609 142311 198643 142327
rect 198945 142361 198979 142377
rect 198945 142311 198979 142327
rect 199281 142361 199315 142377
rect 199281 142311 199315 142327
rect 199617 142361 199651 142377
rect 199617 142311 199651 142327
rect 199953 142361 199987 142377
rect 199953 142311 199987 142327
rect 200289 142361 200323 142377
rect 200289 142311 200323 142327
rect 200625 142361 200659 142377
rect 200625 142311 200659 142327
rect 200961 142361 200995 142377
rect 200961 142311 200995 142327
rect 201297 142361 201331 142377
rect 201297 142311 201331 142327
rect 201633 142361 201667 142377
rect 201633 142311 201667 142327
rect 201969 142361 202003 142377
rect 201969 142311 202003 142327
rect 202305 142361 202339 142377
rect 202305 142311 202339 142327
rect 202641 142361 202675 142377
rect 202641 142311 202675 142327
rect 202977 142361 203011 142377
rect 202977 142311 203011 142327
rect 203313 142361 203347 142377
rect 203313 142311 203347 142327
rect 203649 142361 203683 142377
rect 203649 142311 203683 142327
rect 203985 142361 204019 142377
rect 203985 142311 204019 142327
rect 204321 142361 204355 142377
rect 204321 142311 204355 142327
rect 204657 142361 204691 142377
rect 204657 142311 204691 142327
rect 204993 142361 205027 142377
rect 204993 142311 205027 142327
rect 205329 142361 205363 142377
rect 205329 142311 205363 142327
rect 205665 142361 205699 142377
rect 205665 142311 205699 142327
rect 206001 142361 206035 142377
rect 206001 142311 206035 142327
rect 206337 142361 206371 142377
rect 206337 142311 206371 142327
rect 206673 142361 206707 142377
rect 206673 142311 206707 142327
rect 207009 142361 207043 142377
rect 207009 142311 207043 142327
rect 207345 142361 207379 142377
rect 207345 142311 207379 142327
rect 207681 142361 207715 142377
rect 207681 142311 207715 142327
rect 208017 142361 208051 142377
rect 208017 142311 208051 142327
rect 208353 142361 208387 142377
rect 208353 142311 208387 142327
rect 208689 142361 208723 142377
rect 208689 142311 208723 142327
rect 209025 142361 209059 142377
rect 209025 142311 209059 142327
rect 209361 142361 209395 142377
rect 209361 142311 209395 142327
rect 209697 142361 209731 142377
rect 209697 142311 209731 142327
rect 210033 142361 210067 142377
rect 210033 142311 210067 142327
rect 210369 142361 210403 142377
rect 210369 142311 210403 142327
rect 210705 142361 210739 142377
rect 210705 142311 210739 142327
rect 211041 142361 211075 142377
rect 211041 142311 211075 142327
rect 211377 142361 211411 142377
rect 211377 142311 211411 142327
rect 211713 142361 211747 142377
rect 211713 142311 211747 142327
rect 212049 142361 212083 142377
rect 212049 142311 212083 142327
rect 212385 142361 212419 142377
rect 212385 142311 212419 142327
rect 212721 142361 212755 142377
rect 212721 142311 212755 142327
rect 213057 142361 213091 142377
rect 213057 142311 213091 142327
rect 213393 142361 213427 142377
rect 213393 142311 213427 142327
rect 213729 142361 213763 142377
rect 213729 142311 213763 142327
rect 214065 142361 214099 142377
rect 214065 142311 214099 142327
rect 214401 142361 214435 142377
rect 214401 142311 214435 142327
rect 214737 142361 214771 142377
rect 214737 142311 214771 142327
rect 215073 142361 215107 142377
rect 215073 142311 215107 142327
rect 215409 142361 215443 142377
rect 215409 142311 215443 142327
rect 215745 142361 215779 142377
rect 215745 142311 215779 142327
rect 216081 142361 216115 142377
rect 216081 142311 216115 142327
rect 216417 142361 216451 142377
rect 216417 142311 216451 142327
rect 1713 141977 1747 141993
rect 1713 141927 1747 141943
rect 216919 141977 216953 141993
rect 216919 141927 216953 141943
rect 1713 141641 1747 141657
rect 1713 141591 1747 141607
rect 216919 141641 216953 141657
rect 216919 141591 216953 141607
rect 1713 141305 1747 141321
rect 1713 141255 1747 141271
rect 216919 141305 216953 141321
rect 216919 141255 216953 141271
rect 1713 140969 1747 140985
rect 1713 140919 1747 140935
rect 216919 140969 216953 140985
rect 216919 140919 216953 140935
rect 1713 140633 1747 140649
rect 1713 140583 1747 140599
rect 216919 140633 216953 140649
rect 216919 140583 216953 140599
rect 1713 140297 1747 140313
rect 1713 140247 1747 140263
rect 216919 140297 216953 140313
rect 216919 140247 216953 140263
rect 1713 139961 1747 139977
rect 1713 139911 1747 139927
rect 216919 139961 216953 139977
rect 216919 139911 216953 139927
rect 1713 139625 1747 139641
rect 1713 139575 1747 139591
rect 216919 139625 216953 139641
rect 216919 139575 216953 139591
rect 1713 139289 1747 139305
rect 1713 139239 1747 139255
rect 216919 139289 216953 139305
rect 216919 139239 216953 139255
rect 1713 138953 1747 138969
rect 1713 138903 1747 138919
rect 216919 138953 216953 138969
rect 216919 138903 216953 138919
rect 1713 138617 1747 138633
rect 1713 138567 1747 138583
rect 216919 138617 216953 138633
rect 216919 138567 216953 138583
rect 1713 138281 1747 138297
rect 1713 138231 1747 138247
rect 216919 138281 216953 138297
rect 216919 138231 216953 138247
rect 1713 137945 1747 137961
rect 1713 137895 1747 137911
rect 216919 137945 216953 137961
rect 216919 137895 216953 137911
rect 1713 137609 1747 137625
rect 1713 137559 1747 137575
rect 216919 137609 216953 137625
rect 216919 137559 216953 137575
rect 1713 137273 1747 137289
rect 1713 137223 1747 137239
rect 216919 137273 216953 137289
rect 216919 137223 216953 137239
rect 1713 136937 1747 136953
rect 1713 136887 1747 136903
rect 216919 136937 216953 136953
rect 216919 136887 216953 136903
rect 1713 136601 1747 136617
rect 1713 136551 1747 136567
rect 216919 136601 216953 136617
rect 216919 136551 216953 136567
rect 1713 136265 1747 136281
rect 1713 136215 1747 136231
rect 216919 136265 216953 136281
rect 216919 136215 216953 136231
rect 1713 135929 1747 135945
rect 1713 135879 1747 135895
rect 216919 135929 216953 135945
rect 216919 135879 216953 135895
rect 1713 135593 1747 135609
rect 1713 135543 1747 135559
rect 216919 135593 216953 135609
rect 216919 135543 216953 135559
rect 1713 135257 1747 135273
rect 1713 135207 1747 135223
rect 216919 135257 216953 135273
rect 216919 135207 216953 135223
rect 1713 134921 1747 134937
rect 1713 134871 1747 134887
rect 216919 134921 216953 134937
rect 216919 134871 216953 134887
rect 1713 134585 1747 134601
rect 1713 134535 1747 134551
rect 216919 134585 216953 134601
rect 216919 134535 216953 134551
rect 1713 134249 1747 134265
rect 1713 134199 1747 134215
rect 216919 134249 216953 134265
rect 216919 134199 216953 134215
rect 1713 133913 1747 133929
rect 1713 133863 1747 133879
rect 216919 133913 216953 133929
rect 216919 133863 216953 133879
rect 1713 133577 1747 133593
rect 1713 133527 1747 133543
rect 216919 133577 216953 133593
rect 216919 133527 216953 133543
rect 1713 133241 1747 133257
rect 1713 133191 1747 133207
rect 216919 133241 216953 133257
rect 216919 133191 216953 133207
rect 1713 132905 1747 132921
rect 1713 132855 1747 132871
rect 216919 132905 216953 132921
rect 216919 132855 216953 132871
rect 1713 132569 1747 132585
rect 1713 132519 1747 132535
rect 216919 132569 216953 132585
rect 216919 132519 216953 132535
rect 1713 132233 1747 132249
rect 1713 132183 1747 132199
rect 216919 132233 216953 132249
rect 216919 132183 216953 132199
rect 1713 131897 1747 131913
rect 1713 131847 1747 131863
rect 216919 131897 216953 131913
rect 216919 131847 216953 131863
rect 1713 131561 1747 131577
rect 1713 131511 1747 131527
rect 216919 131561 216953 131577
rect 216919 131511 216953 131527
rect 1713 131225 1747 131241
rect 1713 131175 1747 131191
rect 216919 131225 216953 131241
rect 216919 131175 216953 131191
rect 1713 130889 1747 130905
rect 1713 130839 1747 130855
rect 216919 130889 216953 130905
rect 216919 130839 216953 130855
rect 1713 130553 1747 130569
rect 1713 130503 1747 130519
rect 216919 130553 216953 130569
rect 216919 130503 216953 130519
rect 1713 130217 1747 130233
rect 1713 130167 1747 130183
rect 216919 130217 216953 130233
rect 216919 130167 216953 130183
rect 1713 129881 1747 129897
rect 1713 129831 1747 129847
rect 216919 129881 216953 129897
rect 216919 129831 216953 129847
rect 1713 129545 1747 129561
rect 1713 129495 1747 129511
rect 216919 129545 216953 129561
rect 216919 129495 216953 129511
rect 1713 129209 1747 129225
rect 1713 129159 1747 129175
rect 216919 129209 216953 129225
rect 216919 129159 216953 129175
rect 1713 128873 1747 128889
rect 1713 128823 1747 128839
rect 216919 128873 216953 128889
rect 216919 128823 216953 128839
rect 1713 128537 1747 128553
rect 1713 128487 1747 128503
rect 216919 128537 216953 128553
rect 216919 128487 216953 128503
rect 1713 128201 1747 128217
rect 1713 128151 1747 128167
rect 216919 128201 216953 128217
rect 216919 128151 216953 128167
rect 1713 127865 1747 127881
rect 1713 127815 1747 127831
rect 216919 127865 216953 127881
rect 216919 127815 216953 127831
rect 1713 127529 1747 127545
rect 1713 127479 1747 127495
rect 216919 127529 216953 127545
rect 216919 127479 216953 127495
rect 1713 127193 1747 127209
rect 1713 127143 1747 127159
rect 216919 127193 216953 127209
rect 216919 127143 216953 127159
rect 1713 126857 1747 126873
rect 1713 126807 1747 126823
rect 216919 126857 216953 126873
rect 216919 126807 216953 126823
rect 1713 126521 1747 126537
rect 1713 126471 1747 126487
rect 216919 126521 216953 126537
rect 216919 126471 216953 126487
rect 1713 126185 1747 126201
rect 1713 126135 1747 126151
rect 216919 126185 216953 126201
rect 216919 126135 216953 126151
rect 1713 125849 1747 125865
rect 1713 125799 1747 125815
rect 216919 125849 216953 125865
rect 216919 125799 216953 125815
rect 1713 125513 1747 125529
rect 1713 125463 1747 125479
rect 216919 125513 216953 125529
rect 216919 125463 216953 125479
rect 1713 125177 1747 125193
rect 1713 125127 1747 125143
rect 216919 125177 216953 125193
rect 216919 125127 216953 125143
rect 1713 124841 1747 124857
rect 1713 124791 1747 124807
rect 216919 124841 216953 124857
rect 216919 124791 216953 124807
rect 1713 124505 1747 124521
rect 1713 124455 1747 124471
rect 216919 124505 216953 124521
rect 216919 124455 216953 124471
rect 1713 124169 1747 124185
rect 1713 124119 1747 124135
rect 216919 124169 216953 124185
rect 216919 124119 216953 124135
rect 1713 123833 1747 123849
rect 1713 123783 1747 123799
rect 216919 123833 216953 123849
rect 216919 123783 216953 123799
rect 1713 123497 1747 123513
rect 1713 123447 1747 123463
rect 216919 123497 216953 123513
rect 216919 123447 216953 123463
rect 1713 123161 1747 123177
rect 1713 123111 1747 123127
rect 216919 123161 216953 123177
rect 216919 123111 216953 123127
rect 1713 122825 1747 122841
rect 1713 122775 1747 122791
rect 216919 122825 216953 122841
rect 216919 122775 216953 122791
rect 1713 122489 1747 122505
rect 1713 122439 1747 122455
rect 216919 122489 216953 122505
rect 216919 122439 216953 122455
rect 1713 122153 1747 122169
rect 1713 122103 1747 122119
rect 216919 122153 216953 122169
rect 216919 122103 216953 122119
rect 1713 121817 1747 121833
rect 1713 121767 1747 121783
rect 216919 121817 216953 121833
rect 216919 121767 216953 121783
rect 1713 121481 1747 121497
rect 1713 121431 1747 121447
rect 216919 121481 216953 121497
rect 216919 121431 216953 121447
rect 1713 121145 1747 121161
rect 1713 121095 1747 121111
rect 216919 121145 216953 121161
rect 216919 121095 216953 121111
rect 1713 120809 1747 120825
rect 1713 120759 1747 120775
rect 216919 120809 216953 120825
rect 216919 120759 216953 120775
rect 1713 120473 1747 120489
rect 1713 120423 1747 120439
rect 216919 120473 216953 120489
rect 216919 120423 216953 120439
rect 1713 120137 1747 120153
rect 1713 120087 1747 120103
rect 216919 120137 216953 120153
rect 216919 120087 216953 120103
rect 1713 119801 1747 119817
rect 1713 119751 1747 119767
rect 216919 119801 216953 119817
rect 216919 119751 216953 119767
rect 1713 119465 1747 119481
rect 1713 119415 1747 119431
rect 216919 119465 216953 119481
rect 216919 119415 216953 119431
rect 1713 119129 1747 119145
rect 1713 119079 1747 119095
rect 216919 119129 216953 119145
rect 216919 119079 216953 119095
rect 1713 118793 1747 118809
rect 1713 118743 1747 118759
rect 216919 118793 216953 118809
rect 216919 118743 216953 118759
rect 1713 118457 1747 118473
rect 1713 118407 1747 118423
rect 216919 118457 216953 118473
rect 216919 118407 216953 118423
rect 1713 118121 1747 118137
rect 1713 118071 1747 118087
rect 216919 118121 216953 118137
rect 216919 118071 216953 118087
rect 1713 117785 1747 117801
rect 1713 117735 1747 117751
rect 216919 117785 216953 117801
rect 216919 117735 216953 117751
rect 1713 117449 1747 117465
rect 1713 117399 1747 117415
rect 216919 117449 216953 117465
rect 216919 117399 216953 117415
rect 1713 117113 1747 117129
rect 1713 117063 1747 117079
rect 216919 117113 216953 117129
rect 216919 117063 216953 117079
rect 1713 116777 1747 116793
rect 1713 116727 1747 116743
rect 216919 116777 216953 116793
rect 216919 116727 216953 116743
rect 1713 116441 1747 116457
rect 1713 116391 1747 116407
rect 216919 116441 216953 116457
rect 216919 116391 216953 116407
rect 1713 116105 1747 116121
rect 1713 116055 1747 116071
rect 216919 116105 216953 116121
rect 216919 116055 216953 116071
rect 1713 115769 1747 115785
rect 1713 115719 1747 115735
rect 216919 115769 216953 115785
rect 216919 115719 216953 115735
rect 1713 115433 1747 115449
rect 1713 115383 1747 115399
rect 216919 115433 216953 115449
rect 216919 115383 216953 115399
rect 1713 115097 1747 115113
rect 1713 115047 1747 115063
rect 216919 115097 216953 115113
rect 216919 115047 216953 115063
rect 1713 114761 1747 114777
rect 1713 114711 1747 114727
rect 216919 114761 216953 114777
rect 216919 114711 216953 114727
rect 1713 114425 1747 114441
rect 1713 114375 1747 114391
rect 216919 114425 216953 114441
rect 216919 114375 216953 114391
rect 1713 114089 1747 114105
rect 1713 114039 1747 114055
rect 216919 114089 216953 114105
rect 216919 114039 216953 114055
rect 1713 113753 1747 113769
rect 1713 113703 1747 113719
rect 216919 113753 216953 113769
rect 216919 113703 216953 113719
rect 1713 113417 1747 113433
rect 1713 113367 1747 113383
rect 216919 113417 216953 113433
rect 216919 113367 216953 113383
rect 1713 113081 1747 113097
rect 1713 113031 1747 113047
rect 216919 113081 216953 113097
rect 216919 113031 216953 113047
rect 1713 112745 1747 112761
rect 1713 112695 1747 112711
rect 216919 112745 216953 112761
rect 216919 112695 216953 112711
rect 1713 112409 1747 112425
rect 1713 112359 1747 112375
rect 216919 112409 216953 112425
rect 216919 112359 216953 112375
rect 1713 112073 1747 112089
rect 1713 112023 1747 112039
rect 216919 112073 216953 112089
rect 216919 112023 216953 112039
rect 1713 111737 1747 111753
rect 1713 111687 1747 111703
rect 216919 111737 216953 111753
rect 216919 111687 216953 111703
rect 1713 111401 1747 111417
rect 1713 111351 1747 111367
rect 216919 111401 216953 111417
rect 216919 111351 216953 111367
rect 1713 111065 1747 111081
rect 1713 111015 1747 111031
rect 216919 111065 216953 111081
rect 216919 111015 216953 111031
rect 1713 110729 1747 110745
rect 1713 110679 1747 110695
rect 216919 110729 216953 110745
rect 216919 110679 216953 110695
rect 1713 110393 1747 110409
rect 1713 110343 1747 110359
rect 216919 110393 216953 110409
rect 216919 110343 216953 110359
rect 1713 110057 1747 110073
rect 1713 110007 1747 110023
rect 216919 110057 216953 110073
rect 216919 110007 216953 110023
rect 1713 109721 1747 109737
rect 1713 109671 1747 109687
rect 216919 109721 216953 109737
rect 216919 109671 216953 109687
rect 1713 109385 1747 109401
rect 1713 109335 1747 109351
rect 216919 109385 216953 109401
rect 216919 109335 216953 109351
rect 1713 109049 1747 109065
rect 1713 108999 1747 109015
rect 216919 109049 216953 109065
rect 216919 108999 216953 109015
rect 1713 108713 1747 108729
rect 1713 108663 1747 108679
rect 216919 108713 216953 108729
rect 216919 108663 216953 108679
rect 1713 108377 1747 108393
rect 1713 108327 1747 108343
rect 216919 108377 216953 108393
rect 216919 108327 216953 108343
rect 1713 108041 1747 108057
rect 1713 107991 1747 108007
rect 216919 108041 216953 108057
rect 216919 107991 216953 108007
rect 1713 107705 1747 107721
rect 1713 107655 1747 107671
rect 216919 107705 216953 107721
rect 216919 107655 216953 107671
rect 1713 107369 1747 107385
rect 1713 107319 1747 107335
rect 216919 107369 216953 107385
rect 216919 107319 216953 107335
rect 1713 107033 1747 107049
rect 1713 106983 1747 106999
rect 216919 107033 216953 107049
rect 216919 106983 216953 106999
rect 1713 106697 1747 106713
rect 1713 106647 1747 106663
rect 216919 106697 216953 106713
rect 216919 106647 216953 106663
rect 1713 106361 1747 106377
rect 1713 106311 1747 106327
rect 216919 106361 216953 106377
rect 216919 106311 216953 106327
rect 1713 106025 1747 106041
rect 1713 105975 1747 105991
rect 216919 106025 216953 106041
rect 216919 105975 216953 105991
rect 1713 105689 1747 105705
rect 1713 105639 1747 105655
rect 216919 105689 216953 105705
rect 216919 105639 216953 105655
rect 1713 105353 1747 105369
rect 1713 105303 1747 105319
rect 216919 105353 216953 105369
rect 216919 105303 216953 105319
rect 1713 105017 1747 105033
rect 1713 104967 1747 104983
rect 216919 105017 216953 105033
rect 216919 104967 216953 104983
rect 1713 104681 1747 104697
rect 1713 104631 1747 104647
rect 216919 104681 216953 104697
rect 216919 104631 216953 104647
rect 1713 104345 1747 104361
rect 1713 104295 1747 104311
rect 216919 104345 216953 104361
rect 216919 104295 216953 104311
rect 1713 104009 1747 104025
rect 1713 103959 1747 103975
rect 216919 104009 216953 104025
rect 216919 103959 216953 103975
rect 1713 103673 1747 103689
rect 1713 103623 1747 103639
rect 216919 103673 216953 103689
rect 216919 103623 216953 103639
rect 1713 103337 1747 103353
rect 1713 103287 1747 103303
rect 216919 103337 216953 103353
rect 216919 103287 216953 103303
rect 1713 103001 1747 103017
rect 1713 102951 1747 102967
rect 216919 103001 216953 103017
rect 216919 102951 216953 102967
rect 1713 102665 1747 102681
rect 1713 102615 1747 102631
rect 216919 102665 216953 102681
rect 216919 102615 216953 102631
rect 1713 102329 1747 102345
rect 1713 102279 1747 102295
rect 216919 102329 216953 102345
rect 216919 102279 216953 102295
rect 1713 101993 1747 102009
rect 1713 101943 1747 101959
rect 216919 101993 216953 102009
rect 216919 101943 216953 101959
rect 1713 101657 1747 101673
rect 1713 101607 1747 101623
rect 216919 101657 216953 101673
rect 216919 101607 216953 101623
rect 1713 101321 1747 101337
rect 1713 101271 1747 101287
rect 216919 101321 216953 101337
rect 216919 101271 216953 101287
rect 1713 100985 1747 101001
rect 1713 100935 1747 100951
rect 216919 100985 216953 101001
rect 216919 100935 216953 100951
rect 1713 100649 1747 100665
rect 1713 100599 1747 100615
rect 216919 100649 216953 100665
rect 216919 100599 216953 100615
rect 1713 100313 1747 100329
rect 1713 100263 1747 100279
rect 216919 100313 216953 100329
rect 216919 100263 216953 100279
rect 1713 99977 1747 99993
rect 1713 99927 1747 99943
rect 216919 99977 216953 99993
rect 216919 99927 216953 99943
rect 1713 99641 1747 99657
rect 1713 99591 1747 99607
rect 216919 99641 216953 99657
rect 216919 99591 216953 99607
rect 1713 99305 1747 99321
rect 1713 99255 1747 99271
rect 216919 99305 216953 99321
rect 216919 99255 216953 99271
rect 1713 98969 1747 98985
rect 1713 98919 1747 98935
rect 216919 98969 216953 98985
rect 216919 98919 216953 98935
rect 1713 98633 1747 98649
rect 1713 98583 1747 98599
rect 216919 98633 216953 98649
rect 216919 98583 216953 98599
rect 1713 98297 1747 98313
rect 1713 98247 1747 98263
rect 216919 98297 216953 98313
rect 216919 98247 216953 98263
rect 1713 97961 1747 97977
rect 1713 97911 1747 97927
rect 216919 97961 216953 97977
rect 216919 97911 216953 97927
rect 1713 97625 1747 97641
rect 1713 97575 1747 97591
rect 216919 97625 216953 97641
rect 216919 97575 216953 97591
rect 1713 97289 1747 97305
rect 1713 97239 1747 97255
rect 216919 97289 216953 97305
rect 216919 97239 216953 97255
rect 1713 96953 1747 96969
rect 1713 96903 1747 96919
rect 216919 96953 216953 96969
rect 216919 96903 216953 96919
rect 1713 96617 1747 96633
rect 1713 96567 1747 96583
rect 216919 96617 216953 96633
rect 216919 96567 216953 96583
rect 1713 96281 1747 96297
rect 1713 96231 1747 96247
rect 216919 96281 216953 96297
rect 216919 96231 216953 96247
rect 1713 95945 1747 95961
rect 1713 95895 1747 95911
rect 216919 95945 216953 95961
rect 216919 95895 216953 95911
rect 1713 95609 1747 95625
rect 1713 95559 1747 95575
rect 216919 95609 216953 95625
rect 216919 95559 216953 95575
rect 1713 95273 1747 95289
rect 1713 95223 1747 95239
rect 216919 95273 216953 95289
rect 216919 95223 216953 95239
rect 1713 94937 1747 94953
rect 1713 94887 1747 94903
rect 216919 94937 216953 94953
rect 216919 94887 216953 94903
rect 1713 94601 1747 94617
rect 1713 94551 1747 94567
rect 216919 94601 216953 94617
rect 216919 94551 216953 94567
rect 1713 94265 1747 94281
rect 1713 94215 1747 94231
rect 216919 94265 216953 94281
rect 216919 94215 216953 94231
rect 1713 93929 1747 93945
rect 1713 93879 1747 93895
rect 216919 93929 216953 93945
rect 216919 93879 216953 93895
rect 1713 93593 1747 93609
rect 1713 93543 1747 93559
rect 216919 93593 216953 93609
rect 216919 93543 216953 93559
rect 1713 93257 1747 93273
rect 1713 93207 1747 93223
rect 216919 93257 216953 93273
rect 216919 93207 216953 93223
rect 1713 92921 1747 92937
rect 1713 92871 1747 92887
rect 216919 92921 216953 92937
rect 216919 92871 216953 92887
rect 1713 92585 1747 92601
rect 1713 92535 1747 92551
rect 216919 92585 216953 92601
rect 216919 92535 216953 92551
rect 1713 92249 1747 92265
rect 1713 92199 1747 92215
rect 216919 92249 216953 92265
rect 216919 92199 216953 92215
rect 1713 91913 1747 91929
rect 1713 91863 1747 91879
rect 216919 91913 216953 91929
rect 216919 91863 216953 91879
rect 1713 91577 1747 91593
rect 1713 91527 1747 91543
rect 216919 91577 216953 91593
rect 216919 91527 216953 91543
rect 1713 91241 1747 91257
rect 1713 91191 1747 91207
rect 216919 91241 216953 91257
rect 216919 91191 216953 91207
rect 1713 90905 1747 90921
rect 1713 90855 1747 90871
rect 216919 90905 216953 90921
rect 216919 90855 216953 90871
rect 1713 90569 1747 90585
rect 1713 90519 1747 90535
rect 216919 90569 216953 90585
rect 216919 90519 216953 90535
rect 1713 90233 1747 90249
rect 1713 90183 1747 90199
rect 216919 90233 216953 90249
rect 216919 90183 216953 90199
rect 1713 89897 1747 89913
rect 1713 89847 1747 89863
rect 216919 89897 216953 89913
rect 216919 89847 216953 89863
rect 1713 89561 1747 89577
rect 1713 89511 1747 89527
rect 216919 89561 216953 89577
rect 216919 89511 216953 89527
rect 1713 89225 1747 89241
rect 1713 89175 1747 89191
rect 216919 89225 216953 89241
rect 216919 89175 216953 89191
rect 1713 88889 1747 88905
rect 1713 88839 1747 88855
rect 216919 88889 216953 88905
rect 216919 88839 216953 88855
rect 1713 88553 1747 88569
rect 1713 88503 1747 88519
rect 216919 88553 216953 88569
rect 216919 88503 216953 88519
rect 1713 88217 1747 88233
rect 1713 88167 1747 88183
rect 216919 88217 216953 88233
rect 216919 88167 216953 88183
rect 1713 87881 1747 87897
rect 1713 87831 1747 87847
rect 216919 87881 216953 87897
rect 216919 87831 216953 87847
rect 1713 87545 1747 87561
rect 1713 87495 1747 87511
rect 216919 87545 216953 87561
rect 216919 87495 216953 87511
rect 1713 87209 1747 87225
rect 1713 87159 1747 87175
rect 216919 87209 216953 87225
rect 216919 87159 216953 87175
rect 1713 86873 1747 86889
rect 1713 86823 1747 86839
rect 216919 86873 216953 86889
rect 216919 86823 216953 86839
rect 1713 86537 1747 86553
rect 1713 86487 1747 86503
rect 216919 86537 216953 86553
rect 216919 86487 216953 86503
rect 1713 86201 1747 86217
rect 1713 86151 1747 86167
rect 216919 86201 216953 86217
rect 216919 86151 216953 86167
rect 1713 85865 1747 85881
rect 1713 85815 1747 85831
rect 216919 85865 216953 85881
rect 216919 85815 216953 85831
rect 1713 85529 1747 85545
rect 1713 85479 1747 85495
rect 216919 85529 216953 85545
rect 216919 85479 216953 85495
rect 1713 85193 1747 85209
rect 1713 85143 1747 85159
rect 216919 85193 216953 85209
rect 216919 85143 216953 85159
rect 1713 84857 1747 84873
rect 1713 84807 1747 84823
rect 216919 84857 216953 84873
rect 216919 84807 216953 84823
rect 1713 84521 1747 84537
rect 1713 84471 1747 84487
rect 216919 84521 216953 84537
rect 216919 84471 216953 84487
rect 1713 84185 1747 84201
rect 1713 84135 1747 84151
rect 216919 84185 216953 84201
rect 216919 84135 216953 84151
rect 1713 83849 1747 83865
rect 1713 83799 1747 83815
rect 216919 83849 216953 83865
rect 216919 83799 216953 83815
rect 1713 83513 1747 83529
rect 1713 83463 1747 83479
rect 216919 83513 216953 83529
rect 216919 83463 216953 83479
rect 1713 83177 1747 83193
rect 1713 83127 1747 83143
rect 216919 83177 216953 83193
rect 216919 83127 216953 83143
rect 1713 82841 1747 82857
rect 1713 82791 1747 82807
rect 216919 82841 216953 82857
rect 216919 82791 216953 82807
rect 1713 82505 1747 82521
rect 1713 82455 1747 82471
rect 216919 82505 216953 82521
rect 216919 82455 216953 82471
rect 1713 82169 1747 82185
rect 1713 82119 1747 82135
rect 216919 82169 216953 82185
rect 216919 82119 216953 82135
rect 1713 81833 1747 81849
rect 1713 81783 1747 81799
rect 216919 81833 216953 81849
rect 216919 81783 216953 81799
rect 1713 81497 1747 81513
rect 1713 81447 1747 81463
rect 216919 81497 216953 81513
rect 216919 81447 216953 81463
rect 1713 81161 1747 81177
rect 1713 81111 1747 81127
rect 216919 81161 216953 81177
rect 216919 81111 216953 81127
rect 1713 80825 1747 80841
rect 1713 80775 1747 80791
rect 216919 80825 216953 80841
rect 216919 80775 216953 80791
rect 1713 80489 1747 80505
rect 1713 80439 1747 80455
rect 216919 80489 216953 80505
rect 216919 80439 216953 80455
rect 1713 80153 1747 80169
rect 1713 80103 1747 80119
rect 216919 80153 216953 80169
rect 216919 80103 216953 80119
rect 1713 79817 1747 79833
rect 1713 79767 1747 79783
rect 216919 79817 216953 79833
rect 216919 79767 216953 79783
rect 1713 79481 1747 79497
rect 1713 79431 1747 79447
rect 216919 79481 216953 79497
rect 216919 79431 216953 79447
rect 1713 79145 1747 79161
rect 1713 79095 1747 79111
rect 216919 79145 216953 79161
rect 216919 79095 216953 79111
rect 1713 78809 1747 78825
rect 1713 78759 1747 78775
rect 216919 78809 216953 78825
rect 216919 78759 216953 78775
rect 1713 78473 1747 78489
rect 1713 78423 1747 78439
rect 216919 78473 216953 78489
rect 216919 78423 216953 78439
rect 1713 78137 1747 78153
rect 1713 78087 1747 78103
rect 216919 78137 216953 78153
rect 216919 78087 216953 78103
rect 1713 77801 1747 77817
rect 1713 77751 1747 77767
rect 216919 77801 216953 77817
rect 216919 77751 216953 77767
rect 1713 77465 1747 77481
rect 1713 77415 1747 77431
rect 216919 77465 216953 77481
rect 216919 77415 216953 77431
rect 1713 77129 1747 77145
rect 1713 77079 1747 77095
rect 216919 77129 216953 77145
rect 216919 77079 216953 77095
rect 1713 76793 1747 76809
rect 1713 76743 1747 76759
rect 216919 76793 216953 76809
rect 216919 76743 216953 76759
rect 1713 76457 1747 76473
rect 1713 76407 1747 76423
rect 216919 76457 216953 76473
rect 216919 76407 216953 76423
rect 1713 76121 1747 76137
rect 1713 76071 1747 76087
rect 216919 76121 216953 76137
rect 216919 76071 216953 76087
rect 1713 75785 1747 75801
rect 1713 75735 1747 75751
rect 216919 75785 216953 75801
rect 216919 75735 216953 75751
rect 1713 75449 1747 75465
rect 1713 75399 1747 75415
rect 216919 75449 216953 75465
rect 216919 75399 216953 75415
rect 1713 75113 1747 75129
rect 1713 75063 1747 75079
rect 216919 75113 216953 75129
rect 216919 75063 216953 75079
rect 1713 74777 1747 74793
rect 1713 74727 1747 74743
rect 216919 74777 216953 74793
rect 216919 74727 216953 74743
rect 1713 74441 1747 74457
rect 1713 74391 1747 74407
rect 216919 74441 216953 74457
rect 216919 74391 216953 74407
rect 1713 74105 1747 74121
rect 1713 74055 1747 74071
rect 216919 74105 216953 74121
rect 216919 74055 216953 74071
rect 1713 73769 1747 73785
rect 1713 73719 1747 73735
rect 216919 73769 216953 73785
rect 216919 73719 216953 73735
rect 1713 73433 1747 73449
rect 1713 73383 1747 73399
rect 216919 73433 216953 73449
rect 216919 73383 216953 73399
rect 1713 73097 1747 73113
rect 1713 73047 1747 73063
rect 216919 73097 216953 73113
rect 216919 73047 216953 73063
rect 1713 72761 1747 72777
rect 1713 72711 1747 72727
rect 216919 72761 216953 72777
rect 216919 72711 216953 72727
rect 1713 72425 1747 72441
rect 1713 72375 1747 72391
rect 216919 72425 216953 72441
rect 216919 72375 216953 72391
rect 1713 72089 1747 72105
rect 1713 72039 1747 72055
rect 216919 72089 216953 72105
rect 216919 72039 216953 72055
rect 1713 71753 1747 71769
rect 1713 71703 1747 71719
rect 216919 71753 216953 71769
rect 216919 71703 216953 71719
rect 1713 71417 1747 71433
rect 1713 71367 1747 71383
rect 216919 71417 216953 71433
rect 216919 71367 216953 71383
rect 1713 71081 1747 71097
rect 1713 71031 1747 71047
rect 216919 71081 216953 71097
rect 216919 71031 216953 71047
rect 1713 70745 1747 70761
rect 1713 70695 1747 70711
rect 216919 70745 216953 70761
rect 216919 70695 216953 70711
rect 1713 70409 1747 70425
rect 1713 70359 1747 70375
rect 216919 70409 216953 70425
rect 216919 70359 216953 70375
rect 1713 70073 1747 70089
rect 1713 70023 1747 70039
rect 216919 70073 216953 70089
rect 216919 70023 216953 70039
rect 1713 69737 1747 69753
rect 1713 69687 1747 69703
rect 216919 69737 216953 69753
rect 216919 69687 216953 69703
rect 1713 69401 1747 69417
rect 1713 69351 1747 69367
rect 216919 69401 216953 69417
rect 216919 69351 216953 69367
rect 1713 69065 1747 69081
rect 1713 69015 1747 69031
rect 216919 69065 216953 69081
rect 216919 69015 216953 69031
rect 1713 68729 1747 68745
rect 1713 68679 1747 68695
rect 216919 68729 216953 68745
rect 216919 68679 216953 68695
rect 1713 68393 1747 68409
rect 1713 68343 1747 68359
rect 216919 68393 216953 68409
rect 216919 68343 216953 68359
rect 1713 68057 1747 68073
rect 1713 68007 1747 68023
rect 216919 68057 216953 68073
rect 216919 68007 216953 68023
rect 1713 67721 1747 67737
rect 1713 67671 1747 67687
rect 216919 67721 216953 67737
rect 216919 67671 216953 67687
rect 1713 67385 1747 67401
rect 1713 67335 1747 67351
rect 216919 67385 216953 67401
rect 216919 67335 216953 67351
rect 1713 67049 1747 67065
rect 1713 66999 1747 67015
rect 216919 67049 216953 67065
rect 216919 66999 216953 67015
rect 1713 66713 1747 66729
rect 1713 66663 1747 66679
rect 216919 66713 216953 66729
rect 216919 66663 216953 66679
rect 1713 66377 1747 66393
rect 1713 66327 1747 66343
rect 216919 66377 216953 66393
rect 216919 66327 216953 66343
rect 1713 66041 1747 66057
rect 1713 65991 1747 66007
rect 216919 66041 216953 66057
rect 216919 65991 216953 66007
rect 1713 65705 1747 65721
rect 1713 65655 1747 65671
rect 216919 65705 216953 65721
rect 216919 65655 216953 65671
rect 1713 65369 1747 65385
rect 1713 65319 1747 65335
rect 216919 65369 216953 65385
rect 216919 65319 216953 65335
rect 1713 65033 1747 65049
rect 1713 64983 1747 64999
rect 216919 65033 216953 65049
rect 216919 64983 216953 64999
rect 1713 64697 1747 64713
rect 1713 64647 1747 64663
rect 216919 64697 216953 64713
rect 216919 64647 216953 64663
rect 1713 64361 1747 64377
rect 1713 64311 1747 64327
rect 216919 64361 216953 64377
rect 216919 64311 216953 64327
rect 1713 64025 1747 64041
rect 1713 63975 1747 63991
rect 216919 64025 216953 64041
rect 216919 63975 216953 63991
rect 1713 63689 1747 63705
rect 1713 63639 1747 63655
rect 216919 63689 216953 63705
rect 216919 63639 216953 63655
rect 1713 63353 1747 63369
rect 1713 63303 1747 63319
rect 216919 63353 216953 63369
rect 216919 63303 216953 63319
rect 1713 63017 1747 63033
rect 1713 62967 1747 62983
rect 216919 63017 216953 63033
rect 216919 62967 216953 62983
rect 1713 62681 1747 62697
rect 1713 62631 1747 62647
rect 216919 62681 216953 62697
rect 216919 62631 216953 62647
rect 1713 62345 1747 62361
rect 1713 62295 1747 62311
rect 216919 62345 216953 62361
rect 216919 62295 216953 62311
rect 1713 62009 1747 62025
rect 1713 61959 1747 61975
rect 216919 62009 216953 62025
rect 216919 61959 216953 61975
rect 1713 61673 1747 61689
rect 1713 61623 1747 61639
rect 216919 61673 216953 61689
rect 216919 61623 216953 61639
rect 1713 61337 1747 61353
rect 1713 61287 1747 61303
rect 216919 61337 216953 61353
rect 216919 61287 216953 61303
rect 1713 61001 1747 61017
rect 1713 60951 1747 60967
rect 216919 61001 216953 61017
rect 216919 60951 216953 60967
rect 1713 60665 1747 60681
rect 1713 60615 1747 60631
rect 216919 60665 216953 60681
rect 216919 60615 216953 60631
rect 1713 60329 1747 60345
rect 1713 60279 1747 60295
rect 216919 60329 216953 60345
rect 216919 60279 216953 60295
rect 1713 59993 1747 60009
rect 1713 59943 1747 59959
rect 216919 59993 216953 60009
rect 216919 59943 216953 59959
rect 1713 59657 1747 59673
rect 1713 59607 1747 59623
rect 216919 59657 216953 59673
rect 216919 59607 216953 59623
rect 1713 59321 1747 59337
rect 1713 59271 1747 59287
rect 216919 59321 216953 59337
rect 216919 59271 216953 59287
rect 1713 58985 1747 59001
rect 1713 58935 1747 58951
rect 216919 58985 216953 59001
rect 216919 58935 216953 58951
rect 1713 58649 1747 58665
rect 1713 58599 1747 58615
rect 216919 58649 216953 58665
rect 216919 58599 216953 58615
rect 1713 58313 1747 58329
rect 1713 58263 1747 58279
rect 216919 58313 216953 58329
rect 216919 58263 216953 58279
rect 1713 57977 1747 57993
rect 1713 57927 1747 57943
rect 216919 57977 216953 57993
rect 216919 57927 216953 57943
rect 1713 57641 1747 57657
rect 1713 57591 1747 57607
rect 216919 57641 216953 57657
rect 216919 57591 216953 57607
rect 1713 57305 1747 57321
rect 1713 57255 1747 57271
rect 216919 57305 216953 57321
rect 216919 57255 216953 57271
rect 1713 56969 1747 56985
rect 1713 56919 1747 56935
rect 216919 56969 216953 56985
rect 216919 56919 216953 56935
rect 1713 56633 1747 56649
rect 1713 56583 1747 56599
rect 216919 56633 216953 56649
rect 216919 56583 216953 56599
rect 1713 56297 1747 56313
rect 1713 56247 1747 56263
rect 216919 56297 216953 56313
rect 216919 56247 216953 56263
rect 1713 55961 1747 55977
rect 1713 55911 1747 55927
rect 216919 55961 216953 55977
rect 216919 55911 216953 55927
rect 1713 55625 1747 55641
rect 1713 55575 1747 55591
rect 216919 55625 216953 55641
rect 216919 55575 216953 55591
rect 1713 55289 1747 55305
rect 1713 55239 1747 55255
rect 216919 55289 216953 55305
rect 216919 55239 216953 55255
rect 1713 54953 1747 54969
rect 1713 54903 1747 54919
rect 216919 54953 216953 54969
rect 216919 54903 216953 54919
rect 1713 54617 1747 54633
rect 1713 54567 1747 54583
rect 216919 54617 216953 54633
rect 216919 54567 216953 54583
rect 1713 54281 1747 54297
rect 1713 54231 1747 54247
rect 216919 54281 216953 54297
rect 216919 54231 216953 54247
rect 1713 53945 1747 53961
rect 1713 53895 1747 53911
rect 216919 53945 216953 53961
rect 216919 53895 216953 53911
rect 1713 53609 1747 53625
rect 1713 53559 1747 53575
rect 216919 53609 216953 53625
rect 216919 53559 216953 53575
rect 1713 53273 1747 53289
rect 1713 53223 1747 53239
rect 216919 53273 216953 53289
rect 216919 53223 216953 53239
rect 1713 52937 1747 52953
rect 1713 52887 1747 52903
rect 216919 52937 216953 52953
rect 216919 52887 216953 52903
rect 1713 52601 1747 52617
rect 1713 52551 1747 52567
rect 216919 52601 216953 52617
rect 216919 52551 216953 52567
rect 1713 52265 1747 52281
rect 1713 52215 1747 52231
rect 216919 52265 216953 52281
rect 216919 52215 216953 52231
rect 1713 51929 1747 51945
rect 1713 51879 1747 51895
rect 216919 51929 216953 51945
rect 216919 51879 216953 51895
rect 1713 51593 1747 51609
rect 1713 51543 1747 51559
rect 216919 51593 216953 51609
rect 216919 51543 216953 51559
rect 1713 51257 1747 51273
rect 1713 51207 1747 51223
rect 216919 51257 216953 51273
rect 216919 51207 216953 51223
rect 1713 50921 1747 50937
rect 1713 50871 1747 50887
rect 216919 50921 216953 50937
rect 216919 50871 216953 50887
rect 1713 50585 1747 50601
rect 1713 50535 1747 50551
rect 216919 50585 216953 50601
rect 216919 50535 216953 50551
rect 1713 50249 1747 50265
rect 1713 50199 1747 50215
rect 216919 50249 216953 50265
rect 216919 50199 216953 50215
rect 1713 49913 1747 49929
rect 1713 49863 1747 49879
rect 216919 49913 216953 49929
rect 216919 49863 216953 49879
rect 1713 49577 1747 49593
rect 1713 49527 1747 49543
rect 216919 49577 216953 49593
rect 216919 49527 216953 49543
rect 1713 49241 1747 49257
rect 1713 49191 1747 49207
rect 216919 49241 216953 49257
rect 216919 49191 216953 49207
rect 1713 48905 1747 48921
rect 1713 48855 1747 48871
rect 216919 48905 216953 48921
rect 216919 48855 216953 48871
rect 1713 48569 1747 48585
rect 1713 48519 1747 48535
rect 216919 48569 216953 48585
rect 216919 48519 216953 48535
rect 1713 48233 1747 48249
rect 1713 48183 1747 48199
rect 216919 48233 216953 48249
rect 216919 48183 216953 48199
rect 1713 47897 1747 47913
rect 1713 47847 1747 47863
rect 216919 47897 216953 47913
rect 216919 47847 216953 47863
rect 1713 47561 1747 47577
rect 1713 47511 1747 47527
rect 216919 47561 216953 47577
rect 216919 47511 216953 47527
rect 1713 47225 1747 47241
rect 1713 47175 1747 47191
rect 216919 47225 216953 47241
rect 216919 47175 216953 47191
rect 1713 46889 1747 46905
rect 1713 46839 1747 46855
rect 216919 46889 216953 46905
rect 216919 46839 216953 46855
rect 1713 46553 1747 46569
rect 1713 46503 1747 46519
rect 216919 46553 216953 46569
rect 216919 46503 216953 46519
rect 1713 46217 1747 46233
rect 1713 46167 1747 46183
rect 216919 46217 216953 46233
rect 216919 46167 216953 46183
rect 1713 45881 1747 45897
rect 1713 45831 1747 45847
rect 216919 45881 216953 45897
rect 216919 45831 216953 45847
rect 1713 45545 1747 45561
rect 1713 45495 1747 45511
rect 216919 45545 216953 45561
rect 216919 45495 216953 45511
rect 1713 45209 1747 45225
rect 1713 45159 1747 45175
rect 216919 45209 216953 45225
rect 216919 45159 216953 45175
rect 1713 44873 1747 44889
rect 1713 44823 1747 44839
rect 216919 44873 216953 44889
rect 216919 44823 216953 44839
rect 1713 44537 1747 44553
rect 1713 44487 1747 44503
rect 216919 44537 216953 44553
rect 216919 44487 216953 44503
rect 1713 44201 1747 44217
rect 1713 44151 1747 44167
rect 216919 44201 216953 44217
rect 216919 44151 216953 44167
rect 1713 43865 1747 43881
rect 1713 43815 1747 43831
rect 216919 43865 216953 43881
rect 216919 43815 216953 43831
rect 1713 43529 1747 43545
rect 1713 43479 1747 43495
rect 216919 43529 216953 43545
rect 216919 43479 216953 43495
rect 1713 43193 1747 43209
rect 1713 43143 1747 43159
rect 216919 43193 216953 43209
rect 216919 43143 216953 43159
rect 1713 42857 1747 42873
rect 1713 42807 1747 42823
rect 216919 42857 216953 42873
rect 216919 42807 216953 42823
rect 1713 42521 1747 42537
rect 1713 42471 1747 42487
rect 216919 42521 216953 42537
rect 216919 42471 216953 42487
rect 1713 42185 1747 42201
rect 1713 42135 1747 42151
rect 216919 42185 216953 42201
rect 216919 42135 216953 42151
rect 1713 41849 1747 41865
rect 1713 41799 1747 41815
rect 216919 41849 216953 41865
rect 216919 41799 216953 41815
rect 1713 41513 1747 41529
rect 1713 41463 1747 41479
rect 216919 41513 216953 41529
rect 216919 41463 216953 41479
rect 1713 41177 1747 41193
rect 1713 41127 1747 41143
rect 216919 41177 216953 41193
rect 216919 41127 216953 41143
rect 1713 40841 1747 40857
rect 1713 40791 1747 40807
rect 216919 40841 216953 40857
rect 216919 40791 216953 40807
rect 1713 40505 1747 40521
rect 1713 40455 1747 40471
rect 216919 40505 216953 40521
rect 216919 40455 216953 40471
rect 1713 40169 1747 40185
rect 1713 40119 1747 40135
rect 216919 40169 216953 40185
rect 216919 40119 216953 40135
rect 1713 39833 1747 39849
rect 1713 39783 1747 39799
rect 216919 39833 216953 39849
rect 216919 39783 216953 39799
rect 1713 39497 1747 39513
rect 1713 39447 1747 39463
rect 216919 39497 216953 39513
rect 216919 39447 216953 39463
rect 1713 39161 1747 39177
rect 1713 39111 1747 39127
rect 216919 39161 216953 39177
rect 216919 39111 216953 39127
rect 1713 38825 1747 38841
rect 1713 38775 1747 38791
rect 216919 38825 216953 38841
rect 216919 38775 216953 38791
rect 1713 38489 1747 38505
rect 1713 38439 1747 38455
rect 216919 38489 216953 38505
rect 216919 38439 216953 38455
rect 1713 38153 1747 38169
rect 1713 38103 1747 38119
rect 216919 38153 216953 38169
rect 216919 38103 216953 38119
rect 1713 37817 1747 37833
rect 1713 37767 1747 37783
rect 216919 37817 216953 37833
rect 216919 37767 216953 37783
rect 1713 37481 1747 37497
rect 1713 37431 1747 37447
rect 216919 37481 216953 37497
rect 216919 37431 216953 37447
rect 1713 37145 1747 37161
rect 1713 37095 1747 37111
rect 216919 37145 216953 37161
rect 216919 37095 216953 37111
rect 1713 36809 1747 36825
rect 1713 36759 1747 36775
rect 216919 36809 216953 36825
rect 216919 36759 216953 36775
rect 1713 36473 1747 36489
rect 1713 36423 1747 36439
rect 216919 36473 216953 36489
rect 216919 36423 216953 36439
rect 1713 36137 1747 36153
rect 1713 36087 1747 36103
rect 216919 36137 216953 36153
rect 216919 36087 216953 36103
rect 1713 35801 1747 35817
rect 1713 35751 1747 35767
rect 216919 35801 216953 35817
rect 216919 35751 216953 35767
rect 1713 35465 1747 35481
rect 1713 35415 1747 35431
rect 216919 35465 216953 35481
rect 216919 35415 216953 35431
rect 1713 35129 1747 35145
rect 1713 35079 1747 35095
rect 216919 35129 216953 35145
rect 216919 35079 216953 35095
rect 1713 34793 1747 34809
rect 1713 34743 1747 34759
rect 216919 34793 216953 34809
rect 216919 34743 216953 34759
rect 1713 34457 1747 34473
rect 1713 34407 1747 34423
rect 216919 34457 216953 34473
rect 216919 34407 216953 34423
rect 1713 34121 1747 34137
rect 1713 34071 1747 34087
rect 216919 34121 216953 34137
rect 216919 34071 216953 34087
rect 1713 33785 1747 33801
rect 1713 33735 1747 33751
rect 216919 33785 216953 33801
rect 216919 33735 216953 33751
rect 1713 33449 1747 33465
rect 1713 33399 1747 33415
rect 216919 33449 216953 33465
rect 216919 33399 216953 33415
rect 1713 33113 1747 33129
rect 1713 33063 1747 33079
rect 216919 33113 216953 33129
rect 216919 33063 216953 33079
rect 1713 32777 1747 32793
rect 1713 32727 1747 32743
rect 216919 32777 216953 32793
rect 216919 32727 216953 32743
rect 1713 32441 1747 32457
rect 1713 32391 1747 32407
rect 216919 32441 216953 32457
rect 216919 32391 216953 32407
rect 1713 32105 1747 32121
rect 1713 32055 1747 32071
rect 216919 32105 216953 32121
rect 216919 32055 216953 32071
rect 1713 31769 1747 31785
rect 1713 31719 1747 31735
rect 216919 31769 216953 31785
rect 216919 31719 216953 31735
rect 1713 31433 1747 31449
rect 1713 31383 1747 31399
rect 216919 31433 216953 31449
rect 216919 31383 216953 31399
rect 1713 31097 1747 31113
rect 1713 31047 1747 31063
rect 216919 31097 216953 31113
rect 216919 31047 216953 31063
rect 1713 30761 1747 30777
rect 1713 30711 1747 30727
rect 216919 30761 216953 30777
rect 216919 30711 216953 30727
rect 1713 30425 1747 30441
rect 1713 30375 1747 30391
rect 216919 30425 216953 30441
rect 216919 30375 216953 30391
rect 1713 30089 1747 30105
rect 1713 30039 1747 30055
rect 216919 30089 216953 30105
rect 216919 30039 216953 30055
rect 1713 29753 1747 29769
rect 1713 29703 1747 29719
rect 216919 29753 216953 29769
rect 216919 29703 216953 29719
rect 1713 29417 1747 29433
rect 1713 29367 1747 29383
rect 216919 29417 216953 29433
rect 216919 29367 216953 29383
rect 1713 29081 1747 29097
rect 1713 29031 1747 29047
rect 216919 29081 216953 29097
rect 216919 29031 216953 29047
rect 1713 28745 1747 28761
rect 1713 28695 1747 28711
rect 216919 28745 216953 28761
rect 216919 28695 216953 28711
rect 1713 28409 1747 28425
rect 1713 28359 1747 28375
rect 216919 28409 216953 28425
rect 216919 28359 216953 28375
rect 1713 28073 1747 28089
rect 1713 28023 1747 28039
rect 216919 28073 216953 28089
rect 216919 28023 216953 28039
rect 1713 27737 1747 27753
rect 1713 27687 1747 27703
rect 216919 27737 216953 27753
rect 216919 27687 216953 27703
rect 1713 27401 1747 27417
rect 1713 27351 1747 27367
rect 216919 27401 216953 27417
rect 216919 27351 216953 27367
rect 1713 27065 1747 27081
rect 1713 27015 1747 27031
rect 216919 27065 216953 27081
rect 216919 27015 216953 27031
rect 1713 26729 1747 26745
rect 1713 26679 1747 26695
rect 216919 26729 216953 26745
rect 216919 26679 216953 26695
rect 1713 26393 1747 26409
rect 1713 26343 1747 26359
rect 216919 26393 216953 26409
rect 216919 26343 216953 26359
rect 1713 26057 1747 26073
rect 1713 26007 1747 26023
rect 216919 26057 216953 26073
rect 216919 26007 216953 26023
rect 1713 25721 1747 25737
rect 1713 25671 1747 25687
rect 216919 25721 216953 25737
rect 216919 25671 216953 25687
rect 1713 25385 1747 25401
rect 1713 25335 1747 25351
rect 216919 25385 216953 25401
rect 216919 25335 216953 25351
rect 1713 25049 1747 25065
rect 1713 24999 1747 25015
rect 216919 25049 216953 25065
rect 216919 24999 216953 25015
rect 1713 24713 1747 24729
rect 1713 24663 1747 24679
rect 216919 24713 216953 24729
rect 216919 24663 216953 24679
rect 1713 24377 1747 24393
rect 1713 24327 1747 24343
rect 216919 24377 216953 24393
rect 216919 24327 216953 24343
rect 1713 24041 1747 24057
rect 1713 23991 1747 24007
rect 216919 24041 216953 24057
rect 216919 23991 216953 24007
rect 1713 23705 1747 23721
rect 1713 23655 1747 23671
rect 216919 23705 216953 23721
rect 216919 23655 216953 23671
rect 1713 23369 1747 23385
rect 1713 23319 1747 23335
rect 216919 23369 216953 23385
rect 216919 23319 216953 23335
rect 1713 23033 1747 23049
rect 1713 22983 1747 22999
rect 216919 23033 216953 23049
rect 216919 22983 216953 22999
rect 1713 22697 1747 22713
rect 1713 22647 1747 22663
rect 216919 22697 216953 22713
rect 216919 22647 216953 22663
rect 1713 22361 1747 22377
rect 1713 22311 1747 22327
rect 216919 22361 216953 22377
rect 216919 22311 216953 22327
rect 1713 22025 1747 22041
rect 1713 21975 1747 21991
rect 216919 22025 216953 22041
rect 216919 21975 216953 21991
rect 1713 21689 1747 21705
rect 1713 21639 1747 21655
rect 216919 21689 216953 21705
rect 216919 21639 216953 21655
rect 1713 21353 1747 21369
rect 1713 21303 1747 21319
rect 216919 21353 216953 21369
rect 216919 21303 216953 21319
rect 1713 21017 1747 21033
rect 1713 20967 1747 20983
rect 216919 21017 216953 21033
rect 216919 20967 216953 20983
rect 1713 20681 1747 20697
rect 1713 20631 1747 20647
rect 216919 20681 216953 20697
rect 216919 20631 216953 20647
rect 1713 20345 1747 20361
rect 1713 20295 1747 20311
rect 216919 20345 216953 20361
rect 216919 20295 216953 20311
rect 1713 20009 1747 20025
rect 1713 19959 1747 19975
rect 216919 20009 216953 20025
rect 216919 19959 216953 19975
rect 1713 19673 1747 19689
rect 1713 19623 1747 19639
rect 216919 19673 216953 19689
rect 216919 19623 216953 19639
rect 1713 19337 1747 19353
rect 1713 19287 1747 19303
rect 216919 19337 216953 19353
rect 216919 19287 216953 19303
rect 1713 19001 1747 19017
rect 1713 18951 1747 18967
rect 216919 19001 216953 19017
rect 216919 18951 216953 18967
rect 1713 18665 1747 18681
rect 1713 18615 1747 18631
rect 216919 18665 216953 18681
rect 216919 18615 216953 18631
rect 1713 18329 1747 18345
rect 1713 18279 1747 18295
rect 216919 18329 216953 18345
rect 216919 18279 216953 18295
rect 1713 17993 1747 18009
rect 1713 17943 1747 17959
rect 216919 17993 216953 18009
rect 216919 17943 216953 17959
rect 1713 17657 1747 17673
rect 1713 17607 1747 17623
rect 216919 17657 216953 17673
rect 216919 17607 216953 17623
rect 1713 17321 1747 17337
rect 1713 17271 1747 17287
rect 216919 17321 216953 17337
rect 216919 17271 216953 17287
rect 1713 16985 1747 17001
rect 1713 16935 1747 16951
rect 216919 16985 216953 17001
rect 216919 16935 216953 16951
rect 1713 16649 1747 16665
rect 1713 16599 1747 16615
rect 216919 16649 216953 16665
rect 216919 16599 216953 16615
rect 1713 16313 1747 16329
rect 1713 16263 1747 16279
rect 216919 16313 216953 16329
rect 216919 16263 216953 16279
rect 1713 15977 1747 15993
rect 1713 15927 1747 15943
rect 216919 15977 216953 15993
rect 216919 15927 216953 15943
rect 1713 15641 1747 15657
rect 1713 15591 1747 15607
rect 216919 15641 216953 15657
rect 216919 15591 216953 15607
rect 1713 15305 1747 15321
rect 1713 15255 1747 15271
rect 216919 15305 216953 15321
rect 216919 15255 216953 15271
rect 1713 14969 1747 14985
rect 1713 14919 1747 14935
rect 216919 14969 216953 14985
rect 216919 14919 216953 14935
rect 1713 14633 1747 14649
rect 1713 14583 1747 14599
rect 216919 14633 216953 14649
rect 216919 14583 216953 14599
rect 1713 14297 1747 14313
rect 1713 14247 1747 14263
rect 216919 14297 216953 14313
rect 216919 14247 216953 14263
rect 1713 13961 1747 13977
rect 1713 13911 1747 13927
rect 216919 13961 216953 13977
rect 216919 13911 216953 13927
rect 1713 13625 1747 13641
rect 1713 13575 1747 13591
rect 216919 13625 216953 13641
rect 216919 13575 216953 13591
rect 1713 13289 1747 13305
rect 1713 13239 1747 13255
rect 216919 13289 216953 13305
rect 216919 13239 216953 13255
rect 1713 12953 1747 12969
rect 1713 12903 1747 12919
rect 216919 12953 216953 12969
rect 216919 12903 216953 12919
rect 1713 12617 1747 12633
rect 1713 12567 1747 12583
rect 216919 12617 216953 12633
rect 216919 12567 216953 12583
rect 1713 12281 1747 12297
rect 1713 12231 1747 12247
rect 216919 12281 216953 12297
rect 216919 12231 216953 12247
rect 1713 11945 1747 11961
rect 1713 11895 1747 11911
rect 216919 11945 216953 11961
rect 216919 11895 216953 11911
rect 1713 11609 1747 11625
rect 1713 11559 1747 11575
rect 216919 11609 216953 11625
rect 216919 11559 216953 11575
rect 1713 11273 1747 11289
rect 1713 11223 1747 11239
rect 216919 11273 216953 11289
rect 216919 11223 216953 11239
rect 1713 10937 1747 10953
rect 1713 10887 1747 10903
rect 216919 10937 216953 10953
rect 216919 10887 216953 10903
rect 1713 10601 1747 10617
rect 1713 10551 1747 10567
rect 216919 10601 216953 10617
rect 216919 10551 216953 10567
rect 1713 10265 1747 10281
rect 1713 10215 1747 10231
rect 216919 10265 216953 10281
rect 216919 10215 216953 10231
rect 1713 9929 1747 9945
rect 1713 9879 1747 9895
rect 216919 9929 216953 9945
rect 216919 9879 216953 9895
rect 1713 9593 1747 9609
rect 1713 9543 1747 9559
rect 216919 9593 216953 9609
rect 216919 9543 216953 9559
rect 1713 9257 1747 9273
rect 1713 9207 1747 9223
rect 216919 9257 216953 9273
rect 216919 9207 216953 9223
rect 1713 8921 1747 8937
rect 1713 8871 1747 8887
rect 216919 8921 216953 8937
rect 216919 8871 216953 8887
rect 1713 8585 1747 8601
rect 1713 8535 1747 8551
rect 216919 8585 216953 8601
rect 216919 8535 216953 8551
rect 1713 8249 1747 8265
rect 1713 8199 1747 8215
rect 216919 8249 216953 8265
rect 216919 8199 216953 8215
rect 1713 7913 1747 7929
rect 1713 7863 1747 7879
rect 216919 7913 216953 7929
rect 216919 7863 216953 7879
rect 1713 7577 1747 7593
rect 1713 7527 1747 7543
rect 216919 7577 216953 7593
rect 216919 7527 216953 7543
rect 1713 7241 1747 7257
rect 1713 7191 1747 7207
rect 216919 7241 216953 7257
rect 216919 7191 216953 7207
rect 1713 6905 1747 6921
rect 1713 6855 1747 6871
rect 216919 6905 216953 6921
rect 216919 6855 216953 6871
rect 1713 6569 1747 6585
rect 1713 6519 1747 6535
rect 216919 6569 216953 6585
rect 216919 6519 216953 6535
rect 1713 6233 1747 6249
rect 1713 6183 1747 6199
rect 216919 6233 216953 6249
rect 216919 6183 216953 6199
rect 1713 5897 1747 5913
rect 1713 5847 1747 5863
rect 216919 5897 216953 5913
rect 216919 5847 216953 5863
rect 1713 5561 1747 5577
rect 1713 5511 1747 5527
rect 216919 5561 216953 5577
rect 216919 5511 216953 5527
rect 1713 5225 1747 5241
rect 1713 5175 1747 5191
rect 216919 5225 216953 5241
rect 216919 5175 216953 5191
rect 1713 4889 1747 4905
rect 1713 4839 1747 4855
rect 216919 4889 216953 4905
rect 216919 4839 216953 4855
rect 1713 4553 1747 4569
rect 1713 4503 1747 4519
rect 216919 4553 216953 4569
rect 216919 4503 216953 4519
rect 1713 4217 1747 4233
rect 1713 4167 1747 4183
rect 216919 4217 216953 4233
rect 216919 4167 216953 4183
rect 1713 3881 1747 3897
rect 1713 3831 1747 3847
rect 216919 3881 216953 3897
rect 216919 3831 216953 3847
rect 1713 3545 1747 3561
rect 1713 3495 1747 3511
rect 216919 3545 216953 3561
rect 216919 3495 216953 3511
rect 1713 3209 1747 3225
rect 1713 3159 1747 3175
rect 216919 3209 216953 3225
rect 216919 3159 216953 3175
rect 1713 2873 1747 2889
rect 1713 2823 1747 2839
rect 216919 2873 216953 2889
rect 216919 2823 216953 2839
rect 1713 2537 1747 2553
rect 1713 2487 1747 2503
rect 216919 2537 216953 2553
rect 216919 2487 216953 2503
rect 1713 2201 1747 2217
rect 1713 2151 1747 2167
rect 216919 2201 216953 2217
rect 216919 2151 216953 2167
rect 2049 1865 2083 1881
rect 2049 1815 2083 1831
rect 2385 1865 2419 1881
rect 2385 1815 2419 1831
rect 2721 1865 2755 1881
rect 2721 1815 2755 1831
rect 3057 1865 3091 1881
rect 3057 1815 3091 1831
rect 3393 1865 3427 1881
rect 3393 1815 3427 1831
rect 3729 1865 3763 1881
rect 3729 1815 3763 1831
rect 4065 1865 4099 1881
rect 4065 1815 4099 1831
rect 4401 1865 4435 1881
rect 4401 1815 4435 1831
rect 4737 1865 4771 1881
rect 4737 1815 4771 1831
rect 5073 1865 5107 1881
rect 5073 1815 5107 1831
rect 5409 1865 5443 1881
rect 5409 1815 5443 1831
rect 5745 1865 5779 1881
rect 5745 1815 5779 1831
rect 6081 1865 6115 1881
rect 6081 1815 6115 1831
rect 6417 1865 6451 1881
rect 6417 1815 6451 1831
rect 6753 1865 6787 1881
rect 6753 1815 6787 1831
rect 7089 1865 7123 1881
rect 7089 1815 7123 1831
rect 7425 1865 7459 1881
rect 7425 1815 7459 1831
rect 7761 1865 7795 1881
rect 7761 1815 7795 1831
rect 8097 1865 8131 1881
rect 8097 1815 8131 1831
rect 8433 1865 8467 1881
rect 8433 1815 8467 1831
rect 8769 1865 8803 1881
rect 8769 1815 8803 1831
rect 9105 1865 9139 1881
rect 9105 1815 9139 1831
rect 9441 1865 9475 1881
rect 9441 1815 9475 1831
rect 9777 1865 9811 1881
rect 9777 1815 9811 1831
rect 10113 1865 10147 1881
rect 10113 1815 10147 1831
rect 10449 1865 10483 1881
rect 10449 1815 10483 1831
rect 10785 1865 10819 1881
rect 10785 1815 10819 1831
rect 11121 1865 11155 1881
rect 11121 1815 11155 1831
rect 11457 1865 11491 1881
rect 11457 1815 11491 1831
rect 11793 1865 11827 1881
rect 11793 1815 11827 1831
rect 12129 1865 12163 1881
rect 12129 1815 12163 1831
rect 12465 1865 12499 1881
rect 12465 1815 12499 1831
rect 12801 1865 12835 1881
rect 12801 1815 12835 1831
rect 13137 1865 13171 1881
rect 13137 1815 13171 1831
rect 13473 1865 13507 1881
rect 13473 1815 13507 1831
rect 13809 1865 13843 1881
rect 13809 1815 13843 1831
rect 14145 1865 14179 1881
rect 14145 1815 14179 1831
rect 14481 1865 14515 1881
rect 14481 1815 14515 1831
rect 14817 1865 14851 1881
rect 14817 1815 14851 1831
rect 15153 1865 15187 1881
rect 15153 1815 15187 1831
rect 15489 1865 15523 1881
rect 15489 1815 15523 1831
rect 15825 1865 15859 1881
rect 15825 1815 15859 1831
rect 16161 1865 16195 1881
rect 16161 1815 16195 1831
rect 16497 1865 16531 1881
rect 16497 1815 16531 1831
rect 16833 1865 16867 1881
rect 16833 1815 16867 1831
rect 17169 1865 17203 1881
rect 17169 1815 17203 1831
rect 17505 1865 17539 1881
rect 17505 1815 17539 1831
rect 17841 1865 17875 1881
rect 17841 1815 17875 1831
rect 18177 1865 18211 1881
rect 18177 1815 18211 1831
rect 18513 1865 18547 1881
rect 18513 1815 18547 1831
rect 18849 1865 18883 1881
rect 18849 1815 18883 1831
rect 19185 1865 19219 1881
rect 19185 1815 19219 1831
rect 19521 1865 19555 1881
rect 19521 1815 19555 1831
rect 19857 1865 19891 1881
rect 19857 1815 19891 1831
rect 20193 1865 20227 1881
rect 20193 1815 20227 1831
rect 20529 1865 20563 1881
rect 20529 1815 20563 1831
rect 20865 1865 20899 1881
rect 20865 1815 20899 1831
rect 21201 1865 21235 1881
rect 21201 1815 21235 1831
rect 21537 1865 21571 1881
rect 21537 1815 21571 1831
rect 21873 1865 21907 1881
rect 21873 1815 21907 1831
rect 22209 1865 22243 1881
rect 22209 1815 22243 1831
rect 22545 1865 22579 1881
rect 22545 1815 22579 1831
rect 22881 1865 22915 1881
rect 22881 1815 22915 1831
rect 23217 1865 23251 1881
rect 23217 1815 23251 1831
rect 23553 1865 23587 1881
rect 23553 1815 23587 1831
rect 23889 1865 23923 1881
rect 23889 1815 23923 1831
rect 24225 1865 24259 1881
rect 24225 1815 24259 1831
rect 24561 1865 24595 1881
rect 24561 1815 24595 1831
rect 24897 1865 24931 1881
rect 24897 1815 24931 1831
rect 25233 1865 25267 1881
rect 25233 1815 25267 1831
rect 25569 1865 25603 1881
rect 25569 1815 25603 1831
rect 25905 1865 25939 1881
rect 25905 1815 25939 1831
rect 26241 1865 26275 1881
rect 26241 1815 26275 1831
rect 26577 1865 26611 1881
rect 26577 1815 26611 1831
rect 26913 1865 26947 1881
rect 26913 1815 26947 1831
rect 27249 1865 27283 1881
rect 27249 1815 27283 1831
rect 27585 1865 27619 1881
rect 27585 1815 27619 1831
rect 27921 1865 27955 1881
rect 27921 1815 27955 1831
rect 28257 1865 28291 1881
rect 28257 1815 28291 1831
rect 28593 1865 28627 1881
rect 28593 1815 28627 1831
rect 28929 1865 28963 1881
rect 28929 1815 28963 1831
rect 29265 1865 29299 1881
rect 29265 1815 29299 1831
rect 29601 1865 29635 1881
rect 29601 1815 29635 1831
rect 29937 1865 29971 1881
rect 29937 1815 29971 1831
rect 30273 1865 30307 1881
rect 30273 1815 30307 1831
rect 30609 1865 30643 1881
rect 30609 1815 30643 1831
rect 30945 1865 30979 1881
rect 30945 1815 30979 1831
rect 31281 1865 31315 1881
rect 31281 1815 31315 1831
rect 31617 1865 31651 1881
rect 31617 1815 31651 1831
rect 31953 1865 31987 1881
rect 31953 1815 31987 1831
rect 32289 1865 32323 1881
rect 32289 1815 32323 1831
rect 32625 1865 32659 1881
rect 32625 1815 32659 1831
rect 32961 1865 32995 1881
rect 32961 1815 32995 1831
rect 33297 1865 33331 1881
rect 33297 1815 33331 1831
rect 33633 1865 33667 1881
rect 33633 1815 33667 1831
rect 33969 1865 34003 1881
rect 33969 1815 34003 1831
rect 34305 1865 34339 1881
rect 34305 1815 34339 1831
rect 34641 1865 34675 1881
rect 34641 1815 34675 1831
rect 34977 1865 35011 1881
rect 34977 1815 35011 1831
rect 35313 1865 35347 1881
rect 35313 1815 35347 1831
rect 35649 1865 35683 1881
rect 35649 1815 35683 1831
rect 35985 1865 36019 1881
rect 35985 1815 36019 1831
rect 36321 1865 36355 1881
rect 36321 1815 36355 1831
rect 36657 1865 36691 1881
rect 36657 1815 36691 1831
rect 36993 1865 37027 1881
rect 36993 1815 37027 1831
rect 37329 1865 37363 1881
rect 37329 1815 37363 1831
rect 37665 1865 37699 1881
rect 37665 1815 37699 1831
rect 38001 1865 38035 1881
rect 38001 1815 38035 1831
rect 38337 1865 38371 1881
rect 38337 1815 38371 1831
rect 38673 1865 38707 1881
rect 38673 1815 38707 1831
rect 39009 1865 39043 1881
rect 39009 1815 39043 1831
rect 39345 1865 39379 1881
rect 39345 1815 39379 1831
rect 39681 1865 39715 1881
rect 39681 1815 39715 1831
rect 40017 1865 40051 1881
rect 40017 1815 40051 1831
rect 40353 1865 40387 1881
rect 40353 1815 40387 1831
rect 40689 1865 40723 1881
rect 40689 1815 40723 1831
rect 41025 1865 41059 1881
rect 41025 1815 41059 1831
rect 41361 1865 41395 1881
rect 41361 1815 41395 1831
rect 41697 1865 41731 1881
rect 41697 1815 41731 1831
rect 42033 1865 42067 1881
rect 42033 1815 42067 1831
rect 42369 1865 42403 1881
rect 42369 1815 42403 1831
rect 42705 1865 42739 1881
rect 42705 1815 42739 1831
rect 43041 1865 43075 1881
rect 43041 1815 43075 1831
rect 43377 1865 43411 1881
rect 43377 1815 43411 1831
rect 43713 1865 43747 1881
rect 43713 1815 43747 1831
rect 44049 1865 44083 1881
rect 44049 1815 44083 1831
rect 44385 1865 44419 1881
rect 44385 1815 44419 1831
rect 44721 1865 44755 1881
rect 44721 1815 44755 1831
rect 45057 1865 45091 1881
rect 45057 1815 45091 1831
rect 45393 1865 45427 1881
rect 45393 1815 45427 1831
rect 45729 1865 45763 1881
rect 45729 1815 45763 1831
rect 46065 1865 46099 1881
rect 46065 1815 46099 1831
rect 46401 1865 46435 1881
rect 46401 1815 46435 1831
rect 46737 1865 46771 1881
rect 46737 1815 46771 1831
rect 47073 1865 47107 1881
rect 47073 1815 47107 1831
rect 47409 1865 47443 1881
rect 47409 1815 47443 1831
rect 47745 1865 47779 1881
rect 47745 1815 47779 1831
rect 48081 1865 48115 1881
rect 48081 1815 48115 1831
rect 48417 1865 48451 1881
rect 48417 1815 48451 1831
rect 48753 1865 48787 1881
rect 48753 1815 48787 1831
rect 49089 1865 49123 1881
rect 49089 1815 49123 1831
rect 49425 1865 49459 1881
rect 49425 1815 49459 1831
rect 49761 1865 49795 1881
rect 49761 1815 49795 1831
rect 50097 1865 50131 1881
rect 50097 1815 50131 1831
rect 50433 1865 50467 1881
rect 50433 1815 50467 1831
rect 50769 1865 50803 1881
rect 50769 1815 50803 1831
rect 51105 1865 51139 1881
rect 51105 1815 51139 1831
rect 51441 1865 51475 1881
rect 51441 1815 51475 1831
rect 51777 1865 51811 1881
rect 51777 1815 51811 1831
rect 52113 1865 52147 1881
rect 52113 1815 52147 1831
rect 52449 1865 52483 1881
rect 52449 1815 52483 1831
rect 52785 1865 52819 1881
rect 52785 1815 52819 1831
rect 53121 1865 53155 1881
rect 53121 1815 53155 1831
rect 53457 1865 53491 1881
rect 53457 1815 53491 1831
rect 53793 1865 53827 1881
rect 53793 1815 53827 1831
rect 54129 1865 54163 1881
rect 54129 1815 54163 1831
rect 54465 1865 54499 1881
rect 54465 1815 54499 1831
rect 54801 1865 54835 1881
rect 54801 1815 54835 1831
rect 55137 1865 55171 1881
rect 55137 1815 55171 1831
rect 55473 1865 55507 1881
rect 55473 1815 55507 1831
rect 55809 1865 55843 1881
rect 55809 1815 55843 1831
rect 56145 1865 56179 1881
rect 56145 1815 56179 1831
rect 56481 1865 56515 1881
rect 56481 1815 56515 1831
rect 56817 1865 56851 1881
rect 56817 1815 56851 1831
rect 57153 1865 57187 1881
rect 57153 1815 57187 1831
rect 57489 1865 57523 1881
rect 57489 1815 57523 1831
rect 57825 1865 57859 1881
rect 57825 1815 57859 1831
rect 58161 1865 58195 1881
rect 58161 1815 58195 1831
rect 58497 1865 58531 1881
rect 58497 1815 58531 1831
rect 58833 1865 58867 1881
rect 58833 1815 58867 1831
rect 59169 1865 59203 1881
rect 59169 1815 59203 1831
rect 59505 1865 59539 1881
rect 59505 1815 59539 1831
rect 59841 1865 59875 1881
rect 59841 1815 59875 1831
rect 60177 1865 60211 1881
rect 60177 1815 60211 1831
rect 60513 1865 60547 1881
rect 60513 1815 60547 1831
rect 60849 1865 60883 1881
rect 60849 1815 60883 1831
rect 61185 1865 61219 1881
rect 61185 1815 61219 1831
rect 61521 1865 61555 1881
rect 61521 1815 61555 1831
rect 61857 1865 61891 1881
rect 61857 1815 61891 1831
rect 62193 1865 62227 1881
rect 62193 1815 62227 1831
rect 62529 1865 62563 1881
rect 62529 1815 62563 1831
rect 62865 1865 62899 1881
rect 62865 1815 62899 1831
rect 63201 1865 63235 1881
rect 63201 1815 63235 1831
rect 63537 1865 63571 1881
rect 63537 1815 63571 1831
rect 63873 1865 63907 1881
rect 63873 1815 63907 1831
rect 64209 1865 64243 1881
rect 64209 1815 64243 1831
rect 64545 1865 64579 1881
rect 64545 1815 64579 1831
rect 64881 1865 64915 1881
rect 64881 1815 64915 1831
rect 65217 1865 65251 1881
rect 65217 1815 65251 1831
rect 65553 1865 65587 1881
rect 65553 1815 65587 1831
rect 65889 1865 65923 1881
rect 65889 1815 65923 1831
rect 66225 1865 66259 1881
rect 66225 1815 66259 1831
rect 66561 1865 66595 1881
rect 66561 1815 66595 1831
rect 66897 1865 66931 1881
rect 66897 1815 66931 1831
rect 67233 1865 67267 1881
rect 67233 1815 67267 1831
rect 67569 1865 67603 1881
rect 67569 1815 67603 1831
rect 67905 1865 67939 1881
rect 67905 1815 67939 1831
rect 68241 1865 68275 1881
rect 68241 1815 68275 1831
rect 68577 1865 68611 1881
rect 68577 1815 68611 1831
rect 68913 1865 68947 1881
rect 68913 1815 68947 1831
rect 69249 1865 69283 1881
rect 69249 1815 69283 1831
rect 69585 1865 69619 1881
rect 69585 1815 69619 1831
rect 69921 1865 69955 1881
rect 69921 1815 69955 1831
rect 70257 1865 70291 1881
rect 70257 1815 70291 1831
rect 70593 1865 70627 1881
rect 70593 1815 70627 1831
rect 70929 1865 70963 1881
rect 70929 1815 70963 1831
rect 71265 1865 71299 1881
rect 71265 1815 71299 1831
rect 71601 1865 71635 1881
rect 71601 1815 71635 1831
rect 71937 1865 71971 1881
rect 71937 1815 71971 1831
rect 72273 1865 72307 1881
rect 72273 1815 72307 1831
rect 72609 1865 72643 1881
rect 72609 1815 72643 1831
rect 72945 1865 72979 1881
rect 72945 1815 72979 1831
rect 73281 1865 73315 1881
rect 73281 1815 73315 1831
rect 73617 1865 73651 1881
rect 73617 1815 73651 1831
rect 73953 1865 73987 1881
rect 73953 1815 73987 1831
rect 74289 1865 74323 1881
rect 74289 1815 74323 1831
rect 74625 1865 74659 1881
rect 74625 1815 74659 1831
rect 74961 1865 74995 1881
rect 74961 1815 74995 1831
rect 75297 1865 75331 1881
rect 75297 1815 75331 1831
rect 75633 1865 75667 1881
rect 75633 1815 75667 1831
rect 75969 1865 76003 1881
rect 75969 1815 76003 1831
rect 76305 1865 76339 1881
rect 76305 1815 76339 1831
rect 76641 1865 76675 1881
rect 76641 1815 76675 1831
rect 76977 1865 77011 1881
rect 76977 1815 77011 1831
rect 77313 1865 77347 1881
rect 77313 1815 77347 1831
rect 77649 1865 77683 1881
rect 77649 1815 77683 1831
rect 77985 1865 78019 1881
rect 77985 1815 78019 1831
rect 78321 1865 78355 1881
rect 78321 1815 78355 1831
rect 78657 1865 78691 1881
rect 78657 1815 78691 1831
rect 78993 1865 79027 1881
rect 78993 1815 79027 1831
rect 79329 1865 79363 1881
rect 79329 1815 79363 1831
rect 79665 1865 79699 1881
rect 79665 1815 79699 1831
rect 80001 1865 80035 1881
rect 80001 1815 80035 1831
rect 80337 1865 80371 1881
rect 80337 1815 80371 1831
rect 80673 1865 80707 1881
rect 80673 1815 80707 1831
rect 81009 1865 81043 1881
rect 81009 1815 81043 1831
rect 81345 1865 81379 1881
rect 81345 1815 81379 1831
rect 81681 1865 81715 1881
rect 81681 1815 81715 1831
rect 82017 1865 82051 1881
rect 82017 1815 82051 1831
rect 82353 1865 82387 1881
rect 82353 1815 82387 1831
rect 82689 1865 82723 1881
rect 82689 1815 82723 1831
rect 83025 1865 83059 1881
rect 83025 1815 83059 1831
rect 83361 1865 83395 1881
rect 83361 1815 83395 1831
rect 83697 1865 83731 1881
rect 83697 1815 83731 1831
rect 84033 1865 84067 1881
rect 84033 1815 84067 1831
rect 84369 1865 84403 1881
rect 84369 1815 84403 1831
rect 84705 1865 84739 1881
rect 84705 1815 84739 1831
rect 85041 1865 85075 1881
rect 85041 1815 85075 1831
rect 85377 1865 85411 1881
rect 85377 1815 85411 1831
rect 85713 1865 85747 1881
rect 85713 1815 85747 1831
rect 86049 1865 86083 1881
rect 86049 1815 86083 1831
rect 86385 1865 86419 1881
rect 86385 1815 86419 1831
rect 86721 1865 86755 1881
rect 86721 1815 86755 1831
rect 87057 1865 87091 1881
rect 87057 1815 87091 1831
rect 87393 1865 87427 1881
rect 87393 1815 87427 1831
rect 87729 1865 87763 1881
rect 87729 1815 87763 1831
rect 88065 1865 88099 1881
rect 88065 1815 88099 1831
rect 88401 1865 88435 1881
rect 88401 1815 88435 1831
rect 88737 1865 88771 1881
rect 88737 1815 88771 1831
rect 89073 1865 89107 1881
rect 89073 1815 89107 1831
rect 89409 1865 89443 1881
rect 89409 1815 89443 1831
rect 89745 1865 89779 1881
rect 89745 1815 89779 1831
rect 90081 1865 90115 1881
rect 90081 1815 90115 1831
rect 90417 1865 90451 1881
rect 90417 1815 90451 1831
rect 90753 1865 90787 1881
rect 90753 1815 90787 1831
rect 91089 1865 91123 1881
rect 91089 1815 91123 1831
rect 91425 1865 91459 1881
rect 91425 1815 91459 1831
rect 91761 1865 91795 1881
rect 91761 1815 91795 1831
rect 92097 1865 92131 1881
rect 92097 1815 92131 1831
rect 92433 1865 92467 1881
rect 92433 1815 92467 1831
rect 92769 1865 92803 1881
rect 92769 1815 92803 1831
rect 93105 1865 93139 1881
rect 93105 1815 93139 1831
rect 93441 1865 93475 1881
rect 93441 1815 93475 1831
rect 93777 1865 93811 1881
rect 93777 1815 93811 1831
rect 94113 1865 94147 1881
rect 94113 1815 94147 1831
rect 94449 1865 94483 1881
rect 94449 1815 94483 1831
rect 94785 1865 94819 1881
rect 94785 1815 94819 1831
rect 95121 1865 95155 1881
rect 95121 1815 95155 1831
rect 95457 1865 95491 1881
rect 95457 1815 95491 1831
rect 95793 1865 95827 1881
rect 95793 1815 95827 1831
rect 96129 1865 96163 1881
rect 96129 1815 96163 1831
rect 96465 1865 96499 1881
rect 96465 1815 96499 1831
rect 96801 1865 96835 1881
rect 96801 1815 96835 1831
rect 97137 1865 97171 1881
rect 97137 1815 97171 1831
rect 97473 1865 97507 1881
rect 97473 1815 97507 1831
rect 97809 1865 97843 1881
rect 97809 1815 97843 1831
rect 98145 1865 98179 1881
rect 98145 1815 98179 1831
rect 98481 1865 98515 1881
rect 98481 1815 98515 1831
rect 98817 1865 98851 1881
rect 98817 1815 98851 1831
rect 99153 1865 99187 1881
rect 99153 1815 99187 1831
rect 99489 1865 99523 1881
rect 99489 1815 99523 1831
rect 99825 1865 99859 1881
rect 99825 1815 99859 1831
rect 100161 1865 100195 1881
rect 100161 1815 100195 1831
rect 100497 1865 100531 1881
rect 100497 1815 100531 1831
rect 100833 1865 100867 1881
rect 100833 1815 100867 1831
rect 101169 1865 101203 1881
rect 101169 1815 101203 1831
rect 101505 1865 101539 1881
rect 101505 1815 101539 1831
rect 101841 1865 101875 1881
rect 101841 1815 101875 1831
rect 102177 1865 102211 1881
rect 102177 1815 102211 1831
rect 102513 1865 102547 1881
rect 102513 1815 102547 1831
rect 102849 1865 102883 1881
rect 102849 1815 102883 1831
rect 103185 1865 103219 1881
rect 103185 1815 103219 1831
rect 103521 1865 103555 1881
rect 103521 1815 103555 1831
rect 103857 1865 103891 1881
rect 103857 1815 103891 1831
rect 104193 1865 104227 1881
rect 104193 1815 104227 1831
rect 104529 1865 104563 1881
rect 104529 1815 104563 1831
rect 104865 1865 104899 1881
rect 104865 1815 104899 1831
rect 105201 1865 105235 1881
rect 105201 1815 105235 1831
rect 105537 1865 105571 1881
rect 105537 1815 105571 1831
rect 105873 1865 105907 1881
rect 105873 1815 105907 1831
rect 106209 1865 106243 1881
rect 106209 1815 106243 1831
rect 106545 1865 106579 1881
rect 106545 1815 106579 1831
rect 106881 1865 106915 1881
rect 106881 1815 106915 1831
rect 107217 1865 107251 1881
rect 107217 1815 107251 1831
rect 107553 1865 107587 1881
rect 107553 1815 107587 1831
rect 107889 1865 107923 1881
rect 107889 1815 107923 1831
rect 108225 1865 108259 1881
rect 108225 1815 108259 1831
rect 108561 1865 108595 1881
rect 108561 1815 108595 1831
rect 108897 1865 108931 1881
rect 108897 1815 108931 1831
rect 109233 1865 109267 1881
rect 109233 1815 109267 1831
rect 109569 1865 109603 1881
rect 109569 1815 109603 1831
rect 109905 1865 109939 1881
rect 109905 1815 109939 1831
rect 110241 1865 110275 1881
rect 110241 1815 110275 1831
rect 110577 1865 110611 1881
rect 110577 1815 110611 1831
rect 110913 1865 110947 1881
rect 110913 1815 110947 1831
rect 111249 1865 111283 1881
rect 111249 1815 111283 1831
rect 111585 1865 111619 1881
rect 111585 1815 111619 1831
rect 111921 1865 111955 1881
rect 111921 1815 111955 1831
rect 112257 1865 112291 1881
rect 112257 1815 112291 1831
rect 112593 1865 112627 1881
rect 112593 1815 112627 1831
rect 112929 1865 112963 1881
rect 112929 1815 112963 1831
rect 113265 1865 113299 1881
rect 113265 1815 113299 1831
rect 113601 1865 113635 1881
rect 113601 1815 113635 1831
rect 113937 1865 113971 1881
rect 113937 1815 113971 1831
rect 114273 1865 114307 1881
rect 114273 1815 114307 1831
rect 114609 1865 114643 1881
rect 114609 1815 114643 1831
rect 114945 1865 114979 1881
rect 114945 1815 114979 1831
rect 115281 1865 115315 1881
rect 115281 1815 115315 1831
rect 115617 1865 115651 1881
rect 115617 1815 115651 1831
rect 115953 1865 115987 1881
rect 115953 1815 115987 1831
rect 116289 1865 116323 1881
rect 116289 1815 116323 1831
rect 116625 1865 116659 1881
rect 116625 1815 116659 1831
rect 116961 1865 116995 1881
rect 116961 1815 116995 1831
rect 117297 1865 117331 1881
rect 117297 1815 117331 1831
rect 117633 1865 117667 1881
rect 117633 1815 117667 1831
rect 117969 1865 118003 1881
rect 117969 1815 118003 1831
rect 118305 1865 118339 1881
rect 118305 1815 118339 1831
rect 118641 1865 118675 1881
rect 118641 1815 118675 1831
rect 118977 1865 119011 1881
rect 118977 1815 119011 1831
rect 119313 1865 119347 1881
rect 119313 1815 119347 1831
rect 119649 1865 119683 1881
rect 119649 1815 119683 1831
rect 119985 1865 120019 1881
rect 119985 1815 120019 1831
rect 120321 1865 120355 1881
rect 120321 1815 120355 1831
rect 120657 1865 120691 1881
rect 120657 1815 120691 1831
rect 120993 1865 121027 1881
rect 120993 1815 121027 1831
rect 121329 1865 121363 1881
rect 121329 1815 121363 1831
rect 121665 1865 121699 1881
rect 121665 1815 121699 1831
rect 122001 1865 122035 1881
rect 122001 1815 122035 1831
rect 122337 1865 122371 1881
rect 122337 1815 122371 1831
rect 122673 1865 122707 1881
rect 122673 1815 122707 1831
rect 123009 1865 123043 1881
rect 123009 1815 123043 1831
rect 123345 1865 123379 1881
rect 123345 1815 123379 1831
rect 123681 1865 123715 1881
rect 123681 1815 123715 1831
rect 124017 1865 124051 1881
rect 124017 1815 124051 1831
rect 124353 1865 124387 1881
rect 124353 1815 124387 1831
rect 124689 1865 124723 1881
rect 124689 1815 124723 1831
rect 125025 1865 125059 1881
rect 125025 1815 125059 1831
rect 125361 1865 125395 1881
rect 125361 1815 125395 1831
rect 125697 1865 125731 1881
rect 125697 1815 125731 1831
rect 126033 1865 126067 1881
rect 126033 1815 126067 1831
rect 126369 1865 126403 1881
rect 126369 1815 126403 1831
rect 126705 1865 126739 1881
rect 126705 1815 126739 1831
rect 127041 1865 127075 1881
rect 127041 1815 127075 1831
rect 127377 1865 127411 1881
rect 127377 1815 127411 1831
rect 127713 1865 127747 1881
rect 127713 1815 127747 1831
rect 128049 1865 128083 1881
rect 128049 1815 128083 1831
rect 128385 1865 128419 1881
rect 128385 1815 128419 1831
rect 128721 1865 128755 1881
rect 128721 1815 128755 1831
rect 129057 1865 129091 1881
rect 129057 1815 129091 1831
rect 129393 1865 129427 1881
rect 129393 1815 129427 1831
rect 129729 1865 129763 1881
rect 129729 1815 129763 1831
rect 130065 1865 130099 1881
rect 130065 1815 130099 1831
rect 130401 1865 130435 1881
rect 130401 1815 130435 1831
rect 130737 1865 130771 1881
rect 130737 1815 130771 1831
rect 131073 1865 131107 1881
rect 131073 1815 131107 1831
rect 131409 1865 131443 1881
rect 131409 1815 131443 1831
rect 131745 1865 131779 1881
rect 131745 1815 131779 1831
rect 132081 1865 132115 1881
rect 132081 1815 132115 1831
rect 132417 1865 132451 1881
rect 132417 1815 132451 1831
rect 132753 1865 132787 1881
rect 132753 1815 132787 1831
rect 133089 1865 133123 1881
rect 133089 1815 133123 1831
rect 133425 1865 133459 1881
rect 133425 1815 133459 1831
rect 133761 1865 133795 1881
rect 133761 1815 133795 1831
rect 134097 1865 134131 1881
rect 134097 1815 134131 1831
rect 134433 1865 134467 1881
rect 134433 1815 134467 1831
rect 134769 1865 134803 1881
rect 134769 1815 134803 1831
rect 135105 1865 135139 1881
rect 135105 1815 135139 1831
rect 135441 1865 135475 1881
rect 135441 1815 135475 1831
rect 135777 1865 135811 1881
rect 135777 1815 135811 1831
rect 136113 1865 136147 1881
rect 136113 1815 136147 1831
rect 136449 1865 136483 1881
rect 136449 1815 136483 1831
rect 136785 1865 136819 1881
rect 136785 1815 136819 1831
rect 137121 1865 137155 1881
rect 137121 1815 137155 1831
rect 137457 1865 137491 1881
rect 137457 1815 137491 1831
rect 137793 1865 137827 1881
rect 137793 1815 137827 1831
rect 138129 1865 138163 1881
rect 138129 1815 138163 1831
rect 138465 1865 138499 1881
rect 138465 1815 138499 1831
rect 138801 1865 138835 1881
rect 138801 1815 138835 1831
rect 139137 1865 139171 1881
rect 139137 1815 139171 1831
rect 139473 1865 139507 1881
rect 139473 1815 139507 1831
rect 139809 1865 139843 1881
rect 139809 1815 139843 1831
rect 140145 1865 140179 1881
rect 140145 1815 140179 1831
rect 140481 1865 140515 1881
rect 140481 1815 140515 1831
rect 140817 1865 140851 1881
rect 140817 1815 140851 1831
rect 141153 1865 141187 1881
rect 141153 1815 141187 1831
rect 141489 1865 141523 1881
rect 141489 1815 141523 1831
rect 141825 1865 141859 1881
rect 141825 1815 141859 1831
rect 142161 1865 142195 1881
rect 142161 1815 142195 1831
rect 142497 1865 142531 1881
rect 142497 1815 142531 1831
rect 142833 1865 142867 1881
rect 142833 1815 142867 1831
rect 143169 1865 143203 1881
rect 143169 1815 143203 1831
rect 143505 1865 143539 1881
rect 143505 1815 143539 1831
rect 143841 1865 143875 1881
rect 143841 1815 143875 1831
rect 144177 1865 144211 1881
rect 144177 1815 144211 1831
rect 144513 1865 144547 1881
rect 144513 1815 144547 1831
rect 144849 1865 144883 1881
rect 144849 1815 144883 1831
rect 145185 1865 145219 1881
rect 145185 1815 145219 1831
rect 145521 1865 145555 1881
rect 145521 1815 145555 1831
rect 145857 1865 145891 1881
rect 145857 1815 145891 1831
rect 146193 1865 146227 1881
rect 146193 1815 146227 1831
rect 146529 1865 146563 1881
rect 146529 1815 146563 1831
rect 146865 1865 146899 1881
rect 146865 1815 146899 1831
rect 147201 1865 147235 1881
rect 147201 1815 147235 1831
rect 147537 1865 147571 1881
rect 147537 1815 147571 1831
rect 147873 1865 147907 1881
rect 147873 1815 147907 1831
rect 148209 1865 148243 1881
rect 148209 1815 148243 1831
rect 148545 1865 148579 1881
rect 148545 1815 148579 1831
rect 148881 1865 148915 1881
rect 148881 1815 148915 1831
rect 149217 1865 149251 1881
rect 149217 1815 149251 1831
rect 149553 1865 149587 1881
rect 149553 1815 149587 1831
rect 149889 1865 149923 1881
rect 149889 1815 149923 1831
rect 150225 1865 150259 1881
rect 150225 1815 150259 1831
rect 150561 1865 150595 1881
rect 150561 1815 150595 1831
rect 150897 1865 150931 1881
rect 150897 1815 150931 1831
rect 151233 1865 151267 1881
rect 151233 1815 151267 1831
rect 151569 1865 151603 1881
rect 151569 1815 151603 1831
rect 151905 1865 151939 1881
rect 151905 1815 151939 1831
rect 152241 1865 152275 1881
rect 152241 1815 152275 1831
rect 152577 1865 152611 1881
rect 152577 1815 152611 1831
rect 152913 1865 152947 1881
rect 152913 1815 152947 1831
rect 153249 1865 153283 1881
rect 153249 1815 153283 1831
rect 153585 1865 153619 1881
rect 153585 1815 153619 1831
rect 153921 1865 153955 1881
rect 153921 1815 153955 1831
rect 154257 1865 154291 1881
rect 154257 1815 154291 1831
rect 154593 1865 154627 1881
rect 154593 1815 154627 1831
rect 154929 1865 154963 1881
rect 154929 1815 154963 1831
rect 155265 1865 155299 1881
rect 155265 1815 155299 1831
rect 155601 1865 155635 1881
rect 155601 1815 155635 1831
rect 155937 1865 155971 1881
rect 155937 1815 155971 1831
rect 156273 1865 156307 1881
rect 156273 1815 156307 1831
rect 156609 1865 156643 1881
rect 156609 1815 156643 1831
rect 156945 1865 156979 1881
rect 156945 1815 156979 1831
rect 157281 1865 157315 1881
rect 157281 1815 157315 1831
rect 157617 1865 157651 1881
rect 157617 1815 157651 1831
rect 157953 1865 157987 1881
rect 157953 1815 157987 1831
rect 158289 1865 158323 1881
rect 158289 1815 158323 1831
rect 158625 1865 158659 1881
rect 158625 1815 158659 1831
rect 158961 1865 158995 1881
rect 158961 1815 158995 1831
rect 159297 1865 159331 1881
rect 159297 1815 159331 1831
rect 159633 1865 159667 1881
rect 159633 1815 159667 1831
rect 159969 1865 160003 1881
rect 159969 1815 160003 1831
rect 160305 1865 160339 1881
rect 160305 1815 160339 1831
rect 160641 1865 160675 1881
rect 160641 1815 160675 1831
rect 160977 1865 161011 1881
rect 160977 1815 161011 1831
rect 161313 1865 161347 1881
rect 161313 1815 161347 1831
rect 161649 1865 161683 1881
rect 161649 1815 161683 1831
rect 161985 1865 162019 1881
rect 161985 1815 162019 1831
rect 162321 1865 162355 1881
rect 162321 1815 162355 1831
rect 162657 1865 162691 1881
rect 162657 1815 162691 1831
rect 162993 1865 163027 1881
rect 162993 1815 163027 1831
rect 163329 1865 163363 1881
rect 163329 1815 163363 1831
rect 163665 1865 163699 1881
rect 163665 1815 163699 1831
rect 164001 1865 164035 1881
rect 164001 1815 164035 1831
rect 164337 1865 164371 1881
rect 164337 1815 164371 1831
rect 164673 1865 164707 1881
rect 164673 1815 164707 1831
rect 165009 1865 165043 1881
rect 165009 1815 165043 1831
rect 165345 1865 165379 1881
rect 165345 1815 165379 1831
rect 165681 1865 165715 1881
rect 165681 1815 165715 1831
rect 166017 1865 166051 1881
rect 166017 1815 166051 1831
rect 166353 1865 166387 1881
rect 166353 1815 166387 1831
rect 166689 1865 166723 1881
rect 166689 1815 166723 1831
rect 167025 1865 167059 1881
rect 167025 1815 167059 1831
rect 167361 1865 167395 1881
rect 167361 1815 167395 1831
rect 167697 1865 167731 1881
rect 167697 1815 167731 1831
rect 168033 1865 168067 1881
rect 168033 1815 168067 1831
rect 168369 1865 168403 1881
rect 168369 1815 168403 1831
rect 168705 1865 168739 1881
rect 168705 1815 168739 1831
rect 169041 1865 169075 1881
rect 169041 1815 169075 1831
rect 169377 1865 169411 1881
rect 169377 1815 169411 1831
rect 169713 1865 169747 1881
rect 169713 1815 169747 1831
rect 170049 1865 170083 1881
rect 170049 1815 170083 1831
rect 170385 1865 170419 1881
rect 170385 1815 170419 1831
rect 170721 1865 170755 1881
rect 170721 1815 170755 1831
rect 171057 1865 171091 1881
rect 171057 1815 171091 1831
rect 171393 1865 171427 1881
rect 171393 1815 171427 1831
rect 171729 1865 171763 1881
rect 171729 1815 171763 1831
rect 172065 1865 172099 1881
rect 172065 1815 172099 1831
rect 172401 1865 172435 1881
rect 172401 1815 172435 1831
rect 172737 1865 172771 1881
rect 172737 1815 172771 1831
rect 173073 1865 173107 1881
rect 173073 1815 173107 1831
rect 173409 1865 173443 1881
rect 173409 1815 173443 1831
rect 173745 1865 173779 1881
rect 173745 1815 173779 1831
rect 174081 1865 174115 1881
rect 174081 1815 174115 1831
rect 174417 1865 174451 1881
rect 174417 1815 174451 1831
rect 174753 1865 174787 1881
rect 174753 1815 174787 1831
rect 175089 1865 175123 1881
rect 175089 1815 175123 1831
rect 175425 1865 175459 1881
rect 175425 1815 175459 1831
rect 175761 1865 175795 1881
rect 175761 1815 175795 1831
rect 176097 1865 176131 1881
rect 176097 1815 176131 1831
rect 176433 1865 176467 1881
rect 176433 1815 176467 1831
rect 176769 1865 176803 1881
rect 176769 1815 176803 1831
rect 177105 1865 177139 1881
rect 177105 1815 177139 1831
rect 177441 1865 177475 1881
rect 177441 1815 177475 1831
rect 177777 1865 177811 1881
rect 177777 1815 177811 1831
rect 178113 1865 178147 1881
rect 178113 1815 178147 1831
rect 178449 1865 178483 1881
rect 178449 1815 178483 1831
rect 178785 1865 178819 1881
rect 178785 1815 178819 1831
rect 179121 1865 179155 1881
rect 179121 1815 179155 1831
rect 179457 1865 179491 1881
rect 179457 1815 179491 1831
rect 179793 1865 179827 1881
rect 179793 1815 179827 1831
rect 180129 1865 180163 1881
rect 180129 1815 180163 1831
rect 180465 1865 180499 1881
rect 180465 1815 180499 1831
rect 180801 1865 180835 1881
rect 180801 1815 180835 1831
rect 181137 1865 181171 1881
rect 181137 1815 181171 1831
rect 181473 1865 181507 1881
rect 181473 1815 181507 1831
rect 181809 1865 181843 1881
rect 181809 1815 181843 1831
rect 182145 1865 182179 1881
rect 182145 1815 182179 1831
rect 182481 1865 182515 1881
rect 182481 1815 182515 1831
rect 182817 1865 182851 1881
rect 182817 1815 182851 1831
rect 183153 1865 183187 1881
rect 183153 1815 183187 1831
rect 183489 1865 183523 1881
rect 183489 1815 183523 1831
rect 183825 1865 183859 1881
rect 183825 1815 183859 1831
rect 184161 1865 184195 1881
rect 184161 1815 184195 1831
rect 184497 1865 184531 1881
rect 184497 1815 184531 1831
rect 184833 1865 184867 1881
rect 184833 1815 184867 1831
rect 185169 1865 185203 1881
rect 185169 1815 185203 1831
rect 185505 1865 185539 1881
rect 185505 1815 185539 1831
rect 185841 1865 185875 1881
rect 185841 1815 185875 1831
rect 186177 1865 186211 1881
rect 186177 1815 186211 1831
rect 186513 1865 186547 1881
rect 186513 1815 186547 1831
rect 186849 1865 186883 1881
rect 186849 1815 186883 1831
rect 187185 1865 187219 1881
rect 187185 1815 187219 1831
rect 187521 1865 187555 1881
rect 187521 1815 187555 1831
rect 187857 1865 187891 1881
rect 187857 1815 187891 1831
rect 188193 1865 188227 1881
rect 188193 1815 188227 1831
rect 188529 1865 188563 1881
rect 188529 1815 188563 1831
rect 188865 1865 188899 1881
rect 188865 1815 188899 1831
rect 189201 1865 189235 1881
rect 189201 1815 189235 1831
rect 189537 1865 189571 1881
rect 189537 1815 189571 1831
rect 189873 1865 189907 1881
rect 189873 1815 189907 1831
rect 190209 1865 190243 1881
rect 190209 1815 190243 1831
rect 190545 1865 190579 1881
rect 190545 1815 190579 1831
rect 190881 1865 190915 1881
rect 190881 1815 190915 1831
rect 191217 1865 191251 1881
rect 191217 1815 191251 1831
rect 191553 1865 191587 1881
rect 191553 1815 191587 1831
rect 191889 1865 191923 1881
rect 191889 1815 191923 1831
rect 192225 1865 192259 1881
rect 192225 1815 192259 1831
rect 192561 1865 192595 1881
rect 192561 1815 192595 1831
rect 192897 1865 192931 1881
rect 192897 1815 192931 1831
rect 193233 1865 193267 1881
rect 193233 1815 193267 1831
rect 193569 1865 193603 1881
rect 193569 1815 193603 1831
rect 193905 1865 193939 1881
rect 193905 1815 193939 1831
rect 194241 1865 194275 1881
rect 194241 1815 194275 1831
rect 194577 1865 194611 1881
rect 194577 1815 194611 1831
rect 194913 1865 194947 1881
rect 194913 1815 194947 1831
rect 195249 1865 195283 1881
rect 195249 1815 195283 1831
rect 195585 1865 195619 1881
rect 195585 1815 195619 1831
rect 195921 1865 195955 1881
rect 195921 1815 195955 1831
rect 196257 1865 196291 1881
rect 196257 1815 196291 1831
rect 196593 1865 196627 1881
rect 196593 1815 196627 1831
rect 196929 1865 196963 1881
rect 196929 1815 196963 1831
rect 197265 1865 197299 1881
rect 197265 1815 197299 1831
rect 197601 1865 197635 1881
rect 197601 1815 197635 1831
rect 197937 1865 197971 1881
rect 197937 1815 197971 1831
rect 198273 1865 198307 1881
rect 198273 1815 198307 1831
rect 198609 1865 198643 1881
rect 198609 1815 198643 1831
rect 198945 1865 198979 1881
rect 198945 1815 198979 1831
rect 199281 1865 199315 1881
rect 199281 1815 199315 1831
rect 199617 1865 199651 1881
rect 199617 1815 199651 1831
rect 199953 1865 199987 1881
rect 199953 1815 199987 1831
rect 200289 1865 200323 1881
rect 200289 1815 200323 1831
rect 200625 1865 200659 1881
rect 200625 1815 200659 1831
rect 200961 1865 200995 1881
rect 200961 1815 200995 1831
rect 201297 1865 201331 1881
rect 201297 1815 201331 1831
rect 201633 1865 201667 1881
rect 201633 1815 201667 1831
rect 201969 1865 202003 1881
rect 201969 1815 202003 1831
rect 202305 1865 202339 1881
rect 202305 1815 202339 1831
rect 202641 1865 202675 1881
rect 202641 1815 202675 1831
rect 202977 1865 203011 1881
rect 202977 1815 203011 1831
rect 203313 1865 203347 1881
rect 203313 1815 203347 1831
rect 203649 1865 203683 1881
rect 203649 1815 203683 1831
rect 203985 1865 204019 1881
rect 203985 1815 204019 1831
rect 204321 1865 204355 1881
rect 204321 1815 204355 1831
rect 204657 1865 204691 1881
rect 204657 1815 204691 1831
rect 204993 1865 205027 1881
rect 204993 1815 205027 1831
rect 205329 1865 205363 1881
rect 205329 1815 205363 1831
rect 205665 1865 205699 1881
rect 205665 1815 205699 1831
rect 206001 1865 206035 1881
rect 206001 1815 206035 1831
rect 206337 1865 206371 1881
rect 206337 1815 206371 1831
rect 206673 1865 206707 1881
rect 206673 1815 206707 1831
rect 207009 1865 207043 1881
rect 207009 1815 207043 1831
rect 207345 1865 207379 1881
rect 207345 1815 207379 1831
rect 207681 1865 207715 1881
rect 207681 1815 207715 1831
rect 208017 1865 208051 1881
rect 208017 1815 208051 1831
rect 208353 1865 208387 1881
rect 208353 1815 208387 1831
rect 208689 1865 208723 1881
rect 208689 1815 208723 1831
rect 209025 1865 209059 1881
rect 209025 1815 209059 1831
rect 209361 1865 209395 1881
rect 209361 1815 209395 1831
rect 209697 1865 209731 1881
rect 209697 1815 209731 1831
rect 210033 1865 210067 1881
rect 210033 1815 210067 1831
rect 210369 1865 210403 1881
rect 210369 1815 210403 1831
rect 210705 1865 210739 1881
rect 210705 1815 210739 1831
rect 211041 1865 211075 1881
rect 211041 1815 211075 1831
rect 211377 1865 211411 1881
rect 211377 1815 211411 1831
rect 211713 1865 211747 1881
rect 211713 1815 211747 1831
rect 212049 1865 212083 1881
rect 212049 1815 212083 1831
rect 212385 1865 212419 1881
rect 212385 1815 212419 1831
rect 212721 1865 212755 1881
rect 212721 1815 212755 1831
rect 213057 1865 213091 1881
rect 213057 1815 213091 1831
rect 213393 1865 213427 1881
rect 213393 1815 213427 1831
rect 213729 1865 213763 1881
rect 213729 1815 213763 1831
rect 214065 1865 214099 1881
rect 214065 1815 214099 1831
rect 214401 1865 214435 1881
rect 214401 1815 214435 1831
rect 214737 1865 214771 1881
rect 214737 1815 214771 1831
rect 215073 1865 215107 1881
rect 215073 1815 215107 1831
rect 215409 1865 215443 1881
rect 215409 1815 215443 1831
rect 215745 1865 215779 1881
rect 215745 1815 215779 1831
rect 216081 1865 216115 1881
rect 216081 1815 216115 1831
rect 216417 1865 216451 1881
rect 216417 1815 216451 1831
<< viali >>
rect 2049 142327 2083 142361
rect 2385 142327 2419 142361
rect 2721 142327 2755 142361
rect 3057 142327 3091 142361
rect 3393 142327 3427 142361
rect 3729 142327 3763 142361
rect 4065 142327 4099 142361
rect 4401 142327 4435 142361
rect 4737 142327 4771 142361
rect 5073 142327 5107 142361
rect 5409 142327 5443 142361
rect 5745 142327 5779 142361
rect 6081 142327 6115 142361
rect 6417 142327 6451 142361
rect 6753 142327 6787 142361
rect 7089 142327 7123 142361
rect 7425 142327 7459 142361
rect 7761 142327 7795 142361
rect 8097 142327 8131 142361
rect 8433 142327 8467 142361
rect 8769 142327 8803 142361
rect 9105 142327 9139 142361
rect 9441 142327 9475 142361
rect 9777 142327 9811 142361
rect 10113 142327 10147 142361
rect 10449 142327 10483 142361
rect 10785 142327 10819 142361
rect 11121 142327 11155 142361
rect 11457 142327 11491 142361
rect 11793 142327 11827 142361
rect 12129 142327 12163 142361
rect 12465 142327 12499 142361
rect 12801 142327 12835 142361
rect 13137 142327 13171 142361
rect 13473 142327 13507 142361
rect 13809 142327 13843 142361
rect 14145 142327 14179 142361
rect 14481 142327 14515 142361
rect 14817 142327 14851 142361
rect 15153 142327 15187 142361
rect 15489 142327 15523 142361
rect 15825 142327 15859 142361
rect 16161 142327 16195 142361
rect 16497 142327 16531 142361
rect 16833 142327 16867 142361
rect 17169 142327 17203 142361
rect 17505 142327 17539 142361
rect 17841 142327 17875 142361
rect 18177 142327 18211 142361
rect 18513 142327 18547 142361
rect 18849 142327 18883 142361
rect 19185 142327 19219 142361
rect 19521 142327 19555 142361
rect 19857 142327 19891 142361
rect 20193 142327 20227 142361
rect 20529 142327 20563 142361
rect 20865 142327 20899 142361
rect 21201 142327 21235 142361
rect 21537 142327 21571 142361
rect 21873 142327 21907 142361
rect 22209 142327 22243 142361
rect 22545 142327 22579 142361
rect 22881 142327 22915 142361
rect 23217 142327 23251 142361
rect 23553 142327 23587 142361
rect 23889 142327 23923 142361
rect 24225 142327 24259 142361
rect 24561 142327 24595 142361
rect 24897 142327 24931 142361
rect 25233 142327 25267 142361
rect 25569 142327 25603 142361
rect 25905 142327 25939 142361
rect 26241 142327 26275 142361
rect 26577 142327 26611 142361
rect 26913 142327 26947 142361
rect 27249 142327 27283 142361
rect 27585 142327 27619 142361
rect 27921 142327 27955 142361
rect 28257 142327 28291 142361
rect 28593 142327 28627 142361
rect 28929 142327 28963 142361
rect 29265 142327 29299 142361
rect 29601 142327 29635 142361
rect 29937 142327 29971 142361
rect 30273 142327 30307 142361
rect 30609 142327 30643 142361
rect 30945 142327 30979 142361
rect 31281 142327 31315 142361
rect 31617 142327 31651 142361
rect 31953 142327 31987 142361
rect 32289 142327 32323 142361
rect 32625 142327 32659 142361
rect 32961 142327 32995 142361
rect 33297 142327 33331 142361
rect 33633 142327 33667 142361
rect 33969 142327 34003 142361
rect 34305 142327 34339 142361
rect 34641 142327 34675 142361
rect 34977 142327 35011 142361
rect 35313 142327 35347 142361
rect 35649 142327 35683 142361
rect 35985 142327 36019 142361
rect 36321 142327 36355 142361
rect 36657 142327 36691 142361
rect 36993 142327 37027 142361
rect 37329 142327 37363 142361
rect 37665 142327 37699 142361
rect 38001 142327 38035 142361
rect 38337 142327 38371 142361
rect 38673 142327 38707 142361
rect 39009 142327 39043 142361
rect 39345 142327 39379 142361
rect 39681 142327 39715 142361
rect 40017 142327 40051 142361
rect 40353 142327 40387 142361
rect 40689 142327 40723 142361
rect 41025 142327 41059 142361
rect 41361 142327 41395 142361
rect 41697 142327 41731 142361
rect 42033 142327 42067 142361
rect 42369 142327 42403 142361
rect 42705 142327 42739 142361
rect 43041 142327 43075 142361
rect 43377 142327 43411 142361
rect 43713 142327 43747 142361
rect 44049 142327 44083 142361
rect 44385 142327 44419 142361
rect 44721 142327 44755 142361
rect 45057 142327 45091 142361
rect 45393 142327 45427 142361
rect 45729 142327 45763 142361
rect 46065 142327 46099 142361
rect 46401 142327 46435 142361
rect 46737 142327 46771 142361
rect 47073 142327 47107 142361
rect 47409 142327 47443 142361
rect 47745 142327 47779 142361
rect 48081 142327 48115 142361
rect 48417 142327 48451 142361
rect 48753 142327 48787 142361
rect 49089 142327 49123 142361
rect 49425 142327 49459 142361
rect 49761 142327 49795 142361
rect 50097 142327 50131 142361
rect 50433 142327 50467 142361
rect 50769 142327 50803 142361
rect 51105 142327 51139 142361
rect 51441 142327 51475 142361
rect 51777 142327 51811 142361
rect 52113 142327 52147 142361
rect 52449 142327 52483 142361
rect 52785 142327 52819 142361
rect 53121 142327 53155 142361
rect 53457 142327 53491 142361
rect 53793 142327 53827 142361
rect 54129 142327 54163 142361
rect 54465 142327 54499 142361
rect 54801 142327 54835 142361
rect 55137 142327 55171 142361
rect 55473 142327 55507 142361
rect 55809 142327 55843 142361
rect 56145 142327 56179 142361
rect 56481 142327 56515 142361
rect 56817 142327 56851 142361
rect 57153 142327 57187 142361
rect 57489 142327 57523 142361
rect 57825 142327 57859 142361
rect 58161 142327 58195 142361
rect 58497 142327 58531 142361
rect 58833 142327 58867 142361
rect 59169 142327 59203 142361
rect 59505 142327 59539 142361
rect 59841 142327 59875 142361
rect 60177 142327 60211 142361
rect 60513 142327 60547 142361
rect 60849 142327 60883 142361
rect 61185 142327 61219 142361
rect 61521 142327 61555 142361
rect 61857 142327 61891 142361
rect 62193 142327 62227 142361
rect 62529 142327 62563 142361
rect 62865 142327 62899 142361
rect 63201 142327 63235 142361
rect 63537 142327 63571 142361
rect 63873 142327 63907 142361
rect 64209 142327 64243 142361
rect 64545 142327 64579 142361
rect 64881 142327 64915 142361
rect 65217 142327 65251 142361
rect 65553 142327 65587 142361
rect 65889 142327 65923 142361
rect 66225 142327 66259 142361
rect 66561 142327 66595 142361
rect 66897 142327 66931 142361
rect 67233 142327 67267 142361
rect 67569 142327 67603 142361
rect 67905 142327 67939 142361
rect 68241 142327 68275 142361
rect 68577 142327 68611 142361
rect 68913 142327 68947 142361
rect 69249 142327 69283 142361
rect 69585 142327 69619 142361
rect 69921 142327 69955 142361
rect 70257 142327 70291 142361
rect 70593 142327 70627 142361
rect 70929 142327 70963 142361
rect 71265 142327 71299 142361
rect 71601 142327 71635 142361
rect 71937 142327 71971 142361
rect 72273 142327 72307 142361
rect 72609 142327 72643 142361
rect 72945 142327 72979 142361
rect 73281 142327 73315 142361
rect 73617 142327 73651 142361
rect 73953 142327 73987 142361
rect 74289 142327 74323 142361
rect 74625 142327 74659 142361
rect 74961 142327 74995 142361
rect 75297 142327 75331 142361
rect 75633 142327 75667 142361
rect 75969 142327 76003 142361
rect 76305 142327 76339 142361
rect 76641 142327 76675 142361
rect 76977 142327 77011 142361
rect 77313 142327 77347 142361
rect 77649 142327 77683 142361
rect 77985 142327 78019 142361
rect 78321 142327 78355 142361
rect 78657 142327 78691 142361
rect 78993 142327 79027 142361
rect 79329 142327 79363 142361
rect 79665 142327 79699 142361
rect 80001 142327 80035 142361
rect 80337 142327 80371 142361
rect 80673 142327 80707 142361
rect 81009 142327 81043 142361
rect 81345 142327 81379 142361
rect 81681 142327 81715 142361
rect 82017 142327 82051 142361
rect 82353 142327 82387 142361
rect 82689 142327 82723 142361
rect 83025 142327 83059 142361
rect 83361 142327 83395 142361
rect 83697 142327 83731 142361
rect 84033 142327 84067 142361
rect 84369 142327 84403 142361
rect 84705 142327 84739 142361
rect 85041 142327 85075 142361
rect 85377 142327 85411 142361
rect 85713 142327 85747 142361
rect 86049 142327 86083 142361
rect 86385 142327 86419 142361
rect 86721 142327 86755 142361
rect 87057 142327 87091 142361
rect 87393 142327 87427 142361
rect 87729 142327 87763 142361
rect 88065 142327 88099 142361
rect 88401 142327 88435 142361
rect 88737 142327 88771 142361
rect 89073 142327 89107 142361
rect 89409 142327 89443 142361
rect 89745 142327 89779 142361
rect 90081 142327 90115 142361
rect 90417 142327 90451 142361
rect 90753 142327 90787 142361
rect 91089 142327 91123 142361
rect 91425 142327 91459 142361
rect 91761 142327 91795 142361
rect 92097 142327 92131 142361
rect 92433 142327 92467 142361
rect 92769 142327 92803 142361
rect 93105 142327 93139 142361
rect 93441 142327 93475 142361
rect 93777 142327 93811 142361
rect 94113 142327 94147 142361
rect 94449 142327 94483 142361
rect 94785 142327 94819 142361
rect 95121 142327 95155 142361
rect 95457 142327 95491 142361
rect 95793 142327 95827 142361
rect 96129 142327 96163 142361
rect 96465 142327 96499 142361
rect 96801 142327 96835 142361
rect 97137 142327 97171 142361
rect 97473 142327 97507 142361
rect 97809 142327 97843 142361
rect 98145 142327 98179 142361
rect 98481 142327 98515 142361
rect 98817 142327 98851 142361
rect 99153 142327 99187 142361
rect 99489 142327 99523 142361
rect 99825 142327 99859 142361
rect 100161 142327 100195 142361
rect 100497 142327 100531 142361
rect 100833 142327 100867 142361
rect 101169 142327 101203 142361
rect 101505 142327 101539 142361
rect 101841 142327 101875 142361
rect 102177 142327 102211 142361
rect 102513 142327 102547 142361
rect 102849 142327 102883 142361
rect 103185 142327 103219 142361
rect 103521 142327 103555 142361
rect 103857 142327 103891 142361
rect 104193 142327 104227 142361
rect 104529 142327 104563 142361
rect 104865 142327 104899 142361
rect 105201 142327 105235 142361
rect 105537 142327 105571 142361
rect 105873 142327 105907 142361
rect 106209 142327 106243 142361
rect 106545 142327 106579 142361
rect 106881 142327 106915 142361
rect 107217 142327 107251 142361
rect 107553 142327 107587 142361
rect 107889 142327 107923 142361
rect 108225 142327 108259 142361
rect 108561 142327 108595 142361
rect 108897 142327 108931 142361
rect 109233 142327 109267 142361
rect 109569 142327 109603 142361
rect 109905 142327 109939 142361
rect 110241 142327 110275 142361
rect 110577 142327 110611 142361
rect 110913 142327 110947 142361
rect 111249 142327 111283 142361
rect 111585 142327 111619 142361
rect 111921 142327 111955 142361
rect 112257 142327 112291 142361
rect 112593 142327 112627 142361
rect 112929 142327 112963 142361
rect 113265 142327 113299 142361
rect 113601 142327 113635 142361
rect 113937 142327 113971 142361
rect 114273 142327 114307 142361
rect 114609 142327 114643 142361
rect 114945 142327 114979 142361
rect 115281 142327 115315 142361
rect 115617 142327 115651 142361
rect 115953 142327 115987 142361
rect 116289 142327 116323 142361
rect 116625 142327 116659 142361
rect 116961 142327 116995 142361
rect 117297 142327 117331 142361
rect 117633 142327 117667 142361
rect 117969 142327 118003 142361
rect 118305 142327 118339 142361
rect 118641 142327 118675 142361
rect 118977 142327 119011 142361
rect 119313 142327 119347 142361
rect 119649 142327 119683 142361
rect 119985 142327 120019 142361
rect 120321 142327 120355 142361
rect 120657 142327 120691 142361
rect 120993 142327 121027 142361
rect 121329 142327 121363 142361
rect 121665 142327 121699 142361
rect 122001 142327 122035 142361
rect 122337 142327 122371 142361
rect 122673 142327 122707 142361
rect 123009 142327 123043 142361
rect 123345 142327 123379 142361
rect 123681 142327 123715 142361
rect 124017 142327 124051 142361
rect 124353 142327 124387 142361
rect 124689 142327 124723 142361
rect 125025 142327 125059 142361
rect 125361 142327 125395 142361
rect 125697 142327 125731 142361
rect 126033 142327 126067 142361
rect 126369 142327 126403 142361
rect 126705 142327 126739 142361
rect 127041 142327 127075 142361
rect 127377 142327 127411 142361
rect 127713 142327 127747 142361
rect 128049 142327 128083 142361
rect 128385 142327 128419 142361
rect 128721 142327 128755 142361
rect 129057 142327 129091 142361
rect 129393 142327 129427 142361
rect 129729 142327 129763 142361
rect 130065 142327 130099 142361
rect 130401 142327 130435 142361
rect 130737 142327 130771 142361
rect 131073 142327 131107 142361
rect 131409 142327 131443 142361
rect 131745 142327 131779 142361
rect 132081 142327 132115 142361
rect 132417 142327 132451 142361
rect 132753 142327 132787 142361
rect 133089 142327 133123 142361
rect 133425 142327 133459 142361
rect 133761 142327 133795 142361
rect 134097 142327 134131 142361
rect 134433 142327 134467 142361
rect 134769 142327 134803 142361
rect 135105 142327 135139 142361
rect 135441 142327 135475 142361
rect 135777 142327 135811 142361
rect 136113 142327 136147 142361
rect 136449 142327 136483 142361
rect 136785 142327 136819 142361
rect 137121 142327 137155 142361
rect 137457 142327 137491 142361
rect 137793 142327 137827 142361
rect 138129 142327 138163 142361
rect 138465 142327 138499 142361
rect 138801 142327 138835 142361
rect 139137 142327 139171 142361
rect 139473 142327 139507 142361
rect 139809 142327 139843 142361
rect 140145 142327 140179 142361
rect 140481 142327 140515 142361
rect 140817 142327 140851 142361
rect 141153 142327 141187 142361
rect 141489 142327 141523 142361
rect 141825 142327 141859 142361
rect 142161 142327 142195 142361
rect 142497 142327 142531 142361
rect 142833 142327 142867 142361
rect 143169 142327 143203 142361
rect 143505 142327 143539 142361
rect 143841 142327 143875 142361
rect 144177 142327 144211 142361
rect 144513 142327 144547 142361
rect 144849 142327 144883 142361
rect 145185 142327 145219 142361
rect 145521 142327 145555 142361
rect 145857 142327 145891 142361
rect 146193 142327 146227 142361
rect 146529 142327 146563 142361
rect 146865 142327 146899 142361
rect 147201 142327 147235 142361
rect 147537 142327 147571 142361
rect 147873 142327 147907 142361
rect 148209 142327 148243 142361
rect 148545 142327 148579 142361
rect 148881 142327 148915 142361
rect 149217 142327 149251 142361
rect 149553 142327 149587 142361
rect 149889 142327 149923 142361
rect 150225 142327 150259 142361
rect 150561 142327 150595 142361
rect 150897 142327 150931 142361
rect 151233 142327 151267 142361
rect 151569 142327 151603 142361
rect 151905 142327 151939 142361
rect 152241 142327 152275 142361
rect 152577 142327 152611 142361
rect 152913 142327 152947 142361
rect 153249 142327 153283 142361
rect 153585 142327 153619 142361
rect 153921 142327 153955 142361
rect 154257 142327 154291 142361
rect 154593 142327 154627 142361
rect 154929 142327 154963 142361
rect 155265 142327 155299 142361
rect 155601 142327 155635 142361
rect 155937 142327 155971 142361
rect 156273 142327 156307 142361
rect 156609 142327 156643 142361
rect 156945 142327 156979 142361
rect 157281 142327 157315 142361
rect 157617 142327 157651 142361
rect 157953 142327 157987 142361
rect 158289 142327 158323 142361
rect 158625 142327 158659 142361
rect 158961 142327 158995 142361
rect 159297 142327 159331 142361
rect 159633 142327 159667 142361
rect 159969 142327 160003 142361
rect 160305 142327 160339 142361
rect 160641 142327 160675 142361
rect 160977 142327 161011 142361
rect 161313 142327 161347 142361
rect 161649 142327 161683 142361
rect 161985 142327 162019 142361
rect 162321 142327 162355 142361
rect 162657 142327 162691 142361
rect 162993 142327 163027 142361
rect 163329 142327 163363 142361
rect 163665 142327 163699 142361
rect 164001 142327 164035 142361
rect 164337 142327 164371 142361
rect 164673 142327 164707 142361
rect 165009 142327 165043 142361
rect 165345 142327 165379 142361
rect 165681 142327 165715 142361
rect 166017 142327 166051 142361
rect 166353 142327 166387 142361
rect 166689 142327 166723 142361
rect 167025 142327 167059 142361
rect 167361 142327 167395 142361
rect 167697 142327 167731 142361
rect 168033 142327 168067 142361
rect 168369 142327 168403 142361
rect 168705 142327 168739 142361
rect 169041 142327 169075 142361
rect 169377 142327 169411 142361
rect 169713 142327 169747 142361
rect 170049 142327 170083 142361
rect 170385 142327 170419 142361
rect 170721 142327 170755 142361
rect 171057 142327 171091 142361
rect 171393 142327 171427 142361
rect 171729 142327 171763 142361
rect 172065 142327 172099 142361
rect 172401 142327 172435 142361
rect 172737 142327 172771 142361
rect 173073 142327 173107 142361
rect 173409 142327 173443 142361
rect 173745 142327 173779 142361
rect 174081 142327 174115 142361
rect 174417 142327 174451 142361
rect 174753 142327 174787 142361
rect 175089 142327 175123 142361
rect 175425 142327 175459 142361
rect 175761 142327 175795 142361
rect 176097 142327 176131 142361
rect 176433 142327 176467 142361
rect 176769 142327 176803 142361
rect 177105 142327 177139 142361
rect 177441 142327 177475 142361
rect 177777 142327 177811 142361
rect 178113 142327 178147 142361
rect 178449 142327 178483 142361
rect 178785 142327 178819 142361
rect 179121 142327 179155 142361
rect 179457 142327 179491 142361
rect 179793 142327 179827 142361
rect 180129 142327 180163 142361
rect 180465 142327 180499 142361
rect 180801 142327 180835 142361
rect 181137 142327 181171 142361
rect 181473 142327 181507 142361
rect 181809 142327 181843 142361
rect 182145 142327 182179 142361
rect 182481 142327 182515 142361
rect 182817 142327 182851 142361
rect 183153 142327 183187 142361
rect 183489 142327 183523 142361
rect 183825 142327 183859 142361
rect 184161 142327 184195 142361
rect 184497 142327 184531 142361
rect 184833 142327 184867 142361
rect 185169 142327 185203 142361
rect 185505 142327 185539 142361
rect 185841 142327 185875 142361
rect 186177 142327 186211 142361
rect 186513 142327 186547 142361
rect 186849 142327 186883 142361
rect 187185 142327 187219 142361
rect 187521 142327 187555 142361
rect 187857 142327 187891 142361
rect 188193 142327 188227 142361
rect 188529 142327 188563 142361
rect 188865 142327 188899 142361
rect 189201 142327 189235 142361
rect 189537 142327 189571 142361
rect 189873 142327 189907 142361
rect 190209 142327 190243 142361
rect 190545 142327 190579 142361
rect 190881 142327 190915 142361
rect 191217 142327 191251 142361
rect 191553 142327 191587 142361
rect 191889 142327 191923 142361
rect 192225 142327 192259 142361
rect 192561 142327 192595 142361
rect 192897 142327 192931 142361
rect 193233 142327 193267 142361
rect 193569 142327 193603 142361
rect 193905 142327 193939 142361
rect 194241 142327 194275 142361
rect 194577 142327 194611 142361
rect 194913 142327 194947 142361
rect 195249 142327 195283 142361
rect 195585 142327 195619 142361
rect 195921 142327 195955 142361
rect 196257 142327 196291 142361
rect 196593 142327 196627 142361
rect 196929 142327 196963 142361
rect 197265 142327 197299 142361
rect 197601 142327 197635 142361
rect 197937 142327 197971 142361
rect 198273 142327 198307 142361
rect 198609 142327 198643 142361
rect 198945 142327 198979 142361
rect 199281 142327 199315 142361
rect 199617 142327 199651 142361
rect 199953 142327 199987 142361
rect 200289 142327 200323 142361
rect 200625 142327 200659 142361
rect 200961 142327 200995 142361
rect 201297 142327 201331 142361
rect 201633 142327 201667 142361
rect 201969 142327 202003 142361
rect 202305 142327 202339 142361
rect 202641 142327 202675 142361
rect 202977 142327 203011 142361
rect 203313 142327 203347 142361
rect 203649 142327 203683 142361
rect 203985 142327 204019 142361
rect 204321 142327 204355 142361
rect 204657 142327 204691 142361
rect 204993 142327 205027 142361
rect 205329 142327 205363 142361
rect 205665 142327 205699 142361
rect 206001 142327 206035 142361
rect 206337 142327 206371 142361
rect 206673 142327 206707 142361
rect 207009 142327 207043 142361
rect 207345 142327 207379 142361
rect 207681 142327 207715 142361
rect 208017 142327 208051 142361
rect 208353 142327 208387 142361
rect 208689 142327 208723 142361
rect 209025 142327 209059 142361
rect 209361 142327 209395 142361
rect 209697 142327 209731 142361
rect 210033 142327 210067 142361
rect 210369 142327 210403 142361
rect 210705 142327 210739 142361
rect 211041 142327 211075 142361
rect 211377 142327 211411 142361
rect 211713 142327 211747 142361
rect 212049 142327 212083 142361
rect 212385 142327 212419 142361
rect 212721 142327 212755 142361
rect 213057 142327 213091 142361
rect 213393 142327 213427 142361
rect 213729 142327 213763 142361
rect 214065 142327 214099 142361
rect 214401 142327 214435 142361
rect 214737 142327 214771 142361
rect 215073 142327 215107 142361
rect 215409 142327 215443 142361
rect 215745 142327 215779 142361
rect 216081 142327 216115 142361
rect 216417 142327 216451 142361
rect 1713 141943 1747 141977
rect 216919 141943 216953 141977
rect 1713 141607 1747 141641
rect 216919 141607 216953 141641
rect 1713 141271 1747 141305
rect 216919 141271 216953 141305
rect 1713 140935 1747 140969
rect 216919 140935 216953 140969
rect 1713 140599 1747 140633
rect 216919 140599 216953 140633
rect 1713 140263 1747 140297
rect 216919 140263 216953 140297
rect 1713 139927 1747 139961
rect 216919 139927 216953 139961
rect 1713 139591 1747 139625
rect 216919 139591 216953 139625
rect 1713 139255 1747 139289
rect 216919 139255 216953 139289
rect 1713 138919 1747 138953
rect 216919 138919 216953 138953
rect 1713 138583 1747 138617
rect 216919 138583 216953 138617
rect 1713 138247 1747 138281
rect 216919 138247 216953 138281
rect 1713 137911 1747 137945
rect 216919 137911 216953 137945
rect 1713 137575 1747 137609
rect 216919 137575 216953 137609
rect 1713 137239 1747 137273
rect 216919 137239 216953 137273
rect 1713 136903 1747 136937
rect 216919 136903 216953 136937
rect 1713 136567 1747 136601
rect 216919 136567 216953 136601
rect 1713 136231 1747 136265
rect 216919 136231 216953 136265
rect 1713 135895 1747 135929
rect 216919 135895 216953 135929
rect 1713 135559 1747 135593
rect 216919 135559 216953 135593
rect 1713 135223 1747 135257
rect 216919 135223 216953 135257
rect 1713 134887 1747 134921
rect 216919 134887 216953 134921
rect 1713 134551 1747 134585
rect 216919 134551 216953 134585
rect 1713 134215 1747 134249
rect 216919 134215 216953 134249
rect 1713 133879 1747 133913
rect 216919 133879 216953 133913
rect 1713 133543 1747 133577
rect 216919 133543 216953 133577
rect 1713 133207 1747 133241
rect 216919 133207 216953 133241
rect 1713 132871 1747 132905
rect 216919 132871 216953 132905
rect 1713 132535 1747 132569
rect 216919 132535 216953 132569
rect 1713 132199 1747 132233
rect 216919 132199 216953 132233
rect 1713 131863 1747 131897
rect 216919 131863 216953 131897
rect 1713 131527 1747 131561
rect 216919 131527 216953 131561
rect 1713 131191 1747 131225
rect 216919 131191 216953 131225
rect 1713 130855 1747 130889
rect 216919 130855 216953 130889
rect 1713 130519 1747 130553
rect 216919 130519 216953 130553
rect 1713 130183 1747 130217
rect 216919 130183 216953 130217
rect 1713 129847 1747 129881
rect 216919 129847 216953 129881
rect 1713 129511 1747 129545
rect 216919 129511 216953 129545
rect 1713 129175 1747 129209
rect 216919 129175 216953 129209
rect 1713 128839 1747 128873
rect 216919 128839 216953 128873
rect 1713 128503 1747 128537
rect 216919 128503 216953 128537
rect 1713 128167 1747 128201
rect 216919 128167 216953 128201
rect 1713 127831 1747 127865
rect 216919 127831 216953 127865
rect 1713 127495 1747 127529
rect 216919 127495 216953 127529
rect 1713 127159 1747 127193
rect 216919 127159 216953 127193
rect 1713 126823 1747 126857
rect 216919 126823 216953 126857
rect 1713 126487 1747 126521
rect 216919 126487 216953 126521
rect 1713 126151 1747 126185
rect 216919 126151 216953 126185
rect 1713 125815 1747 125849
rect 216919 125815 216953 125849
rect 1713 125479 1747 125513
rect 216919 125479 216953 125513
rect 1713 125143 1747 125177
rect 216919 125143 216953 125177
rect 1713 124807 1747 124841
rect 216919 124807 216953 124841
rect 1713 124471 1747 124505
rect 216919 124471 216953 124505
rect 1713 124135 1747 124169
rect 216919 124135 216953 124169
rect 1713 123799 1747 123833
rect 216919 123799 216953 123833
rect 1713 123463 1747 123497
rect 216919 123463 216953 123497
rect 1713 123127 1747 123161
rect 216919 123127 216953 123161
rect 1713 122791 1747 122825
rect 216919 122791 216953 122825
rect 1713 122455 1747 122489
rect 216919 122455 216953 122489
rect 1713 122119 1747 122153
rect 216919 122119 216953 122153
rect 1713 121783 1747 121817
rect 216919 121783 216953 121817
rect 1713 121447 1747 121481
rect 216919 121447 216953 121481
rect 1713 121111 1747 121145
rect 216919 121111 216953 121145
rect 1713 120775 1747 120809
rect 216919 120775 216953 120809
rect 1713 120439 1747 120473
rect 216919 120439 216953 120473
rect 1713 120103 1747 120137
rect 216919 120103 216953 120137
rect 1713 119767 1747 119801
rect 216919 119767 216953 119801
rect 1713 119431 1747 119465
rect 216919 119431 216953 119465
rect 1713 119095 1747 119129
rect 216919 119095 216953 119129
rect 1713 118759 1747 118793
rect 216919 118759 216953 118793
rect 1713 118423 1747 118457
rect 216919 118423 216953 118457
rect 1713 118087 1747 118121
rect 216919 118087 216953 118121
rect 1713 117751 1747 117785
rect 216919 117751 216953 117785
rect 1713 117415 1747 117449
rect 216919 117415 216953 117449
rect 1713 117079 1747 117113
rect 216919 117079 216953 117113
rect 1713 116743 1747 116777
rect 216919 116743 216953 116777
rect 1713 116407 1747 116441
rect 216919 116407 216953 116441
rect 1713 116071 1747 116105
rect 216919 116071 216953 116105
rect 1713 115735 1747 115769
rect 216919 115735 216953 115769
rect 1713 115399 1747 115433
rect 216919 115399 216953 115433
rect 1713 115063 1747 115097
rect 216919 115063 216953 115097
rect 1713 114727 1747 114761
rect 216919 114727 216953 114761
rect 1713 114391 1747 114425
rect 216919 114391 216953 114425
rect 1713 114055 1747 114089
rect 216919 114055 216953 114089
rect 1713 113719 1747 113753
rect 216919 113719 216953 113753
rect 1713 113383 1747 113417
rect 216919 113383 216953 113417
rect 1713 113047 1747 113081
rect 216919 113047 216953 113081
rect 1713 112711 1747 112745
rect 216919 112711 216953 112745
rect 1713 112375 1747 112409
rect 216919 112375 216953 112409
rect 1713 112039 1747 112073
rect 216919 112039 216953 112073
rect 1713 111703 1747 111737
rect 216919 111703 216953 111737
rect 1713 111367 1747 111401
rect 216919 111367 216953 111401
rect 1713 111031 1747 111065
rect 216919 111031 216953 111065
rect 1713 110695 1747 110729
rect 216919 110695 216953 110729
rect 1713 110359 1747 110393
rect 216919 110359 216953 110393
rect 1713 110023 1747 110057
rect 216919 110023 216953 110057
rect 1713 109687 1747 109721
rect 216919 109687 216953 109721
rect 1713 109351 1747 109385
rect 216919 109351 216953 109385
rect 1713 109015 1747 109049
rect 216919 109015 216953 109049
rect 1713 108679 1747 108713
rect 216919 108679 216953 108713
rect 1713 108343 1747 108377
rect 216919 108343 216953 108377
rect 1713 108007 1747 108041
rect 216919 108007 216953 108041
rect 1713 107671 1747 107705
rect 216919 107671 216953 107705
rect 1713 107335 1747 107369
rect 216919 107335 216953 107369
rect 1713 106999 1747 107033
rect 216919 106999 216953 107033
rect 1713 106663 1747 106697
rect 216919 106663 216953 106697
rect 1713 106327 1747 106361
rect 216919 106327 216953 106361
rect 1713 105991 1747 106025
rect 216919 105991 216953 106025
rect 1713 105655 1747 105689
rect 216919 105655 216953 105689
rect 1713 105319 1747 105353
rect 216919 105319 216953 105353
rect 1713 104983 1747 105017
rect 216919 104983 216953 105017
rect 1713 104647 1747 104681
rect 216919 104647 216953 104681
rect 1713 104311 1747 104345
rect 216919 104311 216953 104345
rect 1713 103975 1747 104009
rect 216919 103975 216953 104009
rect 1713 103639 1747 103673
rect 216919 103639 216953 103673
rect 1713 103303 1747 103337
rect 216919 103303 216953 103337
rect 1713 102967 1747 103001
rect 216919 102967 216953 103001
rect 1713 102631 1747 102665
rect 216919 102631 216953 102665
rect 1713 102295 1747 102329
rect 216919 102295 216953 102329
rect 1713 101959 1747 101993
rect 216919 101959 216953 101993
rect 1713 101623 1747 101657
rect 216919 101623 216953 101657
rect 1713 101287 1747 101321
rect 216919 101287 216953 101321
rect 1713 100951 1747 100985
rect 216919 100951 216953 100985
rect 1713 100615 1747 100649
rect 216919 100615 216953 100649
rect 1713 100279 1747 100313
rect 216919 100279 216953 100313
rect 1713 99943 1747 99977
rect 216919 99943 216953 99977
rect 1713 99607 1747 99641
rect 216919 99607 216953 99641
rect 1713 99271 1747 99305
rect 216919 99271 216953 99305
rect 1713 98935 1747 98969
rect 216919 98935 216953 98969
rect 1713 98599 1747 98633
rect 216919 98599 216953 98633
rect 1713 98263 1747 98297
rect 216919 98263 216953 98297
rect 1713 97927 1747 97961
rect 216919 97927 216953 97961
rect 1713 97591 1747 97625
rect 216919 97591 216953 97625
rect 1713 97255 1747 97289
rect 216919 97255 216953 97289
rect 1713 96919 1747 96953
rect 216919 96919 216953 96953
rect 1713 96583 1747 96617
rect 216919 96583 216953 96617
rect 1713 96247 1747 96281
rect 216919 96247 216953 96281
rect 1713 95911 1747 95945
rect 216919 95911 216953 95945
rect 1713 95575 1747 95609
rect 216919 95575 216953 95609
rect 1713 95239 1747 95273
rect 216919 95239 216953 95273
rect 1713 94903 1747 94937
rect 216919 94903 216953 94937
rect 1713 94567 1747 94601
rect 216919 94567 216953 94601
rect 1713 94231 1747 94265
rect 216919 94231 216953 94265
rect 1713 93895 1747 93929
rect 216919 93895 216953 93929
rect 1713 93559 1747 93593
rect 216919 93559 216953 93593
rect 1713 93223 1747 93257
rect 216919 93223 216953 93257
rect 1713 92887 1747 92921
rect 216919 92887 216953 92921
rect 1713 92551 1747 92585
rect 216919 92551 216953 92585
rect 1713 92215 1747 92249
rect 216919 92215 216953 92249
rect 1713 91879 1747 91913
rect 216919 91879 216953 91913
rect 1713 91543 1747 91577
rect 216919 91543 216953 91577
rect 1713 91207 1747 91241
rect 216919 91207 216953 91241
rect 1713 90871 1747 90905
rect 216919 90871 216953 90905
rect 1713 90535 1747 90569
rect 216919 90535 216953 90569
rect 1713 90199 1747 90233
rect 216919 90199 216953 90233
rect 1713 89863 1747 89897
rect 216919 89863 216953 89897
rect 1713 89527 1747 89561
rect 216919 89527 216953 89561
rect 1713 89191 1747 89225
rect 216919 89191 216953 89225
rect 1713 88855 1747 88889
rect 216919 88855 216953 88889
rect 1713 88519 1747 88553
rect 216919 88519 216953 88553
rect 1713 88183 1747 88217
rect 216919 88183 216953 88217
rect 1713 87847 1747 87881
rect 216919 87847 216953 87881
rect 1713 87511 1747 87545
rect 216919 87511 216953 87545
rect 1713 87175 1747 87209
rect 216919 87175 216953 87209
rect 1713 86839 1747 86873
rect 216919 86839 216953 86873
rect 1713 86503 1747 86537
rect 216919 86503 216953 86537
rect 1713 86167 1747 86201
rect 216919 86167 216953 86201
rect 1713 85831 1747 85865
rect 216919 85831 216953 85865
rect 1713 85495 1747 85529
rect 216919 85495 216953 85529
rect 1713 85159 1747 85193
rect 216919 85159 216953 85193
rect 1713 84823 1747 84857
rect 216919 84823 216953 84857
rect 1713 84487 1747 84521
rect 216919 84487 216953 84521
rect 1713 84151 1747 84185
rect 216919 84151 216953 84185
rect 1713 83815 1747 83849
rect 216919 83815 216953 83849
rect 1713 83479 1747 83513
rect 216919 83479 216953 83513
rect 1713 83143 1747 83177
rect 216919 83143 216953 83177
rect 1713 82807 1747 82841
rect 216919 82807 216953 82841
rect 1713 82471 1747 82505
rect 216919 82471 216953 82505
rect 1713 82135 1747 82169
rect 216919 82135 216953 82169
rect 1713 81799 1747 81833
rect 216919 81799 216953 81833
rect 1713 81463 1747 81497
rect 216919 81463 216953 81497
rect 1713 81127 1747 81161
rect 216919 81127 216953 81161
rect 1713 80791 1747 80825
rect 216919 80791 216953 80825
rect 1713 80455 1747 80489
rect 216919 80455 216953 80489
rect 1713 80119 1747 80153
rect 216919 80119 216953 80153
rect 1713 79783 1747 79817
rect 216919 79783 216953 79817
rect 1713 79447 1747 79481
rect 216919 79447 216953 79481
rect 1713 79111 1747 79145
rect 216919 79111 216953 79145
rect 1713 78775 1747 78809
rect 216919 78775 216953 78809
rect 1713 78439 1747 78473
rect 216919 78439 216953 78473
rect 1713 78103 1747 78137
rect 216919 78103 216953 78137
rect 1713 77767 1747 77801
rect 216919 77767 216953 77801
rect 1713 77431 1747 77465
rect 216919 77431 216953 77465
rect 1713 77095 1747 77129
rect 216919 77095 216953 77129
rect 1713 76759 1747 76793
rect 216919 76759 216953 76793
rect 1713 76423 1747 76457
rect 216919 76423 216953 76457
rect 1713 76087 1747 76121
rect 216919 76087 216953 76121
rect 1713 75751 1747 75785
rect 216919 75751 216953 75785
rect 1713 75415 1747 75449
rect 216919 75415 216953 75449
rect 1713 75079 1747 75113
rect 216919 75079 216953 75113
rect 1713 74743 1747 74777
rect 216919 74743 216953 74777
rect 1713 74407 1747 74441
rect 216919 74407 216953 74441
rect 1713 74071 1747 74105
rect 216919 74071 216953 74105
rect 1713 73735 1747 73769
rect 216919 73735 216953 73769
rect 1713 73399 1747 73433
rect 216919 73399 216953 73433
rect 1713 73063 1747 73097
rect 216919 73063 216953 73097
rect 1713 72727 1747 72761
rect 216919 72727 216953 72761
rect 1713 72391 1747 72425
rect 216919 72391 216953 72425
rect 1713 72055 1747 72089
rect 216919 72055 216953 72089
rect 1713 71719 1747 71753
rect 216919 71719 216953 71753
rect 1713 71383 1747 71417
rect 216919 71383 216953 71417
rect 1713 71047 1747 71081
rect 216919 71047 216953 71081
rect 1713 70711 1747 70745
rect 216919 70711 216953 70745
rect 1713 70375 1747 70409
rect 216919 70375 216953 70409
rect 1713 70039 1747 70073
rect 216919 70039 216953 70073
rect 1713 69703 1747 69737
rect 216919 69703 216953 69737
rect 1713 69367 1747 69401
rect 216919 69367 216953 69401
rect 1713 69031 1747 69065
rect 216919 69031 216953 69065
rect 1713 68695 1747 68729
rect 216919 68695 216953 68729
rect 1713 68359 1747 68393
rect 216919 68359 216953 68393
rect 1713 68023 1747 68057
rect 216919 68023 216953 68057
rect 1713 67687 1747 67721
rect 216919 67687 216953 67721
rect 1713 67351 1747 67385
rect 216919 67351 216953 67385
rect 1713 67015 1747 67049
rect 216919 67015 216953 67049
rect 1713 66679 1747 66713
rect 216919 66679 216953 66713
rect 1713 66343 1747 66377
rect 216919 66343 216953 66377
rect 1713 66007 1747 66041
rect 216919 66007 216953 66041
rect 1713 65671 1747 65705
rect 216919 65671 216953 65705
rect 1713 65335 1747 65369
rect 216919 65335 216953 65369
rect 1713 64999 1747 65033
rect 216919 64999 216953 65033
rect 1713 64663 1747 64697
rect 216919 64663 216953 64697
rect 1713 64327 1747 64361
rect 216919 64327 216953 64361
rect 1713 63991 1747 64025
rect 216919 63991 216953 64025
rect 1713 63655 1747 63689
rect 216919 63655 216953 63689
rect 1713 63319 1747 63353
rect 216919 63319 216953 63353
rect 1713 62983 1747 63017
rect 216919 62983 216953 63017
rect 1713 62647 1747 62681
rect 216919 62647 216953 62681
rect 1713 62311 1747 62345
rect 216919 62311 216953 62345
rect 1713 61975 1747 62009
rect 216919 61975 216953 62009
rect 1713 61639 1747 61673
rect 216919 61639 216953 61673
rect 1713 61303 1747 61337
rect 216919 61303 216953 61337
rect 1713 60967 1747 61001
rect 216919 60967 216953 61001
rect 1713 60631 1747 60665
rect 216919 60631 216953 60665
rect 1713 60295 1747 60329
rect 216919 60295 216953 60329
rect 1713 59959 1747 59993
rect 216919 59959 216953 59993
rect 1713 59623 1747 59657
rect 216919 59623 216953 59657
rect 1713 59287 1747 59321
rect 216919 59287 216953 59321
rect 1713 58951 1747 58985
rect 216919 58951 216953 58985
rect 1713 58615 1747 58649
rect 216919 58615 216953 58649
rect 1713 58279 1747 58313
rect 216919 58279 216953 58313
rect 1713 57943 1747 57977
rect 216919 57943 216953 57977
rect 1713 57607 1747 57641
rect 216919 57607 216953 57641
rect 1713 57271 1747 57305
rect 216919 57271 216953 57305
rect 1713 56935 1747 56969
rect 216919 56935 216953 56969
rect 1713 56599 1747 56633
rect 216919 56599 216953 56633
rect 1713 56263 1747 56297
rect 216919 56263 216953 56297
rect 1713 55927 1747 55961
rect 216919 55927 216953 55961
rect 1713 55591 1747 55625
rect 216919 55591 216953 55625
rect 1713 55255 1747 55289
rect 216919 55255 216953 55289
rect 1713 54919 1747 54953
rect 216919 54919 216953 54953
rect 1713 54583 1747 54617
rect 216919 54583 216953 54617
rect 1713 54247 1747 54281
rect 216919 54247 216953 54281
rect 1713 53911 1747 53945
rect 216919 53911 216953 53945
rect 1713 53575 1747 53609
rect 216919 53575 216953 53609
rect 1713 53239 1747 53273
rect 216919 53239 216953 53273
rect 1713 52903 1747 52937
rect 216919 52903 216953 52937
rect 1713 52567 1747 52601
rect 216919 52567 216953 52601
rect 1713 52231 1747 52265
rect 216919 52231 216953 52265
rect 1713 51895 1747 51929
rect 216919 51895 216953 51929
rect 1713 51559 1747 51593
rect 216919 51559 216953 51593
rect 1713 51223 1747 51257
rect 216919 51223 216953 51257
rect 1713 50887 1747 50921
rect 216919 50887 216953 50921
rect 1713 50551 1747 50585
rect 216919 50551 216953 50585
rect 1713 50215 1747 50249
rect 216919 50215 216953 50249
rect 1713 49879 1747 49913
rect 216919 49879 216953 49913
rect 1713 49543 1747 49577
rect 216919 49543 216953 49577
rect 1713 49207 1747 49241
rect 216919 49207 216953 49241
rect 1713 48871 1747 48905
rect 216919 48871 216953 48905
rect 1713 48535 1747 48569
rect 216919 48535 216953 48569
rect 1713 48199 1747 48233
rect 216919 48199 216953 48233
rect 1713 47863 1747 47897
rect 216919 47863 216953 47897
rect 1713 47527 1747 47561
rect 216919 47527 216953 47561
rect 1713 47191 1747 47225
rect 216919 47191 216953 47225
rect 1713 46855 1747 46889
rect 216919 46855 216953 46889
rect 1713 46519 1747 46553
rect 216919 46519 216953 46553
rect 1713 46183 1747 46217
rect 216919 46183 216953 46217
rect 1713 45847 1747 45881
rect 216919 45847 216953 45881
rect 1713 45511 1747 45545
rect 216919 45511 216953 45545
rect 1713 45175 1747 45209
rect 216919 45175 216953 45209
rect 1713 44839 1747 44873
rect 216919 44839 216953 44873
rect 1713 44503 1747 44537
rect 216919 44503 216953 44537
rect 1713 44167 1747 44201
rect 216919 44167 216953 44201
rect 1713 43831 1747 43865
rect 216919 43831 216953 43865
rect 1713 43495 1747 43529
rect 216919 43495 216953 43529
rect 1713 43159 1747 43193
rect 216919 43159 216953 43193
rect 1713 42823 1747 42857
rect 216919 42823 216953 42857
rect 1713 42487 1747 42521
rect 216919 42487 216953 42521
rect 1713 42151 1747 42185
rect 216919 42151 216953 42185
rect 1713 41815 1747 41849
rect 216919 41815 216953 41849
rect 1713 41479 1747 41513
rect 216919 41479 216953 41513
rect 1713 41143 1747 41177
rect 216919 41143 216953 41177
rect 1713 40807 1747 40841
rect 216919 40807 216953 40841
rect 1713 40471 1747 40505
rect 216919 40471 216953 40505
rect 1713 40135 1747 40169
rect 216919 40135 216953 40169
rect 1713 39799 1747 39833
rect 216919 39799 216953 39833
rect 1713 39463 1747 39497
rect 216919 39463 216953 39497
rect 1713 39127 1747 39161
rect 216919 39127 216953 39161
rect 1713 38791 1747 38825
rect 216919 38791 216953 38825
rect 1713 38455 1747 38489
rect 216919 38455 216953 38489
rect 1713 38119 1747 38153
rect 216919 38119 216953 38153
rect 1713 37783 1747 37817
rect 216919 37783 216953 37817
rect 1713 37447 1747 37481
rect 216919 37447 216953 37481
rect 1713 37111 1747 37145
rect 216919 37111 216953 37145
rect 1713 36775 1747 36809
rect 216919 36775 216953 36809
rect 1713 36439 1747 36473
rect 216919 36439 216953 36473
rect 1713 36103 1747 36137
rect 216919 36103 216953 36137
rect 1713 35767 1747 35801
rect 216919 35767 216953 35801
rect 1713 35431 1747 35465
rect 216919 35431 216953 35465
rect 1713 35095 1747 35129
rect 216919 35095 216953 35129
rect 1713 34759 1747 34793
rect 216919 34759 216953 34793
rect 1713 34423 1747 34457
rect 216919 34423 216953 34457
rect 1713 34087 1747 34121
rect 216919 34087 216953 34121
rect 1713 33751 1747 33785
rect 216919 33751 216953 33785
rect 1713 33415 1747 33449
rect 216919 33415 216953 33449
rect 1713 33079 1747 33113
rect 216919 33079 216953 33113
rect 1713 32743 1747 32777
rect 216919 32743 216953 32777
rect 1713 32407 1747 32441
rect 216919 32407 216953 32441
rect 1713 32071 1747 32105
rect 216919 32071 216953 32105
rect 1713 31735 1747 31769
rect 216919 31735 216953 31769
rect 1713 31399 1747 31433
rect 216919 31399 216953 31433
rect 1713 31063 1747 31097
rect 216919 31063 216953 31097
rect 1713 30727 1747 30761
rect 216919 30727 216953 30761
rect 1713 30391 1747 30425
rect 216919 30391 216953 30425
rect 1713 30055 1747 30089
rect 216919 30055 216953 30089
rect 1713 29719 1747 29753
rect 216919 29719 216953 29753
rect 1713 29383 1747 29417
rect 216919 29383 216953 29417
rect 1713 29047 1747 29081
rect 216919 29047 216953 29081
rect 1713 28711 1747 28745
rect 216919 28711 216953 28745
rect 1713 28375 1747 28409
rect 216919 28375 216953 28409
rect 1713 28039 1747 28073
rect 216919 28039 216953 28073
rect 1713 27703 1747 27737
rect 216919 27703 216953 27737
rect 1713 27367 1747 27401
rect 216919 27367 216953 27401
rect 1713 27031 1747 27065
rect 216919 27031 216953 27065
rect 1713 26695 1747 26729
rect 216919 26695 216953 26729
rect 1713 26359 1747 26393
rect 216919 26359 216953 26393
rect 1713 26023 1747 26057
rect 216919 26023 216953 26057
rect 1713 25687 1747 25721
rect 216919 25687 216953 25721
rect 1713 25351 1747 25385
rect 216919 25351 216953 25385
rect 1713 25015 1747 25049
rect 216919 25015 216953 25049
rect 1713 24679 1747 24713
rect 216919 24679 216953 24713
rect 1713 24343 1747 24377
rect 216919 24343 216953 24377
rect 1713 24007 1747 24041
rect 216919 24007 216953 24041
rect 1713 23671 1747 23705
rect 216919 23671 216953 23705
rect 1713 23335 1747 23369
rect 216919 23335 216953 23369
rect 1713 22999 1747 23033
rect 216919 22999 216953 23033
rect 1713 22663 1747 22697
rect 216919 22663 216953 22697
rect 1713 22327 1747 22361
rect 216919 22327 216953 22361
rect 1713 21991 1747 22025
rect 216919 21991 216953 22025
rect 1713 21655 1747 21689
rect 216919 21655 216953 21689
rect 1713 21319 1747 21353
rect 216919 21319 216953 21353
rect 1713 20983 1747 21017
rect 216919 20983 216953 21017
rect 1713 20647 1747 20681
rect 216919 20647 216953 20681
rect 1713 20311 1747 20345
rect 216919 20311 216953 20345
rect 1713 19975 1747 20009
rect 216919 19975 216953 20009
rect 1713 19639 1747 19673
rect 216919 19639 216953 19673
rect 1713 19303 1747 19337
rect 216919 19303 216953 19337
rect 1713 18967 1747 19001
rect 216919 18967 216953 19001
rect 1713 18631 1747 18665
rect 216919 18631 216953 18665
rect 1713 18295 1747 18329
rect 216919 18295 216953 18329
rect 1713 17959 1747 17993
rect 216919 17959 216953 17993
rect 1713 17623 1747 17657
rect 216919 17623 216953 17657
rect 1713 17287 1747 17321
rect 216919 17287 216953 17321
rect 1713 16951 1747 16985
rect 216919 16951 216953 16985
rect 1713 16615 1747 16649
rect 216919 16615 216953 16649
rect 1713 16279 1747 16313
rect 216919 16279 216953 16313
rect 1713 15943 1747 15977
rect 216919 15943 216953 15977
rect 1713 15607 1747 15641
rect 216919 15607 216953 15641
rect 1713 15271 1747 15305
rect 216919 15271 216953 15305
rect 1713 14935 1747 14969
rect 216919 14935 216953 14969
rect 1713 14599 1747 14633
rect 216919 14599 216953 14633
rect 1713 14263 1747 14297
rect 216919 14263 216953 14297
rect 1713 13927 1747 13961
rect 216919 13927 216953 13961
rect 1713 13591 1747 13625
rect 216919 13591 216953 13625
rect 1713 13255 1747 13289
rect 216919 13255 216953 13289
rect 1713 12919 1747 12953
rect 216919 12919 216953 12953
rect 1713 12583 1747 12617
rect 216919 12583 216953 12617
rect 1713 12247 1747 12281
rect 216919 12247 216953 12281
rect 1713 11911 1747 11945
rect 216919 11911 216953 11945
rect 1713 11575 1747 11609
rect 216919 11575 216953 11609
rect 1713 11239 1747 11273
rect 216919 11239 216953 11273
rect 1713 10903 1747 10937
rect 216919 10903 216953 10937
rect 1713 10567 1747 10601
rect 216919 10567 216953 10601
rect 1713 10231 1747 10265
rect 216919 10231 216953 10265
rect 1713 9895 1747 9929
rect 216919 9895 216953 9929
rect 1713 9559 1747 9593
rect 216919 9559 216953 9593
rect 1713 9223 1747 9257
rect 216919 9223 216953 9257
rect 1713 8887 1747 8921
rect 216919 8887 216953 8921
rect 1713 8551 1747 8585
rect 216919 8551 216953 8585
rect 1713 8215 1747 8249
rect 216919 8215 216953 8249
rect 1713 7879 1747 7913
rect 216919 7879 216953 7913
rect 1713 7543 1747 7577
rect 216919 7543 216953 7577
rect 1713 7207 1747 7241
rect 216919 7207 216953 7241
rect 1713 6871 1747 6905
rect 216919 6871 216953 6905
rect 1713 6535 1747 6569
rect 216919 6535 216953 6569
rect 1713 6199 1747 6233
rect 216919 6199 216953 6233
rect 1713 5863 1747 5897
rect 216919 5863 216953 5897
rect 1713 5527 1747 5561
rect 216919 5527 216953 5561
rect 1713 5191 1747 5225
rect 216919 5191 216953 5225
rect 1713 4855 1747 4889
rect 216919 4855 216953 4889
rect 1713 4519 1747 4553
rect 216919 4519 216953 4553
rect 1713 4183 1747 4217
rect 216919 4183 216953 4217
rect 1713 3847 1747 3881
rect 216919 3847 216953 3881
rect 1713 3511 1747 3545
rect 216919 3511 216953 3545
rect 1713 3175 1747 3209
rect 216919 3175 216953 3209
rect 1713 2839 1747 2873
rect 216919 2839 216953 2873
rect 1713 2503 1747 2537
rect 216919 2503 216953 2537
rect 1713 2167 1747 2201
rect 216919 2167 216953 2201
rect 2049 1831 2083 1865
rect 2385 1831 2419 1865
rect 2721 1831 2755 1865
rect 3057 1831 3091 1865
rect 3393 1831 3427 1865
rect 3729 1831 3763 1865
rect 4065 1831 4099 1865
rect 4401 1831 4435 1865
rect 4737 1831 4771 1865
rect 5073 1831 5107 1865
rect 5409 1831 5443 1865
rect 5745 1831 5779 1865
rect 6081 1831 6115 1865
rect 6417 1831 6451 1865
rect 6753 1831 6787 1865
rect 7089 1831 7123 1865
rect 7425 1831 7459 1865
rect 7761 1831 7795 1865
rect 8097 1831 8131 1865
rect 8433 1831 8467 1865
rect 8769 1831 8803 1865
rect 9105 1831 9139 1865
rect 9441 1831 9475 1865
rect 9777 1831 9811 1865
rect 10113 1831 10147 1865
rect 10449 1831 10483 1865
rect 10785 1831 10819 1865
rect 11121 1831 11155 1865
rect 11457 1831 11491 1865
rect 11793 1831 11827 1865
rect 12129 1831 12163 1865
rect 12465 1831 12499 1865
rect 12801 1831 12835 1865
rect 13137 1831 13171 1865
rect 13473 1831 13507 1865
rect 13809 1831 13843 1865
rect 14145 1831 14179 1865
rect 14481 1831 14515 1865
rect 14817 1831 14851 1865
rect 15153 1831 15187 1865
rect 15489 1831 15523 1865
rect 15825 1831 15859 1865
rect 16161 1831 16195 1865
rect 16497 1831 16531 1865
rect 16833 1831 16867 1865
rect 17169 1831 17203 1865
rect 17505 1831 17539 1865
rect 17841 1831 17875 1865
rect 18177 1831 18211 1865
rect 18513 1831 18547 1865
rect 18849 1831 18883 1865
rect 19185 1831 19219 1865
rect 19521 1831 19555 1865
rect 19857 1831 19891 1865
rect 20193 1831 20227 1865
rect 20529 1831 20563 1865
rect 20865 1831 20899 1865
rect 21201 1831 21235 1865
rect 21537 1831 21571 1865
rect 21873 1831 21907 1865
rect 22209 1831 22243 1865
rect 22545 1831 22579 1865
rect 22881 1831 22915 1865
rect 23217 1831 23251 1865
rect 23553 1831 23587 1865
rect 23889 1831 23923 1865
rect 24225 1831 24259 1865
rect 24561 1831 24595 1865
rect 24897 1831 24931 1865
rect 25233 1831 25267 1865
rect 25569 1831 25603 1865
rect 25905 1831 25939 1865
rect 26241 1831 26275 1865
rect 26577 1831 26611 1865
rect 26913 1831 26947 1865
rect 27249 1831 27283 1865
rect 27585 1831 27619 1865
rect 27921 1831 27955 1865
rect 28257 1831 28291 1865
rect 28593 1831 28627 1865
rect 28929 1831 28963 1865
rect 29265 1831 29299 1865
rect 29601 1831 29635 1865
rect 29937 1831 29971 1865
rect 30273 1831 30307 1865
rect 30609 1831 30643 1865
rect 30945 1831 30979 1865
rect 31281 1831 31315 1865
rect 31617 1831 31651 1865
rect 31953 1831 31987 1865
rect 32289 1831 32323 1865
rect 32625 1831 32659 1865
rect 32961 1831 32995 1865
rect 33297 1831 33331 1865
rect 33633 1831 33667 1865
rect 33969 1831 34003 1865
rect 34305 1831 34339 1865
rect 34641 1831 34675 1865
rect 34977 1831 35011 1865
rect 35313 1831 35347 1865
rect 35649 1831 35683 1865
rect 35985 1831 36019 1865
rect 36321 1831 36355 1865
rect 36657 1831 36691 1865
rect 36993 1831 37027 1865
rect 37329 1831 37363 1865
rect 37665 1831 37699 1865
rect 38001 1831 38035 1865
rect 38337 1831 38371 1865
rect 38673 1831 38707 1865
rect 39009 1831 39043 1865
rect 39345 1831 39379 1865
rect 39681 1831 39715 1865
rect 40017 1831 40051 1865
rect 40353 1831 40387 1865
rect 40689 1831 40723 1865
rect 41025 1831 41059 1865
rect 41361 1831 41395 1865
rect 41697 1831 41731 1865
rect 42033 1831 42067 1865
rect 42369 1831 42403 1865
rect 42705 1831 42739 1865
rect 43041 1831 43075 1865
rect 43377 1831 43411 1865
rect 43713 1831 43747 1865
rect 44049 1831 44083 1865
rect 44385 1831 44419 1865
rect 44721 1831 44755 1865
rect 45057 1831 45091 1865
rect 45393 1831 45427 1865
rect 45729 1831 45763 1865
rect 46065 1831 46099 1865
rect 46401 1831 46435 1865
rect 46737 1831 46771 1865
rect 47073 1831 47107 1865
rect 47409 1831 47443 1865
rect 47745 1831 47779 1865
rect 48081 1831 48115 1865
rect 48417 1831 48451 1865
rect 48753 1831 48787 1865
rect 49089 1831 49123 1865
rect 49425 1831 49459 1865
rect 49761 1831 49795 1865
rect 50097 1831 50131 1865
rect 50433 1831 50467 1865
rect 50769 1831 50803 1865
rect 51105 1831 51139 1865
rect 51441 1831 51475 1865
rect 51777 1831 51811 1865
rect 52113 1831 52147 1865
rect 52449 1831 52483 1865
rect 52785 1831 52819 1865
rect 53121 1831 53155 1865
rect 53457 1831 53491 1865
rect 53793 1831 53827 1865
rect 54129 1831 54163 1865
rect 54465 1831 54499 1865
rect 54801 1831 54835 1865
rect 55137 1831 55171 1865
rect 55473 1831 55507 1865
rect 55809 1831 55843 1865
rect 56145 1831 56179 1865
rect 56481 1831 56515 1865
rect 56817 1831 56851 1865
rect 57153 1831 57187 1865
rect 57489 1831 57523 1865
rect 57825 1831 57859 1865
rect 58161 1831 58195 1865
rect 58497 1831 58531 1865
rect 58833 1831 58867 1865
rect 59169 1831 59203 1865
rect 59505 1831 59539 1865
rect 59841 1831 59875 1865
rect 60177 1831 60211 1865
rect 60513 1831 60547 1865
rect 60849 1831 60883 1865
rect 61185 1831 61219 1865
rect 61521 1831 61555 1865
rect 61857 1831 61891 1865
rect 62193 1831 62227 1865
rect 62529 1831 62563 1865
rect 62865 1831 62899 1865
rect 63201 1831 63235 1865
rect 63537 1831 63571 1865
rect 63873 1831 63907 1865
rect 64209 1831 64243 1865
rect 64545 1831 64579 1865
rect 64881 1831 64915 1865
rect 65217 1831 65251 1865
rect 65553 1831 65587 1865
rect 65889 1831 65923 1865
rect 66225 1831 66259 1865
rect 66561 1831 66595 1865
rect 66897 1831 66931 1865
rect 67233 1831 67267 1865
rect 67569 1831 67603 1865
rect 67905 1831 67939 1865
rect 68241 1831 68275 1865
rect 68577 1831 68611 1865
rect 68913 1831 68947 1865
rect 69249 1831 69283 1865
rect 69585 1831 69619 1865
rect 69921 1831 69955 1865
rect 70257 1831 70291 1865
rect 70593 1831 70627 1865
rect 70929 1831 70963 1865
rect 71265 1831 71299 1865
rect 71601 1831 71635 1865
rect 71937 1831 71971 1865
rect 72273 1831 72307 1865
rect 72609 1831 72643 1865
rect 72945 1831 72979 1865
rect 73281 1831 73315 1865
rect 73617 1831 73651 1865
rect 73953 1831 73987 1865
rect 74289 1831 74323 1865
rect 74625 1831 74659 1865
rect 74961 1831 74995 1865
rect 75297 1831 75331 1865
rect 75633 1831 75667 1865
rect 75969 1831 76003 1865
rect 76305 1831 76339 1865
rect 76641 1831 76675 1865
rect 76977 1831 77011 1865
rect 77313 1831 77347 1865
rect 77649 1831 77683 1865
rect 77985 1831 78019 1865
rect 78321 1831 78355 1865
rect 78657 1831 78691 1865
rect 78993 1831 79027 1865
rect 79329 1831 79363 1865
rect 79665 1831 79699 1865
rect 80001 1831 80035 1865
rect 80337 1831 80371 1865
rect 80673 1831 80707 1865
rect 81009 1831 81043 1865
rect 81345 1831 81379 1865
rect 81681 1831 81715 1865
rect 82017 1831 82051 1865
rect 82353 1831 82387 1865
rect 82689 1831 82723 1865
rect 83025 1831 83059 1865
rect 83361 1831 83395 1865
rect 83697 1831 83731 1865
rect 84033 1831 84067 1865
rect 84369 1831 84403 1865
rect 84705 1831 84739 1865
rect 85041 1831 85075 1865
rect 85377 1831 85411 1865
rect 85713 1831 85747 1865
rect 86049 1831 86083 1865
rect 86385 1831 86419 1865
rect 86721 1831 86755 1865
rect 87057 1831 87091 1865
rect 87393 1831 87427 1865
rect 87729 1831 87763 1865
rect 88065 1831 88099 1865
rect 88401 1831 88435 1865
rect 88737 1831 88771 1865
rect 89073 1831 89107 1865
rect 89409 1831 89443 1865
rect 89745 1831 89779 1865
rect 90081 1831 90115 1865
rect 90417 1831 90451 1865
rect 90753 1831 90787 1865
rect 91089 1831 91123 1865
rect 91425 1831 91459 1865
rect 91761 1831 91795 1865
rect 92097 1831 92131 1865
rect 92433 1831 92467 1865
rect 92769 1831 92803 1865
rect 93105 1831 93139 1865
rect 93441 1831 93475 1865
rect 93777 1831 93811 1865
rect 94113 1831 94147 1865
rect 94449 1831 94483 1865
rect 94785 1831 94819 1865
rect 95121 1831 95155 1865
rect 95457 1831 95491 1865
rect 95793 1831 95827 1865
rect 96129 1831 96163 1865
rect 96465 1831 96499 1865
rect 96801 1831 96835 1865
rect 97137 1831 97171 1865
rect 97473 1831 97507 1865
rect 97809 1831 97843 1865
rect 98145 1831 98179 1865
rect 98481 1831 98515 1865
rect 98817 1831 98851 1865
rect 99153 1831 99187 1865
rect 99489 1831 99523 1865
rect 99825 1831 99859 1865
rect 100161 1831 100195 1865
rect 100497 1831 100531 1865
rect 100833 1831 100867 1865
rect 101169 1831 101203 1865
rect 101505 1831 101539 1865
rect 101841 1831 101875 1865
rect 102177 1831 102211 1865
rect 102513 1831 102547 1865
rect 102849 1831 102883 1865
rect 103185 1831 103219 1865
rect 103521 1831 103555 1865
rect 103857 1831 103891 1865
rect 104193 1831 104227 1865
rect 104529 1831 104563 1865
rect 104865 1831 104899 1865
rect 105201 1831 105235 1865
rect 105537 1831 105571 1865
rect 105873 1831 105907 1865
rect 106209 1831 106243 1865
rect 106545 1831 106579 1865
rect 106881 1831 106915 1865
rect 107217 1831 107251 1865
rect 107553 1831 107587 1865
rect 107889 1831 107923 1865
rect 108225 1831 108259 1865
rect 108561 1831 108595 1865
rect 108897 1831 108931 1865
rect 109233 1831 109267 1865
rect 109569 1831 109603 1865
rect 109905 1831 109939 1865
rect 110241 1831 110275 1865
rect 110577 1831 110611 1865
rect 110913 1831 110947 1865
rect 111249 1831 111283 1865
rect 111585 1831 111619 1865
rect 111921 1831 111955 1865
rect 112257 1831 112291 1865
rect 112593 1831 112627 1865
rect 112929 1831 112963 1865
rect 113265 1831 113299 1865
rect 113601 1831 113635 1865
rect 113937 1831 113971 1865
rect 114273 1831 114307 1865
rect 114609 1831 114643 1865
rect 114945 1831 114979 1865
rect 115281 1831 115315 1865
rect 115617 1831 115651 1865
rect 115953 1831 115987 1865
rect 116289 1831 116323 1865
rect 116625 1831 116659 1865
rect 116961 1831 116995 1865
rect 117297 1831 117331 1865
rect 117633 1831 117667 1865
rect 117969 1831 118003 1865
rect 118305 1831 118339 1865
rect 118641 1831 118675 1865
rect 118977 1831 119011 1865
rect 119313 1831 119347 1865
rect 119649 1831 119683 1865
rect 119985 1831 120019 1865
rect 120321 1831 120355 1865
rect 120657 1831 120691 1865
rect 120993 1831 121027 1865
rect 121329 1831 121363 1865
rect 121665 1831 121699 1865
rect 122001 1831 122035 1865
rect 122337 1831 122371 1865
rect 122673 1831 122707 1865
rect 123009 1831 123043 1865
rect 123345 1831 123379 1865
rect 123681 1831 123715 1865
rect 124017 1831 124051 1865
rect 124353 1831 124387 1865
rect 124689 1831 124723 1865
rect 125025 1831 125059 1865
rect 125361 1831 125395 1865
rect 125697 1831 125731 1865
rect 126033 1831 126067 1865
rect 126369 1831 126403 1865
rect 126705 1831 126739 1865
rect 127041 1831 127075 1865
rect 127377 1831 127411 1865
rect 127713 1831 127747 1865
rect 128049 1831 128083 1865
rect 128385 1831 128419 1865
rect 128721 1831 128755 1865
rect 129057 1831 129091 1865
rect 129393 1831 129427 1865
rect 129729 1831 129763 1865
rect 130065 1831 130099 1865
rect 130401 1831 130435 1865
rect 130737 1831 130771 1865
rect 131073 1831 131107 1865
rect 131409 1831 131443 1865
rect 131745 1831 131779 1865
rect 132081 1831 132115 1865
rect 132417 1831 132451 1865
rect 132753 1831 132787 1865
rect 133089 1831 133123 1865
rect 133425 1831 133459 1865
rect 133761 1831 133795 1865
rect 134097 1831 134131 1865
rect 134433 1831 134467 1865
rect 134769 1831 134803 1865
rect 135105 1831 135139 1865
rect 135441 1831 135475 1865
rect 135777 1831 135811 1865
rect 136113 1831 136147 1865
rect 136449 1831 136483 1865
rect 136785 1831 136819 1865
rect 137121 1831 137155 1865
rect 137457 1831 137491 1865
rect 137793 1831 137827 1865
rect 138129 1831 138163 1865
rect 138465 1831 138499 1865
rect 138801 1831 138835 1865
rect 139137 1831 139171 1865
rect 139473 1831 139507 1865
rect 139809 1831 139843 1865
rect 140145 1831 140179 1865
rect 140481 1831 140515 1865
rect 140817 1831 140851 1865
rect 141153 1831 141187 1865
rect 141489 1831 141523 1865
rect 141825 1831 141859 1865
rect 142161 1831 142195 1865
rect 142497 1831 142531 1865
rect 142833 1831 142867 1865
rect 143169 1831 143203 1865
rect 143505 1831 143539 1865
rect 143841 1831 143875 1865
rect 144177 1831 144211 1865
rect 144513 1831 144547 1865
rect 144849 1831 144883 1865
rect 145185 1831 145219 1865
rect 145521 1831 145555 1865
rect 145857 1831 145891 1865
rect 146193 1831 146227 1865
rect 146529 1831 146563 1865
rect 146865 1831 146899 1865
rect 147201 1831 147235 1865
rect 147537 1831 147571 1865
rect 147873 1831 147907 1865
rect 148209 1831 148243 1865
rect 148545 1831 148579 1865
rect 148881 1831 148915 1865
rect 149217 1831 149251 1865
rect 149553 1831 149587 1865
rect 149889 1831 149923 1865
rect 150225 1831 150259 1865
rect 150561 1831 150595 1865
rect 150897 1831 150931 1865
rect 151233 1831 151267 1865
rect 151569 1831 151603 1865
rect 151905 1831 151939 1865
rect 152241 1831 152275 1865
rect 152577 1831 152611 1865
rect 152913 1831 152947 1865
rect 153249 1831 153283 1865
rect 153585 1831 153619 1865
rect 153921 1831 153955 1865
rect 154257 1831 154291 1865
rect 154593 1831 154627 1865
rect 154929 1831 154963 1865
rect 155265 1831 155299 1865
rect 155601 1831 155635 1865
rect 155937 1831 155971 1865
rect 156273 1831 156307 1865
rect 156609 1831 156643 1865
rect 156945 1831 156979 1865
rect 157281 1831 157315 1865
rect 157617 1831 157651 1865
rect 157953 1831 157987 1865
rect 158289 1831 158323 1865
rect 158625 1831 158659 1865
rect 158961 1831 158995 1865
rect 159297 1831 159331 1865
rect 159633 1831 159667 1865
rect 159969 1831 160003 1865
rect 160305 1831 160339 1865
rect 160641 1831 160675 1865
rect 160977 1831 161011 1865
rect 161313 1831 161347 1865
rect 161649 1831 161683 1865
rect 161985 1831 162019 1865
rect 162321 1831 162355 1865
rect 162657 1831 162691 1865
rect 162993 1831 163027 1865
rect 163329 1831 163363 1865
rect 163665 1831 163699 1865
rect 164001 1831 164035 1865
rect 164337 1831 164371 1865
rect 164673 1831 164707 1865
rect 165009 1831 165043 1865
rect 165345 1831 165379 1865
rect 165681 1831 165715 1865
rect 166017 1831 166051 1865
rect 166353 1831 166387 1865
rect 166689 1831 166723 1865
rect 167025 1831 167059 1865
rect 167361 1831 167395 1865
rect 167697 1831 167731 1865
rect 168033 1831 168067 1865
rect 168369 1831 168403 1865
rect 168705 1831 168739 1865
rect 169041 1831 169075 1865
rect 169377 1831 169411 1865
rect 169713 1831 169747 1865
rect 170049 1831 170083 1865
rect 170385 1831 170419 1865
rect 170721 1831 170755 1865
rect 171057 1831 171091 1865
rect 171393 1831 171427 1865
rect 171729 1831 171763 1865
rect 172065 1831 172099 1865
rect 172401 1831 172435 1865
rect 172737 1831 172771 1865
rect 173073 1831 173107 1865
rect 173409 1831 173443 1865
rect 173745 1831 173779 1865
rect 174081 1831 174115 1865
rect 174417 1831 174451 1865
rect 174753 1831 174787 1865
rect 175089 1831 175123 1865
rect 175425 1831 175459 1865
rect 175761 1831 175795 1865
rect 176097 1831 176131 1865
rect 176433 1831 176467 1865
rect 176769 1831 176803 1865
rect 177105 1831 177139 1865
rect 177441 1831 177475 1865
rect 177777 1831 177811 1865
rect 178113 1831 178147 1865
rect 178449 1831 178483 1865
rect 178785 1831 178819 1865
rect 179121 1831 179155 1865
rect 179457 1831 179491 1865
rect 179793 1831 179827 1865
rect 180129 1831 180163 1865
rect 180465 1831 180499 1865
rect 180801 1831 180835 1865
rect 181137 1831 181171 1865
rect 181473 1831 181507 1865
rect 181809 1831 181843 1865
rect 182145 1831 182179 1865
rect 182481 1831 182515 1865
rect 182817 1831 182851 1865
rect 183153 1831 183187 1865
rect 183489 1831 183523 1865
rect 183825 1831 183859 1865
rect 184161 1831 184195 1865
rect 184497 1831 184531 1865
rect 184833 1831 184867 1865
rect 185169 1831 185203 1865
rect 185505 1831 185539 1865
rect 185841 1831 185875 1865
rect 186177 1831 186211 1865
rect 186513 1831 186547 1865
rect 186849 1831 186883 1865
rect 187185 1831 187219 1865
rect 187521 1831 187555 1865
rect 187857 1831 187891 1865
rect 188193 1831 188227 1865
rect 188529 1831 188563 1865
rect 188865 1831 188899 1865
rect 189201 1831 189235 1865
rect 189537 1831 189571 1865
rect 189873 1831 189907 1865
rect 190209 1831 190243 1865
rect 190545 1831 190579 1865
rect 190881 1831 190915 1865
rect 191217 1831 191251 1865
rect 191553 1831 191587 1865
rect 191889 1831 191923 1865
rect 192225 1831 192259 1865
rect 192561 1831 192595 1865
rect 192897 1831 192931 1865
rect 193233 1831 193267 1865
rect 193569 1831 193603 1865
rect 193905 1831 193939 1865
rect 194241 1831 194275 1865
rect 194577 1831 194611 1865
rect 194913 1831 194947 1865
rect 195249 1831 195283 1865
rect 195585 1831 195619 1865
rect 195921 1831 195955 1865
rect 196257 1831 196291 1865
rect 196593 1831 196627 1865
rect 196929 1831 196963 1865
rect 197265 1831 197299 1865
rect 197601 1831 197635 1865
rect 197937 1831 197971 1865
rect 198273 1831 198307 1865
rect 198609 1831 198643 1865
rect 198945 1831 198979 1865
rect 199281 1831 199315 1865
rect 199617 1831 199651 1865
rect 199953 1831 199987 1865
rect 200289 1831 200323 1865
rect 200625 1831 200659 1865
rect 200961 1831 200995 1865
rect 201297 1831 201331 1865
rect 201633 1831 201667 1865
rect 201969 1831 202003 1865
rect 202305 1831 202339 1865
rect 202641 1831 202675 1865
rect 202977 1831 203011 1865
rect 203313 1831 203347 1865
rect 203649 1831 203683 1865
rect 203985 1831 204019 1865
rect 204321 1831 204355 1865
rect 204657 1831 204691 1865
rect 204993 1831 205027 1865
rect 205329 1831 205363 1865
rect 205665 1831 205699 1865
rect 206001 1831 206035 1865
rect 206337 1831 206371 1865
rect 206673 1831 206707 1865
rect 207009 1831 207043 1865
rect 207345 1831 207379 1865
rect 207681 1831 207715 1865
rect 208017 1831 208051 1865
rect 208353 1831 208387 1865
rect 208689 1831 208723 1865
rect 209025 1831 209059 1865
rect 209361 1831 209395 1865
rect 209697 1831 209731 1865
rect 210033 1831 210067 1865
rect 210369 1831 210403 1865
rect 210705 1831 210739 1865
rect 211041 1831 211075 1865
rect 211377 1831 211411 1865
rect 211713 1831 211747 1865
rect 212049 1831 212083 1865
rect 212385 1831 212419 1865
rect 212721 1831 212755 1865
rect 213057 1831 213091 1865
rect 213393 1831 213427 1865
rect 213729 1831 213763 1865
rect 214065 1831 214099 1865
rect 214401 1831 214435 1865
rect 214737 1831 214771 1865
rect 215073 1831 215107 1865
rect 215409 1831 215443 1865
rect 215745 1831 215779 1865
rect 216081 1831 216115 1865
rect 216417 1831 216451 1865
<< metal1 >>
rect 1618 142370 217048 142456
rect 1618 142318 2040 142370
rect 2092 142361 3720 142370
rect 3772 142361 5400 142370
rect 5452 142361 7080 142370
rect 7132 142361 8760 142370
rect 8812 142361 10440 142370
rect 10492 142361 12120 142370
rect 12172 142361 13800 142370
rect 13852 142361 15480 142370
rect 15532 142361 17160 142370
rect 17212 142361 18840 142370
rect 18892 142361 20520 142370
rect 20572 142361 22200 142370
rect 22252 142361 23880 142370
rect 23932 142361 25560 142370
rect 25612 142361 27240 142370
rect 27292 142361 28920 142370
rect 28972 142361 30600 142370
rect 30652 142361 32280 142370
rect 32332 142361 33960 142370
rect 34012 142361 35640 142370
rect 35692 142361 37320 142370
rect 37372 142361 39000 142370
rect 39052 142361 40680 142370
rect 40732 142361 42360 142370
rect 42412 142361 44040 142370
rect 44092 142361 45720 142370
rect 45772 142361 47400 142370
rect 47452 142361 49080 142370
rect 49132 142361 50760 142370
rect 50812 142361 52440 142370
rect 52492 142361 54120 142370
rect 54172 142361 55800 142370
rect 55852 142361 57480 142370
rect 57532 142361 59160 142370
rect 59212 142361 60840 142370
rect 60892 142361 62520 142370
rect 62572 142361 64200 142370
rect 64252 142361 65880 142370
rect 65932 142361 67560 142370
rect 67612 142361 69240 142370
rect 69292 142361 70920 142370
rect 70972 142361 72600 142370
rect 72652 142361 74280 142370
rect 74332 142361 75960 142370
rect 76012 142361 77640 142370
rect 77692 142361 79320 142370
rect 79372 142361 81000 142370
rect 81052 142361 82680 142370
rect 82732 142361 84360 142370
rect 84412 142361 86040 142370
rect 86092 142361 87720 142370
rect 87772 142361 89400 142370
rect 89452 142361 91080 142370
rect 91132 142361 92760 142370
rect 92812 142361 94440 142370
rect 94492 142361 96120 142370
rect 96172 142361 97800 142370
rect 97852 142361 99480 142370
rect 99532 142361 101160 142370
rect 101212 142361 102840 142370
rect 102892 142361 104520 142370
rect 104572 142361 106200 142370
rect 106252 142361 107880 142370
rect 107932 142361 109560 142370
rect 109612 142361 111240 142370
rect 111292 142361 112920 142370
rect 112972 142361 114600 142370
rect 114652 142361 116280 142370
rect 116332 142361 117960 142370
rect 118012 142361 119640 142370
rect 119692 142361 121320 142370
rect 121372 142361 123000 142370
rect 123052 142361 124680 142370
rect 124732 142361 126360 142370
rect 126412 142361 128040 142370
rect 128092 142361 129720 142370
rect 129772 142361 131400 142370
rect 131452 142361 133080 142370
rect 133132 142361 134760 142370
rect 134812 142361 136440 142370
rect 136492 142361 138120 142370
rect 138172 142361 139800 142370
rect 139852 142361 141480 142370
rect 141532 142361 143160 142370
rect 143212 142361 144840 142370
rect 144892 142361 146520 142370
rect 146572 142361 148200 142370
rect 148252 142361 149880 142370
rect 149932 142361 151560 142370
rect 151612 142361 153240 142370
rect 153292 142361 154920 142370
rect 154972 142361 156600 142370
rect 156652 142361 158280 142370
rect 158332 142361 159960 142370
rect 160012 142361 161640 142370
rect 161692 142361 163320 142370
rect 163372 142361 165000 142370
rect 165052 142361 166680 142370
rect 166732 142361 168360 142370
rect 168412 142361 170040 142370
rect 170092 142361 171720 142370
rect 171772 142361 173400 142370
rect 173452 142361 175080 142370
rect 175132 142361 176760 142370
rect 176812 142361 178440 142370
rect 178492 142361 180120 142370
rect 180172 142361 181800 142370
rect 181852 142361 183480 142370
rect 183532 142361 185160 142370
rect 185212 142361 186840 142370
rect 186892 142361 188520 142370
rect 188572 142361 190200 142370
rect 190252 142361 191880 142370
rect 191932 142361 193560 142370
rect 193612 142361 195240 142370
rect 195292 142361 196920 142370
rect 196972 142361 198600 142370
rect 198652 142361 200280 142370
rect 200332 142361 201960 142370
rect 202012 142361 203640 142370
rect 203692 142361 205320 142370
rect 205372 142361 207000 142370
rect 207052 142361 208680 142370
rect 208732 142361 210360 142370
rect 210412 142361 212040 142370
rect 212092 142361 213720 142370
rect 213772 142361 215400 142370
rect 215452 142361 217048 142370
rect 2092 142327 2385 142361
rect 2419 142327 2721 142361
rect 2755 142327 3057 142361
rect 3091 142327 3393 142361
rect 3427 142327 3720 142361
rect 3772 142327 4065 142361
rect 4099 142327 4401 142361
rect 4435 142327 4737 142361
rect 4771 142327 5073 142361
rect 5107 142327 5400 142361
rect 5452 142327 5745 142361
rect 5779 142327 6081 142361
rect 6115 142327 6417 142361
rect 6451 142327 6753 142361
rect 6787 142327 7080 142361
rect 7132 142327 7425 142361
rect 7459 142327 7761 142361
rect 7795 142327 8097 142361
rect 8131 142327 8433 142361
rect 8467 142327 8760 142361
rect 8812 142327 9105 142361
rect 9139 142327 9441 142361
rect 9475 142327 9777 142361
rect 9811 142327 10113 142361
rect 10147 142327 10440 142361
rect 10492 142327 10785 142361
rect 10819 142327 11121 142361
rect 11155 142327 11457 142361
rect 11491 142327 11793 142361
rect 11827 142327 12120 142361
rect 12172 142327 12465 142361
rect 12499 142327 12801 142361
rect 12835 142327 13137 142361
rect 13171 142327 13473 142361
rect 13507 142327 13800 142361
rect 13852 142327 14145 142361
rect 14179 142327 14481 142361
rect 14515 142327 14817 142361
rect 14851 142327 15153 142361
rect 15187 142327 15480 142361
rect 15532 142327 15825 142361
rect 15859 142327 16161 142361
rect 16195 142327 16497 142361
rect 16531 142327 16833 142361
rect 16867 142327 17160 142361
rect 17212 142327 17505 142361
rect 17539 142327 17841 142361
rect 17875 142327 18177 142361
rect 18211 142327 18513 142361
rect 18547 142327 18840 142361
rect 18892 142327 19185 142361
rect 19219 142327 19521 142361
rect 19555 142327 19857 142361
rect 19891 142327 20193 142361
rect 20227 142327 20520 142361
rect 20572 142327 20865 142361
rect 20899 142327 21201 142361
rect 21235 142327 21537 142361
rect 21571 142327 21873 142361
rect 21907 142327 22200 142361
rect 22252 142327 22545 142361
rect 22579 142327 22881 142361
rect 22915 142327 23217 142361
rect 23251 142327 23553 142361
rect 23587 142327 23880 142361
rect 23932 142327 24225 142361
rect 24259 142327 24561 142361
rect 24595 142327 24897 142361
rect 24931 142327 25233 142361
rect 25267 142327 25560 142361
rect 25612 142327 25905 142361
rect 25939 142327 26241 142361
rect 26275 142327 26577 142361
rect 26611 142327 26913 142361
rect 26947 142327 27240 142361
rect 27292 142327 27585 142361
rect 27619 142327 27921 142361
rect 27955 142327 28257 142361
rect 28291 142327 28593 142361
rect 28627 142327 28920 142361
rect 28972 142327 29265 142361
rect 29299 142327 29601 142361
rect 29635 142327 29937 142361
rect 29971 142327 30273 142361
rect 30307 142327 30600 142361
rect 30652 142327 30945 142361
rect 30979 142327 31281 142361
rect 31315 142327 31617 142361
rect 31651 142327 31953 142361
rect 31987 142327 32280 142361
rect 32332 142327 32625 142361
rect 32659 142327 32961 142361
rect 32995 142327 33297 142361
rect 33331 142327 33633 142361
rect 33667 142327 33960 142361
rect 34012 142327 34305 142361
rect 34339 142327 34641 142361
rect 34675 142327 34977 142361
rect 35011 142327 35313 142361
rect 35347 142327 35640 142361
rect 35692 142327 35985 142361
rect 36019 142327 36321 142361
rect 36355 142327 36657 142361
rect 36691 142327 36993 142361
rect 37027 142327 37320 142361
rect 37372 142327 37665 142361
rect 37699 142327 38001 142361
rect 38035 142327 38337 142361
rect 38371 142327 38673 142361
rect 38707 142327 39000 142361
rect 39052 142327 39345 142361
rect 39379 142327 39681 142361
rect 39715 142327 40017 142361
rect 40051 142327 40353 142361
rect 40387 142327 40680 142361
rect 40732 142327 41025 142361
rect 41059 142327 41361 142361
rect 41395 142327 41697 142361
rect 41731 142327 42033 142361
rect 42067 142327 42360 142361
rect 42412 142327 42705 142361
rect 42739 142327 43041 142361
rect 43075 142327 43377 142361
rect 43411 142327 43713 142361
rect 43747 142327 44040 142361
rect 44092 142327 44385 142361
rect 44419 142327 44721 142361
rect 44755 142327 45057 142361
rect 45091 142327 45393 142361
rect 45427 142327 45720 142361
rect 45772 142327 46065 142361
rect 46099 142327 46401 142361
rect 46435 142327 46737 142361
rect 46771 142327 47073 142361
rect 47107 142327 47400 142361
rect 47452 142327 47745 142361
rect 47779 142327 48081 142361
rect 48115 142327 48417 142361
rect 48451 142327 48753 142361
rect 48787 142327 49080 142361
rect 49132 142327 49425 142361
rect 49459 142327 49761 142361
rect 49795 142327 50097 142361
rect 50131 142327 50433 142361
rect 50467 142327 50760 142361
rect 50812 142327 51105 142361
rect 51139 142327 51441 142361
rect 51475 142327 51777 142361
rect 51811 142327 52113 142361
rect 52147 142327 52440 142361
rect 52492 142327 52785 142361
rect 52819 142327 53121 142361
rect 53155 142327 53457 142361
rect 53491 142327 53793 142361
rect 53827 142327 54120 142361
rect 54172 142327 54465 142361
rect 54499 142327 54801 142361
rect 54835 142327 55137 142361
rect 55171 142327 55473 142361
rect 55507 142327 55800 142361
rect 55852 142327 56145 142361
rect 56179 142327 56481 142361
rect 56515 142327 56817 142361
rect 56851 142327 57153 142361
rect 57187 142327 57480 142361
rect 57532 142327 57825 142361
rect 57859 142327 58161 142361
rect 58195 142327 58497 142361
rect 58531 142327 58833 142361
rect 58867 142327 59160 142361
rect 59212 142327 59505 142361
rect 59539 142327 59841 142361
rect 59875 142327 60177 142361
rect 60211 142327 60513 142361
rect 60547 142327 60840 142361
rect 60892 142327 61185 142361
rect 61219 142327 61521 142361
rect 61555 142327 61857 142361
rect 61891 142327 62193 142361
rect 62227 142327 62520 142361
rect 62572 142327 62865 142361
rect 62899 142327 63201 142361
rect 63235 142327 63537 142361
rect 63571 142327 63873 142361
rect 63907 142327 64200 142361
rect 64252 142327 64545 142361
rect 64579 142327 64881 142361
rect 64915 142327 65217 142361
rect 65251 142327 65553 142361
rect 65587 142327 65880 142361
rect 65932 142327 66225 142361
rect 66259 142327 66561 142361
rect 66595 142327 66897 142361
rect 66931 142327 67233 142361
rect 67267 142327 67560 142361
rect 67612 142327 67905 142361
rect 67939 142327 68241 142361
rect 68275 142327 68577 142361
rect 68611 142327 68913 142361
rect 68947 142327 69240 142361
rect 69292 142327 69585 142361
rect 69619 142327 69921 142361
rect 69955 142327 70257 142361
rect 70291 142327 70593 142361
rect 70627 142327 70920 142361
rect 70972 142327 71265 142361
rect 71299 142327 71601 142361
rect 71635 142327 71937 142361
rect 71971 142327 72273 142361
rect 72307 142327 72600 142361
rect 72652 142327 72945 142361
rect 72979 142327 73281 142361
rect 73315 142327 73617 142361
rect 73651 142327 73953 142361
rect 73987 142327 74280 142361
rect 74332 142327 74625 142361
rect 74659 142327 74961 142361
rect 74995 142327 75297 142361
rect 75331 142327 75633 142361
rect 75667 142327 75960 142361
rect 76012 142327 76305 142361
rect 76339 142327 76641 142361
rect 76675 142327 76977 142361
rect 77011 142327 77313 142361
rect 77347 142327 77640 142361
rect 77692 142327 77985 142361
rect 78019 142327 78321 142361
rect 78355 142327 78657 142361
rect 78691 142327 78993 142361
rect 79027 142327 79320 142361
rect 79372 142327 79665 142361
rect 79699 142327 80001 142361
rect 80035 142327 80337 142361
rect 80371 142327 80673 142361
rect 80707 142327 81000 142361
rect 81052 142327 81345 142361
rect 81379 142327 81681 142361
rect 81715 142327 82017 142361
rect 82051 142327 82353 142361
rect 82387 142327 82680 142361
rect 82732 142327 83025 142361
rect 83059 142327 83361 142361
rect 83395 142327 83697 142361
rect 83731 142327 84033 142361
rect 84067 142327 84360 142361
rect 84412 142327 84705 142361
rect 84739 142327 85041 142361
rect 85075 142327 85377 142361
rect 85411 142327 85713 142361
rect 85747 142327 86040 142361
rect 86092 142327 86385 142361
rect 86419 142327 86721 142361
rect 86755 142327 87057 142361
rect 87091 142327 87393 142361
rect 87427 142327 87720 142361
rect 87772 142327 88065 142361
rect 88099 142327 88401 142361
rect 88435 142327 88737 142361
rect 88771 142327 89073 142361
rect 89107 142327 89400 142361
rect 89452 142327 89745 142361
rect 89779 142327 90081 142361
rect 90115 142327 90417 142361
rect 90451 142327 90753 142361
rect 90787 142327 91080 142361
rect 91132 142327 91425 142361
rect 91459 142327 91761 142361
rect 91795 142327 92097 142361
rect 92131 142327 92433 142361
rect 92467 142327 92760 142361
rect 92812 142327 93105 142361
rect 93139 142327 93441 142361
rect 93475 142327 93777 142361
rect 93811 142327 94113 142361
rect 94147 142327 94440 142361
rect 94492 142327 94785 142361
rect 94819 142327 95121 142361
rect 95155 142327 95457 142361
rect 95491 142327 95793 142361
rect 95827 142327 96120 142361
rect 96172 142327 96465 142361
rect 96499 142327 96801 142361
rect 96835 142327 97137 142361
rect 97171 142327 97473 142361
rect 97507 142327 97800 142361
rect 97852 142327 98145 142361
rect 98179 142327 98481 142361
rect 98515 142327 98817 142361
rect 98851 142327 99153 142361
rect 99187 142327 99480 142361
rect 99532 142327 99825 142361
rect 99859 142327 100161 142361
rect 100195 142327 100497 142361
rect 100531 142327 100833 142361
rect 100867 142327 101160 142361
rect 101212 142327 101505 142361
rect 101539 142327 101841 142361
rect 101875 142327 102177 142361
rect 102211 142327 102513 142361
rect 102547 142327 102840 142361
rect 102892 142327 103185 142361
rect 103219 142327 103521 142361
rect 103555 142327 103857 142361
rect 103891 142327 104193 142361
rect 104227 142327 104520 142361
rect 104572 142327 104865 142361
rect 104899 142327 105201 142361
rect 105235 142327 105537 142361
rect 105571 142327 105873 142361
rect 105907 142327 106200 142361
rect 106252 142327 106545 142361
rect 106579 142327 106881 142361
rect 106915 142327 107217 142361
rect 107251 142327 107553 142361
rect 107587 142327 107880 142361
rect 107932 142327 108225 142361
rect 108259 142327 108561 142361
rect 108595 142327 108897 142361
rect 108931 142327 109233 142361
rect 109267 142327 109560 142361
rect 109612 142327 109905 142361
rect 109939 142327 110241 142361
rect 110275 142327 110577 142361
rect 110611 142327 110913 142361
rect 110947 142327 111240 142361
rect 111292 142327 111585 142361
rect 111619 142327 111921 142361
rect 111955 142327 112257 142361
rect 112291 142327 112593 142361
rect 112627 142327 112920 142361
rect 112972 142327 113265 142361
rect 113299 142327 113601 142361
rect 113635 142327 113937 142361
rect 113971 142327 114273 142361
rect 114307 142327 114600 142361
rect 114652 142327 114945 142361
rect 114979 142327 115281 142361
rect 115315 142327 115617 142361
rect 115651 142327 115953 142361
rect 115987 142327 116280 142361
rect 116332 142327 116625 142361
rect 116659 142327 116961 142361
rect 116995 142327 117297 142361
rect 117331 142327 117633 142361
rect 117667 142327 117960 142361
rect 118012 142327 118305 142361
rect 118339 142327 118641 142361
rect 118675 142327 118977 142361
rect 119011 142327 119313 142361
rect 119347 142327 119640 142361
rect 119692 142327 119985 142361
rect 120019 142327 120321 142361
rect 120355 142327 120657 142361
rect 120691 142327 120993 142361
rect 121027 142327 121320 142361
rect 121372 142327 121665 142361
rect 121699 142327 122001 142361
rect 122035 142327 122337 142361
rect 122371 142327 122673 142361
rect 122707 142327 123000 142361
rect 123052 142327 123345 142361
rect 123379 142327 123681 142361
rect 123715 142327 124017 142361
rect 124051 142327 124353 142361
rect 124387 142327 124680 142361
rect 124732 142327 125025 142361
rect 125059 142327 125361 142361
rect 125395 142327 125697 142361
rect 125731 142327 126033 142361
rect 126067 142327 126360 142361
rect 126412 142327 126705 142361
rect 126739 142327 127041 142361
rect 127075 142327 127377 142361
rect 127411 142327 127713 142361
rect 127747 142327 128040 142361
rect 128092 142327 128385 142361
rect 128419 142327 128721 142361
rect 128755 142327 129057 142361
rect 129091 142327 129393 142361
rect 129427 142327 129720 142361
rect 129772 142327 130065 142361
rect 130099 142327 130401 142361
rect 130435 142327 130737 142361
rect 130771 142327 131073 142361
rect 131107 142327 131400 142361
rect 131452 142327 131745 142361
rect 131779 142327 132081 142361
rect 132115 142327 132417 142361
rect 132451 142327 132753 142361
rect 132787 142327 133080 142361
rect 133132 142327 133425 142361
rect 133459 142327 133761 142361
rect 133795 142327 134097 142361
rect 134131 142327 134433 142361
rect 134467 142327 134760 142361
rect 134812 142327 135105 142361
rect 135139 142327 135441 142361
rect 135475 142327 135777 142361
rect 135811 142327 136113 142361
rect 136147 142327 136440 142361
rect 136492 142327 136785 142361
rect 136819 142327 137121 142361
rect 137155 142327 137457 142361
rect 137491 142327 137793 142361
rect 137827 142327 138120 142361
rect 138172 142327 138465 142361
rect 138499 142327 138801 142361
rect 138835 142327 139137 142361
rect 139171 142327 139473 142361
rect 139507 142327 139800 142361
rect 139852 142327 140145 142361
rect 140179 142327 140481 142361
rect 140515 142327 140817 142361
rect 140851 142327 141153 142361
rect 141187 142327 141480 142361
rect 141532 142327 141825 142361
rect 141859 142327 142161 142361
rect 142195 142327 142497 142361
rect 142531 142327 142833 142361
rect 142867 142327 143160 142361
rect 143212 142327 143505 142361
rect 143539 142327 143841 142361
rect 143875 142327 144177 142361
rect 144211 142327 144513 142361
rect 144547 142327 144840 142361
rect 144892 142327 145185 142361
rect 145219 142327 145521 142361
rect 145555 142327 145857 142361
rect 145891 142327 146193 142361
rect 146227 142327 146520 142361
rect 146572 142327 146865 142361
rect 146899 142327 147201 142361
rect 147235 142327 147537 142361
rect 147571 142327 147873 142361
rect 147907 142327 148200 142361
rect 148252 142327 148545 142361
rect 148579 142327 148881 142361
rect 148915 142327 149217 142361
rect 149251 142327 149553 142361
rect 149587 142327 149880 142361
rect 149932 142327 150225 142361
rect 150259 142327 150561 142361
rect 150595 142327 150897 142361
rect 150931 142327 151233 142361
rect 151267 142327 151560 142361
rect 151612 142327 151905 142361
rect 151939 142327 152241 142361
rect 152275 142327 152577 142361
rect 152611 142327 152913 142361
rect 152947 142327 153240 142361
rect 153292 142327 153585 142361
rect 153619 142327 153921 142361
rect 153955 142327 154257 142361
rect 154291 142327 154593 142361
rect 154627 142327 154920 142361
rect 154972 142327 155265 142361
rect 155299 142327 155601 142361
rect 155635 142327 155937 142361
rect 155971 142327 156273 142361
rect 156307 142327 156600 142361
rect 156652 142327 156945 142361
rect 156979 142327 157281 142361
rect 157315 142327 157617 142361
rect 157651 142327 157953 142361
rect 157987 142327 158280 142361
rect 158332 142327 158625 142361
rect 158659 142327 158961 142361
rect 158995 142327 159297 142361
rect 159331 142327 159633 142361
rect 159667 142327 159960 142361
rect 160012 142327 160305 142361
rect 160339 142327 160641 142361
rect 160675 142327 160977 142361
rect 161011 142327 161313 142361
rect 161347 142327 161640 142361
rect 161692 142327 161985 142361
rect 162019 142327 162321 142361
rect 162355 142327 162657 142361
rect 162691 142327 162993 142361
rect 163027 142327 163320 142361
rect 163372 142327 163665 142361
rect 163699 142327 164001 142361
rect 164035 142327 164337 142361
rect 164371 142327 164673 142361
rect 164707 142327 165000 142361
rect 165052 142327 165345 142361
rect 165379 142327 165681 142361
rect 165715 142327 166017 142361
rect 166051 142327 166353 142361
rect 166387 142327 166680 142361
rect 166732 142327 167025 142361
rect 167059 142327 167361 142361
rect 167395 142327 167697 142361
rect 167731 142327 168033 142361
rect 168067 142327 168360 142361
rect 168412 142327 168705 142361
rect 168739 142327 169041 142361
rect 169075 142327 169377 142361
rect 169411 142327 169713 142361
rect 169747 142327 170040 142361
rect 170092 142327 170385 142361
rect 170419 142327 170721 142361
rect 170755 142327 171057 142361
rect 171091 142327 171393 142361
rect 171427 142327 171720 142361
rect 171772 142327 172065 142361
rect 172099 142327 172401 142361
rect 172435 142327 172737 142361
rect 172771 142327 173073 142361
rect 173107 142327 173400 142361
rect 173452 142327 173745 142361
rect 173779 142327 174081 142361
rect 174115 142327 174417 142361
rect 174451 142327 174753 142361
rect 174787 142327 175080 142361
rect 175132 142327 175425 142361
rect 175459 142327 175761 142361
rect 175795 142327 176097 142361
rect 176131 142327 176433 142361
rect 176467 142327 176760 142361
rect 176812 142327 177105 142361
rect 177139 142327 177441 142361
rect 177475 142327 177777 142361
rect 177811 142327 178113 142361
rect 178147 142327 178440 142361
rect 178492 142327 178785 142361
rect 178819 142327 179121 142361
rect 179155 142327 179457 142361
rect 179491 142327 179793 142361
rect 179827 142327 180120 142361
rect 180172 142327 180465 142361
rect 180499 142327 180801 142361
rect 180835 142327 181137 142361
rect 181171 142327 181473 142361
rect 181507 142327 181800 142361
rect 181852 142327 182145 142361
rect 182179 142327 182481 142361
rect 182515 142327 182817 142361
rect 182851 142327 183153 142361
rect 183187 142327 183480 142361
rect 183532 142327 183825 142361
rect 183859 142327 184161 142361
rect 184195 142327 184497 142361
rect 184531 142327 184833 142361
rect 184867 142327 185160 142361
rect 185212 142327 185505 142361
rect 185539 142327 185841 142361
rect 185875 142327 186177 142361
rect 186211 142327 186513 142361
rect 186547 142327 186840 142361
rect 186892 142327 187185 142361
rect 187219 142327 187521 142361
rect 187555 142327 187857 142361
rect 187891 142327 188193 142361
rect 188227 142327 188520 142361
rect 188572 142327 188865 142361
rect 188899 142327 189201 142361
rect 189235 142327 189537 142361
rect 189571 142327 189873 142361
rect 189907 142327 190200 142361
rect 190252 142327 190545 142361
rect 190579 142327 190881 142361
rect 190915 142327 191217 142361
rect 191251 142327 191553 142361
rect 191587 142327 191880 142361
rect 191932 142327 192225 142361
rect 192259 142327 192561 142361
rect 192595 142327 192897 142361
rect 192931 142327 193233 142361
rect 193267 142327 193560 142361
rect 193612 142327 193905 142361
rect 193939 142327 194241 142361
rect 194275 142327 194577 142361
rect 194611 142327 194913 142361
rect 194947 142327 195240 142361
rect 195292 142327 195585 142361
rect 195619 142327 195921 142361
rect 195955 142327 196257 142361
rect 196291 142327 196593 142361
rect 196627 142327 196920 142361
rect 196972 142327 197265 142361
rect 197299 142327 197601 142361
rect 197635 142327 197937 142361
rect 197971 142327 198273 142361
rect 198307 142327 198600 142361
rect 198652 142327 198945 142361
rect 198979 142327 199281 142361
rect 199315 142327 199617 142361
rect 199651 142327 199953 142361
rect 199987 142327 200280 142361
rect 200332 142327 200625 142361
rect 200659 142327 200961 142361
rect 200995 142327 201297 142361
rect 201331 142327 201633 142361
rect 201667 142327 201960 142361
rect 202012 142327 202305 142361
rect 202339 142327 202641 142361
rect 202675 142327 202977 142361
rect 203011 142327 203313 142361
rect 203347 142327 203640 142361
rect 203692 142327 203985 142361
rect 204019 142327 204321 142361
rect 204355 142327 204657 142361
rect 204691 142327 204993 142361
rect 205027 142327 205320 142361
rect 205372 142327 205665 142361
rect 205699 142327 206001 142361
rect 206035 142327 206337 142361
rect 206371 142327 206673 142361
rect 206707 142327 207000 142361
rect 207052 142327 207345 142361
rect 207379 142327 207681 142361
rect 207715 142327 208017 142361
rect 208051 142327 208353 142361
rect 208387 142327 208680 142361
rect 208732 142327 209025 142361
rect 209059 142327 209361 142361
rect 209395 142327 209697 142361
rect 209731 142327 210033 142361
rect 210067 142327 210360 142361
rect 210412 142327 210705 142361
rect 210739 142327 211041 142361
rect 211075 142327 211377 142361
rect 211411 142327 211713 142361
rect 211747 142327 212040 142361
rect 212092 142327 212385 142361
rect 212419 142327 212721 142361
rect 212755 142327 213057 142361
rect 213091 142327 213393 142361
rect 213427 142327 213720 142361
rect 213772 142327 214065 142361
rect 214099 142327 214401 142361
rect 214435 142327 214737 142361
rect 214771 142327 215073 142361
rect 215107 142327 215400 142361
rect 215452 142327 215745 142361
rect 215779 142327 216081 142361
rect 216115 142327 216417 142361
rect 216451 142327 217048 142361
rect 2092 142318 3720 142327
rect 3772 142318 5400 142327
rect 5452 142318 7080 142327
rect 7132 142318 8760 142327
rect 8812 142318 10440 142327
rect 10492 142318 12120 142327
rect 12172 142318 13800 142327
rect 13852 142318 15480 142327
rect 15532 142318 17160 142327
rect 17212 142318 18840 142327
rect 18892 142318 20520 142327
rect 20572 142318 22200 142327
rect 22252 142318 23880 142327
rect 23932 142318 25560 142327
rect 25612 142318 27240 142327
rect 27292 142318 28920 142327
rect 28972 142318 30600 142327
rect 30652 142318 32280 142327
rect 32332 142318 33960 142327
rect 34012 142318 35640 142327
rect 35692 142318 37320 142327
rect 37372 142318 39000 142327
rect 39052 142318 40680 142327
rect 40732 142318 42360 142327
rect 42412 142318 44040 142327
rect 44092 142318 45720 142327
rect 45772 142318 47400 142327
rect 47452 142318 49080 142327
rect 49132 142318 50760 142327
rect 50812 142318 52440 142327
rect 52492 142318 54120 142327
rect 54172 142318 55800 142327
rect 55852 142318 57480 142327
rect 57532 142318 59160 142327
rect 59212 142318 60840 142327
rect 60892 142318 62520 142327
rect 62572 142318 64200 142327
rect 64252 142318 65880 142327
rect 65932 142318 67560 142327
rect 67612 142318 69240 142327
rect 69292 142318 70920 142327
rect 70972 142318 72600 142327
rect 72652 142318 74280 142327
rect 74332 142318 75960 142327
rect 76012 142318 77640 142327
rect 77692 142318 79320 142327
rect 79372 142318 81000 142327
rect 81052 142318 82680 142327
rect 82732 142318 84360 142327
rect 84412 142318 86040 142327
rect 86092 142318 87720 142327
rect 87772 142318 89400 142327
rect 89452 142318 91080 142327
rect 91132 142318 92760 142327
rect 92812 142318 94440 142327
rect 94492 142318 96120 142327
rect 96172 142318 97800 142327
rect 97852 142318 99480 142327
rect 99532 142318 101160 142327
rect 101212 142318 102840 142327
rect 102892 142318 104520 142327
rect 104572 142318 106200 142327
rect 106252 142318 107880 142327
rect 107932 142318 109560 142327
rect 109612 142318 111240 142327
rect 111292 142318 112920 142327
rect 112972 142318 114600 142327
rect 114652 142318 116280 142327
rect 116332 142318 117960 142327
rect 118012 142318 119640 142327
rect 119692 142318 121320 142327
rect 121372 142318 123000 142327
rect 123052 142318 124680 142327
rect 124732 142318 126360 142327
rect 126412 142318 128040 142327
rect 128092 142318 129720 142327
rect 129772 142318 131400 142327
rect 131452 142318 133080 142327
rect 133132 142318 134760 142327
rect 134812 142318 136440 142327
rect 136492 142318 138120 142327
rect 138172 142318 139800 142327
rect 139852 142318 141480 142327
rect 141532 142318 143160 142327
rect 143212 142318 144840 142327
rect 144892 142318 146520 142327
rect 146572 142318 148200 142327
rect 148252 142318 149880 142327
rect 149932 142318 151560 142327
rect 151612 142318 153240 142327
rect 153292 142318 154920 142327
rect 154972 142318 156600 142327
rect 156652 142318 158280 142327
rect 158332 142318 159960 142327
rect 160012 142318 161640 142327
rect 161692 142318 163320 142327
rect 163372 142318 165000 142327
rect 165052 142318 166680 142327
rect 166732 142318 168360 142327
rect 168412 142318 170040 142327
rect 170092 142318 171720 142327
rect 171772 142318 173400 142327
rect 173452 142318 175080 142327
rect 175132 142318 176760 142327
rect 176812 142318 178440 142327
rect 178492 142318 180120 142327
rect 180172 142318 181800 142327
rect 181852 142318 183480 142327
rect 183532 142318 185160 142327
rect 185212 142318 186840 142327
rect 186892 142318 188520 142327
rect 188572 142318 190200 142327
rect 190252 142318 191880 142327
rect 191932 142318 193560 142327
rect 193612 142318 195240 142327
rect 195292 142318 196920 142327
rect 196972 142318 198600 142327
rect 198652 142318 200280 142327
rect 200332 142318 201960 142327
rect 202012 142318 203640 142327
rect 203692 142318 205320 142327
rect 205372 142318 207000 142327
rect 207052 142318 208680 142327
rect 208732 142318 210360 142327
rect 210412 142318 212040 142327
rect 212092 142318 213720 142327
rect 213772 142318 215400 142327
rect 215452 142318 217048 142327
rect 1618 142232 217048 142318
rect 1698 141934 1704 141986
rect 1756 141934 1762 141986
rect 216904 141934 216910 141986
rect 216962 141934 216968 141986
rect 1698 141598 1704 141650
rect 1756 141598 1762 141650
rect 216904 141598 216910 141650
rect 216962 141598 216968 141650
rect 1698 141262 1704 141314
rect 1756 141262 1762 141314
rect 216904 141262 216910 141314
rect 216962 141262 216968 141314
rect 1698 140926 1704 140978
rect 1756 140926 1762 140978
rect 216904 140926 216910 140978
rect 216962 140926 216968 140978
rect 1698 140590 1704 140642
rect 1756 140590 1762 140642
rect 216904 140590 216910 140642
rect 216962 140590 216968 140642
rect 1698 140254 1704 140306
rect 1756 140254 1762 140306
rect 216904 140254 216910 140306
rect 216962 140254 216968 140306
rect 1698 139918 1704 139970
rect 1756 139918 1762 139970
rect 216904 139918 216910 139970
rect 216962 139918 216968 139970
rect 1698 139582 1704 139634
rect 1756 139582 1762 139634
rect 216904 139582 216910 139634
rect 216962 139582 216968 139634
rect 1698 139246 1704 139298
rect 1756 139246 1762 139298
rect 216904 139246 216910 139298
rect 216962 139246 216968 139298
rect 1698 138910 1704 138962
rect 1756 138910 1762 138962
rect 216904 138910 216910 138962
rect 216962 138910 216968 138962
rect 1698 138574 1704 138626
rect 1756 138574 1762 138626
rect 216904 138574 216910 138626
rect 216962 138574 216968 138626
rect 1698 138238 1704 138290
rect 1756 138238 1762 138290
rect 216904 138238 216910 138290
rect 216962 138238 216968 138290
rect 1698 137902 1704 137954
rect 1756 137902 1762 137954
rect 216904 137902 216910 137954
rect 216962 137902 216968 137954
rect 1698 137566 1704 137618
rect 1756 137566 1762 137618
rect 216904 137566 216910 137618
rect 216962 137566 216968 137618
rect 1698 137230 1704 137282
rect 1756 137230 1762 137282
rect 216904 137230 216910 137282
rect 216962 137230 216968 137282
rect 1698 136894 1704 136946
rect 1756 136894 1762 136946
rect 216904 136894 216910 136946
rect 216962 136894 216968 136946
rect 1698 136558 1704 136610
rect 1756 136558 1762 136610
rect 216904 136558 216910 136610
rect 216962 136558 216968 136610
rect 1698 136222 1704 136274
rect 1756 136222 1762 136274
rect 216904 136222 216910 136274
rect 216962 136222 216968 136274
rect 1698 135886 1704 135938
rect 1756 135886 1762 135938
rect 216904 135886 216910 135938
rect 216962 135886 216968 135938
rect 1698 135550 1704 135602
rect 1756 135550 1762 135602
rect 216904 135550 216910 135602
rect 216962 135550 216968 135602
rect 1698 135214 1704 135266
rect 1756 135214 1762 135266
rect 216904 135214 216910 135266
rect 216962 135214 216968 135266
rect 1698 134878 1704 134930
rect 1756 134878 1762 134930
rect 216904 134878 216910 134930
rect 216962 134878 216968 134930
rect 1698 134542 1704 134594
rect 1756 134542 1762 134594
rect 216904 134542 216910 134594
rect 216962 134542 216968 134594
rect 1698 134206 1704 134258
rect 1756 134206 1762 134258
rect 216904 134206 216910 134258
rect 216962 134206 216968 134258
rect 1698 133870 1704 133922
rect 1756 133870 1762 133922
rect 216904 133870 216910 133922
rect 216962 133870 216968 133922
rect 1698 133534 1704 133586
rect 1756 133534 1762 133586
rect 216904 133534 216910 133586
rect 216962 133534 216968 133586
rect 1698 133198 1704 133250
rect 1756 133198 1762 133250
rect 216904 133198 216910 133250
rect 216962 133198 216968 133250
rect 29556 133040 29562 133092
rect 29614 133040 29620 133092
rect 34548 133040 34554 133092
rect 34606 133040 34612 133092
rect 39540 133040 39546 133092
rect 39598 133040 39604 133092
rect 44532 133040 44538 133092
rect 44590 133040 44596 133092
rect 49524 133040 49530 133092
rect 49582 133040 49588 133092
rect 54516 133040 54522 133092
rect 54574 133040 54580 133092
rect 59508 133040 59514 133092
rect 59566 133040 59572 133092
rect 64500 133040 64506 133092
rect 64558 133040 64564 133092
rect 69492 133040 69498 133092
rect 69550 133040 69556 133092
rect 74484 133040 74490 133092
rect 74542 133040 74548 133092
rect 79476 133040 79482 133092
rect 79534 133040 79540 133092
rect 84468 133040 84474 133092
rect 84526 133040 84532 133092
rect 89460 133040 89466 133092
rect 89518 133040 89524 133092
rect 94452 133040 94458 133092
rect 94510 133040 94516 133092
rect 99444 133040 99450 133092
rect 99502 133040 99508 133092
rect 104436 133040 104442 133092
rect 104494 133040 104500 133092
rect 109428 133040 109434 133092
rect 109486 133040 109492 133092
rect 114420 133040 114426 133092
rect 114478 133040 114484 133092
rect 119412 133040 119418 133092
rect 119470 133040 119476 133092
rect 124404 133040 124410 133092
rect 124462 133040 124468 133092
rect 129396 133040 129402 133092
rect 129454 133040 129460 133092
rect 134388 133040 134394 133092
rect 134446 133040 134452 133092
rect 139380 133040 139386 133092
rect 139438 133040 139444 133092
rect 144372 133040 144378 133092
rect 144430 133040 144436 133092
rect 149364 133040 149370 133092
rect 149422 133040 149428 133092
rect 154356 133040 154362 133092
rect 154414 133040 154420 133092
rect 159348 133040 159354 133092
rect 159406 133040 159412 133092
rect 164340 133040 164346 133092
rect 164398 133040 164404 133092
rect 169332 133040 169338 133092
rect 169390 133040 169396 133092
rect 174324 133040 174330 133092
rect 174382 133040 174388 133092
rect 179316 133040 179322 133092
rect 179374 133040 179380 133092
rect 184308 133040 184314 133092
rect 184366 133040 184372 133092
rect 1698 132862 1704 132914
rect 1756 132862 1762 132914
rect 216904 132862 216910 132914
rect 216962 132862 216968 132914
rect 1698 132526 1704 132578
rect 1756 132526 1762 132578
rect 216904 132526 216910 132578
rect 216962 132526 216968 132578
rect 1698 132190 1704 132242
rect 1756 132190 1762 132242
rect 216904 132190 216910 132242
rect 216962 132190 216968 132242
rect 1698 131854 1704 131906
rect 1756 131854 1762 131906
rect 216904 131854 216910 131906
rect 216962 131854 216968 131906
rect 1698 131518 1704 131570
rect 1756 131518 1762 131570
rect 216904 131518 216910 131570
rect 216962 131518 216968 131570
rect 1698 131182 1704 131234
rect 1756 131182 1762 131234
rect 216904 131182 216910 131234
rect 216962 131182 216968 131234
rect 1698 130846 1704 130898
rect 1756 130846 1762 130898
rect 216904 130846 216910 130898
rect 216962 130846 216968 130898
rect 1698 130510 1704 130562
rect 1756 130510 1762 130562
rect 216904 130510 216910 130562
rect 216962 130510 216968 130562
rect 1698 130174 1704 130226
rect 1756 130174 1762 130226
rect 216904 130174 216910 130226
rect 216962 130174 216968 130226
rect 1698 129838 1704 129890
rect 1756 129838 1762 129890
rect 216904 129838 216910 129890
rect 216962 129838 216968 129890
rect 1698 129502 1704 129554
rect 1756 129502 1762 129554
rect 216904 129502 216910 129554
rect 216962 129502 216968 129554
rect 1698 129166 1704 129218
rect 1756 129166 1762 129218
rect 216904 129166 216910 129218
rect 216962 129166 216968 129218
rect 1698 128830 1704 128882
rect 1756 128830 1762 128882
rect 216904 128830 216910 128882
rect 216962 128830 216968 128882
rect 1698 128494 1704 128546
rect 1756 128494 1762 128546
rect 216904 128494 216910 128546
rect 216962 128494 216968 128546
rect 1698 128158 1704 128210
rect 1756 128158 1762 128210
rect 216904 128158 216910 128210
rect 216962 128158 216968 128210
rect 1698 127822 1704 127874
rect 1756 127822 1762 127874
rect 216904 127822 216910 127874
rect 216962 127822 216968 127874
rect 1698 127486 1704 127538
rect 1756 127486 1762 127538
rect 216904 127486 216910 127538
rect 216962 127486 216968 127538
rect 1698 127150 1704 127202
rect 1756 127150 1762 127202
rect 216904 127150 216910 127202
rect 216962 127150 216968 127202
rect 1698 126814 1704 126866
rect 1756 126814 1762 126866
rect 216904 126814 216910 126866
rect 216962 126814 216968 126866
rect 1698 126478 1704 126530
rect 1756 126478 1762 126530
rect 216904 126478 216910 126530
rect 216962 126478 216968 126530
rect 1698 126142 1704 126194
rect 1756 126142 1762 126194
rect 216904 126142 216910 126194
rect 216962 126142 216968 126194
rect 1698 125806 1704 125858
rect 1756 125806 1762 125858
rect 216904 125806 216910 125858
rect 216962 125806 216968 125858
rect 1698 125470 1704 125522
rect 1756 125470 1762 125522
rect 216904 125470 216910 125522
rect 216962 125470 216968 125522
rect 1698 125134 1704 125186
rect 1756 125134 1762 125186
rect 216904 125134 216910 125186
rect 216962 125134 216968 125186
rect 1698 124798 1704 124850
rect 1756 124798 1762 124850
rect 216904 124798 216910 124850
rect 216962 124798 216968 124850
rect 1698 124462 1704 124514
rect 1756 124462 1762 124514
rect 216904 124462 216910 124514
rect 216962 124462 216968 124514
rect 1698 124126 1704 124178
rect 1756 124126 1762 124178
rect 216904 124126 216910 124178
rect 216962 124126 216968 124178
rect 1698 123790 1704 123842
rect 1756 123790 1762 123842
rect 216904 123790 216910 123842
rect 216962 123790 216968 123842
rect 1698 123454 1704 123506
rect 1756 123454 1762 123506
rect 216904 123454 216910 123506
rect 216962 123454 216968 123506
rect 1698 123118 1704 123170
rect 1756 123118 1762 123170
rect 216904 123118 216910 123170
rect 216962 123118 216968 123170
rect 1698 122782 1704 122834
rect 1756 122782 1762 122834
rect 216904 122782 216910 122834
rect 216962 122782 216968 122834
rect 1698 122446 1704 122498
rect 1756 122446 1762 122498
rect 216904 122446 216910 122498
rect 216962 122446 216968 122498
rect 1698 122110 1704 122162
rect 1756 122110 1762 122162
rect 216904 122110 216910 122162
rect 216962 122110 216968 122162
rect 1698 121774 1704 121826
rect 1756 121774 1762 121826
rect 216904 121774 216910 121826
rect 216962 121774 216968 121826
rect 1698 121438 1704 121490
rect 1756 121438 1762 121490
rect 216904 121438 216910 121490
rect 216962 121438 216968 121490
rect 1698 121102 1704 121154
rect 1756 121102 1762 121154
rect 216904 121102 216910 121154
rect 216962 121102 216968 121154
rect 1698 120766 1704 120818
rect 1756 120766 1762 120818
rect 216904 120766 216910 120818
rect 216962 120766 216968 120818
rect 1698 120430 1704 120482
rect 1756 120430 1762 120482
rect 216904 120430 216910 120482
rect 216962 120430 216968 120482
rect 1698 120094 1704 120146
rect 1756 120094 1762 120146
rect 216904 120094 216910 120146
rect 216962 120094 216968 120146
rect 1698 119758 1704 119810
rect 1756 119758 1762 119810
rect 216904 119758 216910 119810
rect 216962 119758 216968 119810
rect 1698 119422 1704 119474
rect 1756 119422 1762 119474
rect 216904 119422 216910 119474
rect 216962 119422 216968 119474
rect 1698 119086 1704 119138
rect 1756 119086 1762 119138
rect 216904 119086 216910 119138
rect 216962 119086 216968 119138
rect 1698 118750 1704 118802
rect 1756 118750 1762 118802
rect 216904 118750 216910 118802
rect 216962 118750 216968 118802
rect 1698 118414 1704 118466
rect 1756 118414 1762 118466
rect 216904 118414 216910 118466
rect 216962 118414 216968 118466
rect 1698 118078 1704 118130
rect 1756 118078 1762 118130
rect 216904 118078 216910 118130
rect 216962 118078 216968 118130
rect 1698 117742 1704 117794
rect 1756 117742 1762 117794
rect 216904 117742 216910 117794
rect 216962 117742 216968 117794
rect 1698 117406 1704 117458
rect 1756 117406 1762 117458
rect 216904 117406 216910 117458
rect 216962 117406 216968 117458
rect 1698 117070 1704 117122
rect 1756 117070 1762 117122
rect 216904 117070 216910 117122
rect 216962 117070 216968 117122
rect 1698 116734 1704 116786
rect 1756 116734 1762 116786
rect 216904 116734 216910 116786
rect 216962 116734 216968 116786
rect 1698 116398 1704 116450
rect 1756 116398 1762 116450
rect 216904 116398 216910 116450
rect 216962 116398 216968 116450
rect 1698 116062 1704 116114
rect 1756 116062 1762 116114
rect 216904 116062 216910 116114
rect 216962 116062 216968 116114
rect 1698 115726 1704 115778
rect 1756 115726 1762 115778
rect 216904 115726 216910 115778
rect 216962 115726 216968 115778
rect 1698 115390 1704 115442
rect 1756 115390 1762 115442
rect 216904 115390 216910 115442
rect 216962 115390 216968 115442
rect 1698 115054 1704 115106
rect 1756 115054 1762 115106
rect 216904 115054 216910 115106
rect 216962 115054 216968 115106
rect 1698 114718 1704 114770
rect 1756 114718 1762 114770
rect 216904 114718 216910 114770
rect 216962 114718 216968 114770
rect 1698 114382 1704 114434
rect 1756 114382 1762 114434
rect 216904 114382 216910 114434
rect 216962 114382 216968 114434
rect 1698 114046 1704 114098
rect 1756 114046 1762 114098
rect 216904 114046 216910 114098
rect 216962 114046 216968 114098
rect 1698 113710 1704 113762
rect 1756 113710 1762 113762
rect 216904 113710 216910 113762
rect 216962 113710 216968 113762
rect 1698 113374 1704 113426
rect 1756 113374 1762 113426
rect 216904 113374 216910 113426
rect 216962 113374 216968 113426
rect 1698 113038 1704 113090
rect 1756 113038 1762 113090
rect 216904 113038 216910 113090
rect 216962 113038 216968 113090
rect 1698 112702 1704 112754
rect 1756 112702 1762 112754
rect 216904 112702 216910 112754
rect 216962 112702 216968 112754
rect 1698 112366 1704 112418
rect 1756 112366 1762 112418
rect 216904 112366 216910 112418
rect 216962 112366 216968 112418
rect 1698 112030 1704 112082
rect 1756 112030 1762 112082
rect 216904 112030 216910 112082
rect 216962 112030 216968 112082
rect 1698 111694 1704 111746
rect 1756 111694 1762 111746
rect 216904 111694 216910 111746
rect 216962 111694 216968 111746
rect 1698 111358 1704 111410
rect 1756 111358 1762 111410
rect 216904 111358 216910 111410
rect 216962 111358 216968 111410
rect 1698 111022 1704 111074
rect 1756 111022 1762 111074
rect 216904 111022 216910 111074
rect 216962 111022 216968 111074
rect 1698 110686 1704 110738
rect 1756 110686 1762 110738
rect 216904 110686 216910 110738
rect 216962 110686 216968 110738
rect 1698 110350 1704 110402
rect 1756 110350 1762 110402
rect 216904 110350 216910 110402
rect 216962 110350 216968 110402
rect 1698 110014 1704 110066
rect 1756 110014 1762 110066
rect 216904 110014 216910 110066
rect 216962 110014 216968 110066
rect 1698 109678 1704 109730
rect 1756 109678 1762 109730
rect 216904 109678 216910 109730
rect 216962 109678 216968 109730
rect 1698 109342 1704 109394
rect 1756 109342 1762 109394
rect 216904 109342 216910 109394
rect 216962 109342 216968 109394
rect 1698 109006 1704 109058
rect 1756 109006 1762 109058
rect 216904 109006 216910 109058
rect 216962 109006 216968 109058
rect 1698 108670 1704 108722
rect 1756 108670 1762 108722
rect 216904 108670 216910 108722
rect 216962 108670 216968 108722
rect 1698 108334 1704 108386
rect 1756 108334 1762 108386
rect 216904 108334 216910 108386
rect 216962 108334 216968 108386
rect 1698 107998 1704 108050
rect 1756 107998 1762 108050
rect 216904 107998 216910 108050
rect 216962 107998 216968 108050
rect 1698 107662 1704 107714
rect 1756 107662 1762 107714
rect 216904 107662 216910 107714
rect 216962 107662 216968 107714
rect 1698 107326 1704 107378
rect 1756 107326 1762 107378
rect 216904 107326 216910 107378
rect 216962 107326 216968 107378
rect 1698 106990 1704 107042
rect 1756 106990 1762 107042
rect 216904 106990 216910 107042
rect 216962 106990 216968 107042
rect 1698 106654 1704 106706
rect 1756 106654 1762 106706
rect 216904 106654 216910 106706
rect 216962 106654 216968 106706
rect 1698 106318 1704 106370
rect 1756 106318 1762 106370
rect 216904 106318 216910 106370
rect 216962 106318 216968 106370
rect 1698 105982 1704 106034
rect 1756 105982 1762 106034
rect 216904 105982 216910 106034
rect 216962 105982 216968 106034
rect 1698 105646 1704 105698
rect 1756 105646 1762 105698
rect 216904 105646 216910 105698
rect 216962 105646 216968 105698
rect 1698 105310 1704 105362
rect 1756 105310 1762 105362
rect 216904 105310 216910 105362
rect 216962 105310 216968 105362
rect 1698 104974 1704 105026
rect 1756 104974 1762 105026
rect 216904 104974 216910 105026
rect 216962 104974 216968 105026
rect 1698 104638 1704 104690
rect 1756 104638 1762 104690
rect 216904 104638 216910 104690
rect 216962 104638 216968 104690
rect 1698 104302 1704 104354
rect 1756 104302 1762 104354
rect 216904 104302 216910 104354
rect 216962 104302 216968 104354
rect 1698 103966 1704 104018
rect 1756 103966 1762 104018
rect 216904 103966 216910 104018
rect 216962 103966 216968 104018
rect 1698 103630 1704 103682
rect 1756 103630 1762 103682
rect 216904 103630 216910 103682
rect 216962 103630 216968 103682
rect 1698 103294 1704 103346
rect 1756 103294 1762 103346
rect 216904 103294 216910 103346
rect 216962 103294 216968 103346
rect 1698 102958 1704 103010
rect 1756 102958 1762 103010
rect 216904 102958 216910 103010
rect 216962 102958 216968 103010
rect 1698 102622 1704 102674
rect 1756 102622 1762 102674
rect 216904 102622 216910 102674
rect 216962 102622 216968 102674
rect 1698 102286 1704 102338
rect 1756 102286 1762 102338
rect 216904 102286 216910 102338
rect 216962 102286 216968 102338
rect 1698 101950 1704 102002
rect 1756 101950 1762 102002
rect 216904 101950 216910 102002
rect 216962 101950 216968 102002
rect 1698 101614 1704 101666
rect 1756 101614 1762 101666
rect 216904 101614 216910 101666
rect 216962 101614 216968 101666
rect 1698 101278 1704 101330
rect 1756 101278 1762 101330
rect 216904 101278 216910 101330
rect 216962 101278 216968 101330
rect 1698 100942 1704 100994
rect 1756 100942 1762 100994
rect 216904 100942 216910 100994
rect 216962 100942 216968 100994
rect 1698 100606 1704 100658
rect 1756 100606 1762 100658
rect 216904 100606 216910 100658
rect 216962 100606 216968 100658
rect 1698 100270 1704 100322
rect 1756 100270 1762 100322
rect 216904 100270 216910 100322
rect 216962 100270 216968 100322
rect 1698 99934 1704 99986
rect 1756 99934 1762 99986
rect 216904 99934 216910 99986
rect 216962 99934 216968 99986
rect 1698 99598 1704 99650
rect 1756 99598 1762 99650
rect 216904 99598 216910 99650
rect 216962 99598 216968 99650
rect 1698 99262 1704 99314
rect 1756 99262 1762 99314
rect 216904 99262 216910 99314
rect 216962 99262 216968 99314
rect 1698 98926 1704 98978
rect 1756 98926 1762 98978
rect 216904 98926 216910 98978
rect 216962 98926 216968 98978
rect 1698 98590 1704 98642
rect 1756 98590 1762 98642
rect 216904 98590 216910 98642
rect 216962 98590 216968 98642
rect 1698 98254 1704 98306
rect 1756 98254 1762 98306
rect 216904 98254 216910 98306
rect 216962 98254 216968 98306
rect 1698 97918 1704 97970
rect 1756 97918 1762 97970
rect 216904 97918 216910 97970
rect 216962 97918 216968 97970
rect 1698 97582 1704 97634
rect 1756 97582 1762 97634
rect 216904 97582 216910 97634
rect 216962 97582 216968 97634
rect 1698 97246 1704 97298
rect 1756 97246 1762 97298
rect 216904 97246 216910 97298
rect 216962 97246 216968 97298
rect 1698 96910 1704 96962
rect 1756 96910 1762 96962
rect 216904 96910 216910 96962
rect 216962 96910 216968 96962
rect 1698 96574 1704 96626
rect 1756 96574 1762 96626
rect 216904 96574 216910 96626
rect 216962 96574 216968 96626
rect 1698 96238 1704 96290
rect 1756 96238 1762 96290
rect 216904 96238 216910 96290
rect 216962 96238 216968 96290
rect 1698 95902 1704 95954
rect 1756 95902 1762 95954
rect 216904 95902 216910 95954
rect 216962 95902 216968 95954
rect 1698 95566 1704 95618
rect 1756 95566 1762 95618
rect 216904 95566 216910 95618
rect 216962 95566 216968 95618
rect 1698 95230 1704 95282
rect 1756 95230 1762 95282
rect 216904 95230 216910 95282
rect 216962 95230 216968 95282
rect 1698 94894 1704 94946
rect 1756 94894 1762 94946
rect 216904 94894 216910 94946
rect 216962 94894 216968 94946
rect 1698 94558 1704 94610
rect 1756 94558 1762 94610
rect 216904 94558 216910 94610
rect 216962 94558 216968 94610
rect 1698 94222 1704 94274
rect 1756 94222 1762 94274
rect 216904 94222 216910 94274
rect 216962 94222 216968 94274
rect 1698 93886 1704 93938
rect 1756 93886 1762 93938
rect 216904 93886 216910 93938
rect 216962 93886 216968 93938
rect 1698 93550 1704 93602
rect 1756 93550 1762 93602
rect 216904 93550 216910 93602
rect 216962 93550 216968 93602
rect 1698 93214 1704 93266
rect 1756 93214 1762 93266
rect 216904 93214 216910 93266
rect 216962 93214 216968 93266
rect 1698 92878 1704 92930
rect 1756 92878 1762 92930
rect 216904 92878 216910 92930
rect 216962 92878 216968 92930
rect 1698 92542 1704 92594
rect 1756 92542 1762 92594
rect 216904 92542 216910 92594
rect 216962 92542 216968 92594
rect 1698 92206 1704 92258
rect 1756 92206 1762 92258
rect 216904 92206 216910 92258
rect 216962 92206 216968 92258
rect 1698 91870 1704 91922
rect 1756 91870 1762 91922
rect 216904 91870 216910 91922
rect 216962 91870 216968 91922
rect 1698 91534 1704 91586
rect 1756 91534 1762 91586
rect 216904 91534 216910 91586
rect 216962 91534 216968 91586
rect 1698 91198 1704 91250
rect 1756 91198 1762 91250
rect 216904 91198 216910 91250
rect 216962 91198 216968 91250
rect 1698 90862 1704 90914
rect 1756 90862 1762 90914
rect 216904 90862 216910 90914
rect 216962 90862 216968 90914
rect 1698 90526 1704 90578
rect 1756 90526 1762 90578
rect 216904 90526 216910 90578
rect 216962 90526 216968 90578
rect 1698 90190 1704 90242
rect 1756 90190 1762 90242
rect 216904 90190 216910 90242
rect 216962 90190 216968 90242
rect 1698 89854 1704 89906
rect 1756 89854 1762 89906
rect 216904 89854 216910 89906
rect 216962 89854 216968 89906
rect 1698 89518 1704 89570
rect 1756 89518 1762 89570
rect 216904 89518 216910 89570
rect 216962 89518 216968 89570
rect 1698 89182 1704 89234
rect 1756 89182 1762 89234
rect 216904 89182 216910 89234
rect 216962 89182 216968 89234
rect 1698 88846 1704 88898
rect 1756 88846 1762 88898
rect 216904 88846 216910 88898
rect 216962 88846 216968 88898
rect 1698 88510 1704 88562
rect 1756 88510 1762 88562
rect 216904 88510 216910 88562
rect 216962 88510 216968 88562
rect 1698 88174 1704 88226
rect 1756 88174 1762 88226
rect 216904 88174 216910 88226
rect 216962 88174 216968 88226
rect 1698 87838 1704 87890
rect 1756 87838 1762 87890
rect 216904 87838 216910 87890
rect 216962 87838 216968 87890
rect 1698 87502 1704 87554
rect 1756 87502 1762 87554
rect 216904 87502 216910 87554
rect 216962 87502 216968 87554
rect 1698 87166 1704 87218
rect 1756 87166 1762 87218
rect 216904 87166 216910 87218
rect 216962 87166 216968 87218
rect 1698 86830 1704 86882
rect 1756 86830 1762 86882
rect 216904 86830 216910 86882
rect 216962 86830 216968 86882
rect 1698 86494 1704 86546
rect 1756 86494 1762 86546
rect 216904 86494 216910 86546
rect 216962 86494 216968 86546
rect 1698 86158 1704 86210
rect 1756 86158 1762 86210
rect 216904 86158 216910 86210
rect 216962 86158 216968 86210
rect 1698 85822 1704 85874
rect 1756 85822 1762 85874
rect 216904 85822 216910 85874
rect 216962 85822 216968 85874
rect 1698 85486 1704 85538
rect 1756 85486 1762 85538
rect 216904 85486 216910 85538
rect 216962 85486 216968 85538
rect 1698 85150 1704 85202
rect 1756 85150 1762 85202
rect 216904 85150 216910 85202
rect 216962 85150 216968 85202
rect 1698 84814 1704 84866
rect 1756 84814 1762 84866
rect 216904 84814 216910 84866
rect 216962 84814 216968 84866
rect 1698 84478 1704 84530
rect 1756 84478 1762 84530
rect 216904 84478 216910 84530
rect 216962 84478 216968 84530
rect 1698 84142 1704 84194
rect 1756 84142 1762 84194
rect 216904 84142 216910 84194
rect 216962 84142 216968 84194
rect 1698 83806 1704 83858
rect 1756 83806 1762 83858
rect 216904 83806 216910 83858
rect 216962 83806 216968 83858
rect 1698 83470 1704 83522
rect 1756 83470 1762 83522
rect 216904 83470 216910 83522
rect 216962 83470 216968 83522
rect 1698 83134 1704 83186
rect 1756 83134 1762 83186
rect 216904 83134 216910 83186
rect 216962 83134 216968 83186
rect 1698 82798 1704 82850
rect 1756 82798 1762 82850
rect 216904 82798 216910 82850
rect 216962 82798 216968 82850
rect 1698 82462 1704 82514
rect 1756 82462 1762 82514
rect 216904 82462 216910 82514
rect 216962 82462 216968 82514
rect 1698 82126 1704 82178
rect 1756 82126 1762 82178
rect 216904 82126 216910 82178
rect 216962 82126 216968 82178
rect 1698 81790 1704 81842
rect 1756 81790 1762 81842
rect 216904 81790 216910 81842
rect 216962 81790 216968 81842
rect 1698 81454 1704 81506
rect 1756 81454 1762 81506
rect 216904 81454 216910 81506
rect 216962 81454 216968 81506
rect 1698 81118 1704 81170
rect 1756 81118 1762 81170
rect 216904 81118 216910 81170
rect 216962 81118 216968 81170
rect 1698 80782 1704 80834
rect 1756 80782 1762 80834
rect 216904 80782 216910 80834
rect 216962 80782 216968 80834
rect 1698 80446 1704 80498
rect 1756 80446 1762 80498
rect 216904 80446 216910 80498
rect 216962 80446 216968 80498
rect 1698 80110 1704 80162
rect 1756 80110 1762 80162
rect 216904 80110 216910 80162
rect 216962 80110 216968 80162
rect 1698 79774 1704 79826
rect 1756 79774 1762 79826
rect 216904 79774 216910 79826
rect 216962 79774 216968 79826
rect 1698 79438 1704 79490
rect 1756 79438 1762 79490
rect 216904 79438 216910 79490
rect 216962 79438 216968 79490
rect 1698 79102 1704 79154
rect 1756 79102 1762 79154
rect 216904 79102 216910 79154
rect 216962 79102 216968 79154
rect 1698 78766 1704 78818
rect 1756 78766 1762 78818
rect 216904 78766 216910 78818
rect 216962 78766 216968 78818
rect 1698 78430 1704 78482
rect 1756 78430 1762 78482
rect 216904 78430 216910 78482
rect 216962 78430 216968 78482
rect 1698 78094 1704 78146
rect 1756 78094 1762 78146
rect 216904 78094 216910 78146
rect 216962 78094 216968 78146
rect 1698 77758 1704 77810
rect 1756 77758 1762 77810
rect 216904 77758 216910 77810
rect 216962 77758 216968 77810
rect 1698 77422 1704 77474
rect 1756 77422 1762 77474
rect 216904 77422 216910 77474
rect 216962 77422 216968 77474
rect 1698 77086 1704 77138
rect 1756 77086 1762 77138
rect 216904 77086 216910 77138
rect 216962 77086 216968 77138
rect 1698 76750 1704 76802
rect 1756 76750 1762 76802
rect 216904 76750 216910 76802
rect 216962 76750 216968 76802
rect 1698 76414 1704 76466
rect 1756 76414 1762 76466
rect 216904 76414 216910 76466
rect 216962 76414 216968 76466
rect 1698 76078 1704 76130
rect 1756 76078 1762 76130
rect 216904 76078 216910 76130
rect 216962 76078 216968 76130
rect 1698 75742 1704 75794
rect 1756 75742 1762 75794
rect 216904 75742 216910 75794
rect 216962 75742 216968 75794
rect 1698 75406 1704 75458
rect 1756 75406 1762 75458
rect 216904 75406 216910 75458
rect 216962 75406 216968 75458
rect 1698 75070 1704 75122
rect 1756 75070 1762 75122
rect 216904 75070 216910 75122
rect 216962 75070 216968 75122
rect 1698 74734 1704 74786
rect 1756 74734 1762 74786
rect 216904 74734 216910 74786
rect 216962 74734 216968 74786
rect 1698 74398 1704 74450
rect 1756 74398 1762 74450
rect 216904 74398 216910 74450
rect 216962 74398 216968 74450
rect 1698 74062 1704 74114
rect 1756 74062 1762 74114
rect 216904 74062 216910 74114
rect 216962 74062 216968 74114
rect 1698 73726 1704 73778
rect 1756 73726 1762 73778
rect 216904 73726 216910 73778
rect 216962 73726 216968 73778
rect 1698 73390 1704 73442
rect 1756 73390 1762 73442
rect 216904 73390 216910 73442
rect 216962 73390 216968 73442
rect 1698 73054 1704 73106
rect 1756 73054 1762 73106
rect 216904 73054 216910 73106
rect 216962 73054 216968 73106
rect 1698 72718 1704 72770
rect 1756 72718 1762 72770
rect 216904 72718 216910 72770
rect 216962 72718 216968 72770
rect 1698 72382 1704 72434
rect 1756 72382 1762 72434
rect 216904 72382 216910 72434
rect 216962 72382 216968 72434
rect 1698 72046 1704 72098
rect 1756 72046 1762 72098
rect 216904 72046 216910 72098
rect 216962 72046 216968 72098
rect 1698 71710 1704 71762
rect 1756 71710 1762 71762
rect 216904 71710 216910 71762
rect 216962 71710 216968 71762
rect 1698 71374 1704 71426
rect 1756 71374 1762 71426
rect 216904 71374 216910 71426
rect 216962 71374 216968 71426
rect 1698 71038 1704 71090
rect 1756 71038 1762 71090
rect 216904 71038 216910 71090
rect 216962 71038 216968 71090
rect 1698 70702 1704 70754
rect 1756 70702 1762 70754
rect 216904 70702 216910 70754
rect 216962 70702 216968 70754
rect 1698 70366 1704 70418
rect 1756 70366 1762 70418
rect 216904 70366 216910 70418
rect 216962 70366 216968 70418
rect 1698 70030 1704 70082
rect 1756 70030 1762 70082
rect 216904 70030 216910 70082
rect 216962 70030 216968 70082
rect 1698 69694 1704 69746
rect 1756 69694 1762 69746
rect 216904 69694 216910 69746
rect 216962 69694 216968 69746
rect 1698 69358 1704 69410
rect 1756 69358 1762 69410
rect 216904 69358 216910 69410
rect 216962 69358 216968 69410
rect 1698 69022 1704 69074
rect 1756 69022 1762 69074
rect 216904 69022 216910 69074
rect 216962 69022 216968 69074
rect 1698 68686 1704 68738
rect 1756 68686 1762 68738
rect 216904 68686 216910 68738
rect 216962 68686 216968 68738
rect 1698 68350 1704 68402
rect 1756 68350 1762 68402
rect 216904 68350 216910 68402
rect 216962 68350 216968 68402
rect 1698 68014 1704 68066
rect 1756 68014 1762 68066
rect 216904 68014 216910 68066
rect 216962 68014 216968 68066
rect 1698 67678 1704 67730
rect 1756 67678 1762 67730
rect 216904 67678 216910 67730
rect 216962 67678 216968 67730
rect 1698 67342 1704 67394
rect 1756 67342 1762 67394
rect 216904 67342 216910 67394
rect 216962 67342 216968 67394
rect 1698 67006 1704 67058
rect 1756 67006 1762 67058
rect 216904 67006 216910 67058
rect 216962 67006 216968 67058
rect 1698 66670 1704 66722
rect 1756 66670 1762 66722
rect 216904 66670 216910 66722
rect 216962 66670 216968 66722
rect 1698 66334 1704 66386
rect 1756 66334 1762 66386
rect 216904 66334 216910 66386
rect 216962 66334 216968 66386
rect 1698 65998 1704 66050
rect 1756 65998 1762 66050
rect 216904 65998 216910 66050
rect 216962 65998 216968 66050
rect 1698 65662 1704 65714
rect 1756 65662 1762 65714
rect 216904 65662 216910 65714
rect 216962 65662 216968 65714
rect 1698 65326 1704 65378
rect 1756 65326 1762 65378
rect 216904 65326 216910 65378
rect 216962 65326 216968 65378
rect 1698 64990 1704 65042
rect 1756 64990 1762 65042
rect 216904 64990 216910 65042
rect 216962 64990 216968 65042
rect 1698 64654 1704 64706
rect 1756 64654 1762 64706
rect 216904 64654 216910 64706
rect 216962 64654 216968 64706
rect 1698 64318 1704 64370
rect 1756 64318 1762 64370
rect 216904 64318 216910 64370
rect 216962 64318 216968 64370
rect 1698 63982 1704 64034
rect 1756 63982 1762 64034
rect 216904 63982 216910 64034
rect 216962 63982 216968 64034
rect 1698 63646 1704 63698
rect 1756 63646 1762 63698
rect 216904 63646 216910 63698
rect 216962 63646 216968 63698
rect 1698 63310 1704 63362
rect 1756 63310 1762 63362
rect 216904 63310 216910 63362
rect 216962 63310 216968 63362
rect 1698 62974 1704 63026
rect 1756 62974 1762 63026
rect 216904 62974 216910 63026
rect 216962 62974 216968 63026
rect 1698 62638 1704 62690
rect 1756 62638 1762 62690
rect 216904 62638 216910 62690
rect 216962 62638 216968 62690
rect 1698 62302 1704 62354
rect 1756 62302 1762 62354
rect 216904 62302 216910 62354
rect 216962 62302 216968 62354
rect 1698 61966 1704 62018
rect 1756 61966 1762 62018
rect 216904 61966 216910 62018
rect 216962 61966 216968 62018
rect 1698 61630 1704 61682
rect 1756 61630 1762 61682
rect 216904 61630 216910 61682
rect 216962 61630 216968 61682
rect 1698 61294 1704 61346
rect 1756 61294 1762 61346
rect 216904 61294 216910 61346
rect 216962 61294 216968 61346
rect 1698 60958 1704 61010
rect 1756 60958 1762 61010
rect 216904 60958 216910 61010
rect 216962 60958 216968 61010
rect 1698 60622 1704 60674
rect 1756 60622 1762 60674
rect 216904 60622 216910 60674
rect 216962 60622 216968 60674
rect 1698 60286 1704 60338
rect 1756 60286 1762 60338
rect 216904 60286 216910 60338
rect 216962 60286 216968 60338
rect 1698 59950 1704 60002
rect 1756 59950 1762 60002
rect 216904 59950 216910 60002
rect 216962 59950 216968 60002
rect 1698 59614 1704 59666
rect 1756 59614 1762 59666
rect 216904 59614 216910 59666
rect 216962 59614 216968 59666
rect 1698 59278 1704 59330
rect 1756 59278 1762 59330
rect 216904 59278 216910 59330
rect 216962 59278 216968 59330
rect 1698 58942 1704 58994
rect 1756 58942 1762 58994
rect 216904 58942 216910 58994
rect 216962 58942 216968 58994
rect 1698 58606 1704 58658
rect 1756 58606 1762 58658
rect 216904 58606 216910 58658
rect 216962 58606 216968 58658
rect 1698 58270 1704 58322
rect 1756 58270 1762 58322
rect 216904 58270 216910 58322
rect 216962 58270 216968 58322
rect 1698 57934 1704 57986
rect 1756 57934 1762 57986
rect 216904 57934 216910 57986
rect 216962 57934 216968 57986
rect 1698 57598 1704 57650
rect 1756 57598 1762 57650
rect 216904 57598 216910 57650
rect 216962 57598 216968 57650
rect 1698 57262 1704 57314
rect 1756 57262 1762 57314
rect 216904 57262 216910 57314
rect 216962 57262 216968 57314
rect 1698 56926 1704 56978
rect 1756 56926 1762 56978
rect 216904 56926 216910 56978
rect 216962 56926 216968 56978
rect 1698 56590 1704 56642
rect 1756 56590 1762 56642
rect 216904 56590 216910 56642
rect 216962 56590 216968 56642
rect 1698 56254 1704 56306
rect 1756 56254 1762 56306
rect 216904 56254 216910 56306
rect 216962 56254 216968 56306
rect 1698 55918 1704 55970
rect 1756 55918 1762 55970
rect 216904 55918 216910 55970
rect 216962 55918 216968 55970
rect 1698 55582 1704 55634
rect 1756 55582 1762 55634
rect 216904 55582 216910 55634
rect 216962 55582 216968 55634
rect 1698 55246 1704 55298
rect 1756 55246 1762 55298
rect 216904 55246 216910 55298
rect 216962 55246 216968 55298
rect 1698 54910 1704 54962
rect 1756 54910 1762 54962
rect 216904 54910 216910 54962
rect 216962 54910 216968 54962
rect 1698 54574 1704 54626
rect 1756 54574 1762 54626
rect 216904 54574 216910 54626
rect 216962 54574 216968 54626
rect 1698 54238 1704 54290
rect 1756 54238 1762 54290
rect 216904 54238 216910 54290
rect 216962 54238 216968 54290
rect 1698 53902 1704 53954
rect 1756 53902 1762 53954
rect 216904 53902 216910 53954
rect 216962 53902 216968 53954
rect 1698 53566 1704 53618
rect 1756 53566 1762 53618
rect 216904 53566 216910 53618
rect 216962 53566 216968 53618
rect 1698 53230 1704 53282
rect 1756 53230 1762 53282
rect 216904 53230 216910 53282
rect 216962 53230 216968 53282
rect 1698 52894 1704 52946
rect 1756 52894 1762 52946
rect 216904 52894 216910 52946
rect 216962 52894 216968 52946
rect 1698 52558 1704 52610
rect 1756 52558 1762 52610
rect 216904 52558 216910 52610
rect 216962 52558 216968 52610
rect 1698 52222 1704 52274
rect 1756 52222 1762 52274
rect 216904 52222 216910 52274
rect 216962 52222 216968 52274
rect 1698 51886 1704 51938
rect 1756 51886 1762 51938
rect 216904 51886 216910 51938
rect 216962 51886 216968 51938
rect 1698 51550 1704 51602
rect 1756 51550 1762 51602
rect 216904 51550 216910 51602
rect 216962 51550 216968 51602
rect 1698 51214 1704 51266
rect 1756 51214 1762 51266
rect 216904 51214 216910 51266
rect 216962 51214 216968 51266
rect 1698 50878 1704 50930
rect 1756 50878 1762 50930
rect 216904 50878 216910 50930
rect 216962 50878 216968 50930
rect 1698 50542 1704 50594
rect 1756 50542 1762 50594
rect 216904 50542 216910 50594
rect 216962 50542 216968 50594
rect 1698 50206 1704 50258
rect 1756 50206 1762 50258
rect 216904 50206 216910 50258
rect 216962 50206 216968 50258
rect 1698 49870 1704 49922
rect 1756 49870 1762 49922
rect 216904 49870 216910 49922
rect 216962 49870 216968 49922
rect 1698 49534 1704 49586
rect 1756 49534 1762 49586
rect 216904 49534 216910 49586
rect 216962 49534 216968 49586
rect 1698 49198 1704 49250
rect 1756 49198 1762 49250
rect 216904 49198 216910 49250
rect 216962 49198 216968 49250
rect 1698 48862 1704 48914
rect 1756 48862 1762 48914
rect 216904 48862 216910 48914
rect 216962 48862 216968 48914
rect 1698 48526 1704 48578
rect 1756 48526 1762 48578
rect 216904 48526 216910 48578
rect 216962 48526 216968 48578
rect 1698 48190 1704 48242
rect 1756 48190 1762 48242
rect 216904 48190 216910 48242
rect 216962 48190 216968 48242
rect 1698 47854 1704 47906
rect 1756 47854 1762 47906
rect 216904 47854 216910 47906
rect 216962 47854 216968 47906
rect 1698 47518 1704 47570
rect 1756 47518 1762 47570
rect 216904 47518 216910 47570
rect 216962 47518 216968 47570
rect 1698 47182 1704 47234
rect 1756 47182 1762 47234
rect 216904 47182 216910 47234
rect 216962 47182 216968 47234
rect 1698 46846 1704 46898
rect 1756 46846 1762 46898
rect 216904 46846 216910 46898
rect 216962 46846 216968 46898
rect 1698 46510 1704 46562
rect 1756 46510 1762 46562
rect 216904 46510 216910 46562
rect 216962 46510 216968 46562
rect 1698 46174 1704 46226
rect 1756 46174 1762 46226
rect 216904 46174 216910 46226
rect 216962 46174 216968 46226
rect 1698 45838 1704 45890
rect 1756 45838 1762 45890
rect 216904 45838 216910 45890
rect 216962 45838 216968 45890
rect 1698 45502 1704 45554
rect 1756 45502 1762 45554
rect 216904 45502 216910 45554
rect 216962 45502 216968 45554
rect 1698 45166 1704 45218
rect 1756 45166 1762 45218
rect 216904 45166 216910 45218
rect 216962 45166 216968 45218
rect 15967 44968 15973 45020
rect 16025 44968 16031 45020
rect 1698 44830 1704 44882
rect 1756 44830 1762 44882
rect 1698 44494 1704 44546
rect 1756 44494 1762 44546
rect 1698 44158 1704 44210
rect 1756 44158 1762 44210
rect 1698 43822 1704 43874
rect 1756 43822 1762 43874
rect 1698 43486 1704 43538
rect 1756 43486 1762 43538
rect 15887 43410 15893 43462
rect 15945 43410 15951 43462
rect 1698 43150 1704 43202
rect 1756 43150 1762 43202
rect 1698 42814 1704 42866
rect 1756 42814 1762 42866
rect 1698 42478 1704 42530
rect 1756 42478 1762 42530
rect 1698 42142 1704 42194
rect 1756 42142 1762 42194
rect 15807 42140 15813 42192
rect 15865 42140 15871 42192
rect 1698 41806 1704 41858
rect 1756 41806 1762 41858
rect 1698 41470 1704 41522
rect 1756 41470 1762 41522
rect 1698 41134 1704 41186
rect 1756 41134 1762 41186
rect 1698 40798 1704 40850
rect 1756 40798 1762 40850
rect 15727 40582 15733 40634
rect 15785 40582 15791 40634
rect 1698 40462 1704 40514
rect 1756 40462 1762 40514
rect 1698 40126 1704 40178
rect 1756 40126 1762 40178
rect 1698 39790 1704 39842
rect 1756 39790 1762 39842
rect 1698 39454 1704 39506
rect 1756 39454 1762 39506
rect 15647 39312 15653 39364
rect 15705 39312 15711 39364
rect 1698 39118 1704 39170
rect 1756 39118 1762 39170
rect 1698 38782 1704 38834
rect 1756 38782 1762 38834
rect 1698 38446 1704 38498
rect 1756 38446 1762 38498
rect 1698 38110 1704 38162
rect 1756 38110 1762 38162
rect 1698 37774 1704 37826
rect 1756 37774 1762 37826
rect 15567 37754 15573 37806
rect 15625 37754 15631 37806
rect 1698 37438 1704 37490
rect 1756 37438 1762 37490
rect 1698 37102 1704 37154
rect 1756 37102 1762 37154
rect 1698 36766 1704 36818
rect 1756 36766 1762 36818
rect 15487 36484 15493 36536
rect 15545 36484 15551 36536
rect 1698 36430 1704 36482
rect 1756 36430 1762 36482
rect 1698 36094 1704 36146
rect 1756 36094 1762 36146
rect 1698 35758 1704 35810
rect 1756 35758 1762 35810
rect 1698 35422 1704 35474
rect 1756 35422 1762 35474
rect 1698 35086 1704 35138
rect 1756 35086 1762 35138
rect 15407 34926 15413 34978
rect 15465 34926 15471 34978
rect 1698 34750 1704 34802
rect 1756 34750 1762 34802
rect 1698 34414 1704 34466
rect 1756 34414 1762 34466
rect 1698 34078 1704 34130
rect 1756 34078 1762 34130
rect 1698 33742 1704 33794
rect 1756 33742 1762 33794
rect 1698 33406 1704 33458
rect 1756 33406 1762 33458
rect 1698 33070 1704 33122
rect 1756 33070 1762 33122
rect 1698 32734 1704 32786
rect 1756 32734 1762 32786
rect 1698 32398 1704 32450
rect 1756 32398 1762 32450
rect 1698 32062 1704 32114
rect 1756 32062 1762 32114
rect 1698 31726 1704 31778
rect 1756 31726 1762 31778
rect 1698 31390 1704 31442
rect 1756 31390 1762 31442
rect 1698 31054 1704 31106
rect 1756 31054 1762 31106
rect 1698 30718 1704 30770
rect 1756 30718 1762 30770
rect 1698 30382 1704 30434
rect 1756 30382 1762 30434
rect 1698 30046 1704 30098
rect 1756 30046 1762 30098
rect 1698 29710 1704 29762
rect 1756 29710 1762 29762
rect 15425 29577 15453 34926
rect 15505 29577 15533 36484
rect 15585 29577 15613 37754
rect 15665 29577 15693 39312
rect 15745 29577 15773 40582
rect 15825 29577 15853 42140
rect 15905 29577 15933 43410
rect 15985 29577 16013 44968
rect 216904 44830 216910 44882
rect 216962 44830 216968 44882
rect 216904 44494 216910 44546
rect 216962 44494 216968 44546
rect 216904 44158 216910 44210
rect 216962 44158 216968 44210
rect 216904 43822 216910 43874
rect 216962 43822 216968 43874
rect 216904 43486 216910 43538
rect 216962 43486 216968 43538
rect 216904 43150 216910 43202
rect 216962 43150 216968 43202
rect 216904 42814 216910 42866
rect 216962 42814 216968 42866
rect 216904 42478 216910 42530
rect 216962 42478 216968 42530
rect 216904 42142 216910 42194
rect 216962 42142 216968 42194
rect 216904 41806 216910 41858
rect 216962 41806 216968 41858
rect 216904 41470 216910 41522
rect 216962 41470 216968 41522
rect 216904 41134 216910 41186
rect 216962 41134 216968 41186
rect 216904 40798 216910 40850
rect 216962 40798 216968 40850
rect 216904 40462 216910 40514
rect 216962 40462 216968 40514
rect 216904 40126 216910 40178
rect 216962 40126 216968 40178
rect 216904 39790 216910 39842
rect 216962 39790 216968 39842
rect 216904 39454 216910 39506
rect 216962 39454 216968 39506
rect 216904 39118 216910 39170
rect 216962 39118 216968 39170
rect 216904 38782 216910 38834
rect 216962 38782 216968 38834
rect 216904 38446 216910 38498
rect 216962 38446 216968 38498
rect 216904 38110 216910 38162
rect 216962 38110 216968 38162
rect 216904 37774 216910 37826
rect 216962 37774 216968 37826
rect 216904 37438 216910 37490
rect 216962 37438 216968 37490
rect 216904 37102 216910 37154
rect 216962 37102 216968 37154
rect 216904 36766 216910 36818
rect 216962 36766 216968 36818
rect 216904 36430 216910 36482
rect 216962 36430 216968 36482
rect 216904 36094 216910 36146
rect 216962 36094 216968 36146
rect 216904 35758 216910 35810
rect 216962 35758 216968 35810
rect 216904 35422 216910 35474
rect 216962 35422 216968 35474
rect 216904 35086 216910 35138
rect 216962 35086 216968 35138
rect 216904 34750 216910 34802
rect 216962 34750 216968 34802
rect 216904 34414 216910 34466
rect 216962 34414 216968 34466
rect 216904 34078 216910 34130
rect 216962 34078 216968 34130
rect 216904 33742 216910 33794
rect 216962 33742 216968 33794
rect 216904 33406 216910 33458
rect 216962 33406 216968 33458
rect 216904 33070 216910 33122
rect 216962 33070 216968 33122
rect 216904 32734 216910 32786
rect 216962 32734 216968 32786
rect 216904 32398 216910 32450
rect 216962 32398 216968 32450
rect 216904 32062 216910 32114
rect 216962 32062 216968 32114
rect 216904 31726 216910 31778
rect 216962 31726 216968 31778
rect 216904 31390 216910 31442
rect 216962 31390 216968 31442
rect 216904 31054 216910 31106
rect 216962 31054 216968 31106
rect 216904 30718 216910 30770
rect 216962 30718 216968 30770
rect 216904 30382 216910 30434
rect 216962 30382 216968 30434
rect 216904 30046 216910 30098
rect 216962 30046 216968 30098
rect 216904 29710 216910 29762
rect 216962 29710 216968 29762
rect 1698 29374 1704 29426
rect 1756 29374 1762 29426
rect 1698 29038 1704 29090
rect 1756 29038 1762 29090
rect 1698 28702 1704 28754
rect 1756 28702 1762 28754
rect 1698 28366 1704 28418
rect 1756 28366 1762 28418
rect 1698 28030 1704 28082
rect 1756 28030 1762 28082
rect 1698 27694 1704 27746
rect 1756 27694 1762 27746
rect 1698 27358 1704 27410
rect 1756 27358 1762 27410
rect 1698 27022 1704 27074
rect 1756 27022 1762 27074
rect 1698 26686 1704 26738
rect 1756 26686 1762 26738
rect 1698 26350 1704 26402
rect 1756 26350 1762 26402
rect 1698 26014 1704 26066
rect 1756 26014 1762 26066
rect 1698 25678 1704 25730
rect 1756 25678 1762 25730
rect 1698 25342 1704 25394
rect 1756 25342 1762 25394
rect 1698 25006 1704 25058
rect 1756 25006 1762 25058
rect 1698 24670 1704 24722
rect 1756 24670 1762 24722
rect 1698 24334 1704 24386
rect 1756 24334 1762 24386
rect 1698 23998 1704 24050
rect 1756 23998 1762 24050
rect 1698 23662 1704 23714
rect 1756 23662 1762 23714
rect 1698 23326 1704 23378
rect 1756 23326 1762 23378
rect 1698 22990 1704 23042
rect 1756 22990 1762 23042
rect 1698 22654 1704 22706
rect 1756 22654 1762 22706
rect 1698 22318 1704 22370
rect 1756 22318 1762 22370
rect 1698 21982 1704 22034
rect 1756 21982 1762 22034
rect 1698 21646 1704 21698
rect 1756 21646 1762 21698
rect 1698 21310 1704 21362
rect 1756 21310 1762 21362
rect 1698 20974 1704 21026
rect 1756 20974 1762 21026
rect 1698 20638 1704 20690
rect 1756 20638 1762 20690
rect 1698 20302 1704 20354
rect 1756 20302 1762 20354
rect 1698 19966 1704 20018
rect 1756 19966 1762 20018
rect 1698 19630 1704 19682
rect 1756 19630 1762 19682
rect 1698 19294 1704 19346
rect 1756 19294 1762 19346
rect 1698 18958 1704 19010
rect 1756 18958 1762 19010
rect 1698 18622 1704 18674
rect 1756 18622 1762 18674
rect 1698 18286 1704 18338
rect 1756 18286 1762 18338
rect 1698 17950 1704 18002
rect 1756 17950 1762 18002
rect 29556 17702 29562 17754
rect 29614 17702 29620 17754
rect 34548 17702 34554 17754
rect 34606 17702 34612 17754
rect 39540 17702 39546 17754
rect 39598 17702 39604 17754
rect 44532 17702 44538 17754
rect 44590 17702 44596 17754
rect 49524 17702 49530 17754
rect 49582 17702 49588 17754
rect 54516 17702 54522 17754
rect 54574 17702 54580 17754
rect 59508 17702 59514 17754
rect 59566 17702 59572 17754
rect 64500 17702 64506 17754
rect 64558 17702 64564 17754
rect 69492 17702 69498 17754
rect 69550 17702 69556 17754
rect 74484 17702 74490 17754
rect 74542 17702 74548 17754
rect 79476 17702 79482 17754
rect 79534 17702 79540 17754
rect 84468 17702 84474 17754
rect 84526 17702 84532 17754
rect 89460 17702 89466 17754
rect 89518 17702 89524 17754
rect 94452 17702 94458 17754
rect 94510 17702 94516 17754
rect 99444 17702 99450 17754
rect 99502 17702 99508 17754
rect 104436 17702 104442 17754
rect 104494 17702 104500 17754
rect 109428 17702 109434 17754
rect 109486 17702 109492 17754
rect 114420 17702 114426 17754
rect 114478 17702 114484 17754
rect 119412 17702 119418 17754
rect 119470 17702 119476 17754
rect 124404 17702 124410 17754
rect 124462 17702 124468 17754
rect 129396 17702 129402 17754
rect 129454 17702 129460 17754
rect 134388 17702 134394 17754
rect 134446 17702 134452 17754
rect 139380 17702 139386 17754
rect 139438 17702 139444 17754
rect 144372 17702 144378 17754
rect 144430 17702 144436 17754
rect 149364 17702 149370 17754
rect 149422 17702 149428 17754
rect 154356 17702 154362 17754
rect 154414 17702 154420 17754
rect 159348 17702 159354 17754
rect 159406 17702 159412 17754
rect 164340 17702 164346 17754
rect 164398 17702 164404 17754
rect 169332 17702 169338 17754
rect 169390 17702 169396 17754
rect 174324 17702 174330 17754
rect 174382 17702 174388 17754
rect 179316 17702 179322 17754
rect 179374 17702 179380 17754
rect 184308 17702 184314 17754
rect 184366 17702 184372 17754
rect 1698 17614 1704 17666
rect 1756 17614 1762 17666
rect 1698 17278 1704 17330
rect 1756 17278 1762 17330
rect 1698 16942 1704 16994
rect 1756 16942 1762 16994
rect 1698 16606 1704 16658
rect 1756 16606 1762 16658
rect 1698 16270 1704 16322
rect 1756 16270 1762 16322
rect 1698 15934 1704 15986
rect 1756 15934 1762 15986
rect 1698 15598 1704 15650
rect 1756 15598 1762 15650
rect 1698 15262 1704 15314
rect 1756 15262 1762 15314
rect 1698 14926 1704 14978
rect 1756 14926 1762 14978
rect 1698 14590 1704 14642
rect 1756 14590 1762 14642
rect 1698 14254 1704 14306
rect 1756 14254 1762 14306
rect 202653 14186 202681 29577
rect 202733 15744 202761 29577
rect 202813 17014 202841 29577
rect 202893 18572 202921 29577
rect 202973 19842 203001 29577
rect 203053 21400 203081 29577
rect 203133 22670 203161 29577
rect 203213 24228 203241 29577
rect 216904 29374 216910 29426
rect 216962 29374 216968 29426
rect 216904 29038 216910 29090
rect 216962 29038 216968 29090
rect 216904 28702 216910 28754
rect 216962 28702 216968 28754
rect 216904 28366 216910 28418
rect 216962 28366 216968 28418
rect 216904 28030 216910 28082
rect 216962 28030 216968 28082
rect 216904 27694 216910 27746
rect 216962 27694 216968 27746
rect 216904 27358 216910 27410
rect 216962 27358 216968 27410
rect 216904 27022 216910 27074
rect 216962 27022 216968 27074
rect 216904 26686 216910 26738
rect 216962 26686 216968 26738
rect 216904 26350 216910 26402
rect 216962 26350 216968 26402
rect 216904 26014 216910 26066
rect 216962 26014 216968 26066
rect 216904 25678 216910 25730
rect 216962 25678 216968 25730
rect 216904 25342 216910 25394
rect 216962 25342 216968 25394
rect 216904 25006 216910 25058
rect 216962 25006 216968 25058
rect 216904 24670 216910 24722
rect 216962 24670 216968 24722
rect 216904 24334 216910 24386
rect 216962 24334 216968 24386
rect 203195 24176 203201 24228
rect 203253 24176 203259 24228
rect 216904 23998 216910 24050
rect 216962 23998 216968 24050
rect 216904 23662 216910 23714
rect 216962 23662 216968 23714
rect 216904 23326 216910 23378
rect 216962 23326 216968 23378
rect 216904 22990 216910 23042
rect 216962 22990 216968 23042
rect 203115 22618 203121 22670
rect 203173 22618 203179 22670
rect 216904 22654 216910 22706
rect 216962 22654 216968 22706
rect 216904 22318 216910 22370
rect 216962 22318 216968 22370
rect 216904 21982 216910 22034
rect 216962 21982 216968 22034
rect 216904 21646 216910 21698
rect 216962 21646 216968 21698
rect 203035 21348 203041 21400
rect 203093 21348 203099 21400
rect 216904 21310 216910 21362
rect 216962 21310 216968 21362
rect 216904 20974 216910 21026
rect 216962 20974 216968 21026
rect 216904 20638 216910 20690
rect 216962 20638 216968 20690
rect 216904 20302 216910 20354
rect 216962 20302 216968 20354
rect 216904 19966 216910 20018
rect 216962 19966 216968 20018
rect 202955 19790 202961 19842
rect 203013 19790 203019 19842
rect 216904 19630 216910 19682
rect 216962 19630 216968 19682
rect 216904 19294 216910 19346
rect 216962 19294 216968 19346
rect 216904 18958 216910 19010
rect 216962 18958 216968 19010
rect 216904 18622 216910 18674
rect 216962 18622 216968 18674
rect 202875 18520 202881 18572
rect 202933 18520 202939 18572
rect 216904 18286 216910 18338
rect 216962 18286 216968 18338
rect 216904 17950 216910 18002
rect 216962 17950 216968 18002
rect 216904 17614 216910 17666
rect 216962 17614 216968 17666
rect 216904 17278 216910 17330
rect 216962 17278 216968 17330
rect 202795 16962 202801 17014
rect 202853 16962 202859 17014
rect 216904 16942 216910 16994
rect 216962 16942 216968 16994
rect 216904 16606 216910 16658
rect 216962 16606 216968 16658
rect 216904 16270 216910 16322
rect 216962 16270 216968 16322
rect 216904 15934 216910 15986
rect 216962 15934 216968 15986
rect 202715 15692 202721 15744
rect 202773 15692 202779 15744
rect 216904 15598 216910 15650
rect 216962 15598 216968 15650
rect 216904 15262 216910 15314
rect 216962 15262 216968 15314
rect 216904 14926 216910 14978
rect 216962 14926 216968 14978
rect 216904 14590 216910 14642
rect 216962 14590 216968 14642
rect 216904 14254 216910 14306
rect 216962 14254 216968 14306
rect 202635 14134 202641 14186
rect 202693 14134 202699 14186
rect 1698 13918 1704 13970
rect 1756 13918 1762 13970
rect 216904 13918 216910 13970
rect 216962 13918 216968 13970
rect 1698 13582 1704 13634
rect 1756 13582 1762 13634
rect 216904 13582 216910 13634
rect 216962 13582 216968 13634
rect 1698 13246 1704 13298
rect 1756 13246 1762 13298
rect 216904 13246 216910 13298
rect 216962 13246 216968 13298
rect 1698 12910 1704 12962
rect 1756 12910 1762 12962
rect 216904 12910 216910 12962
rect 216962 12910 216968 12962
rect 1698 12574 1704 12626
rect 1756 12574 1762 12626
rect 216904 12574 216910 12626
rect 216962 12574 216968 12626
rect 1698 12238 1704 12290
rect 1756 12238 1762 12290
rect 216904 12238 216910 12290
rect 216962 12238 216968 12290
rect 1698 11902 1704 11954
rect 1756 11902 1762 11954
rect 216904 11902 216910 11954
rect 216962 11902 216968 11954
rect 1698 11566 1704 11618
rect 1756 11566 1762 11618
rect 216904 11566 216910 11618
rect 216962 11566 216968 11618
rect 1698 11230 1704 11282
rect 1756 11230 1762 11282
rect 216904 11230 216910 11282
rect 216962 11230 216968 11282
rect 1698 10894 1704 10946
rect 1756 10894 1762 10946
rect 216904 10894 216910 10946
rect 216962 10894 216968 10946
rect 1698 10558 1704 10610
rect 1756 10558 1762 10610
rect 216904 10558 216910 10610
rect 216962 10558 216968 10610
rect 1698 10222 1704 10274
rect 1756 10222 1762 10274
rect 216904 10222 216910 10274
rect 216962 10222 216968 10274
rect 1698 9886 1704 9938
rect 1756 9886 1762 9938
rect 216904 9886 216910 9938
rect 216962 9886 216968 9938
rect 1698 9550 1704 9602
rect 1756 9550 1762 9602
rect 216904 9550 216910 9602
rect 216962 9550 216968 9602
rect 1698 9214 1704 9266
rect 1756 9214 1762 9266
rect 216904 9214 216910 9266
rect 216962 9214 216968 9266
rect 1698 8878 1704 8930
rect 1756 8878 1762 8930
rect 216904 8878 216910 8930
rect 216962 8878 216968 8930
rect 1698 8542 1704 8594
rect 1756 8542 1762 8594
rect 216904 8542 216910 8594
rect 216962 8542 216968 8594
rect 1698 8206 1704 8258
rect 1756 8206 1762 8258
rect 216904 8206 216910 8258
rect 216962 8206 216968 8258
rect 1698 7870 1704 7922
rect 1756 7870 1762 7922
rect 216904 7870 216910 7922
rect 216962 7870 216968 7922
rect 1698 7534 1704 7586
rect 1756 7534 1762 7586
rect 216904 7534 216910 7586
rect 216962 7534 216968 7586
rect 1698 7198 1704 7250
rect 1756 7198 1762 7250
rect 216904 7198 216910 7250
rect 216962 7198 216968 7250
rect 1698 6862 1704 6914
rect 1756 6862 1762 6914
rect 216904 6862 216910 6914
rect 216962 6862 216968 6914
rect 1698 6526 1704 6578
rect 1756 6526 1762 6578
rect 216904 6526 216910 6578
rect 216962 6526 216968 6578
rect 1698 6190 1704 6242
rect 1756 6190 1762 6242
rect 216904 6190 216910 6242
rect 216962 6190 216968 6242
rect 1698 5854 1704 5906
rect 1756 5854 1762 5906
rect 216904 5854 216910 5906
rect 216962 5854 216968 5906
rect 1698 5518 1704 5570
rect 1756 5518 1762 5570
rect 216904 5518 216910 5570
rect 216962 5518 216968 5570
rect 1698 5182 1704 5234
rect 1756 5182 1762 5234
rect 216904 5182 216910 5234
rect 216962 5182 216968 5234
rect 1698 4846 1704 4898
rect 1756 4846 1762 4898
rect 216904 4846 216910 4898
rect 216962 4846 216968 4898
rect 1698 4510 1704 4562
rect 1756 4510 1762 4562
rect 216904 4510 216910 4562
rect 216962 4510 216968 4562
rect 1698 4174 1704 4226
rect 1756 4174 1762 4226
rect 216904 4174 216910 4226
rect 216962 4174 216968 4226
rect 1698 3838 1704 3890
rect 1756 3838 1762 3890
rect 216904 3838 216910 3890
rect 216962 3838 216968 3890
rect 1698 3502 1704 3554
rect 1756 3502 1762 3554
rect 216904 3502 216910 3554
rect 216962 3502 216968 3554
rect 1698 3166 1704 3218
rect 1756 3166 1762 3218
rect 216904 3166 216910 3218
rect 216962 3166 216968 3218
rect 1698 2830 1704 2882
rect 1756 2830 1762 2882
rect 216904 2830 216910 2882
rect 216962 2830 216968 2882
rect 1698 2494 1704 2546
rect 1756 2494 1762 2546
rect 216904 2494 216910 2546
rect 216962 2494 216968 2546
rect 1698 2158 1704 2210
rect 1756 2158 1762 2210
rect 216904 2158 216910 2210
rect 216962 2158 216968 2210
rect 1618 1874 217048 1960
rect 1618 1822 2040 1874
rect 2092 1865 3720 1874
rect 3772 1865 5400 1874
rect 5452 1865 7080 1874
rect 7132 1865 8760 1874
rect 8812 1865 10440 1874
rect 10492 1865 12120 1874
rect 12172 1865 13800 1874
rect 13852 1865 15480 1874
rect 15532 1865 17160 1874
rect 17212 1865 18840 1874
rect 18892 1865 20520 1874
rect 20572 1865 22200 1874
rect 22252 1865 23880 1874
rect 23932 1865 25560 1874
rect 25612 1865 27240 1874
rect 27292 1865 28920 1874
rect 28972 1865 30600 1874
rect 30652 1865 32280 1874
rect 32332 1865 33960 1874
rect 34012 1865 35640 1874
rect 35692 1865 37320 1874
rect 37372 1865 39000 1874
rect 39052 1865 40680 1874
rect 40732 1865 42360 1874
rect 42412 1865 44040 1874
rect 44092 1865 45720 1874
rect 45772 1865 47400 1874
rect 47452 1865 49080 1874
rect 49132 1865 50760 1874
rect 50812 1865 52440 1874
rect 52492 1865 54120 1874
rect 54172 1865 55800 1874
rect 55852 1865 57480 1874
rect 57532 1865 59160 1874
rect 59212 1865 60840 1874
rect 60892 1865 62520 1874
rect 62572 1865 64200 1874
rect 64252 1865 65880 1874
rect 65932 1865 67560 1874
rect 67612 1865 69240 1874
rect 69292 1865 70920 1874
rect 70972 1865 72600 1874
rect 72652 1865 74280 1874
rect 74332 1865 75960 1874
rect 76012 1865 77640 1874
rect 77692 1865 79320 1874
rect 79372 1865 81000 1874
rect 81052 1865 82680 1874
rect 82732 1865 84360 1874
rect 84412 1865 86040 1874
rect 86092 1865 87720 1874
rect 87772 1865 89400 1874
rect 89452 1865 91080 1874
rect 91132 1865 92760 1874
rect 92812 1865 94440 1874
rect 94492 1865 96120 1874
rect 96172 1865 97800 1874
rect 97852 1865 99480 1874
rect 99532 1865 101160 1874
rect 101212 1865 102840 1874
rect 102892 1865 104520 1874
rect 104572 1865 106200 1874
rect 106252 1865 107880 1874
rect 107932 1865 109560 1874
rect 109612 1865 111240 1874
rect 111292 1865 112920 1874
rect 112972 1865 114600 1874
rect 114652 1865 116280 1874
rect 116332 1865 117960 1874
rect 118012 1865 119640 1874
rect 119692 1865 121320 1874
rect 121372 1865 123000 1874
rect 123052 1865 124680 1874
rect 124732 1865 126360 1874
rect 126412 1865 128040 1874
rect 128092 1865 129720 1874
rect 129772 1865 131400 1874
rect 131452 1865 133080 1874
rect 133132 1865 134760 1874
rect 134812 1865 136440 1874
rect 136492 1865 138120 1874
rect 138172 1865 139800 1874
rect 139852 1865 141480 1874
rect 141532 1865 143160 1874
rect 143212 1865 144840 1874
rect 144892 1865 146520 1874
rect 146572 1865 148200 1874
rect 148252 1865 149880 1874
rect 149932 1865 151560 1874
rect 151612 1865 153240 1874
rect 153292 1865 154920 1874
rect 154972 1865 156600 1874
rect 156652 1865 158280 1874
rect 158332 1865 159960 1874
rect 160012 1865 161640 1874
rect 161692 1865 163320 1874
rect 163372 1865 165000 1874
rect 165052 1865 166680 1874
rect 166732 1865 168360 1874
rect 168412 1865 170040 1874
rect 170092 1865 171720 1874
rect 171772 1865 173400 1874
rect 173452 1865 175080 1874
rect 175132 1865 176760 1874
rect 176812 1865 178440 1874
rect 178492 1865 180120 1874
rect 180172 1865 181800 1874
rect 181852 1865 183480 1874
rect 183532 1865 185160 1874
rect 185212 1865 186840 1874
rect 186892 1865 188520 1874
rect 188572 1865 190200 1874
rect 190252 1865 191880 1874
rect 191932 1865 193560 1874
rect 193612 1865 195240 1874
rect 195292 1865 196920 1874
rect 196972 1865 198600 1874
rect 198652 1865 200280 1874
rect 200332 1865 201960 1874
rect 202012 1865 203640 1874
rect 203692 1865 205320 1874
rect 205372 1865 207000 1874
rect 207052 1865 208680 1874
rect 208732 1865 210360 1874
rect 210412 1865 212040 1874
rect 212092 1865 213720 1874
rect 213772 1865 215400 1874
rect 215452 1865 217048 1874
rect 2092 1831 2385 1865
rect 2419 1831 2721 1865
rect 2755 1831 3057 1865
rect 3091 1831 3393 1865
rect 3427 1831 3720 1865
rect 3772 1831 4065 1865
rect 4099 1831 4401 1865
rect 4435 1831 4737 1865
rect 4771 1831 5073 1865
rect 5107 1831 5400 1865
rect 5452 1831 5745 1865
rect 5779 1831 6081 1865
rect 6115 1831 6417 1865
rect 6451 1831 6753 1865
rect 6787 1831 7080 1865
rect 7132 1831 7425 1865
rect 7459 1831 7761 1865
rect 7795 1831 8097 1865
rect 8131 1831 8433 1865
rect 8467 1831 8760 1865
rect 8812 1831 9105 1865
rect 9139 1831 9441 1865
rect 9475 1831 9777 1865
rect 9811 1831 10113 1865
rect 10147 1831 10440 1865
rect 10492 1831 10785 1865
rect 10819 1831 11121 1865
rect 11155 1831 11457 1865
rect 11491 1831 11793 1865
rect 11827 1831 12120 1865
rect 12172 1831 12465 1865
rect 12499 1831 12801 1865
rect 12835 1831 13137 1865
rect 13171 1831 13473 1865
rect 13507 1831 13800 1865
rect 13852 1831 14145 1865
rect 14179 1831 14481 1865
rect 14515 1831 14817 1865
rect 14851 1831 15153 1865
rect 15187 1831 15480 1865
rect 15532 1831 15825 1865
rect 15859 1831 16161 1865
rect 16195 1831 16497 1865
rect 16531 1831 16833 1865
rect 16867 1831 17160 1865
rect 17212 1831 17505 1865
rect 17539 1831 17841 1865
rect 17875 1831 18177 1865
rect 18211 1831 18513 1865
rect 18547 1831 18840 1865
rect 18892 1831 19185 1865
rect 19219 1831 19521 1865
rect 19555 1831 19857 1865
rect 19891 1831 20193 1865
rect 20227 1831 20520 1865
rect 20572 1831 20865 1865
rect 20899 1831 21201 1865
rect 21235 1831 21537 1865
rect 21571 1831 21873 1865
rect 21907 1831 22200 1865
rect 22252 1831 22545 1865
rect 22579 1831 22881 1865
rect 22915 1831 23217 1865
rect 23251 1831 23553 1865
rect 23587 1831 23880 1865
rect 23932 1831 24225 1865
rect 24259 1831 24561 1865
rect 24595 1831 24897 1865
rect 24931 1831 25233 1865
rect 25267 1831 25560 1865
rect 25612 1831 25905 1865
rect 25939 1831 26241 1865
rect 26275 1831 26577 1865
rect 26611 1831 26913 1865
rect 26947 1831 27240 1865
rect 27292 1831 27585 1865
rect 27619 1831 27921 1865
rect 27955 1831 28257 1865
rect 28291 1831 28593 1865
rect 28627 1831 28920 1865
rect 28972 1831 29265 1865
rect 29299 1831 29601 1865
rect 29635 1831 29937 1865
rect 29971 1831 30273 1865
rect 30307 1831 30600 1865
rect 30652 1831 30945 1865
rect 30979 1831 31281 1865
rect 31315 1831 31617 1865
rect 31651 1831 31953 1865
rect 31987 1831 32280 1865
rect 32332 1831 32625 1865
rect 32659 1831 32961 1865
rect 32995 1831 33297 1865
rect 33331 1831 33633 1865
rect 33667 1831 33960 1865
rect 34012 1831 34305 1865
rect 34339 1831 34641 1865
rect 34675 1831 34977 1865
rect 35011 1831 35313 1865
rect 35347 1831 35640 1865
rect 35692 1831 35985 1865
rect 36019 1831 36321 1865
rect 36355 1831 36657 1865
rect 36691 1831 36993 1865
rect 37027 1831 37320 1865
rect 37372 1831 37665 1865
rect 37699 1831 38001 1865
rect 38035 1831 38337 1865
rect 38371 1831 38673 1865
rect 38707 1831 39000 1865
rect 39052 1831 39345 1865
rect 39379 1831 39681 1865
rect 39715 1831 40017 1865
rect 40051 1831 40353 1865
rect 40387 1831 40680 1865
rect 40732 1831 41025 1865
rect 41059 1831 41361 1865
rect 41395 1831 41697 1865
rect 41731 1831 42033 1865
rect 42067 1831 42360 1865
rect 42412 1831 42705 1865
rect 42739 1831 43041 1865
rect 43075 1831 43377 1865
rect 43411 1831 43713 1865
rect 43747 1831 44040 1865
rect 44092 1831 44385 1865
rect 44419 1831 44721 1865
rect 44755 1831 45057 1865
rect 45091 1831 45393 1865
rect 45427 1831 45720 1865
rect 45772 1831 46065 1865
rect 46099 1831 46401 1865
rect 46435 1831 46737 1865
rect 46771 1831 47073 1865
rect 47107 1831 47400 1865
rect 47452 1831 47745 1865
rect 47779 1831 48081 1865
rect 48115 1831 48417 1865
rect 48451 1831 48753 1865
rect 48787 1831 49080 1865
rect 49132 1831 49425 1865
rect 49459 1831 49761 1865
rect 49795 1831 50097 1865
rect 50131 1831 50433 1865
rect 50467 1831 50760 1865
rect 50812 1831 51105 1865
rect 51139 1831 51441 1865
rect 51475 1831 51777 1865
rect 51811 1831 52113 1865
rect 52147 1831 52440 1865
rect 52492 1831 52785 1865
rect 52819 1831 53121 1865
rect 53155 1831 53457 1865
rect 53491 1831 53793 1865
rect 53827 1831 54120 1865
rect 54172 1831 54465 1865
rect 54499 1831 54801 1865
rect 54835 1831 55137 1865
rect 55171 1831 55473 1865
rect 55507 1831 55800 1865
rect 55852 1831 56145 1865
rect 56179 1831 56481 1865
rect 56515 1831 56817 1865
rect 56851 1831 57153 1865
rect 57187 1831 57480 1865
rect 57532 1831 57825 1865
rect 57859 1831 58161 1865
rect 58195 1831 58497 1865
rect 58531 1831 58833 1865
rect 58867 1831 59160 1865
rect 59212 1831 59505 1865
rect 59539 1831 59841 1865
rect 59875 1831 60177 1865
rect 60211 1831 60513 1865
rect 60547 1831 60840 1865
rect 60892 1831 61185 1865
rect 61219 1831 61521 1865
rect 61555 1831 61857 1865
rect 61891 1831 62193 1865
rect 62227 1831 62520 1865
rect 62572 1831 62865 1865
rect 62899 1831 63201 1865
rect 63235 1831 63537 1865
rect 63571 1831 63873 1865
rect 63907 1831 64200 1865
rect 64252 1831 64545 1865
rect 64579 1831 64881 1865
rect 64915 1831 65217 1865
rect 65251 1831 65553 1865
rect 65587 1831 65880 1865
rect 65932 1831 66225 1865
rect 66259 1831 66561 1865
rect 66595 1831 66897 1865
rect 66931 1831 67233 1865
rect 67267 1831 67560 1865
rect 67612 1831 67905 1865
rect 67939 1831 68241 1865
rect 68275 1831 68577 1865
rect 68611 1831 68913 1865
rect 68947 1831 69240 1865
rect 69292 1831 69585 1865
rect 69619 1831 69921 1865
rect 69955 1831 70257 1865
rect 70291 1831 70593 1865
rect 70627 1831 70920 1865
rect 70972 1831 71265 1865
rect 71299 1831 71601 1865
rect 71635 1831 71937 1865
rect 71971 1831 72273 1865
rect 72307 1831 72600 1865
rect 72652 1831 72945 1865
rect 72979 1831 73281 1865
rect 73315 1831 73617 1865
rect 73651 1831 73953 1865
rect 73987 1831 74280 1865
rect 74332 1831 74625 1865
rect 74659 1831 74961 1865
rect 74995 1831 75297 1865
rect 75331 1831 75633 1865
rect 75667 1831 75960 1865
rect 76012 1831 76305 1865
rect 76339 1831 76641 1865
rect 76675 1831 76977 1865
rect 77011 1831 77313 1865
rect 77347 1831 77640 1865
rect 77692 1831 77985 1865
rect 78019 1831 78321 1865
rect 78355 1831 78657 1865
rect 78691 1831 78993 1865
rect 79027 1831 79320 1865
rect 79372 1831 79665 1865
rect 79699 1831 80001 1865
rect 80035 1831 80337 1865
rect 80371 1831 80673 1865
rect 80707 1831 81000 1865
rect 81052 1831 81345 1865
rect 81379 1831 81681 1865
rect 81715 1831 82017 1865
rect 82051 1831 82353 1865
rect 82387 1831 82680 1865
rect 82732 1831 83025 1865
rect 83059 1831 83361 1865
rect 83395 1831 83697 1865
rect 83731 1831 84033 1865
rect 84067 1831 84360 1865
rect 84412 1831 84705 1865
rect 84739 1831 85041 1865
rect 85075 1831 85377 1865
rect 85411 1831 85713 1865
rect 85747 1831 86040 1865
rect 86092 1831 86385 1865
rect 86419 1831 86721 1865
rect 86755 1831 87057 1865
rect 87091 1831 87393 1865
rect 87427 1831 87720 1865
rect 87772 1831 88065 1865
rect 88099 1831 88401 1865
rect 88435 1831 88737 1865
rect 88771 1831 89073 1865
rect 89107 1831 89400 1865
rect 89452 1831 89745 1865
rect 89779 1831 90081 1865
rect 90115 1831 90417 1865
rect 90451 1831 90753 1865
rect 90787 1831 91080 1865
rect 91132 1831 91425 1865
rect 91459 1831 91761 1865
rect 91795 1831 92097 1865
rect 92131 1831 92433 1865
rect 92467 1831 92760 1865
rect 92812 1831 93105 1865
rect 93139 1831 93441 1865
rect 93475 1831 93777 1865
rect 93811 1831 94113 1865
rect 94147 1831 94440 1865
rect 94492 1831 94785 1865
rect 94819 1831 95121 1865
rect 95155 1831 95457 1865
rect 95491 1831 95793 1865
rect 95827 1831 96120 1865
rect 96172 1831 96465 1865
rect 96499 1831 96801 1865
rect 96835 1831 97137 1865
rect 97171 1831 97473 1865
rect 97507 1831 97800 1865
rect 97852 1831 98145 1865
rect 98179 1831 98481 1865
rect 98515 1831 98817 1865
rect 98851 1831 99153 1865
rect 99187 1831 99480 1865
rect 99532 1831 99825 1865
rect 99859 1831 100161 1865
rect 100195 1831 100497 1865
rect 100531 1831 100833 1865
rect 100867 1831 101160 1865
rect 101212 1831 101505 1865
rect 101539 1831 101841 1865
rect 101875 1831 102177 1865
rect 102211 1831 102513 1865
rect 102547 1831 102840 1865
rect 102892 1831 103185 1865
rect 103219 1831 103521 1865
rect 103555 1831 103857 1865
rect 103891 1831 104193 1865
rect 104227 1831 104520 1865
rect 104572 1831 104865 1865
rect 104899 1831 105201 1865
rect 105235 1831 105537 1865
rect 105571 1831 105873 1865
rect 105907 1831 106200 1865
rect 106252 1831 106545 1865
rect 106579 1831 106881 1865
rect 106915 1831 107217 1865
rect 107251 1831 107553 1865
rect 107587 1831 107880 1865
rect 107932 1831 108225 1865
rect 108259 1831 108561 1865
rect 108595 1831 108897 1865
rect 108931 1831 109233 1865
rect 109267 1831 109560 1865
rect 109612 1831 109905 1865
rect 109939 1831 110241 1865
rect 110275 1831 110577 1865
rect 110611 1831 110913 1865
rect 110947 1831 111240 1865
rect 111292 1831 111585 1865
rect 111619 1831 111921 1865
rect 111955 1831 112257 1865
rect 112291 1831 112593 1865
rect 112627 1831 112920 1865
rect 112972 1831 113265 1865
rect 113299 1831 113601 1865
rect 113635 1831 113937 1865
rect 113971 1831 114273 1865
rect 114307 1831 114600 1865
rect 114652 1831 114945 1865
rect 114979 1831 115281 1865
rect 115315 1831 115617 1865
rect 115651 1831 115953 1865
rect 115987 1831 116280 1865
rect 116332 1831 116625 1865
rect 116659 1831 116961 1865
rect 116995 1831 117297 1865
rect 117331 1831 117633 1865
rect 117667 1831 117960 1865
rect 118012 1831 118305 1865
rect 118339 1831 118641 1865
rect 118675 1831 118977 1865
rect 119011 1831 119313 1865
rect 119347 1831 119640 1865
rect 119692 1831 119985 1865
rect 120019 1831 120321 1865
rect 120355 1831 120657 1865
rect 120691 1831 120993 1865
rect 121027 1831 121320 1865
rect 121372 1831 121665 1865
rect 121699 1831 122001 1865
rect 122035 1831 122337 1865
rect 122371 1831 122673 1865
rect 122707 1831 123000 1865
rect 123052 1831 123345 1865
rect 123379 1831 123681 1865
rect 123715 1831 124017 1865
rect 124051 1831 124353 1865
rect 124387 1831 124680 1865
rect 124732 1831 125025 1865
rect 125059 1831 125361 1865
rect 125395 1831 125697 1865
rect 125731 1831 126033 1865
rect 126067 1831 126360 1865
rect 126412 1831 126705 1865
rect 126739 1831 127041 1865
rect 127075 1831 127377 1865
rect 127411 1831 127713 1865
rect 127747 1831 128040 1865
rect 128092 1831 128385 1865
rect 128419 1831 128721 1865
rect 128755 1831 129057 1865
rect 129091 1831 129393 1865
rect 129427 1831 129720 1865
rect 129772 1831 130065 1865
rect 130099 1831 130401 1865
rect 130435 1831 130737 1865
rect 130771 1831 131073 1865
rect 131107 1831 131400 1865
rect 131452 1831 131745 1865
rect 131779 1831 132081 1865
rect 132115 1831 132417 1865
rect 132451 1831 132753 1865
rect 132787 1831 133080 1865
rect 133132 1831 133425 1865
rect 133459 1831 133761 1865
rect 133795 1831 134097 1865
rect 134131 1831 134433 1865
rect 134467 1831 134760 1865
rect 134812 1831 135105 1865
rect 135139 1831 135441 1865
rect 135475 1831 135777 1865
rect 135811 1831 136113 1865
rect 136147 1831 136440 1865
rect 136492 1831 136785 1865
rect 136819 1831 137121 1865
rect 137155 1831 137457 1865
rect 137491 1831 137793 1865
rect 137827 1831 138120 1865
rect 138172 1831 138465 1865
rect 138499 1831 138801 1865
rect 138835 1831 139137 1865
rect 139171 1831 139473 1865
rect 139507 1831 139800 1865
rect 139852 1831 140145 1865
rect 140179 1831 140481 1865
rect 140515 1831 140817 1865
rect 140851 1831 141153 1865
rect 141187 1831 141480 1865
rect 141532 1831 141825 1865
rect 141859 1831 142161 1865
rect 142195 1831 142497 1865
rect 142531 1831 142833 1865
rect 142867 1831 143160 1865
rect 143212 1831 143505 1865
rect 143539 1831 143841 1865
rect 143875 1831 144177 1865
rect 144211 1831 144513 1865
rect 144547 1831 144840 1865
rect 144892 1831 145185 1865
rect 145219 1831 145521 1865
rect 145555 1831 145857 1865
rect 145891 1831 146193 1865
rect 146227 1831 146520 1865
rect 146572 1831 146865 1865
rect 146899 1831 147201 1865
rect 147235 1831 147537 1865
rect 147571 1831 147873 1865
rect 147907 1831 148200 1865
rect 148252 1831 148545 1865
rect 148579 1831 148881 1865
rect 148915 1831 149217 1865
rect 149251 1831 149553 1865
rect 149587 1831 149880 1865
rect 149932 1831 150225 1865
rect 150259 1831 150561 1865
rect 150595 1831 150897 1865
rect 150931 1831 151233 1865
rect 151267 1831 151560 1865
rect 151612 1831 151905 1865
rect 151939 1831 152241 1865
rect 152275 1831 152577 1865
rect 152611 1831 152913 1865
rect 152947 1831 153240 1865
rect 153292 1831 153585 1865
rect 153619 1831 153921 1865
rect 153955 1831 154257 1865
rect 154291 1831 154593 1865
rect 154627 1831 154920 1865
rect 154972 1831 155265 1865
rect 155299 1831 155601 1865
rect 155635 1831 155937 1865
rect 155971 1831 156273 1865
rect 156307 1831 156600 1865
rect 156652 1831 156945 1865
rect 156979 1831 157281 1865
rect 157315 1831 157617 1865
rect 157651 1831 157953 1865
rect 157987 1831 158280 1865
rect 158332 1831 158625 1865
rect 158659 1831 158961 1865
rect 158995 1831 159297 1865
rect 159331 1831 159633 1865
rect 159667 1831 159960 1865
rect 160012 1831 160305 1865
rect 160339 1831 160641 1865
rect 160675 1831 160977 1865
rect 161011 1831 161313 1865
rect 161347 1831 161640 1865
rect 161692 1831 161985 1865
rect 162019 1831 162321 1865
rect 162355 1831 162657 1865
rect 162691 1831 162993 1865
rect 163027 1831 163320 1865
rect 163372 1831 163665 1865
rect 163699 1831 164001 1865
rect 164035 1831 164337 1865
rect 164371 1831 164673 1865
rect 164707 1831 165000 1865
rect 165052 1831 165345 1865
rect 165379 1831 165681 1865
rect 165715 1831 166017 1865
rect 166051 1831 166353 1865
rect 166387 1831 166680 1865
rect 166732 1831 167025 1865
rect 167059 1831 167361 1865
rect 167395 1831 167697 1865
rect 167731 1831 168033 1865
rect 168067 1831 168360 1865
rect 168412 1831 168705 1865
rect 168739 1831 169041 1865
rect 169075 1831 169377 1865
rect 169411 1831 169713 1865
rect 169747 1831 170040 1865
rect 170092 1831 170385 1865
rect 170419 1831 170721 1865
rect 170755 1831 171057 1865
rect 171091 1831 171393 1865
rect 171427 1831 171720 1865
rect 171772 1831 172065 1865
rect 172099 1831 172401 1865
rect 172435 1831 172737 1865
rect 172771 1831 173073 1865
rect 173107 1831 173400 1865
rect 173452 1831 173745 1865
rect 173779 1831 174081 1865
rect 174115 1831 174417 1865
rect 174451 1831 174753 1865
rect 174787 1831 175080 1865
rect 175132 1831 175425 1865
rect 175459 1831 175761 1865
rect 175795 1831 176097 1865
rect 176131 1831 176433 1865
rect 176467 1831 176760 1865
rect 176812 1831 177105 1865
rect 177139 1831 177441 1865
rect 177475 1831 177777 1865
rect 177811 1831 178113 1865
rect 178147 1831 178440 1865
rect 178492 1831 178785 1865
rect 178819 1831 179121 1865
rect 179155 1831 179457 1865
rect 179491 1831 179793 1865
rect 179827 1831 180120 1865
rect 180172 1831 180465 1865
rect 180499 1831 180801 1865
rect 180835 1831 181137 1865
rect 181171 1831 181473 1865
rect 181507 1831 181800 1865
rect 181852 1831 182145 1865
rect 182179 1831 182481 1865
rect 182515 1831 182817 1865
rect 182851 1831 183153 1865
rect 183187 1831 183480 1865
rect 183532 1831 183825 1865
rect 183859 1831 184161 1865
rect 184195 1831 184497 1865
rect 184531 1831 184833 1865
rect 184867 1831 185160 1865
rect 185212 1831 185505 1865
rect 185539 1831 185841 1865
rect 185875 1831 186177 1865
rect 186211 1831 186513 1865
rect 186547 1831 186840 1865
rect 186892 1831 187185 1865
rect 187219 1831 187521 1865
rect 187555 1831 187857 1865
rect 187891 1831 188193 1865
rect 188227 1831 188520 1865
rect 188572 1831 188865 1865
rect 188899 1831 189201 1865
rect 189235 1831 189537 1865
rect 189571 1831 189873 1865
rect 189907 1831 190200 1865
rect 190252 1831 190545 1865
rect 190579 1831 190881 1865
rect 190915 1831 191217 1865
rect 191251 1831 191553 1865
rect 191587 1831 191880 1865
rect 191932 1831 192225 1865
rect 192259 1831 192561 1865
rect 192595 1831 192897 1865
rect 192931 1831 193233 1865
rect 193267 1831 193560 1865
rect 193612 1831 193905 1865
rect 193939 1831 194241 1865
rect 194275 1831 194577 1865
rect 194611 1831 194913 1865
rect 194947 1831 195240 1865
rect 195292 1831 195585 1865
rect 195619 1831 195921 1865
rect 195955 1831 196257 1865
rect 196291 1831 196593 1865
rect 196627 1831 196920 1865
rect 196972 1831 197265 1865
rect 197299 1831 197601 1865
rect 197635 1831 197937 1865
rect 197971 1831 198273 1865
rect 198307 1831 198600 1865
rect 198652 1831 198945 1865
rect 198979 1831 199281 1865
rect 199315 1831 199617 1865
rect 199651 1831 199953 1865
rect 199987 1831 200280 1865
rect 200332 1831 200625 1865
rect 200659 1831 200961 1865
rect 200995 1831 201297 1865
rect 201331 1831 201633 1865
rect 201667 1831 201960 1865
rect 202012 1831 202305 1865
rect 202339 1831 202641 1865
rect 202675 1831 202977 1865
rect 203011 1831 203313 1865
rect 203347 1831 203640 1865
rect 203692 1831 203985 1865
rect 204019 1831 204321 1865
rect 204355 1831 204657 1865
rect 204691 1831 204993 1865
rect 205027 1831 205320 1865
rect 205372 1831 205665 1865
rect 205699 1831 206001 1865
rect 206035 1831 206337 1865
rect 206371 1831 206673 1865
rect 206707 1831 207000 1865
rect 207052 1831 207345 1865
rect 207379 1831 207681 1865
rect 207715 1831 208017 1865
rect 208051 1831 208353 1865
rect 208387 1831 208680 1865
rect 208732 1831 209025 1865
rect 209059 1831 209361 1865
rect 209395 1831 209697 1865
rect 209731 1831 210033 1865
rect 210067 1831 210360 1865
rect 210412 1831 210705 1865
rect 210739 1831 211041 1865
rect 211075 1831 211377 1865
rect 211411 1831 211713 1865
rect 211747 1831 212040 1865
rect 212092 1831 212385 1865
rect 212419 1831 212721 1865
rect 212755 1831 213057 1865
rect 213091 1831 213393 1865
rect 213427 1831 213720 1865
rect 213772 1831 214065 1865
rect 214099 1831 214401 1865
rect 214435 1831 214737 1865
rect 214771 1831 215073 1865
rect 215107 1831 215400 1865
rect 215452 1831 215745 1865
rect 215779 1831 216081 1865
rect 216115 1831 216417 1865
rect 216451 1831 217048 1865
rect 2092 1822 3720 1831
rect 3772 1822 5400 1831
rect 5452 1822 7080 1831
rect 7132 1822 8760 1831
rect 8812 1822 10440 1831
rect 10492 1822 12120 1831
rect 12172 1822 13800 1831
rect 13852 1822 15480 1831
rect 15532 1822 17160 1831
rect 17212 1822 18840 1831
rect 18892 1822 20520 1831
rect 20572 1822 22200 1831
rect 22252 1822 23880 1831
rect 23932 1822 25560 1831
rect 25612 1822 27240 1831
rect 27292 1822 28920 1831
rect 28972 1822 30600 1831
rect 30652 1822 32280 1831
rect 32332 1822 33960 1831
rect 34012 1822 35640 1831
rect 35692 1822 37320 1831
rect 37372 1822 39000 1831
rect 39052 1822 40680 1831
rect 40732 1822 42360 1831
rect 42412 1822 44040 1831
rect 44092 1822 45720 1831
rect 45772 1822 47400 1831
rect 47452 1822 49080 1831
rect 49132 1822 50760 1831
rect 50812 1822 52440 1831
rect 52492 1822 54120 1831
rect 54172 1822 55800 1831
rect 55852 1822 57480 1831
rect 57532 1822 59160 1831
rect 59212 1822 60840 1831
rect 60892 1822 62520 1831
rect 62572 1822 64200 1831
rect 64252 1822 65880 1831
rect 65932 1822 67560 1831
rect 67612 1822 69240 1831
rect 69292 1822 70920 1831
rect 70972 1822 72600 1831
rect 72652 1822 74280 1831
rect 74332 1822 75960 1831
rect 76012 1822 77640 1831
rect 77692 1822 79320 1831
rect 79372 1822 81000 1831
rect 81052 1822 82680 1831
rect 82732 1822 84360 1831
rect 84412 1822 86040 1831
rect 86092 1822 87720 1831
rect 87772 1822 89400 1831
rect 89452 1822 91080 1831
rect 91132 1822 92760 1831
rect 92812 1822 94440 1831
rect 94492 1822 96120 1831
rect 96172 1822 97800 1831
rect 97852 1822 99480 1831
rect 99532 1822 101160 1831
rect 101212 1822 102840 1831
rect 102892 1822 104520 1831
rect 104572 1822 106200 1831
rect 106252 1822 107880 1831
rect 107932 1822 109560 1831
rect 109612 1822 111240 1831
rect 111292 1822 112920 1831
rect 112972 1822 114600 1831
rect 114652 1822 116280 1831
rect 116332 1822 117960 1831
rect 118012 1822 119640 1831
rect 119692 1822 121320 1831
rect 121372 1822 123000 1831
rect 123052 1822 124680 1831
rect 124732 1822 126360 1831
rect 126412 1822 128040 1831
rect 128092 1822 129720 1831
rect 129772 1822 131400 1831
rect 131452 1822 133080 1831
rect 133132 1822 134760 1831
rect 134812 1822 136440 1831
rect 136492 1822 138120 1831
rect 138172 1822 139800 1831
rect 139852 1822 141480 1831
rect 141532 1822 143160 1831
rect 143212 1822 144840 1831
rect 144892 1822 146520 1831
rect 146572 1822 148200 1831
rect 148252 1822 149880 1831
rect 149932 1822 151560 1831
rect 151612 1822 153240 1831
rect 153292 1822 154920 1831
rect 154972 1822 156600 1831
rect 156652 1822 158280 1831
rect 158332 1822 159960 1831
rect 160012 1822 161640 1831
rect 161692 1822 163320 1831
rect 163372 1822 165000 1831
rect 165052 1822 166680 1831
rect 166732 1822 168360 1831
rect 168412 1822 170040 1831
rect 170092 1822 171720 1831
rect 171772 1822 173400 1831
rect 173452 1822 175080 1831
rect 175132 1822 176760 1831
rect 176812 1822 178440 1831
rect 178492 1822 180120 1831
rect 180172 1822 181800 1831
rect 181852 1822 183480 1831
rect 183532 1822 185160 1831
rect 185212 1822 186840 1831
rect 186892 1822 188520 1831
rect 188572 1822 190200 1831
rect 190252 1822 191880 1831
rect 191932 1822 193560 1831
rect 193612 1822 195240 1831
rect 195292 1822 196920 1831
rect 196972 1822 198600 1831
rect 198652 1822 200280 1831
rect 200332 1822 201960 1831
rect 202012 1822 203640 1831
rect 203692 1822 205320 1831
rect 205372 1822 207000 1831
rect 207052 1822 208680 1831
rect 208732 1822 210360 1831
rect 210412 1822 212040 1831
rect 212092 1822 213720 1831
rect 213772 1822 215400 1831
rect 215452 1822 217048 1831
rect 1618 1736 217048 1822
<< via1 >>
rect 2040 142361 2092 142370
rect 3720 142361 3772 142370
rect 5400 142361 5452 142370
rect 7080 142361 7132 142370
rect 8760 142361 8812 142370
rect 10440 142361 10492 142370
rect 12120 142361 12172 142370
rect 13800 142361 13852 142370
rect 15480 142361 15532 142370
rect 17160 142361 17212 142370
rect 18840 142361 18892 142370
rect 20520 142361 20572 142370
rect 22200 142361 22252 142370
rect 23880 142361 23932 142370
rect 25560 142361 25612 142370
rect 27240 142361 27292 142370
rect 28920 142361 28972 142370
rect 30600 142361 30652 142370
rect 32280 142361 32332 142370
rect 33960 142361 34012 142370
rect 35640 142361 35692 142370
rect 37320 142361 37372 142370
rect 39000 142361 39052 142370
rect 40680 142361 40732 142370
rect 42360 142361 42412 142370
rect 44040 142361 44092 142370
rect 45720 142361 45772 142370
rect 47400 142361 47452 142370
rect 49080 142361 49132 142370
rect 50760 142361 50812 142370
rect 52440 142361 52492 142370
rect 54120 142361 54172 142370
rect 55800 142361 55852 142370
rect 57480 142361 57532 142370
rect 59160 142361 59212 142370
rect 60840 142361 60892 142370
rect 62520 142361 62572 142370
rect 64200 142361 64252 142370
rect 65880 142361 65932 142370
rect 67560 142361 67612 142370
rect 69240 142361 69292 142370
rect 70920 142361 70972 142370
rect 72600 142361 72652 142370
rect 74280 142361 74332 142370
rect 75960 142361 76012 142370
rect 77640 142361 77692 142370
rect 79320 142361 79372 142370
rect 81000 142361 81052 142370
rect 82680 142361 82732 142370
rect 84360 142361 84412 142370
rect 86040 142361 86092 142370
rect 87720 142361 87772 142370
rect 89400 142361 89452 142370
rect 91080 142361 91132 142370
rect 92760 142361 92812 142370
rect 94440 142361 94492 142370
rect 96120 142361 96172 142370
rect 97800 142361 97852 142370
rect 99480 142361 99532 142370
rect 101160 142361 101212 142370
rect 102840 142361 102892 142370
rect 104520 142361 104572 142370
rect 106200 142361 106252 142370
rect 107880 142361 107932 142370
rect 109560 142361 109612 142370
rect 111240 142361 111292 142370
rect 112920 142361 112972 142370
rect 114600 142361 114652 142370
rect 116280 142361 116332 142370
rect 117960 142361 118012 142370
rect 119640 142361 119692 142370
rect 121320 142361 121372 142370
rect 123000 142361 123052 142370
rect 124680 142361 124732 142370
rect 126360 142361 126412 142370
rect 128040 142361 128092 142370
rect 129720 142361 129772 142370
rect 131400 142361 131452 142370
rect 133080 142361 133132 142370
rect 134760 142361 134812 142370
rect 136440 142361 136492 142370
rect 138120 142361 138172 142370
rect 139800 142361 139852 142370
rect 141480 142361 141532 142370
rect 143160 142361 143212 142370
rect 144840 142361 144892 142370
rect 146520 142361 146572 142370
rect 148200 142361 148252 142370
rect 149880 142361 149932 142370
rect 151560 142361 151612 142370
rect 153240 142361 153292 142370
rect 154920 142361 154972 142370
rect 156600 142361 156652 142370
rect 158280 142361 158332 142370
rect 159960 142361 160012 142370
rect 161640 142361 161692 142370
rect 163320 142361 163372 142370
rect 165000 142361 165052 142370
rect 166680 142361 166732 142370
rect 168360 142361 168412 142370
rect 170040 142361 170092 142370
rect 171720 142361 171772 142370
rect 173400 142361 173452 142370
rect 175080 142361 175132 142370
rect 176760 142361 176812 142370
rect 178440 142361 178492 142370
rect 180120 142361 180172 142370
rect 181800 142361 181852 142370
rect 183480 142361 183532 142370
rect 185160 142361 185212 142370
rect 186840 142361 186892 142370
rect 188520 142361 188572 142370
rect 190200 142361 190252 142370
rect 191880 142361 191932 142370
rect 193560 142361 193612 142370
rect 195240 142361 195292 142370
rect 196920 142361 196972 142370
rect 198600 142361 198652 142370
rect 200280 142361 200332 142370
rect 201960 142361 202012 142370
rect 203640 142361 203692 142370
rect 205320 142361 205372 142370
rect 207000 142361 207052 142370
rect 208680 142361 208732 142370
rect 210360 142361 210412 142370
rect 212040 142361 212092 142370
rect 213720 142361 213772 142370
rect 215400 142361 215452 142370
rect 2040 142327 2049 142361
rect 2049 142327 2083 142361
rect 2083 142327 2092 142361
rect 3720 142327 3729 142361
rect 3729 142327 3763 142361
rect 3763 142327 3772 142361
rect 5400 142327 5409 142361
rect 5409 142327 5443 142361
rect 5443 142327 5452 142361
rect 7080 142327 7089 142361
rect 7089 142327 7123 142361
rect 7123 142327 7132 142361
rect 8760 142327 8769 142361
rect 8769 142327 8803 142361
rect 8803 142327 8812 142361
rect 10440 142327 10449 142361
rect 10449 142327 10483 142361
rect 10483 142327 10492 142361
rect 12120 142327 12129 142361
rect 12129 142327 12163 142361
rect 12163 142327 12172 142361
rect 13800 142327 13809 142361
rect 13809 142327 13843 142361
rect 13843 142327 13852 142361
rect 15480 142327 15489 142361
rect 15489 142327 15523 142361
rect 15523 142327 15532 142361
rect 17160 142327 17169 142361
rect 17169 142327 17203 142361
rect 17203 142327 17212 142361
rect 18840 142327 18849 142361
rect 18849 142327 18883 142361
rect 18883 142327 18892 142361
rect 20520 142327 20529 142361
rect 20529 142327 20563 142361
rect 20563 142327 20572 142361
rect 22200 142327 22209 142361
rect 22209 142327 22243 142361
rect 22243 142327 22252 142361
rect 23880 142327 23889 142361
rect 23889 142327 23923 142361
rect 23923 142327 23932 142361
rect 25560 142327 25569 142361
rect 25569 142327 25603 142361
rect 25603 142327 25612 142361
rect 27240 142327 27249 142361
rect 27249 142327 27283 142361
rect 27283 142327 27292 142361
rect 28920 142327 28929 142361
rect 28929 142327 28963 142361
rect 28963 142327 28972 142361
rect 30600 142327 30609 142361
rect 30609 142327 30643 142361
rect 30643 142327 30652 142361
rect 32280 142327 32289 142361
rect 32289 142327 32323 142361
rect 32323 142327 32332 142361
rect 33960 142327 33969 142361
rect 33969 142327 34003 142361
rect 34003 142327 34012 142361
rect 35640 142327 35649 142361
rect 35649 142327 35683 142361
rect 35683 142327 35692 142361
rect 37320 142327 37329 142361
rect 37329 142327 37363 142361
rect 37363 142327 37372 142361
rect 39000 142327 39009 142361
rect 39009 142327 39043 142361
rect 39043 142327 39052 142361
rect 40680 142327 40689 142361
rect 40689 142327 40723 142361
rect 40723 142327 40732 142361
rect 42360 142327 42369 142361
rect 42369 142327 42403 142361
rect 42403 142327 42412 142361
rect 44040 142327 44049 142361
rect 44049 142327 44083 142361
rect 44083 142327 44092 142361
rect 45720 142327 45729 142361
rect 45729 142327 45763 142361
rect 45763 142327 45772 142361
rect 47400 142327 47409 142361
rect 47409 142327 47443 142361
rect 47443 142327 47452 142361
rect 49080 142327 49089 142361
rect 49089 142327 49123 142361
rect 49123 142327 49132 142361
rect 50760 142327 50769 142361
rect 50769 142327 50803 142361
rect 50803 142327 50812 142361
rect 52440 142327 52449 142361
rect 52449 142327 52483 142361
rect 52483 142327 52492 142361
rect 54120 142327 54129 142361
rect 54129 142327 54163 142361
rect 54163 142327 54172 142361
rect 55800 142327 55809 142361
rect 55809 142327 55843 142361
rect 55843 142327 55852 142361
rect 57480 142327 57489 142361
rect 57489 142327 57523 142361
rect 57523 142327 57532 142361
rect 59160 142327 59169 142361
rect 59169 142327 59203 142361
rect 59203 142327 59212 142361
rect 60840 142327 60849 142361
rect 60849 142327 60883 142361
rect 60883 142327 60892 142361
rect 62520 142327 62529 142361
rect 62529 142327 62563 142361
rect 62563 142327 62572 142361
rect 64200 142327 64209 142361
rect 64209 142327 64243 142361
rect 64243 142327 64252 142361
rect 65880 142327 65889 142361
rect 65889 142327 65923 142361
rect 65923 142327 65932 142361
rect 67560 142327 67569 142361
rect 67569 142327 67603 142361
rect 67603 142327 67612 142361
rect 69240 142327 69249 142361
rect 69249 142327 69283 142361
rect 69283 142327 69292 142361
rect 70920 142327 70929 142361
rect 70929 142327 70963 142361
rect 70963 142327 70972 142361
rect 72600 142327 72609 142361
rect 72609 142327 72643 142361
rect 72643 142327 72652 142361
rect 74280 142327 74289 142361
rect 74289 142327 74323 142361
rect 74323 142327 74332 142361
rect 75960 142327 75969 142361
rect 75969 142327 76003 142361
rect 76003 142327 76012 142361
rect 77640 142327 77649 142361
rect 77649 142327 77683 142361
rect 77683 142327 77692 142361
rect 79320 142327 79329 142361
rect 79329 142327 79363 142361
rect 79363 142327 79372 142361
rect 81000 142327 81009 142361
rect 81009 142327 81043 142361
rect 81043 142327 81052 142361
rect 82680 142327 82689 142361
rect 82689 142327 82723 142361
rect 82723 142327 82732 142361
rect 84360 142327 84369 142361
rect 84369 142327 84403 142361
rect 84403 142327 84412 142361
rect 86040 142327 86049 142361
rect 86049 142327 86083 142361
rect 86083 142327 86092 142361
rect 87720 142327 87729 142361
rect 87729 142327 87763 142361
rect 87763 142327 87772 142361
rect 89400 142327 89409 142361
rect 89409 142327 89443 142361
rect 89443 142327 89452 142361
rect 91080 142327 91089 142361
rect 91089 142327 91123 142361
rect 91123 142327 91132 142361
rect 92760 142327 92769 142361
rect 92769 142327 92803 142361
rect 92803 142327 92812 142361
rect 94440 142327 94449 142361
rect 94449 142327 94483 142361
rect 94483 142327 94492 142361
rect 96120 142327 96129 142361
rect 96129 142327 96163 142361
rect 96163 142327 96172 142361
rect 97800 142327 97809 142361
rect 97809 142327 97843 142361
rect 97843 142327 97852 142361
rect 99480 142327 99489 142361
rect 99489 142327 99523 142361
rect 99523 142327 99532 142361
rect 101160 142327 101169 142361
rect 101169 142327 101203 142361
rect 101203 142327 101212 142361
rect 102840 142327 102849 142361
rect 102849 142327 102883 142361
rect 102883 142327 102892 142361
rect 104520 142327 104529 142361
rect 104529 142327 104563 142361
rect 104563 142327 104572 142361
rect 106200 142327 106209 142361
rect 106209 142327 106243 142361
rect 106243 142327 106252 142361
rect 107880 142327 107889 142361
rect 107889 142327 107923 142361
rect 107923 142327 107932 142361
rect 109560 142327 109569 142361
rect 109569 142327 109603 142361
rect 109603 142327 109612 142361
rect 111240 142327 111249 142361
rect 111249 142327 111283 142361
rect 111283 142327 111292 142361
rect 112920 142327 112929 142361
rect 112929 142327 112963 142361
rect 112963 142327 112972 142361
rect 114600 142327 114609 142361
rect 114609 142327 114643 142361
rect 114643 142327 114652 142361
rect 116280 142327 116289 142361
rect 116289 142327 116323 142361
rect 116323 142327 116332 142361
rect 117960 142327 117969 142361
rect 117969 142327 118003 142361
rect 118003 142327 118012 142361
rect 119640 142327 119649 142361
rect 119649 142327 119683 142361
rect 119683 142327 119692 142361
rect 121320 142327 121329 142361
rect 121329 142327 121363 142361
rect 121363 142327 121372 142361
rect 123000 142327 123009 142361
rect 123009 142327 123043 142361
rect 123043 142327 123052 142361
rect 124680 142327 124689 142361
rect 124689 142327 124723 142361
rect 124723 142327 124732 142361
rect 126360 142327 126369 142361
rect 126369 142327 126403 142361
rect 126403 142327 126412 142361
rect 128040 142327 128049 142361
rect 128049 142327 128083 142361
rect 128083 142327 128092 142361
rect 129720 142327 129729 142361
rect 129729 142327 129763 142361
rect 129763 142327 129772 142361
rect 131400 142327 131409 142361
rect 131409 142327 131443 142361
rect 131443 142327 131452 142361
rect 133080 142327 133089 142361
rect 133089 142327 133123 142361
rect 133123 142327 133132 142361
rect 134760 142327 134769 142361
rect 134769 142327 134803 142361
rect 134803 142327 134812 142361
rect 136440 142327 136449 142361
rect 136449 142327 136483 142361
rect 136483 142327 136492 142361
rect 138120 142327 138129 142361
rect 138129 142327 138163 142361
rect 138163 142327 138172 142361
rect 139800 142327 139809 142361
rect 139809 142327 139843 142361
rect 139843 142327 139852 142361
rect 141480 142327 141489 142361
rect 141489 142327 141523 142361
rect 141523 142327 141532 142361
rect 143160 142327 143169 142361
rect 143169 142327 143203 142361
rect 143203 142327 143212 142361
rect 144840 142327 144849 142361
rect 144849 142327 144883 142361
rect 144883 142327 144892 142361
rect 146520 142327 146529 142361
rect 146529 142327 146563 142361
rect 146563 142327 146572 142361
rect 148200 142327 148209 142361
rect 148209 142327 148243 142361
rect 148243 142327 148252 142361
rect 149880 142327 149889 142361
rect 149889 142327 149923 142361
rect 149923 142327 149932 142361
rect 151560 142327 151569 142361
rect 151569 142327 151603 142361
rect 151603 142327 151612 142361
rect 153240 142327 153249 142361
rect 153249 142327 153283 142361
rect 153283 142327 153292 142361
rect 154920 142327 154929 142361
rect 154929 142327 154963 142361
rect 154963 142327 154972 142361
rect 156600 142327 156609 142361
rect 156609 142327 156643 142361
rect 156643 142327 156652 142361
rect 158280 142327 158289 142361
rect 158289 142327 158323 142361
rect 158323 142327 158332 142361
rect 159960 142327 159969 142361
rect 159969 142327 160003 142361
rect 160003 142327 160012 142361
rect 161640 142327 161649 142361
rect 161649 142327 161683 142361
rect 161683 142327 161692 142361
rect 163320 142327 163329 142361
rect 163329 142327 163363 142361
rect 163363 142327 163372 142361
rect 165000 142327 165009 142361
rect 165009 142327 165043 142361
rect 165043 142327 165052 142361
rect 166680 142327 166689 142361
rect 166689 142327 166723 142361
rect 166723 142327 166732 142361
rect 168360 142327 168369 142361
rect 168369 142327 168403 142361
rect 168403 142327 168412 142361
rect 170040 142327 170049 142361
rect 170049 142327 170083 142361
rect 170083 142327 170092 142361
rect 171720 142327 171729 142361
rect 171729 142327 171763 142361
rect 171763 142327 171772 142361
rect 173400 142327 173409 142361
rect 173409 142327 173443 142361
rect 173443 142327 173452 142361
rect 175080 142327 175089 142361
rect 175089 142327 175123 142361
rect 175123 142327 175132 142361
rect 176760 142327 176769 142361
rect 176769 142327 176803 142361
rect 176803 142327 176812 142361
rect 178440 142327 178449 142361
rect 178449 142327 178483 142361
rect 178483 142327 178492 142361
rect 180120 142327 180129 142361
rect 180129 142327 180163 142361
rect 180163 142327 180172 142361
rect 181800 142327 181809 142361
rect 181809 142327 181843 142361
rect 181843 142327 181852 142361
rect 183480 142327 183489 142361
rect 183489 142327 183523 142361
rect 183523 142327 183532 142361
rect 185160 142327 185169 142361
rect 185169 142327 185203 142361
rect 185203 142327 185212 142361
rect 186840 142327 186849 142361
rect 186849 142327 186883 142361
rect 186883 142327 186892 142361
rect 188520 142327 188529 142361
rect 188529 142327 188563 142361
rect 188563 142327 188572 142361
rect 190200 142327 190209 142361
rect 190209 142327 190243 142361
rect 190243 142327 190252 142361
rect 191880 142327 191889 142361
rect 191889 142327 191923 142361
rect 191923 142327 191932 142361
rect 193560 142327 193569 142361
rect 193569 142327 193603 142361
rect 193603 142327 193612 142361
rect 195240 142327 195249 142361
rect 195249 142327 195283 142361
rect 195283 142327 195292 142361
rect 196920 142327 196929 142361
rect 196929 142327 196963 142361
rect 196963 142327 196972 142361
rect 198600 142327 198609 142361
rect 198609 142327 198643 142361
rect 198643 142327 198652 142361
rect 200280 142327 200289 142361
rect 200289 142327 200323 142361
rect 200323 142327 200332 142361
rect 201960 142327 201969 142361
rect 201969 142327 202003 142361
rect 202003 142327 202012 142361
rect 203640 142327 203649 142361
rect 203649 142327 203683 142361
rect 203683 142327 203692 142361
rect 205320 142327 205329 142361
rect 205329 142327 205363 142361
rect 205363 142327 205372 142361
rect 207000 142327 207009 142361
rect 207009 142327 207043 142361
rect 207043 142327 207052 142361
rect 208680 142327 208689 142361
rect 208689 142327 208723 142361
rect 208723 142327 208732 142361
rect 210360 142327 210369 142361
rect 210369 142327 210403 142361
rect 210403 142327 210412 142361
rect 212040 142327 212049 142361
rect 212049 142327 212083 142361
rect 212083 142327 212092 142361
rect 213720 142327 213729 142361
rect 213729 142327 213763 142361
rect 213763 142327 213772 142361
rect 215400 142327 215409 142361
rect 215409 142327 215443 142361
rect 215443 142327 215452 142361
rect 2040 142318 2092 142327
rect 3720 142318 3772 142327
rect 5400 142318 5452 142327
rect 7080 142318 7132 142327
rect 8760 142318 8812 142327
rect 10440 142318 10492 142327
rect 12120 142318 12172 142327
rect 13800 142318 13852 142327
rect 15480 142318 15532 142327
rect 17160 142318 17212 142327
rect 18840 142318 18892 142327
rect 20520 142318 20572 142327
rect 22200 142318 22252 142327
rect 23880 142318 23932 142327
rect 25560 142318 25612 142327
rect 27240 142318 27292 142327
rect 28920 142318 28972 142327
rect 30600 142318 30652 142327
rect 32280 142318 32332 142327
rect 33960 142318 34012 142327
rect 35640 142318 35692 142327
rect 37320 142318 37372 142327
rect 39000 142318 39052 142327
rect 40680 142318 40732 142327
rect 42360 142318 42412 142327
rect 44040 142318 44092 142327
rect 45720 142318 45772 142327
rect 47400 142318 47452 142327
rect 49080 142318 49132 142327
rect 50760 142318 50812 142327
rect 52440 142318 52492 142327
rect 54120 142318 54172 142327
rect 55800 142318 55852 142327
rect 57480 142318 57532 142327
rect 59160 142318 59212 142327
rect 60840 142318 60892 142327
rect 62520 142318 62572 142327
rect 64200 142318 64252 142327
rect 65880 142318 65932 142327
rect 67560 142318 67612 142327
rect 69240 142318 69292 142327
rect 70920 142318 70972 142327
rect 72600 142318 72652 142327
rect 74280 142318 74332 142327
rect 75960 142318 76012 142327
rect 77640 142318 77692 142327
rect 79320 142318 79372 142327
rect 81000 142318 81052 142327
rect 82680 142318 82732 142327
rect 84360 142318 84412 142327
rect 86040 142318 86092 142327
rect 87720 142318 87772 142327
rect 89400 142318 89452 142327
rect 91080 142318 91132 142327
rect 92760 142318 92812 142327
rect 94440 142318 94492 142327
rect 96120 142318 96172 142327
rect 97800 142318 97852 142327
rect 99480 142318 99532 142327
rect 101160 142318 101212 142327
rect 102840 142318 102892 142327
rect 104520 142318 104572 142327
rect 106200 142318 106252 142327
rect 107880 142318 107932 142327
rect 109560 142318 109612 142327
rect 111240 142318 111292 142327
rect 112920 142318 112972 142327
rect 114600 142318 114652 142327
rect 116280 142318 116332 142327
rect 117960 142318 118012 142327
rect 119640 142318 119692 142327
rect 121320 142318 121372 142327
rect 123000 142318 123052 142327
rect 124680 142318 124732 142327
rect 126360 142318 126412 142327
rect 128040 142318 128092 142327
rect 129720 142318 129772 142327
rect 131400 142318 131452 142327
rect 133080 142318 133132 142327
rect 134760 142318 134812 142327
rect 136440 142318 136492 142327
rect 138120 142318 138172 142327
rect 139800 142318 139852 142327
rect 141480 142318 141532 142327
rect 143160 142318 143212 142327
rect 144840 142318 144892 142327
rect 146520 142318 146572 142327
rect 148200 142318 148252 142327
rect 149880 142318 149932 142327
rect 151560 142318 151612 142327
rect 153240 142318 153292 142327
rect 154920 142318 154972 142327
rect 156600 142318 156652 142327
rect 158280 142318 158332 142327
rect 159960 142318 160012 142327
rect 161640 142318 161692 142327
rect 163320 142318 163372 142327
rect 165000 142318 165052 142327
rect 166680 142318 166732 142327
rect 168360 142318 168412 142327
rect 170040 142318 170092 142327
rect 171720 142318 171772 142327
rect 173400 142318 173452 142327
rect 175080 142318 175132 142327
rect 176760 142318 176812 142327
rect 178440 142318 178492 142327
rect 180120 142318 180172 142327
rect 181800 142318 181852 142327
rect 183480 142318 183532 142327
rect 185160 142318 185212 142327
rect 186840 142318 186892 142327
rect 188520 142318 188572 142327
rect 190200 142318 190252 142327
rect 191880 142318 191932 142327
rect 193560 142318 193612 142327
rect 195240 142318 195292 142327
rect 196920 142318 196972 142327
rect 198600 142318 198652 142327
rect 200280 142318 200332 142327
rect 201960 142318 202012 142327
rect 203640 142318 203692 142327
rect 205320 142318 205372 142327
rect 207000 142318 207052 142327
rect 208680 142318 208732 142327
rect 210360 142318 210412 142327
rect 212040 142318 212092 142327
rect 213720 142318 213772 142327
rect 215400 142318 215452 142327
rect 1704 141977 1756 141986
rect 1704 141943 1713 141977
rect 1713 141943 1747 141977
rect 1747 141943 1756 141977
rect 1704 141934 1756 141943
rect 216910 141977 216962 141986
rect 216910 141943 216919 141977
rect 216919 141943 216953 141977
rect 216953 141943 216962 141977
rect 216910 141934 216962 141943
rect 1704 141641 1756 141650
rect 1704 141607 1713 141641
rect 1713 141607 1747 141641
rect 1747 141607 1756 141641
rect 1704 141598 1756 141607
rect 216910 141641 216962 141650
rect 216910 141607 216919 141641
rect 216919 141607 216953 141641
rect 216953 141607 216962 141641
rect 216910 141598 216962 141607
rect 1704 141305 1756 141314
rect 1704 141271 1713 141305
rect 1713 141271 1747 141305
rect 1747 141271 1756 141305
rect 1704 141262 1756 141271
rect 216910 141305 216962 141314
rect 216910 141271 216919 141305
rect 216919 141271 216953 141305
rect 216953 141271 216962 141305
rect 216910 141262 216962 141271
rect 1704 140969 1756 140978
rect 1704 140935 1713 140969
rect 1713 140935 1747 140969
rect 1747 140935 1756 140969
rect 1704 140926 1756 140935
rect 216910 140969 216962 140978
rect 216910 140935 216919 140969
rect 216919 140935 216953 140969
rect 216953 140935 216962 140969
rect 216910 140926 216962 140935
rect 1704 140633 1756 140642
rect 1704 140599 1713 140633
rect 1713 140599 1747 140633
rect 1747 140599 1756 140633
rect 1704 140590 1756 140599
rect 216910 140633 216962 140642
rect 216910 140599 216919 140633
rect 216919 140599 216953 140633
rect 216953 140599 216962 140633
rect 216910 140590 216962 140599
rect 1704 140297 1756 140306
rect 1704 140263 1713 140297
rect 1713 140263 1747 140297
rect 1747 140263 1756 140297
rect 1704 140254 1756 140263
rect 216910 140297 216962 140306
rect 216910 140263 216919 140297
rect 216919 140263 216953 140297
rect 216953 140263 216962 140297
rect 216910 140254 216962 140263
rect 1704 139961 1756 139970
rect 1704 139927 1713 139961
rect 1713 139927 1747 139961
rect 1747 139927 1756 139961
rect 1704 139918 1756 139927
rect 216910 139961 216962 139970
rect 216910 139927 216919 139961
rect 216919 139927 216953 139961
rect 216953 139927 216962 139961
rect 216910 139918 216962 139927
rect 1704 139625 1756 139634
rect 1704 139591 1713 139625
rect 1713 139591 1747 139625
rect 1747 139591 1756 139625
rect 1704 139582 1756 139591
rect 216910 139625 216962 139634
rect 216910 139591 216919 139625
rect 216919 139591 216953 139625
rect 216953 139591 216962 139625
rect 216910 139582 216962 139591
rect 1704 139289 1756 139298
rect 1704 139255 1713 139289
rect 1713 139255 1747 139289
rect 1747 139255 1756 139289
rect 1704 139246 1756 139255
rect 216910 139289 216962 139298
rect 216910 139255 216919 139289
rect 216919 139255 216953 139289
rect 216953 139255 216962 139289
rect 216910 139246 216962 139255
rect 1704 138953 1756 138962
rect 1704 138919 1713 138953
rect 1713 138919 1747 138953
rect 1747 138919 1756 138953
rect 1704 138910 1756 138919
rect 216910 138953 216962 138962
rect 216910 138919 216919 138953
rect 216919 138919 216953 138953
rect 216953 138919 216962 138953
rect 216910 138910 216962 138919
rect 1704 138617 1756 138626
rect 1704 138583 1713 138617
rect 1713 138583 1747 138617
rect 1747 138583 1756 138617
rect 1704 138574 1756 138583
rect 216910 138617 216962 138626
rect 216910 138583 216919 138617
rect 216919 138583 216953 138617
rect 216953 138583 216962 138617
rect 216910 138574 216962 138583
rect 1704 138281 1756 138290
rect 1704 138247 1713 138281
rect 1713 138247 1747 138281
rect 1747 138247 1756 138281
rect 1704 138238 1756 138247
rect 216910 138281 216962 138290
rect 216910 138247 216919 138281
rect 216919 138247 216953 138281
rect 216953 138247 216962 138281
rect 216910 138238 216962 138247
rect 1704 137945 1756 137954
rect 1704 137911 1713 137945
rect 1713 137911 1747 137945
rect 1747 137911 1756 137945
rect 1704 137902 1756 137911
rect 216910 137945 216962 137954
rect 216910 137911 216919 137945
rect 216919 137911 216953 137945
rect 216953 137911 216962 137945
rect 216910 137902 216962 137911
rect 1704 137609 1756 137618
rect 1704 137575 1713 137609
rect 1713 137575 1747 137609
rect 1747 137575 1756 137609
rect 1704 137566 1756 137575
rect 216910 137609 216962 137618
rect 216910 137575 216919 137609
rect 216919 137575 216953 137609
rect 216953 137575 216962 137609
rect 216910 137566 216962 137575
rect 1704 137273 1756 137282
rect 1704 137239 1713 137273
rect 1713 137239 1747 137273
rect 1747 137239 1756 137273
rect 1704 137230 1756 137239
rect 216910 137273 216962 137282
rect 216910 137239 216919 137273
rect 216919 137239 216953 137273
rect 216953 137239 216962 137273
rect 216910 137230 216962 137239
rect 1704 136937 1756 136946
rect 1704 136903 1713 136937
rect 1713 136903 1747 136937
rect 1747 136903 1756 136937
rect 1704 136894 1756 136903
rect 216910 136937 216962 136946
rect 216910 136903 216919 136937
rect 216919 136903 216953 136937
rect 216953 136903 216962 136937
rect 216910 136894 216962 136903
rect 1704 136601 1756 136610
rect 1704 136567 1713 136601
rect 1713 136567 1747 136601
rect 1747 136567 1756 136601
rect 1704 136558 1756 136567
rect 216910 136601 216962 136610
rect 216910 136567 216919 136601
rect 216919 136567 216953 136601
rect 216953 136567 216962 136601
rect 216910 136558 216962 136567
rect 1704 136265 1756 136274
rect 1704 136231 1713 136265
rect 1713 136231 1747 136265
rect 1747 136231 1756 136265
rect 1704 136222 1756 136231
rect 216910 136265 216962 136274
rect 216910 136231 216919 136265
rect 216919 136231 216953 136265
rect 216953 136231 216962 136265
rect 216910 136222 216962 136231
rect 1704 135929 1756 135938
rect 1704 135895 1713 135929
rect 1713 135895 1747 135929
rect 1747 135895 1756 135929
rect 1704 135886 1756 135895
rect 216910 135929 216962 135938
rect 216910 135895 216919 135929
rect 216919 135895 216953 135929
rect 216953 135895 216962 135929
rect 216910 135886 216962 135895
rect 1704 135593 1756 135602
rect 1704 135559 1713 135593
rect 1713 135559 1747 135593
rect 1747 135559 1756 135593
rect 1704 135550 1756 135559
rect 216910 135593 216962 135602
rect 216910 135559 216919 135593
rect 216919 135559 216953 135593
rect 216953 135559 216962 135593
rect 216910 135550 216962 135559
rect 1704 135257 1756 135266
rect 1704 135223 1713 135257
rect 1713 135223 1747 135257
rect 1747 135223 1756 135257
rect 1704 135214 1756 135223
rect 216910 135257 216962 135266
rect 216910 135223 216919 135257
rect 216919 135223 216953 135257
rect 216953 135223 216962 135257
rect 216910 135214 216962 135223
rect 1704 134921 1756 134930
rect 1704 134887 1713 134921
rect 1713 134887 1747 134921
rect 1747 134887 1756 134921
rect 1704 134878 1756 134887
rect 216910 134921 216962 134930
rect 216910 134887 216919 134921
rect 216919 134887 216953 134921
rect 216953 134887 216962 134921
rect 216910 134878 216962 134887
rect 1704 134585 1756 134594
rect 1704 134551 1713 134585
rect 1713 134551 1747 134585
rect 1747 134551 1756 134585
rect 1704 134542 1756 134551
rect 216910 134585 216962 134594
rect 216910 134551 216919 134585
rect 216919 134551 216953 134585
rect 216953 134551 216962 134585
rect 216910 134542 216962 134551
rect 1704 134249 1756 134258
rect 1704 134215 1713 134249
rect 1713 134215 1747 134249
rect 1747 134215 1756 134249
rect 1704 134206 1756 134215
rect 216910 134249 216962 134258
rect 216910 134215 216919 134249
rect 216919 134215 216953 134249
rect 216953 134215 216962 134249
rect 216910 134206 216962 134215
rect 1704 133913 1756 133922
rect 1704 133879 1713 133913
rect 1713 133879 1747 133913
rect 1747 133879 1756 133913
rect 1704 133870 1756 133879
rect 216910 133913 216962 133922
rect 216910 133879 216919 133913
rect 216919 133879 216953 133913
rect 216953 133879 216962 133913
rect 216910 133870 216962 133879
rect 1704 133577 1756 133586
rect 1704 133543 1713 133577
rect 1713 133543 1747 133577
rect 1747 133543 1756 133577
rect 1704 133534 1756 133543
rect 216910 133577 216962 133586
rect 216910 133543 216919 133577
rect 216919 133543 216953 133577
rect 216953 133543 216962 133577
rect 216910 133534 216962 133543
rect 1704 133241 1756 133250
rect 1704 133207 1713 133241
rect 1713 133207 1747 133241
rect 1747 133207 1756 133241
rect 1704 133198 1756 133207
rect 216910 133241 216962 133250
rect 216910 133207 216919 133241
rect 216919 133207 216953 133241
rect 216953 133207 216962 133241
rect 216910 133198 216962 133207
rect 29562 133040 29614 133092
rect 34554 133040 34606 133092
rect 39546 133040 39598 133092
rect 44538 133040 44590 133092
rect 49530 133040 49582 133092
rect 54522 133040 54574 133092
rect 59514 133040 59566 133092
rect 64506 133040 64558 133092
rect 69498 133040 69550 133092
rect 74490 133040 74542 133092
rect 79482 133040 79534 133092
rect 84474 133040 84526 133092
rect 89466 133040 89518 133092
rect 94458 133040 94510 133092
rect 99450 133040 99502 133092
rect 104442 133040 104494 133092
rect 109434 133040 109486 133092
rect 114426 133040 114478 133092
rect 119418 133040 119470 133092
rect 124410 133040 124462 133092
rect 129402 133040 129454 133092
rect 134394 133040 134446 133092
rect 139386 133040 139438 133092
rect 144378 133040 144430 133092
rect 149370 133040 149422 133092
rect 154362 133040 154414 133092
rect 159354 133040 159406 133092
rect 164346 133040 164398 133092
rect 169338 133040 169390 133092
rect 174330 133040 174382 133092
rect 179322 133040 179374 133092
rect 184314 133040 184366 133092
rect 1704 132905 1756 132914
rect 1704 132871 1713 132905
rect 1713 132871 1747 132905
rect 1747 132871 1756 132905
rect 1704 132862 1756 132871
rect 216910 132905 216962 132914
rect 216910 132871 216919 132905
rect 216919 132871 216953 132905
rect 216953 132871 216962 132905
rect 216910 132862 216962 132871
rect 1704 132569 1756 132578
rect 1704 132535 1713 132569
rect 1713 132535 1747 132569
rect 1747 132535 1756 132569
rect 1704 132526 1756 132535
rect 216910 132569 216962 132578
rect 216910 132535 216919 132569
rect 216919 132535 216953 132569
rect 216953 132535 216962 132569
rect 216910 132526 216962 132535
rect 1704 132233 1756 132242
rect 1704 132199 1713 132233
rect 1713 132199 1747 132233
rect 1747 132199 1756 132233
rect 1704 132190 1756 132199
rect 216910 132233 216962 132242
rect 216910 132199 216919 132233
rect 216919 132199 216953 132233
rect 216953 132199 216962 132233
rect 216910 132190 216962 132199
rect 1704 131897 1756 131906
rect 1704 131863 1713 131897
rect 1713 131863 1747 131897
rect 1747 131863 1756 131897
rect 1704 131854 1756 131863
rect 216910 131897 216962 131906
rect 216910 131863 216919 131897
rect 216919 131863 216953 131897
rect 216953 131863 216962 131897
rect 216910 131854 216962 131863
rect 1704 131561 1756 131570
rect 1704 131527 1713 131561
rect 1713 131527 1747 131561
rect 1747 131527 1756 131561
rect 1704 131518 1756 131527
rect 216910 131561 216962 131570
rect 216910 131527 216919 131561
rect 216919 131527 216953 131561
rect 216953 131527 216962 131561
rect 216910 131518 216962 131527
rect 1704 131225 1756 131234
rect 1704 131191 1713 131225
rect 1713 131191 1747 131225
rect 1747 131191 1756 131225
rect 1704 131182 1756 131191
rect 216910 131225 216962 131234
rect 216910 131191 216919 131225
rect 216919 131191 216953 131225
rect 216953 131191 216962 131225
rect 216910 131182 216962 131191
rect 1704 130889 1756 130898
rect 1704 130855 1713 130889
rect 1713 130855 1747 130889
rect 1747 130855 1756 130889
rect 1704 130846 1756 130855
rect 216910 130889 216962 130898
rect 216910 130855 216919 130889
rect 216919 130855 216953 130889
rect 216953 130855 216962 130889
rect 216910 130846 216962 130855
rect 1704 130553 1756 130562
rect 1704 130519 1713 130553
rect 1713 130519 1747 130553
rect 1747 130519 1756 130553
rect 1704 130510 1756 130519
rect 216910 130553 216962 130562
rect 216910 130519 216919 130553
rect 216919 130519 216953 130553
rect 216953 130519 216962 130553
rect 216910 130510 216962 130519
rect 1704 130217 1756 130226
rect 1704 130183 1713 130217
rect 1713 130183 1747 130217
rect 1747 130183 1756 130217
rect 1704 130174 1756 130183
rect 216910 130217 216962 130226
rect 216910 130183 216919 130217
rect 216919 130183 216953 130217
rect 216953 130183 216962 130217
rect 216910 130174 216962 130183
rect 1704 129881 1756 129890
rect 1704 129847 1713 129881
rect 1713 129847 1747 129881
rect 1747 129847 1756 129881
rect 1704 129838 1756 129847
rect 216910 129881 216962 129890
rect 216910 129847 216919 129881
rect 216919 129847 216953 129881
rect 216953 129847 216962 129881
rect 216910 129838 216962 129847
rect 1704 129545 1756 129554
rect 1704 129511 1713 129545
rect 1713 129511 1747 129545
rect 1747 129511 1756 129545
rect 1704 129502 1756 129511
rect 216910 129545 216962 129554
rect 216910 129511 216919 129545
rect 216919 129511 216953 129545
rect 216953 129511 216962 129545
rect 216910 129502 216962 129511
rect 1704 129209 1756 129218
rect 1704 129175 1713 129209
rect 1713 129175 1747 129209
rect 1747 129175 1756 129209
rect 1704 129166 1756 129175
rect 216910 129209 216962 129218
rect 216910 129175 216919 129209
rect 216919 129175 216953 129209
rect 216953 129175 216962 129209
rect 216910 129166 216962 129175
rect 1704 128873 1756 128882
rect 1704 128839 1713 128873
rect 1713 128839 1747 128873
rect 1747 128839 1756 128873
rect 1704 128830 1756 128839
rect 216910 128873 216962 128882
rect 216910 128839 216919 128873
rect 216919 128839 216953 128873
rect 216953 128839 216962 128873
rect 216910 128830 216962 128839
rect 1704 128537 1756 128546
rect 1704 128503 1713 128537
rect 1713 128503 1747 128537
rect 1747 128503 1756 128537
rect 1704 128494 1756 128503
rect 216910 128537 216962 128546
rect 216910 128503 216919 128537
rect 216919 128503 216953 128537
rect 216953 128503 216962 128537
rect 216910 128494 216962 128503
rect 1704 128201 1756 128210
rect 1704 128167 1713 128201
rect 1713 128167 1747 128201
rect 1747 128167 1756 128201
rect 1704 128158 1756 128167
rect 216910 128201 216962 128210
rect 216910 128167 216919 128201
rect 216919 128167 216953 128201
rect 216953 128167 216962 128201
rect 216910 128158 216962 128167
rect 1704 127865 1756 127874
rect 1704 127831 1713 127865
rect 1713 127831 1747 127865
rect 1747 127831 1756 127865
rect 1704 127822 1756 127831
rect 216910 127865 216962 127874
rect 216910 127831 216919 127865
rect 216919 127831 216953 127865
rect 216953 127831 216962 127865
rect 216910 127822 216962 127831
rect 1704 127529 1756 127538
rect 1704 127495 1713 127529
rect 1713 127495 1747 127529
rect 1747 127495 1756 127529
rect 1704 127486 1756 127495
rect 216910 127529 216962 127538
rect 216910 127495 216919 127529
rect 216919 127495 216953 127529
rect 216953 127495 216962 127529
rect 216910 127486 216962 127495
rect 1704 127193 1756 127202
rect 1704 127159 1713 127193
rect 1713 127159 1747 127193
rect 1747 127159 1756 127193
rect 1704 127150 1756 127159
rect 216910 127193 216962 127202
rect 216910 127159 216919 127193
rect 216919 127159 216953 127193
rect 216953 127159 216962 127193
rect 216910 127150 216962 127159
rect 1704 126857 1756 126866
rect 1704 126823 1713 126857
rect 1713 126823 1747 126857
rect 1747 126823 1756 126857
rect 1704 126814 1756 126823
rect 216910 126857 216962 126866
rect 216910 126823 216919 126857
rect 216919 126823 216953 126857
rect 216953 126823 216962 126857
rect 216910 126814 216962 126823
rect 1704 126521 1756 126530
rect 1704 126487 1713 126521
rect 1713 126487 1747 126521
rect 1747 126487 1756 126521
rect 1704 126478 1756 126487
rect 216910 126521 216962 126530
rect 216910 126487 216919 126521
rect 216919 126487 216953 126521
rect 216953 126487 216962 126521
rect 216910 126478 216962 126487
rect 1704 126185 1756 126194
rect 1704 126151 1713 126185
rect 1713 126151 1747 126185
rect 1747 126151 1756 126185
rect 1704 126142 1756 126151
rect 216910 126185 216962 126194
rect 216910 126151 216919 126185
rect 216919 126151 216953 126185
rect 216953 126151 216962 126185
rect 216910 126142 216962 126151
rect 1704 125849 1756 125858
rect 1704 125815 1713 125849
rect 1713 125815 1747 125849
rect 1747 125815 1756 125849
rect 1704 125806 1756 125815
rect 216910 125849 216962 125858
rect 216910 125815 216919 125849
rect 216919 125815 216953 125849
rect 216953 125815 216962 125849
rect 216910 125806 216962 125815
rect 1704 125513 1756 125522
rect 1704 125479 1713 125513
rect 1713 125479 1747 125513
rect 1747 125479 1756 125513
rect 1704 125470 1756 125479
rect 216910 125513 216962 125522
rect 216910 125479 216919 125513
rect 216919 125479 216953 125513
rect 216953 125479 216962 125513
rect 216910 125470 216962 125479
rect 1704 125177 1756 125186
rect 1704 125143 1713 125177
rect 1713 125143 1747 125177
rect 1747 125143 1756 125177
rect 1704 125134 1756 125143
rect 216910 125177 216962 125186
rect 216910 125143 216919 125177
rect 216919 125143 216953 125177
rect 216953 125143 216962 125177
rect 216910 125134 216962 125143
rect 1704 124841 1756 124850
rect 1704 124807 1713 124841
rect 1713 124807 1747 124841
rect 1747 124807 1756 124841
rect 1704 124798 1756 124807
rect 216910 124841 216962 124850
rect 216910 124807 216919 124841
rect 216919 124807 216953 124841
rect 216953 124807 216962 124841
rect 216910 124798 216962 124807
rect 1704 124505 1756 124514
rect 1704 124471 1713 124505
rect 1713 124471 1747 124505
rect 1747 124471 1756 124505
rect 1704 124462 1756 124471
rect 216910 124505 216962 124514
rect 216910 124471 216919 124505
rect 216919 124471 216953 124505
rect 216953 124471 216962 124505
rect 216910 124462 216962 124471
rect 1704 124169 1756 124178
rect 1704 124135 1713 124169
rect 1713 124135 1747 124169
rect 1747 124135 1756 124169
rect 1704 124126 1756 124135
rect 216910 124169 216962 124178
rect 216910 124135 216919 124169
rect 216919 124135 216953 124169
rect 216953 124135 216962 124169
rect 216910 124126 216962 124135
rect 1704 123833 1756 123842
rect 1704 123799 1713 123833
rect 1713 123799 1747 123833
rect 1747 123799 1756 123833
rect 1704 123790 1756 123799
rect 216910 123833 216962 123842
rect 216910 123799 216919 123833
rect 216919 123799 216953 123833
rect 216953 123799 216962 123833
rect 216910 123790 216962 123799
rect 1704 123497 1756 123506
rect 1704 123463 1713 123497
rect 1713 123463 1747 123497
rect 1747 123463 1756 123497
rect 1704 123454 1756 123463
rect 216910 123497 216962 123506
rect 216910 123463 216919 123497
rect 216919 123463 216953 123497
rect 216953 123463 216962 123497
rect 216910 123454 216962 123463
rect 1704 123161 1756 123170
rect 1704 123127 1713 123161
rect 1713 123127 1747 123161
rect 1747 123127 1756 123161
rect 1704 123118 1756 123127
rect 216910 123161 216962 123170
rect 216910 123127 216919 123161
rect 216919 123127 216953 123161
rect 216953 123127 216962 123161
rect 216910 123118 216962 123127
rect 1704 122825 1756 122834
rect 1704 122791 1713 122825
rect 1713 122791 1747 122825
rect 1747 122791 1756 122825
rect 1704 122782 1756 122791
rect 216910 122825 216962 122834
rect 216910 122791 216919 122825
rect 216919 122791 216953 122825
rect 216953 122791 216962 122825
rect 216910 122782 216962 122791
rect 1704 122489 1756 122498
rect 1704 122455 1713 122489
rect 1713 122455 1747 122489
rect 1747 122455 1756 122489
rect 1704 122446 1756 122455
rect 216910 122489 216962 122498
rect 216910 122455 216919 122489
rect 216919 122455 216953 122489
rect 216953 122455 216962 122489
rect 216910 122446 216962 122455
rect 1704 122153 1756 122162
rect 1704 122119 1713 122153
rect 1713 122119 1747 122153
rect 1747 122119 1756 122153
rect 1704 122110 1756 122119
rect 216910 122153 216962 122162
rect 216910 122119 216919 122153
rect 216919 122119 216953 122153
rect 216953 122119 216962 122153
rect 216910 122110 216962 122119
rect 1704 121817 1756 121826
rect 1704 121783 1713 121817
rect 1713 121783 1747 121817
rect 1747 121783 1756 121817
rect 1704 121774 1756 121783
rect 216910 121817 216962 121826
rect 216910 121783 216919 121817
rect 216919 121783 216953 121817
rect 216953 121783 216962 121817
rect 216910 121774 216962 121783
rect 1704 121481 1756 121490
rect 1704 121447 1713 121481
rect 1713 121447 1747 121481
rect 1747 121447 1756 121481
rect 1704 121438 1756 121447
rect 216910 121481 216962 121490
rect 216910 121447 216919 121481
rect 216919 121447 216953 121481
rect 216953 121447 216962 121481
rect 216910 121438 216962 121447
rect 1704 121145 1756 121154
rect 1704 121111 1713 121145
rect 1713 121111 1747 121145
rect 1747 121111 1756 121145
rect 1704 121102 1756 121111
rect 216910 121145 216962 121154
rect 216910 121111 216919 121145
rect 216919 121111 216953 121145
rect 216953 121111 216962 121145
rect 216910 121102 216962 121111
rect 1704 120809 1756 120818
rect 1704 120775 1713 120809
rect 1713 120775 1747 120809
rect 1747 120775 1756 120809
rect 1704 120766 1756 120775
rect 216910 120809 216962 120818
rect 216910 120775 216919 120809
rect 216919 120775 216953 120809
rect 216953 120775 216962 120809
rect 216910 120766 216962 120775
rect 1704 120473 1756 120482
rect 1704 120439 1713 120473
rect 1713 120439 1747 120473
rect 1747 120439 1756 120473
rect 1704 120430 1756 120439
rect 216910 120473 216962 120482
rect 216910 120439 216919 120473
rect 216919 120439 216953 120473
rect 216953 120439 216962 120473
rect 216910 120430 216962 120439
rect 1704 120137 1756 120146
rect 1704 120103 1713 120137
rect 1713 120103 1747 120137
rect 1747 120103 1756 120137
rect 1704 120094 1756 120103
rect 216910 120137 216962 120146
rect 216910 120103 216919 120137
rect 216919 120103 216953 120137
rect 216953 120103 216962 120137
rect 216910 120094 216962 120103
rect 1704 119801 1756 119810
rect 1704 119767 1713 119801
rect 1713 119767 1747 119801
rect 1747 119767 1756 119801
rect 1704 119758 1756 119767
rect 216910 119801 216962 119810
rect 216910 119767 216919 119801
rect 216919 119767 216953 119801
rect 216953 119767 216962 119801
rect 216910 119758 216962 119767
rect 1704 119465 1756 119474
rect 1704 119431 1713 119465
rect 1713 119431 1747 119465
rect 1747 119431 1756 119465
rect 1704 119422 1756 119431
rect 216910 119465 216962 119474
rect 216910 119431 216919 119465
rect 216919 119431 216953 119465
rect 216953 119431 216962 119465
rect 216910 119422 216962 119431
rect 1704 119129 1756 119138
rect 1704 119095 1713 119129
rect 1713 119095 1747 119129
rect 1747 119095 1756 119129
rect 1704 119086 1756 119095
rect 216910 119129 216962 119138
rect 216910 119095 216919 119129
rect 216919 119095 216953 119129
rect 216953 119095 216962 119129
rect 216910 119086 216962 119095
rect 1704 118793 1756 118802
rect 1704 118759 1713 118793
rect 1713 118759 1747 118793
rect 1747 118759 1756 118793
rect 1704 118750 1756 118759
rect 216910 118793 216962 118802
rect 216910 118759 216919 118793
rect 216919 118759 216953 118793
rect 216953 118759 216962 118793
rect 216910 118750 216962 118759
rect 1704 118457 1756 118466
rect 1704 118423 1713 118457
rect 1713 118423 1747 118457
rect 1747 118423 1756 118457
rect 1704 118414 1756 118423
rect 216910 118457 216962 118466
rect 216910 118423 216919 118457
rect 216919 118423 216953 118457
rect 216953 118423 216962 118457
rect 216910 118414 216962 118423
rect 1704 118121 1756 118130
rect 1704 118087 1713 118121
rect 1713 118087 1747 118121
rect 1747 118087 1756 118121
rect 1704 118078 1756 118087
rect 216910 118121 216962 118130
rect 216910 118087 216919 118121
rect 216919 118087 216953 118121
rect 216953 118087 216962 118121
rect 216910 118078 216962 118087
rect 1704 117785 1756 117794
rect 1704 117751 1713 117785
rect 1713 117751 1747 117785
rect 1747 117751 1756 117785
rect 1704 117742 1756 117751
rect 216910 117785 216962 117794
rect 216910 117751 216919 117785
rect 216919 117751 216953 117785
rect 216953 117751 216962 117785
rect 216910 117742 216962 117751
rect 1704 117449 1756 117458
rect 1704 117415 1713 117449
rect 1713 117415 1747 117449
rect 1747 117415 1756 117449
rect 1704 117406 1756 117415
rect 216910 117449 216962 117458
rect 216910 117415 216919 117449
rect 216919 117415 216953 117449
rect 216953 117415 216962 117449
rect 216910 117406 216962 117415
rect 1704 117113 1756 117122
rect 1704 117079 1713 117113
rect 1713 117079 1747 117113
rect 1747 117079 1756 117113
rect 1704 117070 1756 117079
rect 216910 117113 216962 117122
rect 216910 117079 216919 117113
rect 216919 117079 216953 117113
rect 216953 117079 216962 117113
rect 216910 117070 216962 117079
rect 1704 116777 1756 116786
rect 1704 116743 1713 116777
rect 1713 116743 1747 116777
rect 1747 116743 1756 116777
rect 1704 116734 1756 116743
rect 216910 116777 216962 116786
rect 216910 116743 216919 116777
rect 216919 116743 216953 116777
rect 216953 116743 216962 116777
rect 216910 116734 216962 116743
rect 1704 116441 1756 116450
rect 1704 116407 1713 116441
rect 1713 116407 1747 116441
rect 1747 116407 1756 116441
rect 1704 116398 1756 116407
rect 216910 116441 216962 116450
rect 216910 116407 216919 116441
rect 216919 116407 216953 116441
rect 216953 116407 216962 116441
rect 216910 116398 216962 116407
rect 1704 116105 1756 116114
rect 1704 116071 1713 116105
rect 1713 116071 1747 116105
rect 1747 116071 1756 116105
rect 1704 116062 1756 116071
rect 216910 116105 216962 116114
rect 216910 116071 216919 116105
rect 216919 116071 216953 116105
rect 216953 116071 216962 116105
rect 216910 116062 216962 116071
rect 1704 115769 1756 115778
rect 1704 115735 1713 115769
rect 1713 115735 1747 115769
rect 1747 115735 1756 115769
rect 1704 115726 1756 115735
rect 216910 115769 216962 115778
rect 216910 115735 216919 115769
rect 216919 115735 216953 115769
rect 216953 115735 216962 115769
rect 216910 115726 216962 115735
rect 1704 115433 1756 115442
rect 1704 115399 1713 115433
rect 1713 115399 1747 115433
rect 1747 115399 1756 115433
rect 1704 115390 1756 115399
rect 216910 115433 216962 115442
rect 216910 115399 216919 115433
rect 216919 115399 216953 115433
rect 216953 115399 216962 115433
rect 216910 115390 216962 115399
rect 1704 115097 1756 115106
rect 1704 115063 1713 115097
rect 1713 115063 1747 115097
rect 1747 115063 1756 115097
rect 1704 115054 1756 115063
rect 216910 115097 216962 115106
rect 216910 115063 216919 115097
rect 216919 115063 216953 115097
rect 216953 115063 216962 115097
rect 216910 115054 216962 115063
rect 1704 114761 1756 114770
rect 1704 114727 1713 114761
rect 1713 114727 1747 114761
rect 1747 114727 1756 114761
rect 1704 114718 1756 114727
rect 216910 114761 216962 114770
rect 216910 114727 216919 114761
rect 216919 114727 216953 114761
rect 216953 114727 216962 114761
rect 216910 114718 216962 114727
rect 1704 114425 1756 114434
rect 1704 114391 1713 114425
rect 1713 114391 1747 114425
rect 1747 114391 1756 114425
rect 1704 114382 1756 114391
rect 216910 114425 216962 114434
rect 216910 114391 216919 114425
rect 216919 114391 216953 114425
rect 216953 114391 216962 114425
rect 216910 114382 216962 114391
rect 1704 114089 1756 114098
rect 1704 114055 1713 114089
rect 1713 114055 1747 114089
rect 1747 114055 1756 114089
rect 1704 114046 1756 114055
rect 216910 114089 216962 114098
rect 216910 114055 216919 114089
rect 216919 114055 216953 114089
rect 216953 114055 216962 114089
rect 216910 114046 216962 114055
rect 1704 113753 1756 113762
rect 1704 113719 1713 113753
rect 1713 113719 1747 113753
rect 1747 113719 1756 113753
rect 1704 113710 1756 113719
rect 216910 113753 216962 113762
rect 216910 113719 216919 113753
rect 216919 113719 216953 113753
rect 216953 113719 216962 113753
rect 216910 113710 216962 113719
rect 1704 113417 1756 113426
rect 1704 113383 1713 113417
rect 1713 113383 1747 113417
rect 1747 113383 1756 113417
rect 1704 113374 1756 113383
rect 216910 113417 216962 113426
rect 216910 113383 216919 113417
rect 216919 113383 216953 113417
rect 216953 113383 216962 113417
rect 216910 113374 216962 113383
rect 1704 113081 1756 113090
rect 1704 113047 1713 113081
rect 1713 113047 1747 113081
rect 1747 113047 1756 113081
rect 1704 113038 1756 113047
rect 216910 113081 216962 113090
rect 216910 113047 216919 113081
rect 216919 113047 216953 113081
rect 216953 113047 216962 113081
rect 216910 113038 216962 113047
rect 1704 112745 1756 112754
rect 1704 112711 1713 112745
rect 1713 112711 1747 112745
rect 1747 112711 1756 112745
rect 1704 112702 1756 112711
rect 216910 112745 216962 112754
rect 216910 112711 216919 112745
rect 216919 112711 216953 112745
rect 216953 112711 216962 112745
rect 216910 112702 216962 112711
rect 1704 112409 1756 112418
rect 1704 112375 1713 112409
rect 1713 112375 1747 112409
rect 1747 112375 1756 112409
rect 1704 112366 1756 112375
rect 216910 112409 216962 112418
rect 216910 112375 216919 112409
rect 216919 112375 216953 112409
rect 216953 112375 216962 112409
rect 216910 112366 216962 112375
rect 1704 112073 1756 112082
rect 1704 112039 1713 112073
rect 1713 112039 1747 112073
rect 1747 112039 1756 112073
rect 1704 112030 1756 112039
rect 216910 112073 216962 112082
rect 216910 112039 216919 112073
rect 216919 112039 216953 112073
rect 216953 112039 216962 112073
rect 216910 112030 216962 112039
rect 1704 111737 1756 111746
rect 1704 111703 1713 111737
rect 1713 111703 1747 111737
rect 1747 111703 1756 111737
rect 1704 111694 1756 111703
rect 216910 111737 216962 111746
rect 216910 111703 216919 111737
rect 216919 111703 216953 111737
rect 216953 111703 216962 111737
rect 216910 111694 216962 111703
rect 1704 111401 1756 111410
rect 1704 111367 1713 111401
rect 1713 111367 1747 111401
rect 1747 111367 1756 111401
rect 1704 111358 1756 111367
rect 216910 111401 216962 111410
rect 216910 111367 216919 111401
rect 216919 111367 216953 111401
rect 216953 111367 216962 111401
rect 216910 111358 216962 111367
rect 1704 111065 1756 111074
rect 1704 111031 1713 111065
rect 1713 111031 1747 111065
rect 1747 111031 1756 111065
rect 1704 111022 1756 111031
rect 216910 111065 216962 111074
rect 216910 111031 216919 111065
rect 216919 111031 216953 111065
rect 216953 111031 216962 111065
rect 216910 111022 216962 111031
rect 1704 110729 1756 110738
rect 1704 110695 1713 110729
rect 1713 110695 1747 110729
rect 1747 110695 1756 110729
rect 1704 110686 1756 110695
rect 216910 110729 216962 110738
rect 216910 110695 216919 110729
rect 216919 110695 216953 110729
rect 216953 110695 216962 110729
rect 216910 110686 216962 110695
rect 1704 110393 1756 110402
rect 1704 110359 1713 110393
rect 1713 110359 1747 110393
rect 1747 110359 1756 110393
rect 1704 110350 1756 110359
rect 216910 110393 216962 110402
rect 216910 110359 216919 110393
rect 216919 110359 216953 110393
rect 216953 110359 216962 110393
rect 216910 110350 216962 110359
rect 1704 110057 1756 110066
rect 1704 110023 1713 110057
rect 1713 110023 1747 110057
rect 1747 110023 1756 110057
rect 1704 110014 1756 110023
rect 216910 110057 216962 110066
rect 216910 110023 216919 110057
rect 216919 110023 216953 110057
rect 216953 110023 216962 110057
rect 216910 110014 216962 110023
rect 1704 109721 1756 109730
rect 1704 109687 1713 109721
rect 1713 109687 1747 109721
rect 1747 109687 1756 109721
rect 1704 109678 1756 109687
rect 216910 109721 216962 109730
rect 216910 109687 216919 109721
rect 216919 109687 216953 109721
rect 216953 109687 216962 109721
rect 216910 109678 216962 109687
rect 1704 109385 1756 109394
rect 1704 109351 1713 109385
rect 1713 109351 1747 109385
rect 1747 109351 1756 109385
rect 1704 109342 1756 109351
rect 216910 109385 216962 109394
rect 216910 109351 216919 109385
rect 216919 109351 216953 109385
rect 216953 109351 216962 109385
rect 216910 109342 216962 109351
rect 1704 109049 1756 109058
rect 1704 109015 1713 109049
rect 1713 109015 1747 109049
rect 1747 109015 1756 109049
rect 1704 109006 1756 109015
rect 216910 109049 216962 109058
rect 216910 109015 216919 109049
rect 216919 109015 216953 109049
rect 216953 109015 216962 109049
rect 216910 109006 216962 109015
rect 1704 108713 1756 108722
rect 1704 108679 1713 108713
rect 1713 108679 1747 108713
rect 1747 108679 1756 108713
rect 1704 108670 1756 108679
rect 216910 108713 216962 108722
rect 216910 108679 216919 108713
rect 216919 108679 216953 108713
rect 216953 108679 216962 108713
rect 216910 108670 216962 108679
rect 1704 108377 1756 108386
rect 1704 108343 1713 108377
rect 1713 108343 1747 108377
rect 1747 108343 1756 108377
rect 1704 108334 1756 108343
rect 216910 108377 216962 108386
rect 216910 108343 216919 108377
rect 216919 108343 216953 108377
rect 216953 108343 216962 108377
rect 216910 108334 216962 108343
rect 1704 108041 1756 108050
rect 1704 108007 1713 108041
rect 1713 108007 1747 108041
rect 1747 108007 1756 108041
rect 1704 107998 1756 108007
rect 216910 108041 216962 108050
rect 216910 108007 216919 108041
rect 216919 108007 216953 108041
rect 216953 108007 216962 108041
rect 216910 107998 216962 108007
rect 1704 107705 1756 107714
rect 1704 107671 1713 107705
rect 1713 107671 1747 107705
rect 1747 107671 1756 107705
rect 1704 107662 1756 107671
rect 216910 107705 216962 107714
rect 216910 107671 216919 107705
rect 216919 107671 216953 107705
rect 216953 107671 216962 107705
rect 216910 107662 216962 107671
rect 1704 107369 1756 107378
rect 1704 107335 1713 107369
rect 1713 107335 1747 107369
rect 1747 107335 1756 107369
rect 1704 107326 1756 107335
rect 216910 107369 216962 107378
rect 216910 107335 216919 107369
rect 216919 107335 216953 107369
rect 216953 107335 216962 107369
rect 216910 107326 216962 107335
rect 1704 107033 1756 107042
rect 1704 106999 1713 107033
rect 1713 106999 1747 107033
rect 1747 106999 1756 107033
rect 1704 106990 1756 106999
rect 216910 107033 216962 107042
rect 216910 106999 216919 107033
rect 216919 106999 216953 107033
rect 216953 106999 216962 107033
rect 216910 106990 216962 106999
rect 1704 106697 1756 106706
rect 1704 106663 1713 106697
rect 1713 106663 1747 106697
rect 1747 106663 1756 106697
rect 1704 106654 1756 106663
rect 216910 106697 216962 106706
rect 216910 106663 216919 106697
rect 216919 106663 216953 106697
rect 216953 106663 216962 106697
rect 216910 106654 216962 106663
rect 1704 106361 1756 106370
rect 1704 106327 1713 106361
rect 1713 106327 1747 106361
rect 1747 106327 1756 106361
rect 1704 106318 1756 106327
rect 216910 106361 216962 106370
rect 216910 106327 216919 106361
rect 216919 106327 216953 106361
rect 216953 106327 216962 106361
rect 216910 106318 216962 106327
rect 1704 106025 1756 106034
rect 1704 105991 1713 106025
rect 1713 105991 1747 106025
rect 1747 105991 1756 106025
rect 1704 105982 1756 105991
rect 216910 106025 216962 106034
rect 216910 105991 216919 106025
rect 216919 105991 216953 106025
rect 216953 105991 216962 106025
rect 216910 105982 216962 105991
rect 1704 105689 1756 105698
rect 1704 105655 1713 105689
rect 1713 105655 1747 105689
rect 1747 105655 1756 105689
rect 1704 105646 1756 105655
rect 216910 105689 216962 105698
rect 216910 105655 216919 105689
rect 216919 105655 216953 105689
rect 216953 105655 216962 105689
rect 216910 105646 216962 105655
rect 1704 105353 1756 105362
rect 1704 105319 1713 105353
rect 1713 105319 1747 105353
rect 1747 105319 1756 105353
rect 1704 105310 1756 105319
rect 216910 105353 216962 105362
rect 216910 105319 216919 105353
rect 216919 105319 216953 105353
rect 216953 105319 216962 105353
rect 216910 105310 216962 105319
rect 1704 105017 1756 105026
rect 1704 104983 1713 105017
rect 1713 104983 1747 105017
rect 1747 104983 1756 105017
rect 1704 104974 1756 104983
rect 216910 105017 216962 105026
rect 216910 104983 216919 105017
rect 216919 104983 216953 105017
rect 216953 104983 216962 105017
rect 216910 104974 216962 104983
rect 1704 104681 1756 104690
rect 1704 104647 1713 104681
rect 1713 104647 1747 104681
rect 1747 104647 1756 104681
rect 1704 104638 1756 104647
rect 216910 104681 216962 104690
rect 216910 104647 216919 104681
rect 216919 104647 216953 104681
rect 216953 104647 216962 104681
rect 216910 104638 216962 104647
rect 1704 104345 1756 104354
rect 1704 104311 1713 104345
rect 1713 104311 1747 104345
rect 1747 104311 1756 104345
rect 1704 104302 1756 104311
rect 216910 104345 216962 104354
rect 216910 104311 216919 104345
rect 216919 104311 216953 104345
rect 216953 104311 216962 104345
rect 216910 104302 216962 104311
rect 1704 104009 1756 104018
rect 1704 103975 1713 104009
rect 1713 103975 1747 104009
rect 1747 103975 1756 104009
rect 1704 103966 1756 103975
rect 216910 104009 216962 104018
rect 216910 103975 216919 104009
rect 216919 103975 216953 104009
rect 216953 103975 216962 104009
rect 216910 103966 216962 103975
rect 1704 103673 1756 103682
rect 1704 103639 1713 103673
rect 1713 103639 1747 103673
rect 1747 103639 1756 103673
rect 1704 103630 1756 103639
rect 216910 103673 216962 103682
rect 216910 103639 216919 103673
rect 216919 103639 216953 103673
rect 216953 103639 216962 103673
rect 216910 103630 216962 103639
rect 1704 103337 1756 103346
rect 1704 103303 1713 103337
rect 1713 103303 1747 103337
rect 1747 103303 1756 103337
rect 1704 103294 1756 103303
rect 216910 103337 216962 103346
rect 216910 103303 216919 103337
rect 216919 103303 216953 103337
rect 216953 103303 216962 103337
rect 216910 103294 216962 103303
rect 1704 103001 1756 103010
rect 1704 102967 1713 103001
rect 1713 102967 1747 103001
rect 1747 102967 1756 103001
rect 1704 102958 1756 102967
rect 216910 103001 216962 103010
rect 216910 102967 216919 103001
rect 216919 102967 216953 103001
rect 216953 102967 216962 103001
rect 216910 102958 216962 102967
rect 1704 102665 1756 102674
rect 1704 102631 1713 102665
rect 1713 102631 1747 102665
rect 1747 102631 1756 102665
rect 1704 102622 1756 102631
rect 216910 102665 216962 102674
rect 216910 102631 216919 102665
rect 216919 102631 216953 102665
rect 216953 102631 216962 102665
rect 216910 102622 216962 102631
rect 1704 102329 1756 102338
rect 1704 102295 1713 102329
rect 1713 102295 1747 102329
rect 1747 102295 1756 102329
rect 1704 102286 1756 102295
rect 216910 102329 216962 102338
rect 216910 102295 216919 102329
rect 216919 102295 216953 102329
rect 216953 102295 216962 102329
rect 216910 102286 216962 102295
rect 1704 101993 1756 102002
rect 1704 101959 1713 101993
rect 1713 101959 1747 101993
rect 1747 101959 1756 101993
rect 1704 101950 1756 101959
rect 216910 101993 216962 102002
rect 216910 101959 216919 101993
rect 216919 101959 216953 101993
rect 216953 101959 216962 101993
rect 216910 101950 216962 101959
rect 1704 101657 1756 101666
rect 1704 101623 1713 101657
rect 1713 101623 1747 101657
rect 1747 101623 1756 101657
rect 1704 101614 1756 101623
rect 216910 101657 216962 101666
rect 216910 101623 216919 101657
rect 216919 101623 216953 101657
rect 216953 101623 216962 101657
rect 216910 101614 216962 101623
rect 1704 101321 1756 101330
rect 1704 101287 1713 101321
rect 1713 101287 1747 101321
rect 1747 101287 1756 101321
rect 1704 101278 1756 101287
rect 216910 101321 216962 101330
rect 216910 101287 216919 101321
rect 216919 101287 216953 101321
rect 216953 101287 216962 101321
rect 216910 101278 216962 101287
rect 1704 100985 1756 100994
rect 1704 100951 1713 100985
rect 1713 100951 1747 100985
rect 1747 100951 1756 100985
rect 1704 100942 1756 100951
rect 216910 100985 216962 100994
rect 216910 100951 216919 100985
rect 216919 100951 216953 100985
rect 216953 100951 216962 100985
rect 216910 100942 216962 100951
rect 1704 100649 1756 100658
rect 1704 100615 1713 100649
rect 1713 100615 1747 100649
rect 1747 100615 1756 100649
rect 1704 100606 1756 100615
rect 216910 100649 216962 100658
rect 216910 100615 216919 100649
rect 216919 100615 216953 100649
rect 216953 100615 216962 100649
rect 216910 100606 216962 100615
rect 1704 100313 1756 100322
rect 1704 100279 1713 100313
rect 1713 100279 1747 100313
rect 1747 100279 1756 100313
rect 1704 100270 1756 100279
rect 216910 100313 216962 100322
rect 216910 100279 216919 100313
rect 216919 100279 216953 100313
rect 216953 100279 216962 100313
rect 216910 100270 216962 100279
rect 1704 99977 1756 99986
rect 1704 99943 1713 99977
rect 1713 99943 1747 99977
rect 1747 99943 1756 99977
rect 1704 99934 1756 99943
rect 216910 99977 216962 99986
rect 216910 99943 216919 99977
rect 216919 99943 216953 99977
rect 216953 99943 216962 99977
rect 216910 99934 216962 99943
rect 1704 99641 1756 99650
rect 1704 99607 1713 99641
rect 1713 99607 1747 99641
rect 1747 99607 1756 99641
rect 1704 99598 1756 99607
rect 216910 99641 216962 99650
rect 216910 99607 216919 99641
rect 216919 99607 216953 99641
rect 216953 99607 216962 99641
rect 216910 99598 216962 99607
rect 1704 99305 1756 99314
rect 1704 99271 1713 99305
rect 1713 99271 1747 99305
rect 1747 99271 1756 99305
rect 1704 99262 1756 99271
rect 216910 99305 216962 99314
rect 216910 99271 216919 99305
rect 216919 99271 216953 99305
rect 216953 99271 216962 99305
rect 216910 99262 216962 99271
rect 1704 98969 1756 98978
rect 1704 98935 1713 98969
rect 1713 98935 1747 98969
rect 1747 98935 1756 98969
rect 1704 98926 1756 98935
rect 216910 98969 216962 98978
rect 216910 98935 216919 98969
rect 216919 98935 216953 98969
rect 216953 98935 216962 98969
rect 216910 98926 216962 98935
rect 1704 98633 1756 98642
rect 1704 98599 1713 98633
rect 1713 98599 1747 98633
rect 1747 98599 1756 98633
rect 1704 98590 1756 98599
rect 216910 98633 216962 98642
rect 216910 98599 216919 98633
rect 216919 98599 216953 98633
rect 216953 98599 216962 98633
rect 216910 98590 216962 98599
rect 1704 98297 1756 98306
rect 1704 98263 1713 98297
rect 1713 98263 1747 98297
rect 1747 98263 1756 98297
rect 1704 98254 1756 98263
rect 216910 98297 216962 98306
rect 216910 98263 216919 98297
rect 216919 98263 216953 98297
rect 216953 98263 216962 98297
rect 216910 98254 216962 98263
rect 1704 97961 1756 97970
rect 1704 97927 1713 97961
rect 1713 97927 1747 97961
rect 1747 97927 1756 97961
rect 1704 97918 1756 97927
rect 216910 97961 216962 97970
rect 216910 97927 216919 97961
rect 216919 97927 216953 97961
rect 216953 97927 216962 97961
rect 216910 97918 216962 97927
rect 1704 97625 1756 97634
rect 1704 97591 1713 97625
rect 1713 97591 1747 97625
rect 1747 97591 1756 97625
rect 1704 97582 1756 97591
rect 216910 97625 216962 97634
rect 216910 97591 216919 97625
rect 216919 97591 216953 97625
rect 216953 97591 216962 97625
rect 216910 97582 216962 97591
rect 1704 97289 1756 97298
rect 1704 97255 1713 97289
rect 1713 97255 1747 97289
rect 1747 97255 1756 97289
rect 1704 97246 1756 97255
rect 216910 97289 216962 97298
rect 216910 97255 216919 97289
rect 216919 97255 216953 97289
rect 216953 97255 216962 97289
rect 216910 97246 216962 97255
rect 1704 96953 1756 96962
rect 1704 96919 1713 96953
rect 1713 96919 1747 96953
rect 1747 96919 1756 96953
rect 1704 96910 1756 96919
rect 216910 96953 216962 96962
rect 216910 96919 216919 96953
rect 216919 96919 216953 96953
rect 216953 96919 216962 96953
rect 216910 96910 216962 96919
rect 1704 96617 1756 96626
rect 1704 96583 1713 96617
rect 1713 96583 1747 96617
rect 1747 96583 1756 96617
rect 1704 96574 1756 96583
rect 216910 96617 216962 96626
rect 216910 96583 216919 96617
rect 216919 96583 216953 96617
rect 216953 96583 216962 96617
rect 216910 96574 216962 96583
rect 1704 96281 1756 96290
rect 1704 96247 1713 96281
rect 1713 96247 1747 96281
rect 1747 96247 1756 96281
rect 1704 96238 1756 96247
rect 216910 96281 216962 96290
rect 216910 96247 216919 96281
rect 216919 96247 216953 96281
rect 216953 96247 216962 96281
rect 216910 96238 216962 96247
rect 1704 95945 1756 95954
rect 1704 95911 1713 95945
rect 1713 95911 1747 95945
rect 1747 95911 1756 95945
rect 1704 95902 1756 95911
rect 216910 95945 216962 95954
rect 216910 95911 216919 95945
rect 216919 95911 216953 95945
rect 216953 95911 216962 95945
rect 216910 95902 216962 95911
rect 1704 95609 1756 95618
rect 1704 95575 1713 95609
rect 1713 95575 1747 95609
rect 1747 95575 1756 95609
rect 1704 95566 1756 95575
rect 216910 95609 216962 95618
rect 216910 95575 216919 95609
rect 216919 95575 216953 95609
rect 216953 95575 216962 95609
rect 216910 95566 216962 95575
rect 1704 95273 1756 95282
rect 1704 95239 1713 95273
rect 1713 95239 1747 95273
rect 1747 95239 1756 95273
rect 1704 95230 1756 95239
rect 216910 95273 216962 95282
rect 216910 95239 216919 95273
rect 216919 95239 216953 95273
rect 216953 95239 216962 95273
rect 216910 95230 216962 95239
rect 1704 94937 1756 94946
rect 1704 94903 1713 94937
rect 1713 94903 1747 94937
rect 1747 94903 1756 94937
rect 1704 94894 1756 94903
rect 216910 94937 216962 94946
rect 216910 94903 216919 94937
rect 216919 94903 216953 94937
rect 216953 94903 216962 94937
rect 216910 94894 216962 94903
rect 1704 94601 1756 94610
rect 1704 94567 1713 94601
rect 1713 94567 1747 94601
rect 1747 94567 1756 94601
rect 1704 94558 1756 94567
rect 216910 94601 216962 94610
rect 216910 94567 216919 94601
rect 216919 94567 216953 94601
rect 216953 94567 216962 94601
rect 216910 94558 216962 94567
rect 1704 94265 1756 94274
rect 1704 94231 1713 94265
rect 1713 94231 1747 94265
rect 1747 94231 1756 94265
rect 1704 94222 1756 94231
rect 216910 94265 216962 94274
rect 216910 94231 216919 94265
rect 216919 94231 216953 94265
rect 216953 94231 216962 94265
rect 216910 94222 216962 94231
rect 1704 93929 1756 93938
rect 1704 93895 1713 93929
rect 1713 93895 1747 93929
rect 1747 93895 1756 93929
rect 1704 93886 1756 93895
rect 216910 93929 216962 93938
rect 216910 93895 216919 93929
rect 216919 93895 216953 93929
rect 216953 93895 216962 93929
rect 216910 93886 216962 93895
rect 1704 93593 1756 93602
rect 1704 93559 1713 93593
rect 1713 93559 1747 93593
rect 1747 93559 1756 93593
rect 1704 93550 1756 93559
rect 216910 93593 216962 93602
rect 216910 93559 216919 93593
rect 216919 93559 216953 93593
rect 216953 93559 216962 93593
rect 216910 93550 216962 93559
rect 1704 93257 1756 93266
rect 1704 93223 1713 93257
rect 1713 93223 1747 93257
rect 1747 93223 1756 93257
rect 1704 93214 1756 93223
rect 216910 93257 216962 93266
rect 216910 93223 216919 93257
rect 216919 93223 216953 93257
rect 216953 93223 216962 93257
rect 216910 93214 216962 93223
rect 1704 92921 1756 92930
rect 1704 92887 1713 92921
rect 1713 92887 1747 92921
rect 1747 92887 1756 92921
rect 1704 92878 1756 92887
rect 216910 92921 216962 92930
rect 216910 92887 216919 92921
rect 216919 92887 216953 92921
rect 216953 92887 216962 92921
rect 216910 92878 216962 92887
rect 1704 92585 1756 92594
rect 1704 92551 1713 92585
rect 1713 92551 1747 92585
rect 1747 92551 1756 92585
rect 1704 92542 1756 92551
rect 216910 92585 216962 92594
rect 216910 92551 216919 92585
rect 216919 92551 216953 92585
rect 216953 92551 216962 92585
rect 216910 92542 216962 92551
rect 1704 92249 1756 92258
rect 1704 92215 1713 92249
rect 1713 92215 1747 92249
rect 1747 92215 1756 92249
rect 1704 92206 1756 92215
rect 216910 92249 216962 92258
rect 216910 92215 216919 92249
rect 216919 92215 216953 92249
rect 216953 92215 216962 92249
rect 216910 92206 216962 92215
rect 1704 91913 1756 91922
rect 1704 91879 1713 91913
rect 1713 91879 1747 91913
rect 1747 91879 1756 91913
rect 1704 91870 1756 91879
rect 216910 91913 216962 91922
rect 216910 91879 216919 91913
rect 216919 91879 216953 91913
rect 216953 91879 216962 91913
rect 216910 91870 216962 91879
rect 1704 91577 1756 91586
rect 1704 91543 1713 91577
rect 1713 91543 1747 91577
rect 1747 91543 1756 91577
rect 1704 91534 1756 91543
rect 216910 91577 216962 91586
rect 216910 91543 216919 91577
rect 216919 91543 216953 91577
rect 216953 91543 216962 91577
rect 216910 91534 216962 91543
rect 1704 91241 1756 91250
rect 1704 91207 1713 91241
rect 1713 91207 1747 91241
rect 1747 91207 1756 91241
rect 1704 91198 1756 91207
rect 216910 91241 216962 91250
rect 216910 91207 216919 91241
rect 216919 91207 216953 91241
rect 216953 91207 216962 91241
rect 216910 91198 216962 91207
rect 1704 90905 1756 90914
rect 1704 90871 1713 90905
rect 1713 90871 1747 90905
rect 1747 90871 1756 90905
rect 1704 90862 1756 90871
rect 216910 90905 216962 90914
rect 216910 90871 216919 90905
rect 216919 90871 216953 90905
rect 216953 90871 216962 90905
rect 216910 90862 216962 90871
rect 1704 90569 1756 90578
rect 1704 90535 1713 90569
rect 1713 90535 1747 90569
rect 1747 90535 1756 90569
rect 1704 90526 1756 90535
rect 216910 90569 216962 90578
rect 216910 90535 216919 90569
rect 216919 90535 216953 90569
rect 216953 90535 216962 90569
rect 216910 90526 216962 90535
rect 1704 90233 1756 90242
rect 1704 90199 1713 90233
rect 1713 90199 1747 90233
rect 1747 90199 1756 90233
rect 1704 90190 1756 90199
rect 216910 90233 216962 90242
rect 216910 90199 216919 90233
rect 216919 90199 216953 90233
rect 216953 90199 216962 90233
rect 216910 90190 216962 90199
rect 1704 89897 1756 89906
rect 1704 89863 1713 89897
rect 1713 89863 1747 89897
rect 1747 89863 1756 89897
rect 1704 89854 1756 89863
rect 216910 89897 216962 89906
rect 216910 89863 216919 89897
rect 216919 89863 216953 89897
rect 216953 89863 216962 89897
rect 216910 89854 216962 89863
rect 1704 89561 1756 89570
rect 1704 89527 1713 89561
rect 1713 89527 1747 89561
rect 1747 89527 1756 89561
rect 1704 89518 1756 89527
rect 216910 89561 216962 89570
rect 216910 89527 216919 89561
rect 216919 89527 216953 89561
rect 216953 89527 216962 89561
rect 216910 89518 216962 89527
rect 1704 89225 1756 89234
rect 1704 89191 1713 89225
rect 1713 89191 1747 89225
rect 1747 89191 1756 89225
rect 1704 89182 1756 89191
rect 216910 89225 216962 89234
rect 216910 89191 216919 89225
rect 216919 89191 216953 89225
rect 216953 89191 216962 89225
rect 216910 89182 216962 89191
rect 1704 88889 1756 88898
rect 1704 88855 1713 88889
rect 1713 88855 1747 88889
rect 1747 88855 1756 88889
rect 1704 88846 1756 88855
rect 216910 88889 216962 88898
rect 216910 88855 216919 88889
rect 216919 88855 216953 88889
rect 216953 88855 216962 88889
rect 216910 88846 216962 88855
rect 1704 88553 1756 88562
rect 1704 88519 1713 88553
rect 1713 88519 1747 88553
rect 1747 88519 1756 88553
rect 1704 88510 1756 88519
rect 216910 88553 216962 88562
rect 216910 88519 216919 88553
rect 216919 88519 216953 88553
rect 216953 88519 216962 88553
rect 216910 88510 216962 88519
rect 1704 88217 1756 88226
rect 1704 88183 1713 88217
rect 1713 88183 1747 88217
rect 1747 88183 1756 88217
rect 1704 88174 1756 88183
rect 216910 88217 216962 88226
rect 216910 88183 216919 88217
rect 216919 88183 216953 88217
rect 216953 88183 216962 88217
rect 216910 88174 216962 88183
rect 1704 87881 1756 87890
rect 1704 87847 1713 87881
rect 1713 87847 1747 87881
rect 1747 87847 1756 87881
rect 1704 87838 1756 87847
rect 216910 87881 216962 87890
rect 216910 87847 216919 87881
rect 216919 87847 216953 87881
rect 216953 87847 216962 87881
rect 216910 87838 216962 87847
rect 1704 87545 1756 87554
rect 1704 87511 1713 87545
rect 1713 87511 1747 87545
rect 1747 87511 1756 87545
rect 1704 87502 1756 87511
rect 216910 87545 216962 87554
rect 216910 87511 216919 87545
rect 216919 87511 216953 87545
rect 216953 87511 216962 87545
rect 216910 87502 216962 87511
rect 1704 87209 1756 87218
rect 1704 87175 1713 87209
rect 1713 87175 1747 87209
rect 1747 87175 1756 87209
rect 1704 87166 1756 87175
rect 216910 87209 216962 87218
rect 216910 87175 216919 87209
rect 216919 87175 216953 87209
rect 216953 87175 216962 87209
rect 216910 87166 216962 87175
rect 1704 86873 1756 86882
rect 1704 86839 1713 86873
rect 1713 86839 1747 86873
rect 1747 86839 1756 86873
rect 1704 86830 1756 86839
rect 216910 86873 216962 86882
rect 216910 86839 216919 86873
rect 216919 86839 216953 86873
rect 216953 86839 216962 86873
rect 216910 86830 216962 86839
rect 1704 86537 1756 86546
rect 1704 86503 1713 86537
rect 1713 86503 1747 86537
rect 1747 86503 1756 86537
rect 1704 86494 1756 86503
rect 216910 86537 216962 86546
rect 216910 86503 216919 86537
rect 216919 86503 216953 86537
rect 216953 86503 216962 86537
rect 216910 86494 216962 86503
rect 1704 86201 1756 86210
rect 1704 86167 1713 86201
rect 1713 86167 1747 86201
rect 1747 86167 1756 86201
rect 1704 86158 1756 86167
rect 216910 86201 216962 86210
rect 216910 86167 216919 86201
rect 216919 86167 216953 86201
rect 216953 86167 216962 86201
rect 216910 86158 216962 86167
rect 1704 85865 1756 85874
rect 1704 85831 1713 85865
rect 1713 85831 1747 85865
rect 1747 85831 1756 85865
rect 1704 85822 1756 85831
rect 216910 85865 216962 85874
rect 216910 85831 216919 85865
rect 216919 85831 216953 85865
rect 216953 85831 216962 85865
rect 216910 85822 216962 85831
rect 1704 85529 1756 85538
rect 1704 85495 1713 85529
rect 1713 85495 1747 85529
rect 1747 85495 1756 85529
rect 1704 85486 1756 85495
rect 216910 85529 216962 85538
rect 216910 85495 216919 85529
rect 216919 85495 216953 85529
rect 216953 85495 216962 85529
rect 216910 85486 216962 85495
rect 1704 85193 1756 85202
rect 1704 85159 1713 85193
rect 1713 85159 1747 85193
rect 1747 85159 1756 85193
rect 1704 85150 1756 85159
rect 216910 85193 216962 85202
rect 216910 85159 216919 85193
rect 216919 85159 216953 85193
rect 216953 85159 216962 85193
rect 216910 85150 216962 85159
rect 1704 84857 1756 84866
rect 1704 84823 1713 84857
rect 1713 84823 1747 84857
rect 1747 84823 1756 84857
rect 1704 84814 1756 84823
rect 216910 84857 216962 84866
rect 216910 84823 216919 84857
rect 216919 84823 216953 84857
rect 216953 84823 216962 84857
rect 216910 84814 216962 84823
rect 1704 84521 1756 84530
rect 1704 84487 1713 84521
rect 1713 84487 1747 84521
rect 1747 84487 1756 84521
rect 1704 84478 1756 84487
rect 216910 84521 216962 84530
rect 216910 84487 216919 84521
rect 216919 84487 216953 84521
rect 216953 84487 216962 84521
rect 216910 84478 216962 84487
rect 1704 84185 1756 84194
rect 1704 84151 1713 84185
rect 1713 84151 1747 84185
rect 1747 84151 1756 84185
rect 1704 84142 1756 84151
rect 216910 84185 216962 84194
rect 216910 84151 216919 84185
rect 216919 84151 216953 84185
rect 216953 84151 216962 84185
rect 216910 84142 216962 84151
rect 1704 83849 1756 83858
rect 1704 83815 1713 83849
rect 1713 83815 1747 83849
rect 1747 83815 1756 83849
rect 1704 83806 1756 83815
rect 216910 83849 216962 83858
rect 216910 83815 216919 83849
rect 216919 83815 216953 83849
rect 216953 83815 216962 83849
rect 216910 83806 216962 83815
rect 1704 83513 1756 83522
rect 1704 83479 1713 83513
rect 1713 83479 1747 83513
rect 1747 83479 1756 83513
rect 1704 83470 1756 83479
rect 216910 83513 216962 83522
rect 216910 83479 216919 83513
rect 216919 83479 216953 83513
rect 216953 83479 216962 83513
rect 216910 83470 216962 83479
rect 1704 83177 1756 83186
rect 1704 83143 1713 83177
rect 1713 83143 1747 83177
rect 1747 83143 1756 83177
rect 1704 83134 1756 83143
rect 216910 83177 216962 83186
rect 216910 83143 216919 83177
rect 216919 83143 216953 83177
rect 216953 83143 216962 83177
rect 216910 83134 216962 83143
rect 1704 82841 1756 82850
rect 1704 82807 1713 82841
rect 1713 82807 1747 82841
rect 1747 82807 1756 82841
rect 1704 82798 1756 82807
rect 216910 82841 216962 82850
rect 216910 82807 216919 82841
rect 216919 82807 216953 82841
rect 216953 82807 216962 82841
rect 216910 82798 216962 82807
rect 1704 82505 1756 82514
rect 1704 82471 1713 82505
rect 1713 82471 1747 82505
rect 1747 82471 1756 82505
rect 1704 82462 1756 82471
rect 216910 82505 216962 82514
rect 216910 82471 216919 82505
rect 216919 82471 216953 82505
rect 216953 82471 216962 82505
rect 216910 82462 216962 82471
rect 1704 82169 1756 82178
rect 1704 82135 1713 82169
rect 1713 82135 1747 82169
rect 1747 82135 1756 82169
rect 1704 82126 1756 82135
rect 216910 82169 216962 82178
rect 216910 82135 216919 82169
rect 216919 82135 216953 82169
rect 216953 82135 216962 82169
rect 216910 82126 216962 82135
rect 1704 81833 1756 81842
rect 1704 81799 1713 81833
rect 1713 81799 1747 81833
rect 1747 81799 1756 81833
rect 1704 81790 1756 81799
rect 216910 81833 216962 81842
rect 216910 81799 216919 81833
rect 216919 81799 216953 81833
rect 216953 81799 216962 81833
rect 216910 81790 216962 81799
rect 1704 81497 1756 81506
rect 1704 81463 1713 81497
rect 1713 81463 1747 81497
rect 1747 81463 1756 81497
rect 1704 81454 1756 81463
rect 216910 81497 216962 81506
rect 216910 81463 216919 81497
rect 216919 81463 216953 81497
rect 216953 81463 216962 81497
rect 216910 81454 216962 81463
rect 1704 81161 1756 81170
rect 1704 81127 1713 81161
rect 1713 81127 1747 81161
rect 1747 81127 1756 81161
rect 1704 81118 1756 81127
rect 216910 81161 216962 81170
rect 216910 81127 216919 81161
rect 216919 81127 216953 81161
rect 216953 81127 216962 81161
rect 216910 81118 216962 81127
rect 1704 80825 1756 80834
rect 1704 80791 1713 80825
rect 1713 80791 1747 80825
rect 1747 80791 1756 80825
rect 1704 80782 1756 80791
rect 216910 80825 216962 80834
rect 216910 80791 216919 80825
rect 216919 80791 216953 80825
rect 216953 80791 216962 80825
rect 216910 80782 216962 80791
rect 1704 80489 1756 80498
rect 1704 80455 1713 80489
rect 1713 80455 1747 80489
rect 1747 80455 1756 80489
rect 1704 80446 1756 80455
rect 216910 80489 216962 80498
rect 216910 80455 216919 80489
rect 216919 80455 216953 80489
rect 216953 80455 216962 80489
rect 216910 80446 216962 80455
rect 1704 80153 1756 80162
rect 1704 80119 1713 80153
rect 1713 80119 1747 80153
rect 1747 80119 1756 80153
rect 1704 80110 1756 80119
rect 216910 80153 216962 80162
rect 216910 80119 216919 80153
rect 216919 80119 216953 80153
rect 216953 80119 216962 80153
rect 216910 80110 216962 80119
rect 1704 79817 1756 79826
rect 1704 79783 1713 79817
rect 1713 79783 1747 79817
rect 1747 79783 1756 79817
rect 1704 79774 1756 79783
rect 216910 79817 216962 79826
rect 216910 79783 216919 79817
rect 216919 79783 216953 79817
rect 216953 79783 216962 79817
rect 216910 79774 216962 79783
rect 1704 79481 1756 79490
rect 1704 79447 1713 79481
rect 1713 79447 1747 79481
rect 1747 79447 1756 79481
rect 1704 79438 1756 79447
rect 216910 79481 216962 79490
rect 216910 79447 216919 79481
rect 216919 79447 216953 79481
rect 216953 79447 216962 79481
rect 216910 79438 216962 79447
rect 1704 79145 1756 79154
rect 1704 79111 1713 79145
rect 1713 79111 1747 79145
rect 1747 79111 1756 79145
rect 1704 79102 1756 79111
rect 216910 79145 216962 79154
rect 216910 79111 216919 79145
rect 216919 79111 216953 79145
rect 216953 79111 216962 79145
rect 216910 79102 216962 79111
rect 1704 78809 1756 78818
rect 1704 78775 1713 78809
rect 1713 78775 1747 78809
rect 1747 78775 1756 78809
rect 1704 78766 1756 78775
rect 216910 78809 216962 78818
rect 216910 78775 216919 78809
rect 216919 78775 216953 78809
rect 216953 78775 216962 78809
rect 216910 78766 216962 78775
rect 1704 78473 1756 78482
rect 1704 78439 1713 78473
rect 1713 78439 1747 78473
rect 1747 78439 1756 78473
rect 1704 78430 1756 78439
rect 216910 78473 216962 78482
rect 216910 78439 216919 78473
rect 216919 78439 216953 78473
rect 216953 78439 216962 78473
rect 216910 78430 216962 78439
rect 1704 78137 1756 78146
rect 1704 78103 1713 78137
rect 1713 78103 1747 78137
rect 1747 78103 1756 78137
rect 1704 78094 1756 78103
rect 216910 78137 216962 78146
rect 216910 78103 216919 78137
rect 216919 78103 216953 78137
rect 216953 78103 216962 78137
rect 216910 78094 216962 78103
rect 1704 77801 1756 77810
rect 1704 77767 1713 77801
rect 1713 77767 1747 77801
rect 1747 77767 1756 77801
rect 1704 77758 1756 77767
rect 216910 77801 216962 77810
rect 216910 77767 216919 77801
rect 216919 77767 216953 77801
rect 216953 77767 216962 77801
rect 216910 77758 216962 77767
rect 1704 77465 1756 77474
rect 1704 77431 1713 77465
rect 1713 77431 1747 77465
rect 1747 77431 1756 77465
rect 1704 77422 1756 77431
rect 216910 77465 216962 77474
rect 216910 77431 216919 77465
rect 216919 77431 216953 77465
rect 216953 77431 216962 77465
rect 216910 77422 216962 77431
rect 1704 77129 1756 77138
rect 1704 77095 1713 77129
rect 1713 77095 1747 77129
rect 1747 77095 1756 77129
rect 1704 77086 1756 77095
rect 216910 77129 216962 77138
rect 216910 77095 216919 77129
rect 216919 77095 216953 77129
rect 216953 77095 216962 77129
rect 216910 77086 216962 77095
rect 1704 76793 1756 76802
rect 1704 76759 1713 76793
rect 1713 76759 1747 76793
rect 1747 76759 1756 76793
rect 1704 76750 1756 76759
rect 216910 76793 216962 76802
rect 216910 76759 216919 76793
rect 216919 76759 216953 76793
rect 216953 76759 216962 76793
rect 216910 76750 216962 76759
rect 1704 76457 1756 76466
rect 1704 76423 1713 76457
rect 1713 76423 1747 76457
rect 1747 76423 1756 76457
rect 1704 76414 1756 76423
rect 216910 76457 216962 76466
rect 216910 76423 216919 76457
rect 216919 76423 216953 76457
rect 216953 76423 216962 76457
rect 216910 76414 216962 76423
rect 1704 76121 1756 76130
rect 1704 76087 1713 76121
rect 1713 76087 1747 76121
rect 1747 76087 1756 76121
rect 1704 76078 1756 76087
rect 216910 76121 216962 76130
rect 216910 76087 216919 76121
rect 216919 76087 216953 76121
rect 216953 76087 216962 76121
rect 216910 76078 216962 76087
rect 1704 75785 1756 75794
rect 1704 75751 1713 75785
rect 1713 75751 1747 75785
rect 1747 75751 1756 75785
rect 1704 75742 1756 75751
rect 216910 75785 216962 75794
rect 216910 75751 216919 75785
rect 216919 75751 216953 75785
rect 216953 75751 216962 75785
rect 216910 75742 216962 75751
rect 1704 75449 1756 75458
rect 1704 75415 1713 75449
rect 1713 75415 1747 75449
rect 1747 75415 1756 75449
rect 1704 75406 1756 75415
rect 216910 75449 216962 75458
rect 216910 75415 216919 75449
rect 216919 75415 216953 75449
rect 216953 75415 216962 75449
rect 216910 75406 216962 75415
rect 1704 75113 1756 75122
rect 1704 75079 1713 75113
rect 1713 75079 1747 75113
rect 1747 75079 1756 75113
rect 1704 75070 1756 75079
rect 216910 75113 216962 75122
rect 216910 75079 216919 75113
rect 216919 75079 216953 75113
rect 216953 75079 216962 75113
rect 216910 75070 216962 75079
rect 1704 74777 1756 74786
rect 1704 74743 1713 74777
rect 1713 74743 1747 74777
rect 1747 74743 1756 74777
rect 1704 74734 1756 74743
rect 216910 74777 216962 74786
rect 216910 74743 216919 74777
rect 216919 74743 216953 74777
rect 216953 74743 216962 74777
rect 216910 74734 216962 74743
rect 1704 74441 1756 74450
rect 1704 74407 1713 74441
rect 1713 74407 1747 74441
rect 1747 74407 1756 74441
rect 1704 74398 1756 74407
rect 216910 74441 216962 74450
rect 216910 74407 216919 74441
rect 216919 74407 216953 74441
rect 216953 74407 216962 74441
rect 216910 74398 216962 74407
rect 1704 74105 1756 74114
rect 1704 74071 1713 74105
rect 1713 74071 1747 74105
rect 1747 74071 1756 74105
rect 1704 74062 1756 74071
rect 216910 74105 216962 74114
rect 216910 74071 216919 74105
rect 216919 74071 216953 74105
rect 216953 74071 216962 74105
rect 216910 74062 216962 74071
rect 1704 73769 1756 73778
rect 1704 73735 1713 73769
rect 1713 73735 1747 73769
rect 1747 73735 1756 73769
rect 1704 73726 1756 73735
rect 216910 73769 216962 73778
rect 216910 73735 216919 73769
rect 216919 73735 216953 73769
rect 216953 73735 216962 73769
rect 216910 73726 216962 73735
rect 1704 73433 1756 73442
rect 1704 73399 1713 73433
rect 1713 73399 1747 73433
rect 1747 73399 1756 73433
rect 1704 73390 1756 73399
rect 216910 73433 216962 73442
rect 216910 73399 216919 73433
rect 216919 73399 216953 73433
rect 216953 73399 216962 73433
rect 216910 73390 216962 73399
rect 1704 73097 1756 73106
rect 1704 73063 1713 73097
rect 1713 73063 1747 73097
rect 1747 73063 1756 73097
rect 1704 73054 1756 73063
rect 216910 73097 216962 73106
rect 216910 73063 216919 73097
rect 216919 73063 216953 73097
rect 216953 73063 216962 73097
rect 216910 73054 216962 73063
rect 1704 72761 1756 72770
rect 1704 72727 1713 72761
rect 1713 72727 1747 72761
rect 1747 72727 1756 72761
rect 1704 72718 1756 72727
rect 216910 72761 216962 72770
rect 216910 72727 216919 72761
rect 216919 72727 216953 72761
rect 216953 72727 216962 72761
rect 216910 72718 216962 72727
rect 1704 72425 1756 72434
rect 1704 72391 1713 72425
rect 1713 72391 1747 72425
rect 1747 72391 1756 72425
rect 1704 72382 1756 72391
rect 216910 72425 216962 72434
rect 216910 72391 216919 72425
rect 216919 72391 216953 72425
rect 216953 72391 216962 72425
rect 216910 72382 216962 72391
rect 1704 72089 1756 72098
rect 1704 72055 1713 72089
rect 1713 72055 1747 72089
rect 1747 72055 1756 72089
rect 1704 72046 1756 72055
rect 216910 72089 216962 72098
rect 216910 72055 216919 72089
rect 216919 72055 216953 72089
rect 216953 72055 216962 72089
rect 216910 72046 216962 72055
rect 1704 71753 1756 71762
rect 1704 71719 1713 71753
rect 1713 71719 1747 71753
rect 1747 71719 1756 71753
rect 1704 71710 1756 71719
rect 216910 71753 216962 71762
rect 216910 71719 216919 71753
rect 216919 71719 216953 71753
rect 216953 71719 216962 71753
rect 216910 71710 216962 71719
rect 1704 71417 1756 71426
rect 1704 71383 1713 71417
rect 1713 71383 1747 71417
rect 1747 71383 1756 71417
rect 1704 71374 1756 71383
rect 216910 71417 216962 71426
rect 216910 71383 216919 71417
rect 216919 71383 216953 71417
rect 216953 71383 216962 71417
rect 216910 71374 216962 71383
rect 1704 71081 1756 71090
rect 1704 71047 1713 71081
rect 1713 71047 1747 71081
rect 1747 71047 1756 71081
rect 1704 71038 1756 71047
rect 216910 71081 216962 71090
rect 216910 71047 216919 71081
rect 216919 71047 216953 71081
rect 216953 71047 216962 71081
rect 216910 71038 216962 71047
rect 1704 70745 1756 70754
rect 1704 70711 1713 70745
rect 1713 70711 1747 70745
rect 1747 70711 1756 70745
rect 1704 70702 1756 70711
rect 216910 70745 216962 70754
rect 216910 70711 216919 70745
rect 216919 70711 216953 70745
rect 216953 70711 216962 70745
rect 216910 70702 216962 70711
rect 1704 70409 1756 70418
rect 1704 70375 1713 70409
rect 1713 70375 1747 70409
rect 1747 70375 1756 70409
rect 1704 70366 1756 70375
rect 216910 70409 216962 70418
rect 216910 70375 216919 70409
rect 216919 70375 216953 70409
rect 216953 70375 216962 70409
rect 216910 70366 216962 70375
rect 1704 70073 1756 70082
rect 1704 70039 1713 70073
rect 1713 70039 1747 70073
rect 1747 70039 1756 70073
rect 1704 70030 1756 70039
rect 216910 70073 216962 70082
rect 216910 70039 216919 70073
rect 216919 70039 216953 70073
rect 216953 70039 216962 70073
rect 216910 70030 216962 70039
rect 1704 69737 1756 69746
rect 1704 69703 1713 69737
rect 1713 69703 1747 69737
rect 1747 69703 1756 69737
rect 1704 69694 1756 69703
rect 216910 69737 216962 69746
rect 216910 69703 216919 69737
rect 216919 69703 216953 69737
rect 216953 69703 216962 69737
rect 216910 69694 216962 69703
rect 1704 69401 1756 69410
rect 1704 69367 1713 69401
rect 1713 69367 1747 69401
rect 1747 69367 1756 69401
rect 1704 69358 1756 69367
rect 216910 69401 216962 69410
rect 216910 69367 216919 69401
rect 216919 69367 216953 69401
rect 216953 69367 216962 69401
rect 216910 69358 216962 69367
rect 1704 69065 1756 69074
rect 1704 69031 1713 69065
rect 1713 69031 1747 69065
rect 1747 69031 1756 69065
rect 1704 69022 1756 69031
rect 216910 69065 216962 69074
rect 216910 69031 216919 69065
rect 216919 69031 216953 69065
rect 216953 69031 216962 69065
rect 216910 69022 216962 69031
rect 1704 68729 1756 68738
rect 1704 68695 1713 68729
rect 1713 68695 1747 68729
rect 1747 68695 1756 68729
rect 1704 68686 1756 68695
rect 216910 68729 216962 68738
rect 216910 68695 216919 68729
rect 216919 68695 216953 68729
rect 216953 68695 216962 68729
rect 216910 68686 216962 68695
rect 1704 68393 1756 68402
rect 1704 68359 1713 68393
rect 1713 68359 1747 68393
rect 1747 68359 1756 68393
rect 1704 68350 1756 68359
rect 216910 68393 216962 68402
rect 216910 68359 216919 68393
rect 216919 68359 216953 68393
rect 216953 68359 216962 68393
rect 216910 68350 216962 68359
rect 1704 68057 1756 68066
rect 1704 68023 1713 68057
rect 1713 68023 1747 68057
rect 1747 68023 1756 68057
rect 1704 68014 1756 68023
rect 216910 68057 216962 68066
rect 216910 68023 216919 68057
rect 216919 68023 216953 68057
rect 216953 68023 216962 68057
rect 216910 68014 216962 68023
rect 1704 67721 1756 67730
rect 1704 67687 1713 67721
rect 1713 67687 1747 67721
rect 1747 67687 1756 67721
rect 1704 67678 1756 67687
rect 216910 67721 216962 67730
rect 216910 67687 216919 67721
rect 216919 67687 216953 67721
rect 216953 67687 216962 67721
rect 216910 67678 216962 67687
rect 1704 67385 1756 67394
rect 1704 67351 1713 67385
rect 1713 67351 1747 67385
rect 1747 67351 1756 67385
rect 1704 67342 1756 67351
rect 216910 67385 216962 67394
rect 216910 67351 216919 67385
rect 216919 67351 216953 67385
rect 216953 67351 216962 67385
rect 216910 67342 216962 67351
rect 1704 67049 1756 67058
rect 1704 67015 1713 67049
rect 1713 67015 1747 67049
rect 1747 67015 1756 67049
rect 1704 67006 1756 67015
rect 216910 67049 216962 67058
rect 216910 67015 216919 67049
rect 216919 67015 216953 67049
rect 216953 67015 216962 67049
rect 216910 67006 216962 67015
rect 1704 66713 1756 66722
rect 1704 66679 1713 66713
rect 1713 66679 1747 66713
rect 1747 66679 1756 66713
rect 1704 66670 1756 66679
rect 216910 66713 216962 66722
rect 216910 66679 216919 66713
rect 216919 66679 216953 66713
rect 216953 66679 216962 66713
rect 216910 66670 216962 66679
rect 1704 66377 1756 66386
rect 1704 66343 1713 66377
rect 1713 66343 1747 66377
rect 1747 66343 1756 66377
rect 1704 66334 1756 66343
rect 216910 66377 216962 66386
rect 216910 66343 216919 66377
rect 216919 66343 216953 66377
rect 216953 66343 216962 66377
rect 216910 66334 216962 66343
rect 1704 66041 1756 66050
rect 1704 66007 1713 66041
rect 1713 66007 1747 66041
rect 1747 66007 1756 66041
rect 1704 65998 1756 66007
rect 216910 66041 216962 66050
rect 216910 66007 216919 66041
rect 216919 66007 216953 66041
rect 216953 66007 216962 66041
rect 216910 65998 216962 66007
rect 1704 65705 1756 65714
rect 1704 65671 1713 65705
rect 1713 65671 1747 65705
rect 1747 65671 1756 65705
rect 1704 65662 1756 65671
rect 216910 65705 216962 65714
rect 216910 65671 216919 65705
rect 216919 65671 216953 65705
rect 216953 65671 216962 65705
rect 216910 65662 216962 65671
rect 1704 65369 1756 65378
rect 1704 65335 1713 65369
rect 1713 65335 1747 65369
rect 1747 65335 1756 65369
rect 1704 65326 1756 65335
rect 216910 65369 216962 65378
rect 216910 65335 216919 65369
rect 216919 65335 216953 65369
rect 216953 65335 216962 65369
rect 216910 65326 216962 65335
rect 1704 65033 1756 65042
rect 1704 64999 1713 65033
rect 1713 64999 1747 65033
rect 1747 64999 1756 65033
rect 1704 64990 1756 64999
rect 216910 65033 216962 65042
rect 216910 64999 216919 65033
rect 216919 64999 216953 65033
rect 216953 64999 216962 65033
rect 216910 64990 216962 64999
rect 1704 64697 1756 64706
rect 1704 64663 1713 64697
rect 1713 64663 1747 64697
rect 1747 64663 1756 64697
rect 1704 64654 1756 64663
rect 216910 64697 216962 64706
rect 216910 64663 216919 64697
rect 216919 64663 216953 64697
rect 216953 64663 216962 64697
rect 216910 64654 216962 64663
rect 1704 64361 1756 64370
rect 1704 64327 1713 64361
rect 1713 64327 1747 64361
rect 1747 64327 1756 64361
rect 1704 64318 1756 64327
rect 216910 64361 216962 64370
rect 216910 64327 216919 64361
rect 216919 64327 216953 64361
rect 216953 64327 216962 64361
rect 216910 64318 216962 64327
rect 1704 64025 1756 64034
rect 1704 63991 1713 64025
rect 1713 63991 1747 64025
rect 1747 63991 1756 64025
rect 1704 63982 1756 63991
rect 216910 64025 216962 64034
rect 216910 63991 216919 64025
rect 216919 63991 216953 64025
rect 216953 63991 216962 64025
rect 216910 63982 216962 63991
rect 1704 63689 1756 63698
rect 1704 63655 1713 63689
rect 1713 63655 1747 63689
rect 1747 63655 1756 63689
rect 1704 63646 1756 63655
rect 216910 63689 216962 63698
rect 216910 63655 216919 63689
rect 216919 63655 216953 63689
rect 216953 63655 216962 63689
rect 216910 63646 216962 63655
rect 1704 63353 1756 63362
rect 1704 63319 1713 63353
rect 1713 63319 1747 63353
rect 1747 63319 1756 63353
rect 1704 63310 1756 63319
rect 216910 63353 216962 63362
rect 216910 63319 216919 63353
rect 216919 63319 216953 63353
rect 216953 63319 216962 63353
rect 216910 63310 216962 63319
rect 1704 63017 1756 63026
rect 1704 62983 1713 63017
rect 1713 62983 1747 63017
rect 1747 62983 1756 63017
rect 1704 62974 1756 62983
rect 216910 63017 216962 63026
rect 216910 62983 216919 63017
rect 216919 62983 216953 63017
rect 216953 62983 216962 63017
rect 216910 62974 216962 62983
rect 1704 62681 1756 62690
rect 1704 62647 1713 62681
rect 1713 62647 1747 62681
rect 1747 62647 1756 62681
rect 1704 62638 1756 62647
rect 216910 62681 216962 62690
rect 216910 62647 216919 62681
rect 216919 62647 216953 62681
rect 216953 62647 216962 62681
rect 216910 62638 216962 62647
rect 1704 62345 1756 62354
rect 1704 62311 1713 62345
rect 1713 62311 1747 62345
rect 1747 62311 1756 62345
rect 1704 62302 1756 62311
rect 216910 62345 216962 62354
rect 216910 62311 216919 62345
rect 216919 62311 216953 62345
rect 216953 62311 216962 62345
rect 216910 62302 216962 62311
rect 1704 62009 1756 62018
rect 1704 61975 1713 62009
rect 1713 61975 1747 62009
rect 1747 61975 1756 62009
rect 1704 61966 1756 61975
rect 216910 62009 216962 62018
rect 216910 61975 216919 62009
rect 216919 61975 216953 62009
rect 216953 61975 216962 62009
rect 216910 61966 216962 61975
rect 1704 61673 1756 61682
rect 1704 61639 1713 61673
rect 1713 61639 1747 61673
rect 1747 61639 1756 61673
rect 1704 61630 1756 61639
rect 216910 61673 216962 61682
rect 216910 61639 216919 61673
rect 216919 61639 216953 61673
rect 216953 61639 216962 61673
rect 216910 61630 216962 61639
rect 1704 61337 1756 61346
rect 1704 61303 1713 61337
rect 1713 61303 1747 61337
rect 1747 61303 1756 61337
rect 1704 61294 1756 61303
rect 216910 61337 216962 61346
rect 216910 61303 216919 61337
rect 216919 61303 216953 61337
rect 216953 61303 216962 61337
rect 216910 61294 216962 61303
rect 1704 61001 1756 61010
rect 1704 60967 1713 61001
rect 1713 60967 1747 61001
rect 1747 60967 1756 61001
rect 1704 60958 1756 60967
rect 216910 61001 216962 61010
rect 216910 60967 216919 61001
rect 216919 60967 216953 61001
rect 216953 60967 216962 61001
rect 216910 60958 216962 60967
rect 1704 60665 1756 60674
rect 1704 60631 1713 60665
rect 1713 60631 1747 60665
rect 1747 60631 1756 60665
rect 1704 60622 1756 60631
rect 216910 60665 216962 60674
rect 216910 60631 216919 60665
rect 216919 60631 216953 60665
rect 216953 60631 216962 60665
rect 216910 60622 216962 60631
rect 1704 60329 1756 60338
rect 1704 60295 1713 60329
rect 1713 60295 1747 60329
rect 1747 60295 1756 60329
rect 1704 60286 1756 60295
rect 216910 60329 216962 60338
rect 216910 60295 216919 60329
rect 216919 60295 216953 60329
rect 216953 60295 216962 60329
rect 216910 60286 216962 60295
rect 1704 59993 1756 60002
rect 1704 59959 1713 59993
rect 1713 59959 1747 59993
rect 1747 59959 1756 59993
rect 1704 59950 1756 59959
rect 216910 59993 216962 60002
rect 216910 59959 216919 59993
rect 216919 59959 216953 59993
rect 216953 59959 216962 59993
rect 216910 59950 216962 59959
rect 1704 59657 1756 59666
rect 1704 59623 1713 59657
rect 1713 59623 1747 59657
rect 1747 59623 1756 59657
rect 1704 59614 1756 59623
rect 216910 59657 216962 59666
rect 216910 59623 216919 59657
rect 216919 59623 216953 59657
rect 216953 59623 216962 59657
rect 216910 59614 216962 59623
rect 1704 59321 1756 59330
rect 1704 59287 1713 59321
rect 1713 59287 1747 59321
rect 1747 59287 1756 59321
rect 1704 59278 1756 59287
rect 216910 59321 216962 59330
rect 216910 59287 216919 59321
rect 216919 59287 216953 59321
rect 216953 59287 216962 59321
rect 216910 59278 216962 59287
rect 1704 58985 1756 58994
rect 1704 58951 1713 58985
rect 1713 58951 1747 58985
rect 1747 58951 1756 58985
rect 1704 58942 1756 58951
rect 216910 58985 216962 58994
rect 216910 58951 216919 58985
rect 216919 58951 216953 58985
rect 216953 58951 216962 58985
rect 216910 58942 216962 58951
rect 1704 58649 1756 58658
rect 1704 58615 1713 58649
rect 1713 58615 1747 58649
rect 1747 58615 1756 58649
rect 1704 58606 1756 58615
rect 216910 58649 216962 58658
rect 216910 58615 216919 58649
rect 216919 58615 216953 58649
rect 216953 58615 216962 58649
rect 216910 58606 216962 58615
rect 1704 58313 1756 58322
rect 1704 58279 1713 58313
rect 1713 58279 1747 58313
rect 1747 58279 1756 58313
rect 1704 58270 1756 58279
rect 216910 58313 216962 58322
rect 216910 58279 216919 58313
rect 216919 58279 216953 58313
rect 216953 58279 216962 58313
rect 216910 58270 216962 58279
rect 1704 57977 1756 57986
rect 1704 57943 1713 57977
rect 1713 57943 1747 57977
rect 1747 57943 1756 57977
rect 1704 57934 1756 57943
rect 216910 57977 216962 57986
rect 216910 57943 216919 57977
rect 216919 57943 216953 57977
rect 216953 57943 216962 57977
rect 216910 57934 216962 57943
rect 1704 57641 1756 57650
rect 1704 57607 1713 57641
rect 1713 57607 1747 57641
rect 1747 57607 1756 57641
rect 1704 57598 1756 57607
rect 216910 57641 216962 57650
rect 216910 57607 216919 57641
rect 216919 57607 216953 57641
rect 216953 57607 216962 57641
rect 216910 57598 216962 57607
rect 1704 57305 1756 57314
rect 1704 57271 1713 57305
rect 1713 57271 1747 57305
rect 1747 57271 1756 57305
rect 1704 57262 1756 57271
rect 216910 57305 216962 57314
rect 216910 57271 216919 57305
rect 216919 57271 216953 57305
rect 216953 57271 216962 57305
rect 216910 57262 216962 57271
rect 1704 56969 1756 56978
rect 1704 56935 1713 56969
rect 1713 56935 1747 56969
rect 1747 56935 1756 56969
rect 1704 56926 1756 56935
rect 216910 56969 216962 56978
rect 216910 56935 216919 56969
rect 216919 56935 216953 56969
rect 216953 56935 216962 56969
rect 216910 56926 216962 56935
rect 1704 56633 1756 56642
rect 1704 56599 1713 56633
rect 1713 56599 1747 56633
rect 1747 56599 1756 56633
rect 1704 56590 1756 56599
rect 216910 56633 216962 56642
rect 216910 56599 216919 56633
rect 216919 56599 216953 56633
rect 216953 56599 216962 56633
rect 216910 56590 216962 56599
rect 1704 56297 1756 56306
rect 1704 56263 1713 56297
rect 1713 56263 1747 56297
rect 1747 56263 1756 56297
rect 1704 56254 1756 56263
rect 216910 56297 216962 56306
rect 216910 56263 216919 56297
rect 216919 56263 216953 56297
rect 216953 56263 216962 56297
rect 216910 56254 216962 56263
rect 1704 55961 1756 55970
rect 1704 55927 1713 55961
rect 1713 55927 1747 55961
rect 1747 55927 1756 55961
rect 1704 55918 1756 55927
rect 216910 55961 216962 55970
rect 216910 55927 216919 55961
rect 216919 55927 216953 55961
rect 216953 55927 216962 55961
rect 216910 55918 216962 55927
rect 1704 55625 1756 55634
rect 1704 55591 1713 55625
rect 1713 55591 1747 55625
rect 1747 55591 1756 55625
rect 1704 55582 1756 55591
rect 216910 55625 216962 55634
rect 216910 55591 216919 55625
rect 216919 55591 216953 55625
rect 216953 55591 216962 55625
rect 216910 55582 216962 55591
rect 1704 55289 1756 55298
rect 1704 55255 1713 55289
rect 1713 55255 1747 55289
rect 1747 55255 1756 55289
rect 1704 55246 1756 55255
rect 216910 55289 216962 55298
rect 216910 55255 216919 55289
rect 216919 55255 216953 55289
rect 216953 55255 216962 55289
rect 216910 55246 216962 55255
rect 1704 54953 1756 54962
rect 1704 54919 1713 54953
rect 1713 54919 1747 54953
rect 1747 54919 1756 54953
rect 1704 54910 1756 54919
rect 216910 54953 216962 54962
rect 216910 54919 216919 54953
rect 216919 54919 216953 54953
rect 216953 54919 216962 54953
rect 216910 54910 216962 54919
rect 1704 54617 1756 54626
rect 1704 54583 1713 54617
rect 1713 54583 1747 54617
rect 1747 54583 1756 54617
rect 1704 54574 1756 54583
rect 216910 54617 216962 54626
rect 216910 54583 216919 54617
rect 216919 54583 216953 54617
rect 216953 54583 216962 54617
rect 216910 54574 216962 54583
rect 1704 54281 1756 54290
rect 1704 54247 1713 54281
rect 1713 54247 1747 54281
rect 1747 54247 1756 54281
rect 1704 54238 1756 54247
rect 216910 54281 216962 54290
rect 216910 54247 216919 54281
rect 216919 54247 216953 54281
rect 216953 54247 216962 54281
rect 216910 54238 216962 54247
rect 1704 53945 1756 53954
rect 1704 53911 1713 53945
rect 1713 53911 1747 53945
rect 1747 53911 1756 53945
rect 1704 53902 1756 53911
rect 216910 53945 216962 53954
rect 216910 53911 216919 53945
rect 216919 53911 216953 53945
rect 216953 53911 216962 53945
rect 216910 53902 216962 53911
rect 1704 53609 1756 53618
rect 1704 53575 1713 53609
rect 1713 53575 1747 53609
rect 1747 53575 1756 53609
rect 1704 53566 1756 53575
rect 216910 53609 216962 53618
rect 216910 53575 216919 53609
rect 216919 53575 216953 53609
rect 216953 53575 216962 53609
rect 216910 53566 216962 53575
rect 1704 53273 1756 53282
rect 1704 53239 1713 53273
rect 1713 53239 1747 53273
rect 1747 53239 1756 53273
rect 1704 53230 1756 53239
rect 216910 53273 216962 53282
rect 216910 53239 216919 53273
rect 216919 53239 216953 53273
rect 216953 53239 216962 53273
rect 216910 53230 216962 53239
rect 1704 52937 1756 52946
rect 1704 52903 1713 52937
rect 1713 52903 1747 52937
rect 1747 52903 1756 52937
rect 1704 52894 1756 52903
rect 216910 52937 216962 52946
rect 216910 52903 216919 52937
rect 216919 52903 216953 52937
rect 216953 52903 216962 52937
rect 216910 52894 216962 52903
rect 1704 52601 1756 52610
rect 1704 52567 1713 52601
rect 1713 52567 1747 52601
rect 1747 52567 1756 52601
rect 1704 52558 1756 52567
rect 216910 52601 216962 52610
rect 216910 52567 216919 52601
rect 216919 52567 216953 52601
rect 216953 52567 216962 52601
rect 216910 52558 216962 52567
rect 1704 52265 1756 52274
rect 1704 52231 1713 52265
rect 1713 52231 1747 52265
rect 1747 52231 1756 52265
rect 1704 52222 1756 52231
rect 216910 52265 216962 52274
rect 216910 52231 216919 52265
rect 216919 52231 216953 52265
rect 216953 52231 216962 52265
rect 216910 52222 216962 52231
rect 1704 51929 1756 51938
rect 1704 51895 1713 51929
rect 1713 51895 1747 51929
rect 1747 51895 1756 51929
rect 1704 51886 1756 51895
rect 216910 51929 216962 51938
rect 216910 51895 216919 51929
rect 216919 51895 216953 51929
rect 216953 51895 216962 51929
rect 216910 51886 216962 51895
rect 1704 51593 1756 51602
rect 1704 51559 1713 51593
rect 1713 51559 1747 51593
rect 1747 51559 1756 51593
rect 1704 51550 1756 51559
rect 216910 51593 216962 51602
rect 216910 51559 216919 51593
rect 216919 51559 216953 51593
rect 216953 51559 216962 51593
rect 216910 51550 216962 51559
rect 1704 51257 1756 51266
rect 1704 51223 1713 51257
rect 1713 51223 1747 51257
rect 1747 51223 1756 51257
rect 1704 51214 1756 51223
rect 216910 51257 216962 51266
rect 216910 51223 216919 51257
rect 216919 51223 216953 51257
rect 216953 51223 216962 51257
rect 216910 51214 216962 51223
rect 1704 50921 1756 50930
rect 1704 50887 1713 50921
rect 1713 50887 1747 50921
rect 1747 50887 1756 50921
rect 1704 50878 1756 50887
rect 216910 50921 216962 50930
rect 216910 50887 216919 50921
rect 216919 50887 216953 50921
rect 216953 50887 216962 50921
rect 216910 50878 216962 50887
rect 1704 50585 1756 50594
rect 1704 50551 1713 50585
rect 1713 50551 1747 50585
rect 1747 50551 1756 50585
rect 1704 50542 1756 50551
rect 216910 50585 216962 50594
rect 216910 50551 216919 50585
rect 216919 50551 216953 50585
rect 216953 50551 216962 50585
rect 216910 50542 216962 50551
rect 1704 50249 1756 50258
rect 1704 50215 1713 50249
rect 1713 50215 1747 50249
rect 1747 50215 1756 50249
rect 1704 50206 1756 50215
rect 216910 50249 216962 50258
rect 216910 50215 216919 50249
rect 216919 50215 216953 50249
rect 216953 50215 216962 50249
rect 216910 50206 216962 50215
rect 1704 49913 1756 49922
rect 1704 49879 1713 49913
rect 1713 49879 1747 49913
rect 1747 49879 1756 49913
rect 1704 49870 1756 49879
rect 216910 49913 216962 49922
rect 216910 49879 216919 49913
rect 216919 49879 216953 49913
rect 216953 49879 216962 49913
rect 216910 49870 216962 49879
rect 1704 49577 1756 49586
rect 1704 49543 1713 49577
rect 1713 49543 1747 49577
rect 1747 49543 1756 49577
rect 1704 49534 1756 49543
rect 216910 49577 216962 49586
rect 216910 49543 216919 49577
rect 216919 49543 216953 49577
rect 216953 49543 216962 49577
rect 216910 49534 216962 49543
rect 1704 49241 1756 49250
rect 1704 49207 1713 49241
rect 1713 49207 1747 49241
rect 1747 49207 1756 49241
rect 1704 49198 1756 49207
rect 216910 49241 216962 49250
rect 216910 49207 216919 49241
rect 216919 49207 216953 49241
rect 216953 49207 216962 49241
rect 216910 49198 216962 49207
rect 1704 48905 1756 48914
rect 1704 48871 1713 48905
rect 1713 48871 1747 48905
rect 1747 48871 1756 48905
rect 1704 48862 1756 48871
rect 216910 48905 216962 48914
rect 216910 48871 216919 48905
rect 216919 48871 216953 48905
rect 216953 48871 216962 48905
rect 216910 48862 216962 48871
rect 1704 48569 1756 48578
rect 1704 48535 1713 48569
rect 1713 48535 1747 48569
rect 1747 48535 1756 48569
rect 1704 48526 1756 48535
rect 216910 48569 216962 48578
rect 216910 48535 216919 48569
rect 216919 48535 216953 48569
rect 216953 48535 216962 48569
rect 216910 48526 216962 48535
rect 1704 48233 1756 48242
rect 1704 48199 1713 48233
rect 1713 48199 1747 48233
rect 1747 48199 1756 48233
rect 1704 48190 1756 48199
rect 216910 48233 216962 48242
rect 216910 48199 216919 48233
rect 216919 48199 216953 48233
rect 216953 48199 216962 48233
rect 216910 48190 216962 48199
rect 1704 47897 1756 47906
rect 1704 47863 1713 47897
rect 1713 47863 1747 47897
rect 1747 47863 1756 47897
rect 1704 47854 1756 47863
rect 216910 47897 216962 47906
rect 216910 47863 216919 47897
rect 216919 47863 216953 47897
rect 216953 47863 216962 47897
rect 216910 47854 216962 47863
rect 1704 47561 1756 47570
rect 1704 47527 1713 47561
rect 1713 47527 1747 47561
rect 1747 47527 1756 47561
rect 1704 47518 1756 47527
rect 216910 47561 216962 47570
rect 216910 47527 216919 47561
rect 216919 47527 216953 47561
rect 216953 47527 216962 47561
rect 216910 47518 216962 47527
rect 1704 47225 1756 47234
rect 1704 47191 1713 47225
rect 1713 47191 1747 47225
rect 1747 47191 1756 47225
rect 1704 47182 1756 47191
rect 216910 47225 216962 47234
rect 216910 47191 216919 47225
rect 216919 47191 216953 47225
rect 216953 47191 216962 47225
rect 216910 47182 216962 47191
rect 1704 46889 1756 46898
rect 1704 46855 1713 46889
rect 1713 46855 1747 46889
rect 1747 46855 1756 46889
rect 1704 46846 1756 46855
rect 216910 46889 216962 46898
rect 216910 46855 216919 46889
rect 216919 46855 216953 46889
rect 216953 46855 216962 46889
rect 216910 46846 216962 46855
rect 1704 46553 1756 46562
rect 1704 46519 1713 46553
rect 1713 46519 1747 46553
rect 1747 46519 1756 46553
rect 1704 46510 1756 46519
rect 216910 46553 216962 46562
rect 216910 46519 216919 46553
rect 216919 46519 216953 46553
rect 216953 46519 216962 46553
rect 216910 46510 216962 46519
rect 1704 46217 1756 46226
rect 1704 46183 1713 46217
rect 1713 46183 1747 46217
rect 1747 46183 1756 46217
rect 1704 46174 1756 46183
rect 216910 46217 216962 46226
rect 216910 46183 216919 46217
rect 216919 46183 216953 46217
rect 216953 46183 216962 46217
rect 216910 46174 216962 46183
rect 1704 45881 1756 45890
rect 1704 45847 1713 45881
rect 1713 45847 1747 45881
rect 1747 45847 1756 45881
rect 1704 45838 1756 45847
rect 216910 45881 216962 45890
rect 216910 45847 216919 45881
rect 216919 45847 216953 45881
rect 216953 45847 216962 45881
rect 216910 45838 216962 45847
rect 1704 45545 1756 45554
rect 1704 45511 1713 45545
rect 1713 45511 1747 45545
rect 1747 45511 1756 45545
rect 1704 45502 1756 45511
rect 216910 45545 216962 45554
rect 216910 45511 216919 45545
rect 216919 45511 216953 45545
rect 216953 45511 216962 45545
rect 216910 45502 216962 45511
rect 1704 45209 1756 45218
rect 1704 45175 1713 45209
rect 1713 45175 1747 45209
rect 1747 45175 1756 45209
rect 1704 45166 1756 45175
rect 216910 45209 216962 45218
rect 216910 45175 216919 45209
rect 216919 45175 216953 45209
rect 216953 45175 216962 45209
rect 216910 45166 216962 45175
rect 15973 44968 16025 45020
rect 1704 44873 1756 44882
rect 1704 44839 1713 44873
rect 1713 44839 1747 44873
rect 1747 44839 1756 44873
rect 1704 44830 1756 44839
rect 1704 44537 1756 44546
rect 1704 44503 1713 44537
rect 1713 44503 1747 44537
rect 1747 44503 1756 44537
rect 1704 44494 1756 44503
rect 1704 44201 1756 44210
rect 1704 44167 1713 44201
rect 1713 44167 1747 44201
rect 1747 44167 1756 44201
rect 1704 44158 1756 44167
rect 1704 43865 1756 43874
rect 1704 43831 1713 43865
rect 1713 43831 1747 43865
rect 1747 43831 1756 43865
rect 1704 43822 1756 43831
rect 1704 43529 1756 43538
rect 1704 43495 1713 43529
rect 1713 43495 1747 43529
rect 1747 43495 1756 43529
rect 1704 43486 1756 43495
rect 15893 43410 15945 43462
rect 1704 43193 1756 43202
rect 1704 43159 1713 43193
rect 1713 43159 1747 43193
rect 1747 43159 1756 43193
rect 1704 43150 1756 43159
rect 1704 42857 1756 42866
rect 1704 42823 1713 42857
rect 1713 42823 1747 42857
rect 1747 42823 1756 42857
rect 1704 42814 1756 42823
rect 1704 42521 1756 42530
rect 1704 42487 1713 42521
rect 1713 42487 1747 42521
rect 1747 42487 1756 42521
rect 1704 42478 1756 42487
rect 1704 42185 1756 42194
rect 1704 42151 1713 42185
rect 1713 42151 1747 42185
rect 1747 42151 1756 42185
rect 1704 42142 1756 42151
rect 15813 42140 15865 42192
rect 1704 41849 1756 41858
rect 1704 41815 1713 41849
rect 1713 41815 1747 41849
rect 1747 41815 1756 41849
rect 1704 41806 1756 41815
rect 1704 41513 1756 41522
rect 1704 41479 1713 41513
rect 1713 41479 1747 41513
rect 1747 41479 1756 41513
rect 1704 41470 1756 41479
rect 1704 41177 1756 41186
rect 1704 41143 1713 41177
rect 1713 41143 1747 41177
rect 1747 41143 1756 41177
rect 1704 41134 1756 41143
rect 1704 40841 1756 40850
rect 1704 40807 1713 40841
rect 1713 40807 1747 40841
rect 1747 40807 1756 40841
rect 1704 40798 1756 40807
rect 15733 40582 15785 40634
rect 1704 40505 1756 40514
rect 1704 40471 1713 40505
rect 1713 40471 1747 40505
rect 1747 40471 1756 40505
rect 1704 40462 1756 40471
rect 1704 40169 1756 40178
rect 1704 40135 1713 40169
rect 1713 40135 1747 40169
rect 1747 40135 1756 40169
rect 1704 40126 1756 40135
rect 1704 39833 1756 39842
rect 1704 39799 1713 39833
rect 1713 39799 1747 39833
rect 1747 39799 1756 39833
rect 1704 39790 1756 39799
rect 1704 39497 1756 39506
rect 1704 39463 1713 39497
rect 1713 39463 1747 39497
rect 1747 39463 1756 39497
rect 1704 39454 1756 39463
rect 15653 39312 15705 39364
rect 1704 39161 1756 39170
rect 1704 39127 1713 39161
rect 1713 39127 1747 39161
rect 1747 39127 1756 39161
rect 1704 39118 1756 39127
rect 1704 38825 1756 38834
rect 1704 38791 1713 38825
rect 1713 38791 1747 38825
rect 1747 38791 1756 38825
rect 1704 38782 1756 38791
rect 1704 38489 1756 38498
rect 1704 38455 1713 38489
rect 1713 38455 1747 38489
rect 1747 38455 1756 38489
rect 1704 38446 1756 38455
rect 1704 38153 1756 38162
rect 1704 38119 1713 38153
rect 1713 38119 1747 38153
rect 1747 38119 1756 38153
rect 1704 38110 1756 38119
rect 1704 37817 1756 37826
rect 1704 37783 1713 37817
rect 1713 37783 1747 37817
rect 1747 37783 1756 37817
rect 1704 37774 1756 37783
rect 15573 37754 15625 37806
rect 1704 37481 1756 37490
rect 1704 37447 1713 37481
rect 1713 37447 1747 37481
rect 1747 37447 1756 37481
rect 1704 37438 1756 37447
rect 1704 37145 1756 37154
rect 1704 37111 1713 37145
rect 1713 37111 1747 37145
rect 1747 37111 1756 37145
rect 1704 37102 1756 37111
rect 1704 36809 1756 36818
rect 1704 36775 1713 36809
rect 1713 36775 1747 36809
rect 1747 36775 1756 36809
rect 1704 36766 1756 36775
rect 15493 36484 15545 36536
rect 1704 36473 1756 36482
rect 1704 36439 1713 36473
rect 1713 36439 1747 36473
rect 1747 36439 1756 36473
rect 1704 36430 1756 36439
rect 1704 36137 1756 36146
rect 1704 36103 1713 36137
rect 1713 36103 1747 36137
rect 1747 36103 1756 36137
rect 1704 36094 1756 36103
rect 1704 35801 1756 35810
rect 1704 35767 1713 35801
rect 1713 35767 1747 35801
rect 1747 35767 1756 35801
rect 1704 35758 1756 35767
rect 1704 35465 1756 35474
rect 1704 35431 1713 35465
rect 1713 35431 1747 35465
rect 1747 35431 1756 35465
rect 1704 35422 1756 35431
rect 1704 35129 1756 35138
rect 1704 35095 1713 35129
rect 1713 35095 1747 35129
rect 1747 35095 1756 35129
rect 1704 35086 1756 35095
rect 15413 34926 15465 34978
rect 1704 34793 1756 34802
rect 1704 34759 1713 34793
rect 1713 34759 1747 34793
rect 1747 34759 1756 34793
rect 1704 34750 1756 34759
rect 1704 34457 1756 34466
rect 1704 34423 1713 34457
rect 1713 34423 1747 34457
rect 1747 34423 1756 34457
rect 1704 34414 1756 34423
rect 1704 34121 1756 34130
rect 1704 34087 1713 34121
rect 1713 34087 1747 34121
rect 1747 34087 1756 34121
rect 1704 34078 1756 34087
rect 1704 33785 1756 33794
rect 1704 33751 1713 33785
rect 1713 33751 1747 33785
rect 1747 33751 1756 33785
rect 1704 33742 1756 33751
rect 1704 33449 1756 33458
rect 1704 33415 1713 33449
rect 1713 33415 1747 33449
rect 1747 33415 1756 33449
rect 1704 33406 1756 33415
rect 1704 33113 1756 33122
rect 1704 33079 1713 33113
rect 1713 33079 1747 33113
rect 1747 33079 1756 33113
rect 1704 33070 1756 33079
rect 1704 32777 1756 32786
rect 1704 32743 1713 32777
rect 1713 32743 1747 32777
rect 1747 32743 1756 32777
rect 1704 32734 1756 32743
rect 1704 32441 1756 32450
rect 1704 32407 1713 32441
rect 1713 32407 1747 32441
rect 1747 32407 1756 32441
rect 1704 32398 1756 32407
rect 1704 32105 1756 32114
rect 1704 32071 1713 32105
rect 1713 32071 1747 32105
rect 1747 32071 1756 32105
rect 1704 32062 1756 32071
rect 1704 31769 1756 31778
rect 1704 31735 1713 31769
rect 1713 31735 1747 31769
rect 1747 31735 1756 31769
rect 1704 31726 1756 31735
rect 1704 31433 1756 31442
rect 1704 31399 1713 31433
rect 1713 31399 1747 31433
rect 1747 31399 1756 31433
rect 1704 31390 1756 31399
rect 1704 31097 1756 31106
rect 1704 31063 1713 31097
rect 1713 31063 1747 31097
rect 1747 31063 1756 31097
rect 1704 31054 1756 31063
rect 1704 30761 1756 30770
rect 1704 30727 1713 30761
rect 1713 30727 1747 30761
rect 1747 30727 1756 30761
rect 1704 30718 1756 30727
rect 1704 30425 1756 30434
rect 1704 30391 1713 30425
rect 1713 30391 1747 30425
rect 1747 30391 1756 30425
rect 1704 30382 1756 30391
rect 1704 30089 1756 30098
rect 1704 30055 1713 30089
rect 1713 30055 1747 30089
rect 1747 30055 1756 30089
rect 1704 30046 1756 30055
rect 1704 29753 1756 29762
rect 1704 29719 1713 29753
rect 1713 29719 1747 29753
rect 1747 29719 1756 29753
rect 1704 29710 1756 29719
rect 216910 44873 216962 44882
rect 216910 44839 216919 44873
rect 216919 44839 216953 44873
rect 216953 44839 216962 44873
rect 216910 44830 216962 44839
rect 216910 44537 216962 44546
rect 216910 44503 216919 44537
rect 216919 44503 216953 44537
rect 216953 44503 216962 44537
rect 216910 44494 216962 44503
rect 216910 44201 216962 44210
rect 216910 44167 216919 44201
rect 216919 44167 216953 44201
rect 216953 44167 216962 44201
rect 216910 44158 216962 44167
rect 216910 43865 216962 43874
rect 216910 43831 216919 43865
rect 216919 43831 216953 43865
rect 216953 43831 216962 43865
rect 216910 43822 216962 43831
rect 216910 43529 216962 43538
rect 216910 43495 216919 43529
rect 216919 43495 216953 43529
rect 216953 43495 216962 43529
rect 216910 43486 216962 43495
rect 216910 43193 216962 43202
rect 216910 43159 216919 43193
rect 216919 43159 216953 43193
rect 216953 43159 216962 43193
rect 216910 43150 216962 43159
rect 216910 42857 216962 42866
rect 216910 42823 216919 42857
rect 216919 42823 216953 42857
rect 216953 42823 216962 42857
rect 216910 42814 216962 42823
rect 216910 42521 216962 42530
rect 216910 42487 216919 42521
rect 216919 42487 216953 42521
rect 216953 42487 216962 42521
rect 216910 42478 216962 42487
rect 216910 42185 216962 42194
rect 216910 42151 216919 42185
rect 216919 42151 216953 42185
rect 216953 42151 216962 42185
rect 216910 42142 216962 42151
rect 216910 41849 216962 41858
rect 216910 41815 216919 41849
rect 216919 41815 216953 41849
rect 216953 41815 216962 41849
rect 216910 41806 216962 41815
rect 216910 41513 216962 41522
rect 216910 41479 216919 41513
rect 216919 41479 216953 41513
rect 216953 41479 216962 41513
rect 216910 41470 216962 41479
rect 216910 41177 216962 41186
rect 216910 41143 216919 41177
rect 216919 41143 216953 41177
rect 216953 41143 216962 41177
rect 216910 41134 216962 41143
rect 216910 40841 216962 40850
rect 216910 40807 216919 40841
rect 216919 40807 216953 40841
rect 216953 40807 216962 40841
rect 216910 40798 216962 40807
rect 216910 40505 216962 40514
rect 216910 40471 216919 40505
rect 216919 40471 216953 40505
rect 216953 40471 216962 40505
rect 216910 40462 216962 40471
rect 216910 40169 216962 40178
rect 216910 40135 216919 40169
rect 216919 40135 216953 40169
rect 216953 40135 216962 40169
rect 216910 40126 216962 40135
rect 216910 39833 216962 39842
rect 216910 39799 216919 39833
rect 216919 39799 216953 39833
rect 216953 39799 216962 39833
rect 216910 39790 216962 39799
rect 216910 39497 216962 39506
rect 216910 39463 216919 39497
rect 216919 39463 216953 39497
rect 216953 39463 216962 39497
rect 216910 39454 216962 39463
rect 216910 39161 216962 39170
rect 216910 39127 216919 39161
rect 216919 39127 216953 39161
rect 216953 39127 216962 39161
rect 216910 39118 216962 39127
rect 216910 38825 216962 38834
rect 216910 38791 216919 38825
rect 216919 38791 216953 38825
rect 216953 38791 216962 38825
rect 216910 38782 216962 38791
rect 216910 38489 216962 38498
rect 216910 38455 216919 38489
rect 216919 38455 216953 38489
rect 216953 38455 216962 38489
rect 216910 38446 216962 38455
rect 216910 38153 216962 38162
rect 216910 38119 216919 38153
rect 216919 38119 216953 38153
rect 216953 38119 216962 38153
rect 216910 38110 216962 38119
rect 216910 37817 216962 37826
rect 216910 37783 216919 37817
rect 216919 37783 216953 37817
rect 216953 37783 216962 37817
rect 216910 37774 216962 37783
rect 216910 37481 216962 37490
rect 216910 37447 216919 37481
rect 216919 37447 216953 37481
rect 216953 37447 216962 37481
rect 216910 37438 216962 37447
rect 216910 37145 216962 37154
rect 216910 37111 216919 37145
rect 216919 37111 216953 37145
rect 216953 37111 216962 37145
rect 216910 37102 216962 37111
rect 216910 36809 216962 36818
rect 216910 36775 216919 36809
rect 216919 36775 216953 36809
rect 216953 36775 216962 36809
rect 216910 36766 216962 36775
rect 216910 36473 216962 36482
rect 216910 36439 216919 36473
rect 216919 36439 216953 36473
rect 216953 36439 216962 36473
rect 216910 36430 216962 36439
rect 216910 36137 216962 36146
rect 216910 36103 216919 36137
rect 216919 36103 216953 36137
rect 216953 36103 216962 36137
rect 216910 36094 216962 36103
rect 216910 35801 216962 35810
rect 216910 35767 216919 35801
rect 216919 35767 216953 35801
rect 216953 35767 216962 35801
rect 216910 35758 216962 35767
rect 216910 35465 216962 35474
rect 216910 35431 216919 35465
rect 216919 35431 216953 35465
rect 216953 35431 216962 35465
rect 216910 35422 216962 35431
rect 216910 35129 216962 35138
rect 216910 35095 216919 35129
rect 216919 35095 216953 35129
rect 216953 35095 216962 35129
rect 216910 35086 216962 35095
rect 216910 34793 216962 34802
rect 216910 34759 216919 34793
rect 216919 34759 216953 34793
rect 216953 34759 216962 34793
rect 216910 34750 216962 34759
rect 216910 34457 216962 34466
rect 216910 34423 216919 34457
rect 216919 34423 216953 34457
rect 216953 34423 216962 34457
rect 216910 34414 216962 34423
rect 216910 34121 216962 34130
rect 216910 34087 216919 34121
rect 216919 34087 216953 34121
rect 216953 34087 216962 34121
rect 216910 34078 216962 34087
rect 216910 33785 216962 33794
rect 216910 33751 216919 33785
rect 216919 33751 216953 33785
rect 216953 33751 216962 33785
rect 216910 33742 216962 33751
rect 216910 33449 216962 33458
rect 216910 33415 216919 33449
rect 216919 33415 216953 33449
rect 216953 33415 216962 33449
rect 216910 33406 216962 33415
rect 216910 33113 216962 33122
rect 216910 33079 216919 33113
rect 216919 33079 216953 33113
rect 216953 33079 216962 33113
rect 216910 33070 216962 33079
rect 216910 32777 216962 32786
rect 216910 32743 216919 32777
rect 216919 32743 216953 32777
rect 216953 32743 216962 32777
rect 216910 32734 216962 32743
rect 216910 32441 216962 32450
rect 216910 32407 216919 32441
rect 216919 32407 216953 32441
rect 216953 32407 216962 32441
rect 216910 32398 216962 32407
rect 216910 32105 216962 32114
rect 216910 32071 216919 32105
rect 216919 32071 216953 32105
rect 216953 32071 216962 32105
rect 216910 32062 216962 32071
rect 216910 31769 216962 31778
rect 216910 31735 216919 31769
rect 216919 31735 216953 31769
rect 216953 31735 216962 31769
rect 216910 31726 216962 31735
rect 216910 31433 216962 31442
rect 216910 31399 216919 31433
rect 216919 31399 216953 31433
rect 216953 31399 216962 31433
rect 216910 31390 216962 31399
rect 216910 31097 216962 31106
rect 216910 31063 216919 31097
rect 216919 31063 216953 31097
rect 216953 31063 216962 31097
rect 216910 31054 216962 31063
rect 216910 30761 216962 30770
rect 216910 30727 216919 30761
rect 216919 30727 216953 30761
rect 216953 30727 216962 30761
rect 216910 30718 216962 30727
rect 216910 30425 216962 30434
rect 216910 30391 216919 30425
rect 216919 30391 216953 30425
rect 216953 30391 216962 30425
rect 216910 30382 216962 30391
rect 216910 30089 216962 30098
rect 216910 30055 216919 30089
rect 216919 30055 216953 30089
rect 216953 30055 216962 30089
rect 216910 30046 216962 30055
rect 216910 29753 216962 29762
rect 216910 29719 216919 29753
rect 216919 29719 216953 29753
rect 216953 29719 216962 29753
rect 216910 29710 216962 29719
rect 1704 29417 1756 29426
rect 1704 29383 1713 29417
rect 1713 29383 1747 29417
rect 1747 29383 1756 29417
rect 1704 29374 1756 29383
rect 1704 29081 1756 29090
rect 1704 29047 1713 29081
rect 1713 29047 1747 29081
rect 1747 29047 1756 29081
rect 1704 29038 1756 29047
rect 1704 28745 1756 28754
rect 1704 28711 1713 28745
rect 1713 28711 1747 28745
rect 1747 28711 1756 28745
rect 1704 28702 1756 28711
rect 1704 28409 1756 28418
rect 1704 28375 1713 28409
rect 1713 28375 1747 28409
rect 1747 28375 1756 28409
rect 1704 28366 1756 28375
rect 1704 28073 1756 28082
rect 1704 28039 1713 28073
rect 1713 28039 1747 28073
rect 1747 28039 1756 28073
rect 1704 28030 1756 28039
rect 1704 27737 1756 27746
rect 1704 27703 1713 27737
rect 1713 27703 1747 27737
rect 1747 27703 1756 27737
rect 1704 27694 1756 27703
rect 1704 27401 1756 27410
rect 1704 27367 1713 27401
rect 1713 27367 1747 27401
rect 1747 27367 1756 27401
rect 1704 27358 1756 27367
rect 1704 27065 1756 27074
rect 1704 27031 1713 27065
rect 1713 27031 1747 27065
rect 1747 27031 1756 27065
rect 1704 27022 1756 27031
rect 1704 26729 1756 26738
rect 1704 26695 1713 26729
rect 1713 26695 1747 26729
rect 1747 26695 1756 26729
rect 1704 26686 1756 26695
rect 1704 26393 1756 26402
rect 1704 26359 1713 26393
rect 1713 26359 1747 26393
rect 1747 26359 1756 26393
rect 1704 26350 1756 26359
rect 1704 26057 1756 26066
rect 1704 26023 1713 26057
rect 1713 26023 1747 26057
rect 1747 26023 1756 26057
rect 1704 26014 1756 26023
rect 1704 25721 1756 25730
rect 1704 25687 1713 25721
rect 1713 25687 1747 25721
rect 1747 25687 1756 25721
rect 1704 25678 1756 25687
rect 1704 25385 1756 25394
rect 1704 25351 1713 25385
rect 1713 25351 1747 25385
rect 1747 25351 1756 25385
rect 1704 25342 1756 25351
rect 1704 25049 1756 25058
rect 1704 25015 1713 25049
rect 1713 25015 1747 25049
rect 1747 25015 1756 25049
rect 1704 25006 1756 25015
rect 1704 24713 1756 24722
rect 1704 24679 1713 24713
rect 1713 24679 1747 24713
rect 1747 24679 1756 24713
rect 1704 24670 1756 24679
rect 1704 24377 1756 24386
rect 1704 24343 1713 24377
rect 1713 24343 1747 24377
rect 1747 24343 1756 24377
rect 1704 24334 1756 24343
rect 1704 24041 1756 24050
rect 1704 24007 1713 24041
rect 1713 24007 1747 24041
rect 1747 24007 1756 24041
rect 1704 23998 1756 24007
rect 1704 23705 1756 23714
rect 1704 23671 1713 23705
rect 1713 23671 1747 23705
rect 1747 23671 1756 23705
rect 1704 23662 1756 23671
rect 1704 23369 1756 23378
rect 1704 23335 1713 23369
rect 1713 23335 1747 23369
rect 1747 23335 1756 23369
rect 1704 23326 1756 23335
rect 1704 23033 1756 23042
rect 1704 22999 1713 23033
rect 1713 22999 1747 23033
rect 1747 22999 1756 23033
rect 1704 22990 1756 22999
rect 1704 22697 1756 22706
rect 1704 22663 1713 22697
rect 1713 22663 1747 22697
rect 1747 22663 1756 22697
rect 1704 22654 1756 22663
rect 1704 22361 1756 22370
rect 1704 22327 1713 22361
rect 1713 22327 1747 22361
rect 1747 22327 1756 22361
rect 1704 22318 1756 22327
rect 1704 22025 1756 22034
rect 1704 21991 1713 22025
rect 1713 21991 1747 22025
rect 1747 21991 1756 22025
rect 1704 21982 1756 21991
rect 1704 21689 1756 21698
rect 1704 21655 1713 21689
rect 1713 21655 1747 21689
rect 1747 21655 1756 21689
rect 1704 21646 1756 21655
rect 1704 21353 1756 21362
rect 1704 21319 1713 21353
rect 1713 21319 1747 21353
rect 1747 21319 1756 21353
rect 1704 21310 1756 21319
rect 1704 21017 1756 21026
rect 1704 20983 1713 21017
rect 1713 20983 1747 21017
rect 1747 20983 1756 21017
rect 1704 20974 1756 20983
rect 1704 20681 1756 20690
rect 1704 20647 1713 20681
rect 1713 20647 1747 20681
rect 1747 20647 1756 20681
rect 1704 20638 1756 20647
rect 1704 20345 1756 20354
rect 1704 20311 1713 20345
rect 1713 20311 1747 20345
rect 1747 20311 1756 20345
rect 1704 20302 1756 20311
rect 1704 20009 1756 20018
rect 1704 19975 1713 20009
rect 1713 19975 1747 20009
rect 1747 19975 1756 20009
rect 1704 19966 1756 19975
rect 1704 19673 1756 19682
rect 1704 19639 1713 19673
rect 1713 19639 1747 19673
rect 1747 19639 1756 19673
rect 1704 19630 1756 19639
rect 1704 19337 1756 19346
rect 1704 19303 1713 19337
rect 1713 19303 1747 19337
rect 1747 19303 1756 19337
rect 1704 19294 1756 19303
rect 1704 19001 1756 19010
rect 1704 18967 1713 19001
rect 1713 18967 1747 19001
rect 1747 18967 1756 19001
rect 1704 18958 1756 18967
rect 1704 18665 1756 18674
rect 1704 18631 1713 18665
rect 1713 18631 1747 18665
rect 1747 18631 1756 18665
rect 1704 18622 1756 18631
rect 1704 18329 1756 18338
rect 1704 18295 1713 18329
rect 1713 18295 1747 18329
rect 1747 18295 1756 18329
rect 1704 18286 1756 18295
rect 1704 17993 1756 18002
rect 1704 17959 1713 17993
rect 1713 17959 1747 17993
rect 1747 17959 1756 17993
rect 1704 17950 1756 17959
rect 29562 17702 29614 17754
rect 34554 17702 34606 17754
rect 39546 17702 39598 17754
rect 44538 17702 44590 17754
rect 49530 17702 49582 17754
rect 54522 17702 54574 17754
rect 59514 17702 59566 17754
rect 64506 17702 64558 17754
rect 69498 17702 69550 17754
rect 74490 17702 74542 17754
rect 79482 17702 79534 17754
rect 84474 17702 84526 17754
rect 89466 17702 89518 17754
rect 94458 17702 94510 17754
rect 99450 17702 99502 17754
rect 104442 17702 104494 17754
rect 109434 17702 109486 17754
rect 114426 17702 114478 17754
rect 119418 17702 119470 17754
rect 124410 17702 124462 17754
rect 129402 17702 129454 17754
rect 134394 17702 134446 17754
rect 139386 17702 139438 17754
rect 144378 17702 144430 17754
rect 149370 17702 149422 17754
rect 154362 17702 154414 17754
rect 159354 17702 159406 17754
rect 164346 17702 164398 17754
rect 169338 17702 169390 17754
rect 174330 17702 174382 17754
rect 179322 17702 179374 17754
rect 184314 17702 184366 17754
rect 1704 17657 1756 17666
rect 1704 17623 1713 17657
rect 1713 17623 1747 17657
rect 1747 17623 1756 17657
rect 1704 17614 1756 17623
rect 1704 17321 1756 17330
rect 1704 17287 1713 17321
rect 1713 17287 1747 17321
rect 1747 17287 1756 17321
rect 1704 17278 1756 17287
rect 1704 16985 1756 16994
rect 1704 16951 1713 16985
rect 1713 16951 1747 16985
rect 1747 16951 1756 16985
rect 1704 16942 1756 16951
rect 1704 16649 1756 16658
rect 1704 16615 1713 16649
rect 1713 16615 1747 16649
rect 1747 16615 1756 16649
rect 1704 16606 1756 16615
rect 1704 16313 1756 16322
rect 1704 16279 1713 16313
rect 1713 16279 1747 16313
rect 1747 16279 1756 16313
rect 1704 16270 1756 16279
rect 1704 15977 1756 15986
rect 1704 15943 1713 15977
rect 1713 15943 1747 15977
rect 1747 15943 1756 15977
rect 1704 15934 1756 15943
rect 1704 15641 1756 15650
rect 1704 15607 1713 15641
rect 1713 15607 1747 15641
rect 1747 15607 1756 15641
rect 1704 15598 1756 15607
rect 1704 15305 1756 15314
rect 1704 15271 1713 15305
rect 1713 15271 1747 15305
rect 1747 15271 1756 15305
rect 1704 15262 1756 15271
rect 1704 14969 1756 14978
rect 1704 14935 1713 14969
rect 1713 14935 1747 14969
rect 1747 14935 1756 14969
rect 1704 14926 1756 14935
rect 1704 14633 1756 14642
rect 1704 14599 1713 14633
rect 1713 14599 1747 14633
rect 1747 14599 1756 14633
rect 1704 14590 1756 14599
rect 1704 14297 1756 14306
rect 1704 14263 1713 14297
rect 1713 14263 1747 14297
rect 1747 14263 1756 14297
rect 1704 14254 1756 14263
rect 216910 29417 216962 29426
rect 216910 29383 216919 29417
rect 216919 29383 216953 29417
rect 216953 29383 216962 29417
rect 216910 29374 216962 29383
rect 216910 29081 216962 29090
rect 216910 29047 216919 29081
rect 216919 29047 216953 29081
rect 216953 29047 216962 29081
rect 216910 29038 216962 29047
rect 216910 28745 216962 28754
rect 216910 28711 216919 28745
rect 216919 28711 216953 28745
rect 216953 28711 216962 28745
rect 216910 28702 216962 28711
rect 216910 28409 216962 28418
rect 216910 28375 216919 28409
rect 216919 28375 216953 28409
rect 216953 28375 216962 28409
rect 216910 28366 216962 28375
rect 216910 28073 216962 28082
rect 216910 28039 216919 28073
rect 216919 28039 216953 28073
rect 216953 28039 216962 28073
rect 216910 28030 216962 28039
rect 216910 27737 216962 27746
rect 216910 27703 216919 27737
rect 216919 27703 216953 27737
rect 216953 27703 216962 27737
rect 216910 27694 216962 27703
rect 216910 27401 216962 27410
rect 216910 27367 216919 27401
rect 216919 27367 216953 27401
rect 216953 27367 216962 27401
rect 216910 27358 216962 27367
rect 216910 27065 216962 27074
rect 216910 27031 216919 27065
rect 216919 27031 216953 27065
rect 216953 27031 216962 27065
rect 216910 27022 216962 27031
rect 216910 26729 216962 26738
rect 216910 26695 216919 26729
rect 216919 26695 216953 26729
rect 216953 26695 216962 26729
rect 216910 26686 216962 26695
rect 216910 26393 216962 26402
rect 216910 26359 216919 26393
rect 216919 26359 216953 26393
rect 216953 26359 216962 26393
rect 216910 26350 216962 26359
rect 216910 26057 216962 26066
rect 216910 26023 216919 26057
rect 216919 26023 216953 26057
rect 216953 26023 216962 26057
rect 216910 26014 216962 26023
rect 216910 25721 216962 25730
rect 216910 25687 216919 25721
rect 216919 25687 216953 25721
rect 216953 25687 216962 25721
rect 216910 25678 216962 25687
rect 216910 25385 216962 25394
rect 216910 25351 216919 25385
rect 216919 25351 216953 25385
rect 216953 25351 216962 25385
rect 216910 25342 216962 25351
rect 216910 25049 216962 25058
rect 216910 25015 216919 25049
rect 216919 25015 216953 25049
rect 216953 25015 216962 25049
rect 216910 25006 216962 25015
rect 216910 24713 216962 24722
rect 216910 24679 216919 24713
rect 216919 24679 216953 24713
rect 216953 24679 216962 24713
rect 216910 24670 216962 24679
rect 216910 24377 216962 24386
rect 216910 24343 216919 24377
rect 216919 24343 216953 24377
rect 216953 24343 216962 24377
rect 216910 24334 216962 24343
rect 203201 24176 203253 24228
rect 216910 24041 216962 24050
rect 216910 24007 216919 24041
rect 216919 24007 216953 24041
rect 216953 24007 216962 24041
rect 216910 23998 216962 24007
rect 216910 23705 216962 23714
rect 216910 23671 216919 23705
rect 216919 23671 216953 23705
rect 216953 23671 216962 23705
rect 216910 23662 216962 23671
rect 216910 23369 216962 23378
rect 216910 23335 216919 23369
rect 216919 23335 216953 23369
rect 216953 23335 216962 23369
rect 216910 23326 216962 23335
rect 216910 23033 216962 23042
rect 216910 22999 216919 23033
rect 216919 22999 216953 23033
rect 216953 22999 216962 23033
rect 216910 22990 216962 22999
rect 203121 22618 203173 22670
rect 216910 22697 216962 22706
rect 216910 22663 216919 22697
rect 216919 22663 216953 22697
rect 216953 22663 216962 22697
rect 216910 22654 216962 22663
rect 216910 22361 216962 22370
rect 216910 22327 216919 22361
rect 216919 22327 216953 22361
rect 216953 22327 216962 22361
rect 216910 22318 216962 22327
rect 216910 22025 216962 22034
rect 216910 21991 216919 22025
rect 216919 21991 216953 22025
rect 216953 21991 216962 22025
rect 216910 21982 216962 21991
rect 216910 21689 216962 21698
rect 216910 21655 216919 21689
rect 216919 21655 216953 21689
rect 216953 21655 216962 21689
rect 216910 21646 216962 21655
rect 203041 21348 203093 21400
rect 216910 21353 216962 21362
rect 216910 21319 216919 21353
rect 216919 21319 216953 21353
rect 216953 21319 216962 21353
rect 216910 21310 216962 21319
rect 216910 21017 216962 21026
rect 216910 20983 216919 21017
rect 216919 20983 216953 21017
rect 216953 20983 216962 21017
rect 216910 20974 216962 20983
rect 216910 20681 216962 20690
rect 216910 20647 216919 20681
rect 216919 20647 216953 20681
rect 216953 20647 216962 20681
rect 216910 20638 216962 20647
rect 216910 20345 216962 20354
rect 216910 20311 216919 20345
rect 216919 20311 216953 20345
rect 216953 20311 216962 20345
rect 216910 20302 216962 20311
rect 216910 20009 216962 20018
rect 216910 19975 216919 20009
rect 216919 19975 216953 20009
rect 216953 19975 216962 20009
rect 216910 19966 216962 19975
rect 202961 19790 203013 19842
rect 216910 19673 216962 19682
rect 216910 19639 216919 19673
rect 216919 19639 216953 19673
rect 216953 19639 216962 19673
rect 216910 19630 216962 19639
rect 216910 19337 216962 19346
rect 216910 19303 216919 19337
rect 216919 19303 216953 19337
rect 216953 19303 216962 19337
rect 216910 19294 216962 19303
rect 216910 19001 216962 19010
rect 216910 18967 216919 19001
rect 216919 18967 216953 19001
rect 216953 18967 216962 19001
rect 216910 18958 216962 18967
rect 216910 18665 216962 18674
rect 216910 18631 216919 18665
rect 216919 18631 216953 18665
rect 216953 18631 216962 18665
rect 216910 18622 216962 18631
rect 202881 18520 202933 18572
rect 216910 18329 216962 18338
rect 216910 18295 216919 18329
rect 216919 18295 216953 18329
rect 216953 18295 216962 18329
rect 216910 18286 216962 18295
rect 216910 17993 216962 18002
rect 216910 17959 216919 17993
rect 216919 17959 216953 17993
rect 216953 17959 216962 17993
rect 216910 17950 216962 17959
rect 216910 17657 216962 17666
rect 216910 17623 216919 17657
rect 216919 17623 216953 17657
rect 216953 17623 216962 17657
rect 216910 17614 216962 17623
rect 216910 17321 216962 17330
rect 216910 17287 216919 17321
rect 216919 17287 216953 17321
rect 216953 17287 216962 17321
rect 216910 17278 216962 17287
rect 202801 16962 202853 17014
rect 216910 16985 216962 16994
rect 216910 16951 216919 16985
rect 216919 16951 216953 16985
rect 216953 16951 216962 16985
rect 216910 16942 216962 16951
rect 216910 16649 216962 16658
rect 216910 16615 216919 16649
rect 216919 16615 216953 16649
rect 216953 16615 216962 16649
rect 216910 16606 216962 16615
rect 216910 16313 216962 16322
rect 216910 16279 216919 16313
rect 216919 16279 216953 16313
rect 216953 16279 216962 16313
rect 216910 16270 216962 16279
rect 216910 15977 216962 15986
rect 216910 15943 216919 15977
rect 216919 15943 216953 15977
rect 216953 15943 216962 15977
rect 216910 15934 216962 15943
rect 202721 15692 202773 15744
rect 216910 15641 216962 15650
rect 216910 15607 216919 15641
rect 216919 15607 216953 15641
rect 216953 15607 216962 15641
rect 216910 15598 216962 15607
rect 216910 15305 216962 15314
rect 216910 15271 216919 15305
rect 216919 15271 216953 15305
rect 216953 15271 216962 15305
rect 216910 15262 216962 15271
rect 216910 14969 216962 14978
rect 216910 14935 216919 14969
rect 216919 14935 216953 14969
rect 216953 14935 216962 14969
rect 216910 14926 216962 14935
rect 216910 14633 216962 14642
rect 216910 14599 216919 14633
rect 216919 14599 216953 14633
rect 216953 14599 216962 14633
rect 216910 14590 216962 14599
rect 216910 14297 216962 14306
rect 216910 14263 216919 14297
rect 216919 14263 216953 14297
rect 216953 14263 216962 14297
rect 216910 14254 216962 14263
rect 202641 14134 202693 14186
rect 1704 13961 1756 13970
rect 1704 13927 1713 13961
rect 1713 13927 1747 13961
rect 1747 13927 1756 13961
rect 1704 13918 1756 13927
rect 216910 13961 216962 13970
rect 216910 13927 216919 13961
rect 216919 13927 216953 13961
rect 216953 13927 216962 13961
rect 216910 13918 216962 13927
rect 1704 13625 1756 13634
rect 1704 13591 1713 13625
rect 1713 13591 1747 13625
rect 1747 13591 1756 13625
rect 1704 13582 1756 13591
rect 216910 13625 216962 13634
rect 216910 13591 216919 13625
rect 216919 13591 216953 13625
rect 216953 13591 216962 13625
rect 216910 13582 216962 13591
rect 1704 13289 1756 13298
rect 1704 13255 1713 13289
rect 1713 13255 1747 13289
rect 1747 13255 1756 13289
rect 1704 13246 1756 13255
rect 216910 13289 216962 13298
rect 216910 13255 216919 13289
rect 216919 13255 216953 13289
rect 216953 13255 216962 13289
rect 216910 13246 216962 13255
rect 1704 12953 1756 12962
rect 1704 12919 1713 12953
rect 1713 12919 1747 12953
rect 1747 12919 1756 12953
rect 1704 12910 1756 12919
rect 216910 12953 216962 12962
rect 216910 12919 216919 12953
rect 216919 12919 216953 12953
rect 216953 12919 216962 12953
rect 216910 12910 216962 12919
rect 1704 12617 1756 12626
rect 1704 12583 1713 12617
rect 1713 12583 1747 12617
rect 1747 12583 1756 12617
rect 1704 12574 1756 12583
rect 216910 12617 216962 12626
rect 216910 12583 216919 12617
rect 216919 12583 216953 12617
rect 216953 12583 216962 12617
rect 216910 12574 216962 12583
rect 1704 12281 1756 12290
rect 1704 12247 1713 12281
rect 1713 12247 1747 12281
rect 1747 12247 1756 12281
rect 1704 12238 1756 12247
rect 216910 12281 216962 12290
rect 216910 12247 216919 12281
rect 216919 12247 216953 12281
rect 216953 12247 216962 12281
rect 216910 12238 216962 12247
rect 1704 11945 1756 11954
rect 1704 11911 1713 11945
rect 1713 11911 1747 11945
rect 1747 11911 1756 11945
rect 1704 11902 1756 11911
rect 216910 11945 216962 11954
rect 216910 11911 216919 11945
rect 216919 11911 216953 11945
rect 216953 11911 216962 11945
rect 216910 11902 216962 11911
rect 1704 11609 1756 11618
rect 1704 11575 1713 11609
rect 1713 11575 1747 11609
rect 1747 11575 1756 11609
rect 1704 11566 1756 11575
rect 216910 11609 216962 11618
rect 216910 11575 216919 11609
rect 216919 11575 216953 11609
rect 216953 11575 216962 11609
rect 216910 11566 216962 11575
rect 1704 11273 1756 11282
rect 1704 11239 1713 11273
rect 1713 11239 1747 11273
rect 1747 11239 1756 11273
rect 1704 11230 1756 11239
rect 216910 11273 216962 11282
rect 216910 11239 216919 11273
rect 216919 11239 216953 11273
rect 216953 11239 216962 11273
rect 216910 11230 216962 11239
rect 1704 10937 1756 10946
rect 1704 10903 1713 10937
rect 1713 10903 1747 10937
rect 1747 10903 1756 10937
rect 1704 10894 1756 10903
rect 216910 10937 216962 10946
rect 216910 10903 216919 10937
rect 216919 10903 216953 10937
rect 216953 10903 216962 10937
rect 216910 10894 216962 10903
rect 1704 10601 1756 10610
rect 1704 10567 1713 10601
rect 1713 10567 1747 10601
rect 1747 10567 1756 10601
rect 1704 10558 1756 10567
rect 216910 10601 216962 10610
rect 216910 10567 216919 10601
rect 216919 10567 216953 10601
rect 216953 10567 216962 10601
rect 216910 10558 216962 10567
rect 1704 10265 1756 10274
rect 1704 10231 1713 10265
rect 1713 10231 1747 10265
rect 1747 10231 1756 10265
rect 1704 10222 1756 10231
rect 216910 10265 216962 10274
rect 216910 10231 216919 10265
rect 216919 10231 216953 10265
rect 216953 10231 216962 10265
rect 216910 10222 216962 10231
rect 1704 9929 1756 9938
rect 1704 9895 1713 9929
rect 1713 9895 1747 9929
rect 1747 9895 1756 9929
rect 1704 9886 1756 9895
rect 216910 9929 216962 9938
rect 216910 9895 216919 9929
rect 216919 9895 216953 9929
rect 216953 9895 216962 9929
rect 216910 9886 216962 9895
rect 1704 9593 1756 9602
rect 1704 9559 1713 9593
rect 1713 9559 1747 9593
rect 1747 9559 1756 9593
rect 1704 9550 1756 9559
rect 216910 9593 216962 9602
rect 216910 9559 216919 9593
rect 216919 9559 216953 9593
rect 216953 9559 216962 9593
rect 216910 9550 216962 9559
rect 1704 9257 1756 9266
rect 1704 9223 1713 9257
rect 1713 9223 1747 9257
rect 1747 9223 1756 9257
rect 1704 9214 1756 9223
rect 216910 9257 216962 9266
rect 216910 9223 216919 9257
rect 216919 9223 216953 9257
rect 216953 9223 216962 9257
rect 216910 9214 216962 9223
rect 1704 8921 1756 8930
rect 1704 8887 1713 8921
rect 1713 8887 1747 8921
rect 1747 8887 1756 8921
rect 1704 8878 1756 8887
rect 216910 8921 216962 8930
rect 216910 8887 216919 8921
rect 216919 8887 216953 8921
rect 216953 8887 216962 8921
rect 216910 8878 216962 8887
rect 1704 8585 1756 8594
rect 1704 8551 1713 8585
rect 1713 8551 1747 8585
rect 1747 8551 1756 8585
rect 1704 8542 1756 8551
rect 216910 8585 216962 8594
rect 216910 8551 216919 8585
rect 216919 8551 216953 8585
rect 216953 8551 216962 8585
rect 216910 8542 216962 8551
rect 1704 8249 1756 8258
rect 1704 8215 1713 8249
rect 1713 8215 1747 8249
rect 1747 8215 1756 8249
rect 1704 8206 1756 8215
rect 216910 8249 216962 8258
rect 216910 8215 216919 8249
rect 216919 8215 216953 8249
rect 216953 8215 216962 8249
rect 216910 8206 216962 8215
rect 1704 7913 1756 7922
rect 1704 7879 1713 7913
rect 1713 7879 1747 7913
rect 1747 7879 1756 7913
rect 1704 7870 1756 7879
rect 216910 7913 216962 7922
rect 216910 7879 216919 7913
rect 216919 7879 216953 7913
rect 216953 7879 216962 7913
rect 216910 7870 216962 7879
rect 1704 7577 1756 7586
rect 1704 7543 1713 7577
rect 1713 7543 1747 7577
rect 1747 7543 1756 7577
rect 1704 7534 1756 7543
rect 216910 7577 216962 7586
rect 216910 7543 216919 7577
rect 216919 7543 216953 7577
rect 216953 7543 216962 7577
rect 216910 7534 216962 7543
rect 1704 7241 1756 7250
rect 1704 7207 1713 7241
rect 1713 7207 1747 7241
rect 1747 7207 1756 7241
rect 1704 7198 1756 7207
rect 216910 7241 216962 7250
rect 216910 7207 216919 7241
rect 216919 7207 216953 7241
rect 216953 7207 216962 7241
rect 216910 7198 216962 7207
rect 1704 6905 1756 6914
rect 1704 6871 1713 6905
rect 1713 6871 1747 6905
rect 1747 6871 1756 6905
rect 1704 6862 1756 6871
rect 216910 6905 216962 6914
rect 216910 6871 216919 6905
rect 216919 6871 216953 6905
rect 216953 6871 216962 6905
rect 216910 6862 216962 6871
rect 1704 6569 1756 6578
rect 1704 6535 1713 6569
rect 1713 6535 1747 6569
rect 1747 6535 1756 6569
rect 1704 6526 1756 6535
rect 216910 6569 216962 6578
rect 216910 6535 216919 6569
rect 216919 6535 216953 6569
rect 216953 6535 216962 6569
rect 216910 6526 216962 6535
rect 1704 6233 1756 6242
rect 1704 6199 1713 6233
rect 1713 6199 1747 6233
rect 1747 6199 1756 6233
rect 1704 6190 1756 6199
rect 216910 6233 216962 6242
rect 216910 6199 216919 6233
rect 216919 6199 216953 6233
rect 216953 6199 216962 6233
rect 216910 6190 216962 6199
rect 1704 5897 1756 5906
rect 1704 5863 1713 5897
rect 1713 5863 1747 5897
rect 1747 5863 1756 5897
rect 1704 5854 1756 5863
rect 216910 5897 216962 5906
rect 216910 5863 216919 5897
rect 216919 5863 216953 5897
rect 216953 5863 216962 5897
rect 216910 5854 216962 5863
rect 1704 5561 1756 5570
rect 1704 5527 1713 5561
rect 1713 5527 1747 5561
rect 1747 5527 1756 5561
rect 1704 5518 1756 5527
rect 216910 5561 216962 5570
rect 216910 5527 216919 5561
rect 216919 5527 216953 5561
rect 216953 5527 216962 5561
rect 216910 5518 216962 5527
rect 1704 5225 1756 5234
rect 1704 5191 1713 5225
rect 1713 5191 1747 5225
rect 1747 5191 1756 5225
rect 1704 5182 1756 5191
rect 216910 5225 216962 5234
rect 216910 5191 216919 5225
rect 216919 5191 216953 5225
rect 216953 5191 216962 5225
rect 216910 5182 216962 5191
rect 1704 4889 1756 4898
rect 1704 4855 1713 4889
rect 1713 4855 1747 4889
rect 1747 4855 1756 4889
rect 1704 4846 1756 4855
rect 216910 4889 216962 4898
rect 216910 4855 216919 4889
rect 216919 4855 216953 4889
rect 216953 4855 216962 4889
rect 216910 4846 216962 4855
rect 1704 4553 1756 4562
rect 1704 4519 1713 4553
rect 1713 4519 1747 4553
rect 1747 4519 1756 4553
rect 1704 4510 1756 4519
rect 216910 4553 216962 4562
rect 216910 4519 216919 4553
rect 216919 4519 216953 4553
rect 216953 4519 216962 4553
rect 216910 4510 216962 4519
rect 1704 4217 1756 4226
rect 1704 4183 1713 4217
rect 1713 4183 1747 4217
rect 1747 4183 1756 4217
rect 1704 4174 1756 4183
rect 216910 4217 216962 4226
rect 216910 4183 216919 4217
rect 216919 4183 216953 4217
rect 216953 4183 216962 4217
rect 216910 4174 216962 4183
rect 1704 3881 1756 3890
rect 1704 3847 1713 3881
rect 1713 3847 1747 3881
rect 1747 3847 1756 3881
rect 1704 3838 1756 3847
rect 216910 3881 216962 3890
rect 216910 3847 216919 3881
rect 216919 3847 216953 3881
rect 216953 3847 216962 3881
rect 216910 3838 216962 3847
rect 1704 3545 1756 3554
rect 1704 3511 1713 3545
rect 1713 3511 1747 3545
rect 1747 3511 1756 3545
rect 1704 3502 1756 3511
rect 216910 3545 216962 3554
rect 216910 3511 216919 3545
rect 216919 3511 216953 3545
rect 216953 3511 216962 3545
rect 216910 3502 216962 3511
rect 1704 3209 1756 3218
rect 1704 3175 1713 3209
rect 1713 3175 1747 3209
rect 1747 3175 1756 3209
rect 1704 3166 1756 3175
rect 216910 3209 216962 3218
rect 216910 3175 216919 3209
rect 216919 3175 216953 3209
rect 216953 3175 216962 3209
rect 216910 3166 216962 3175
rect 1704 2873 1756 2882
rect 1704 2839 1713 2873
rect 1713 2839 1747 2873
rect 1747 2839 1756 2873
rect 1704 2830 1756 2839
rect 216910 2873 216962 2882
rect 216910 2839 216919 2873
rect 216919 2839 216953 2873
rect 216953 2839 216962 2873
rect 216910 2830 216962 2839
rect 1704 2537 1756 2546
rect 1704 2503 1713 2537
rect 1713 2503 1747 2537
rect 1747 2503 1756 2537
rect 1704 2494 1756 2503
rect 216910 2537 216962 2546
rect 216910 2503 216919 2537
rect 216919 2503 216953 2537
rect 216953 2503 216962 2537
rect 216910 2494 216962 2503
rect 1704 2201 1756 2210
rect 1704 2167 1713 2201
rect 1713 2167 1747 2201
rect 1747 2167 1756 2201
rect 1704 2158 1756 2167
rect 216910 2201 216962 2210
rect 216910 2167 216919 2201
rect 216919 2167 216953 2201
rect 216953 2167 216962 2201
rect 216910 2158 216962 2167
rect 2040 1865 2092 1874
rect 3720 1865 3772 1874
rect 5400 1865 5452 1874
rect 7080 1865 7132 1874
rect 8760 1865 8812 1874
rect 10440 1865 10492 1874
rect 12120 1865 12172 1874
rect 13800 1865 13852 1874
rect 15480 1865 15532 1874
rect 17160 1865 17212 1874
rect 18840 1865 18892 1874
rect 20520 1865 20572 1874
rect 22200 1865 22252 1874
rect 23880 1865 23932 1874
rect 25560 1865 25612 1874
rect 27240 1865 27292 1874
rect 28920 1865 28972 1874
rect 30600 1865 30652 1874
rect 32280 1865 32332 1874
rect 33960 1865 34012 1874
rect 35640 1865 35692 1874
rect 37320 1865 37372 1874
rect 39000 1865 39052 1874
rect 40680 1865 40732 1874
rect 42360 1865 42412 1874
rect 44040 1865 44092 1874
rect 45720 1865 45772 1874
rect 47400 1865 47452 1874
rect 49080 1865 49132 1874
rect 50760 1865 50812 1874
rect 52440 1865 52492 1874
rect 54120 1865 54172 1874
rect 55800 1865 55852 1874
rect 57480 1865 57532 1874
rect 59160 1865 59212 1874
rect 60840 1865 60892 1874
rect 62520 1865 62572 1874
rect 64200 1865 64252 1874
rect 65880 1865 65932 1874
rect 67560 1865 67612 1874
rect 69240 1865 69292 1874
rect 70920 1865 70972 1874
rect 72600 1865 72652 1874
rect 74280 1865 74332 1874
rect 75960 1865 76012 1874
rect 77640 1865 77692 1874
rect 79320 1865 79372 1874
rect 81000 1865 81052 1874
rect 82680 1865 82732 1874
rect 84360 1865 84412 1874
rect 86040 1865 86092 1874
rect 87720 1865 87772 1874
rect 89400 1865 89452 1874
rect 91080 1865 91132 1874
rect 92760 1865 92812 1874
rect 94440 1865 94492 1874
rect 96120 1865 96172 1874
rect 97800 1865 97852 1874
rect 99480 1865 99532 1874
rect 101160 1865 101212 1874
rect 102840 1865 102892 1874
rect 104520 1865 104572 1874
rect 106200 1865 106252 1874
rect 107880 1865 107932 1874
rect 109560 1865 109612 1874
rect 111240 1865 111292 1874
rect 112920 1865 112972 1874
rect 114600 1865 114652 1874
rect 116280 1865 116332 1874
rect 117960 1865 118012 1874
rect 119640 1865 119692 1874
rect 121320 1865 121372 1874
rect 123000 1865 123052 1874
rect 124680 1865 124732 1874
rect 126360 1865 126412 1874
rect 128040 1865 128092 1874
rect 129720 1865 129772 1874
rect 131400 1865 131452 1874
rect 133080 1865 133132 1874
rect 134760 1865 134812 1874
rect 136440 1865 136492 1874
rect 138120 1865 138172 1874
rect 139800 1865 139852 1874
rect 141480 1865 141532 1874
rect 143160 1865 143212 1874
rect 144840 1865 144892 1874
rect 146520 1865 146572 1874
rect 148200 1865 148252 1874
rect 149880 1865 149932 1874
rect 151560 1865 151612 1874
rect 153240 1865 153292 1874
rect 154920 1865 154972 1874
rect 156600 1865 156652 1874
rect 158280 1865 158332 1874
rect 159960 1865 160012 1874
rect 161640 1865 161692 1874
rect 163320 1865 163372 1874
rect 165000 1865 165052 1874
rect 166680 1865 166732 1874
rect 168360 1865 168412 1874
rect 170040 1865 170092 1874
rect 171720 1865 171772 1874
rect 173400 1865 173452 1874
rect 175080 1865 175132 1874
rect 176760 1865 176812 1874
rect 178440 1865 178492 1874
rect 180120 1865 180172 1874
rect 181800 1865 181852 1874
rect 183480 1865 183532 1874
rect 185160 1865 185212 1874
rect 186840 1865 186892 1874
rect 188520 1865 188572 1874
rect 190200 1865 190252 1874
rect 191880 1865 191932 1874
rect 193560 1865 193612 1874
rect 195240 1865 195292 1874
rect 196920 1865 196972 1874
rect 198600 1865 198652 1874
rect 200280 1865 200332 1874
rect 201960 1865 202012 1874
rect 203640 1865 203692 1874
rect 205320 1865 205372 1874
rect 207000 1865 207052 1874
rect 208680 1865 208732 1874
rect 210360 1865 210412 1874
rect 212040 1865 212092 1874
rect 213720 1865 213772 1874
rect 215400 1865 215452 1874
rect 2040 1831 2049 1865
rect 2049 1831 2083 1865
rect 2083 1831 2092 1865
rect 3720 1831 3729 1865
rect 3729 1831 3763 1865
rect 3763 1831 3772 1865
rect 5400 1831 5409 1865
rect 5409 1831 5443 1865
rect 5443 1831 5452 1865
rect 7080 1831 7089 1865
rect 7089 1831 7123 1865
rect 7123 1831 7132 1865
rect 8760 1831 8769 1865
rect 8769 1831 8803 1865
rect 8803 1831 8812 1865
rect 10440 1831 10449 1865
rect 10449 1831 10483 1865
rect 10483 1831 10492 1865
rect 12120 1831 12129 1865
rect 12129 1831 12163 1865
rect 12163 1831 12172 1865
rect 13800 1831 13809 1865
rect 13809 1831 13843 1865
rect 13843 1831 13852 1865
rect 15480 1831 15489 1865
rect 15489 1831 15523 1865
rect 15523 1831 15532 1865
rect 17160 1831 17169 1865
rect 17169 1831 17203 1865
rect 17203 1831 17212 1865
rect 18840 1831 18849 1865
rect 18849 1831 18883 1865
rect 18883 1831 18892 1865
rect 20520 1831 20529 1865
rect 20529 1831 20563 1865
rect 20563 1831 20572 1865
rect 22200 1831 22209 1865
rect 22209 1831 22243 1865
rect 22243 1831 22252 1865
rect 23880 1831 23889 1865
rect 23889 1831 23923 1865
rect 23923 1831 23932 1865
rect 25560 1831 25569 1865
rect 25569 1831 25603 1865
rect 25603 1831 25612 1865
rect 27240 1831 27249 1865
rect 27249 1831 27283 1865
rect 27283 1831 27292 1865
rect 28920 1831 28929 1865
rect 28929 1831 28963 1865
rect 28963 1831 28972 1865
rect 30600 1831 30609 1865
rect 30609 1831 30643 1865
rect 30643 1831 30652 1865
rect 32280 1831 32289 1865
rect 32289 1831 32323 1865
rect 32323 1831 32332 1865
rect 33960 1831 33969 1865
rect 33969 1831 34003 1865
rect 34003 1831 34012 1865
rect 35640 1831 35649 1865
rect 35649 1831 35683 1865
rect 35683 1831 35692 1865
rect 37320 1831 37329 1865
rect 37329 1831 37363 1865
rect 37363 1831 37372 1865
rect 39000 1831 39009 1865
rect 39009 1831 39043 1865
rect 39043 1831 39052 1865
rect 40680 1831 40689 1865
rect 40689 1831 40723 1865
rect 40723 1831 40732 1865
rect 42360 1831 42369 1865
rect 42369 1831 42403 1865
rect 42403 1831 42412 1865
rect 44040 1831 44049 1865
rect 44049 1831 44083 1865
rect 44083 1831 44092 1865
rect 45720 1831 45729 1865
rect 45729 1831 45763 1865
rect 45763 1831 45772 1865
rect 47400 1831 47409 1865
rect 47409 1831 47443 1865
rect 47443 1831 47452 1865
rect 49080 1831 49089 1865
rect 49089 1831 49123 1865
rect 49123 1831 49132 1865
rect 50760 1831 50769 1865
rect 50769 1831 50803 1865
rect 50803 1831 50812 1865
rect 52440 1831 52449 1865
rect 52449 1831 52483 1865
rect 52483 1831 52492 1865
rect 54120 1831 54129 1865
rect 54129 1831 54163 1865
rect 54163 1831 54172 1865
rect 55800 1831 55809 1865
rect 55809 1831 55843 1865
rect 55843 1831 55852 1865
rect 57480 1831 57489 1865
rect 57489 1831 57523 1865
rect 57523 1831 57532 1865
rect 59160 1831 59169 1865
rect 59169 1831 59203 1865
rect 59203 1831 59212 1865
rect 60840 1831 60849 1865
rect 60849 1831 60883 1865
rect 60883 1831 60892 1865
rect 62520 1831 62529 1865
rect 62529 1831 62563 1865
rect 62563 1831 62572 1865
rect 64200 1831 64209 1865
rect 64209 1831 64243 1865
rect 64243 1831 64252 1865
rect 65880 1831 65889 1865
rect 65889 1831 65923 1865
rect 65923 1831 65932 1865
rect 67560 1831 67569 1865
rect 67569 1831 67603 1865
rect 67603 1831 67612 1865
rect 69240 1831 69249 1865
rect 69249 1831 69283 1865
rect 69283 1831 69292 1865
rect 70920 1831 70929 1865
rect 70929 1831 70963 1865
rect 70963 1831 70972 1865
rect 72600 1831 72609 1865
rect 72609 1831 72643 1865
rect 72643 1831 72652 1865
rect 74280 1831 74289 1865
rect 74289 1831 74323 1865
rect 74323 1831 74332 1865
rect 75960 1831 75969 1865
rect 75969 1831 76003 1865
rect 76003 1831 76012 1865
rect 77640 1831 77649 1865
rect 77649 1831 77683 1865
rect 77683 1831 77692 1865
rect 79320 1831 79329 1865
rect 79329 1831 79363 1865
rect 79363 1831 79372 1865
rect 81000 1831 81009 1865
rect 81009 1831 81043 1865
rect 81043 1831 81052 1865
rect 82680 1831 82689 1865
rect 82689 1831 82723 1865
rect 82723 1831 82732 1865
rect 84360 1831 84369 1865
rect 84369 1831 84403 1865
rect 84403 1831 84412 1865
rect 86040 1831 86049 1865
rect 86049 1831 86083 1865
rect 86083 1831 86092 1865
rect 87720 1831 87729 1865
rect 87729 1831 87763 1865
rect 87763 1831 87772 1865
rect 89400 1831 89409 1865
rect 89409 1831 89443 1865
rect 89443 1831 89452 1865
rect 91080 1831 91089 1865
rect 91089 1831 91123 1865
rect 91123 1831 91132 1865
rect 92760 1831 92769 1865
rect 92769 1831 92803 1865
rect 92803 1831 92812 1865
rect 94440 1831 94449 1865
rect 94449 1831 94483 1865
rect 94483 1831 94492 1865
rect 96120 1831 96129 1865
rect 96129 1831 96163 1865
rect 96163 1831 96172 1865
rect 97800 1831 97809 1865
rect 97809 1831 97843 1865
rect 97843 1831 97852 1865
rect 99480 1831 99489 1865
rect 99489 1831 99523 1865
rect 99523 1831 99532 1865
rect 101160 1831 101169 1865
rect 101169 1831 101203 1865
rect 101203 1831 101212 1865
rect 102840 1831 102849 1865
rect 102849 1831 102883 1865
rect 102883 1831 102892 1865
rect 104520 1831 104529 1865
rect 104529 1831 104563 1865
rect 104563 1831 104572 1865
rect 106200 1831 106209 1865
rect 106209 1831 106243 1865
rect 106243 1831 106252 1865
rect 107880 1831 107889 1865
rect 107889 1831 107923 1865
rect 107923 1831 107932 1865
rect 109560 1831 109569 1865
rect 109569 1831 109603 1865
rect 109603 1831 109612 1865
rect 111240 1831 111249 1865
rect 111249 1831 111283 1865
rect 111283 1831 111292 1865
rect 112920 1831 112929 1865
rect 112929 1831 112963 1865
rect 112963 1831 112972 1865
rect 114600 1831 114609 1865
rect 114609 1831 114643 1865
rect 114643 1831 114652 1865
rect 116280 1831 116289 1865
rect 116289 1831 116323 1865
rect 116323 1831 116332 1865
rect 117960 1831 117969 1865
rect 117969 1831 118003 1865
rect 118003 1831 118012 1865
rect 119640 1831 119649 1865
rect 119649 1831 119683 1865
rect 119683 1831 119692 1865
rect 121320 1831 121329 1865
rect 121329 1831 121363 1865
rect 121363 1831 121372 1865
rect 123000 1831 123009 1865
rect 123009 1831 123043 1865
rect 123043 1831 123052 1865
rect 124680 1831 124689 1865
rect 124689 1831 124723 1865
rect 124723 1831 124732 1865
rect 126360 1831 126369 1865
rect 126369 1831 126403 1865
rect 126403 1831 126412 1865
rect 128040 1831 128049 1865
rect 128049 1831 128083 1865
rect 128083 1831 128092 1865
rect 129720 1831 129729 1865
rect 129729 1831 129763 1865
rect 129763 1831 129772 1865
rect 131400 1831 131409 1865
rect 131409 1831 131443 1865
rect 131443 1831 131452 1865
rect 133080 1831 133089 1865
rect 133089 1831 133123 1865
rect 133123 1831 133132 1865
rect 134760 1831 134769 1865
rect 134769 1831 134803 1865
rect 134803 1831 134812 1865
rect 136440 1831 136449 1865
rect 136449 1831 136483 1865
rect 136483 1831 136492 1865
rect 138120 1831 138129 1865
rect 138129 1831 138163 1865
rect 138163 1831 138172 1865
rect 139800 1831 139809 1865
rect 139809 1831 139843 1865
rect 139843 1831 139852 1865
rect 141480 1831 141489 1865
rect 141489 1831 141523 1865
rect 141523 1831 141532 1865
rect 143160 1831 143169 1865
rect 143169 1831 143203 1865
rect 143203 1831 143212 1865
rect 144840 1831 144849 1865
rect 144849 1831 144883 1865
rect 144883 1831 144892 1865
rect 146520 1831 146529 1865
rect 146529 1831 146563 1865
rect 146563 1831 146572 1865
rect 148200 1831 148209 1865
rect 148209 1831 148243 1865
rect 148243 1831 148252 1865
rect 149880 1831 149889 1865
rect 149889 1831 149923 1865
rect 149923 1831 149932 1865
rect 151560 1831 151569 1865
rect 151569 1831 151603 1865
rect 151603 1831 151612 1865
rect 153240 1831 153249 1865
rect 153249 1831 153283 1865
rect 153283 1831 153292 1865
rect 154920 1831 154929 1865
rect 154929 1831 154963 1865
rect 154963 1831 154972 1865
rect 156600 1831 156609 1865
rect 156609 1831 156643 1865
rect 156643 1831 156652 1865
rect 158280 1831 158289 1865
rect 158289 1831 158323 1865
rect 158323 1831 158332 1865
rect 159960 1831 159969 1865
rect 159969 1831 160003 1865
rect 160003 1831 160012 1865
rect 161640 1831 161649 1865
rect 161649 1831 161683 1865
rect 161683 1831 161692 1865
rect 163320 1831 163329 1865
rect 163329 1831 163363 1865
rect 163363 1831 163372 1865
rect 165000 1831 165009 1865
rect 165009 1831 165043 1865
rect 165043 1831 165052 1865
rect 166680 1831 166689 1865
rect 166689 1831 166723 1865
rect 166723 1831 166732 1865
rect 168360 1831 168369 1865
rect 168369 1831 168403 1865
rect 168403 1831 168412 1865
rect 170040 1831 170049 1865
rect 170049 1831 170083 1865
rect 170083 1831 170092 1865
rect 171720 1831 171729 1865
rect 171729 1831 171763 1865
rect 171763 1831 171772 1865
rect 173400 1831 173409 1865
rect 173409 1831 173443 1865
rect 173443 1831 173452 1865
rect 175080 1831 175089 1865
rect 175089 1831 175123 1865
rect 175123 1831 175132 1865
rect 176760 1831 176769 1865
rect 176769 1831 176803 1865
rect 176803 1831 176812 1865
rect 178440 1831 178449 1865
rect 178449 1831 178483 1865
rect 178483 1831 178492 1865
rect 180120 1831 180129 1865
rect 180129 1831 180163 1865
rect 180163 1831 180172 1865
rect 181800 1831 181809 1865
rect 181809 1831 181843 1865
rect 181843 1831 181852 1865
rect 183480 1831 183489 1865
rect 183489 1831 183523 1865
rect 183523 1831 183532 1865
rect 185160 1831 185169 1865
rect 185169 1831 185203 1865
rect 185203 1831 185212 1865
rect 186840 1831 186849 1865
rect 186849 1831 186883 1865
rect 186883 1831 186892 1865
rect 188520 1831 188529 1865
rect 188529 1831 188563 1865
rect 188563 1831 188572 1865
rect 190200 1831 190209 1865
rect 190209 1831 190243 1865
rect 190243 1831 190252 1865
rect 191880 1831 191889 1865
rect 191889 1831 191923 1865
rect 191923 1831 191932 1865
rect 193560 1831 193569 1865
rect 193569 1831 193603 1865
rect 193603 1831 193612 1865
rect 195240 1831 195249 1865
rect 195249 1831 195283 1865
rect 195283 1831 195292 1865
rect 196920 1831 196929 1865
rect 196929 1831 196963 1865
rect 196963 1831 196972 1865
rect 198600 1831 198609 1865
rect 198609 1831 198643 1865
rect 198643 1831 198652 1865
rect 200280 1831 200289 1865
rect 200289 1831 200323 1865
rect 200323 1831 200332 1865
rect 201960 1831 201969 1865
rect 201969 1831 202003 1865
rect 202003 1831 202012 1865
rect 203640 1831 203649 1865
rect 203649 1831 203683 1865
rect 203683 1831 203692 1865
rect 205320 1831 205329 1865
rect 205329 1831 205363 1865
rect 205363 1831 205372 1865
rect 207000 1831 207009 1865
rect 207009 1831 207043 1865
rect 207043 1831 207052 1865
rect 208680 1831 208689 1865
rect 208689 1831 208723 1865
rect 208723 1831 208732 1865
rect 210360 1831 210369 1865
rect 210369 1831 210403 1865
rect 210403 1831 210412 1865
rect 212040 1831 212049 1865
rect 212049 1831 212083 1865
rect 212083 1831 212092 1865
rect 213720 1831 213729 1865
rect 213729 1831 213763 1865
rect 213763 1831 213772 1865
rect 215400 1831 215409 1865
rect 215409 1831 215443 1865
rect 215443 1831 215452 1865
rect 2040 1822 2092 1831
rect 3720 1822 3772 1831
rect 5400 1822 5452 1831
rect 7080 1822 7132 1831
rect 8760 1822 8812 1831
rect 10440 1822 10492 1831
rect 12120 1822 12172 1831
rect 13800 1822 13852 1831
rect 15480 1822 15532 1831
rect 17160 1822 17212 1831
rect 18840 1822 18892 1831
rect 20520 1822 20572 1831
rect 22200 1822 22252 1831
rect 23880 1822 23932 1831
rect 25560 1822 25612 1831
rect 27240 1822 27292 1831
rect 28920 1822 28972 1831
rect 30600 1822 30652 1831
rect 32280 1822 32332 1831
rect 33960 1822 34012 1831
rect 35640 1822 35692 1831
rect 37320 1822 37372 1831
rect 39000 1822 39052 1831
rect 40680 1822 40732 1831
rect 42360 1822 42412 1831
rect 44040 1822 44092 1831
rect 45720 1822 45772 1831
rect 47400 1822 47452 1831
rect 49080 1822 49132 1831
rect 50760 1822 50812 1831
rect 52440 1822 52492 1831
rect 54120 1822 54172 1831
rect 55800 1822 55852 1831
rect 57480 1822 57532 1831
rect 59160 1822 59212 1831
rect 60840 1822 60892 1831
rect 62520 1822 62572 1831
rect 64200 1822 64252 1831
rect 65880 1822 65932 1831
rect 67560 1822 67612 1831
rect 69240 1822 69292 1831
rect 70920 1822 70972 1831
rect 72600 1822 72652 1831
rect 74280 1822 74332 1831
rect 75960 1822 76012 1831
rect 77640 1822 77692 1831
rect 79320 1822 79372 1831
rect 81000 1822 81052 1831
rect 82680 1822 82732 1831
rect 84360 1822 84412 1831
rect 86040 1822 86092 1831
rect 87720 1822 87772 1831
rect 89400 1822 89452 1831
rect 91080 1822 91132 1831
rect 92760 1822 92812 1831
rect 94440 1822 94492 1831
rect 96120 1822 96172 1831
rect 97800 1822 97852 1831
rect 99480 1822 99532 1831
rect 101160 1822 101212 1831
rect 102840 1822 102892 1831
rect 104520 1822 104572 1831
rect 106200 1822 106252 1831
rect 107880 1822 107932 1831
rect 109560 1822 109612 1831
rect 111240 1822 111292 1831
rect 112920 1822 112972 1831
rect 114600 1822 114652 1831
rect 116280 1822 116332 1831
rect 117960 1822 118012 1831
rect 119640 1822 119692 1831
rect 121320 1822 121372 1831
rect 123000 1822 123052 1831
rect 124680 1822 124732 1831
rect 126360 1822 126412 1831
rect 128040 1822 128092 1831
rect 129720 1822 129772 1831
rect 131400 1822 131452 1831
rect 133080 1822 133132 1831
rect 134760 1822 134812 1831
rect 136440 1822 136492 1831
rect 138120 1822 138172 1831
rect 139800 1822 139852 1831
rect 141480 1822 141532 1831
rect 143160 1822 143212 1831
rect 144840 1822 144892 1831
rect 146520 1822 146572 1831
rect 148200 1822 148252 1831
rect 149880 1822 149932 1831
rect 151560 1822 151612 1831
rect 153240 1822 153292 1831
rect 154920 1822 154972 1831
rect 156600 1822 156652 1831
rect 158280 1822 158332 1831
rect 159960 1822 160012 1831
rect 161640 1822 161692 1831
rect 163320 1822 163372 1831
rect 165000 1822 165052 1831
rect 166680 1822 166732 1831
rect 168360 1822 168412 1831
rect 170040 1822 170092 1831
rect 171720 1822 171772 1831
rect 173400 1822 173452 1831
rect 175080 1822 175132 1831
rect 176760 1822 176812 1831
rect 178440 1822 178492 1831
rect 180120 1822 180172 1831
rect 181800 1822 181852 1831
rect 183480 1822 183532 1831
rect 185160 1822 185212 1831
rect 186840 1822 186892 1831
rect 188520 1822 188572 1831
rect 190200 1822 190252 1831
rect 191880 1822 191932 1831
rect 193560 1822 193612 1831
rect 195240 1822 195292 1831
rect 196920 1822 196972 1831
rect 198600 1822 198652 1831
rect 200280 1822 200332 1831
rect 201960 1822 202012 1831
rect 203640 1822 203692 1831
rect 205320 1822 205372 1831
rect 207000 1822 207052 1831
rect 208680 1822 208732 1831
rect 210360 1822 210412 1831
rect 212040 1822 212092 1831
rect 213720 1822 213772 1831
rect 215400 1822 215452 1831
<< metal2 >>
rect 1618 141986 1842 142456
rect 2038 142372 2094 142381
rect 2038 142307 2094 142316
rect 3718 142372 3774 142381
rect 3718 142307 3774 142316
rect 5398 142372 5454 142381
rect 5398 142307 5454 142316
rect 7078 142372 7134 142381
rect 7078 142307 7134 142316
rect 8758 142372 8814 142381
rect 8758 142307 8814 142316
rect 10438 142372 10494 142381
rect 10438 142307 10494 142316
rect 12118 142372 12174 142381
rect 12118 142307 12174 142316
rect 13798 142372 13854 142381
rect 13798 142307 13854 142316
rect 15478 142372 15534 142381
rect 15478 142307 15534 142316
rect 17158 142372 17214 142381
rect 17158 142307 17214 142316
rect 18838 142372 18894 142381
rect 18838 142307 18894 142316
rect 20518 142372 20574 142381
rect 20518 142307 20574 142316
rect 22198 142372 22254 142381
rect 22198 142307 22254 142316
rect 23878 142372 23934 142381
rect 23878 142307 23934 142316
rect 25558 142372 25614 142381
rect 25558 142307 25614 142316
rect 27238 142372 27294 142381
rect 27238 142307 27294 142316
rect 28918 142372 28974 142381
rect 28918 142307 28974 142316
rect 30598 142372 30654 142381
rect 30598 142307 30654 142316
rect 32278 142372 32334 142381
rect 32278 142307 32334 142316
rect 33958 142372 34014 142381
rect 33958 142307 34014 142316
rect 35638 142372 35694 142381
rect 35638 142307 35694 142316
rect 37318 142372 37374 142381
rect 37318 142307 37374 142316
rect 38998 142372 39054 142381
rect 38998 142307 39054 142316
rect 40678 142372 40734 142381
rect 40678 142307 40734 142316
rect 42358 142372 42414 142381
rect 42358 142307 42414 142316
rect 44038 142372 44094 142381
rect 44038 142307 44094 142316
rect 45718 142372 45774 142381
rect 45718 142307 45774 142316
rect 47398 142372 47454 142381
rect 47398 142307 47454 142316
rect 49078 142372 49134 142381
rect 49078 142307 49134 142316
rect 50758 142372 50814 142381
rect 50758 142307 50814 142316
rect 52438 142372 52494 142381
rect 52438 142307 52494 142316
rect 54118 142372 54174 142381
rect 54118 142307 54174 142316
rect 55798 142372 55854 142381
rect 55798 142307 55854 142316
rect 57478 142372 57534 142381
rect 57478 142307 57534 142316
rect 59158 142372 59214 142381
rect 59158 142307 59214 142316
rect 60838 142372 60894 142381
rect 60838 142307 60894 142316
rect 62518 142372 62574 142381
rect 62518 142307 62574 142316
rect 64198 142372 64254 142381
rect 64198 142307 64254 142316
rect 65878 142372 65934 142381
rect 65878 142307 65934 142316
rect 67558 142372 67614 142381
rect 67558 142307 67614 142316
rect 69238 142372 69294 142381
rect 69238 142307 69294 142316
rect 70918 142372 70974 142381
rect 70918 142307 70974 142316
rect 72598 142372 72654 142381
rect 72598 142307 72654 142316
rect 74278 142372 74334 142381
rect 74278 142307 74334 142316
rect 75958 142372 76014 142381
rect 75958 142307 76014 142316
rect 77638 142372 77694 142381
rect 77638 142307 77694 142316
rect 79318 142372 79374 142381
rect 79318 142307 79374 142316
rect 80998 142372 81054 142381
rect 80998 142307 81054 142316
rect 82678 142372 82734 142381
rect 82678 142307 82734 142316
rect 84358 142372 84414 142381
rect 84358 142307 84414 142316
rect 86038 142372 86094 142381
rect 86038 142307 86094 142316
rect 87718 142372 87774 142381
rect 87718 142307 87774 142316
rect 89398 142372 89454 142381
rect 89398 142307 89454 142316
rect 91078 142372 91134 142381
rect 91078 142307 91134 142316
rect 92758 142372 92814 142381
rect 92758 142307 92814 142316
rect 94438 142372 94494 142381
rect 94438 142307 94494 142316
rect 96118 142372 96174 142381
rect 96118 142307 96174 142316
rect 97798 142372 97854 142381
rect 97798 142307 97854 142316
rect 99478 142372 99534 142381
rect 99478 142307 99534 142316
rect 101158 142372 101214 142381
rect 101158 142307 101214 142316
rect 102838 142372 102894 142381
rect 102838 142307 102894 142316
rect 104518 142372 104574 142381
rect 104518 142307 104574 142316
rect 106198 142372 106254 142381
rect 106198 142307 106254 142316
rect 107878 142372 107934 142381
rect 107878 142307 107934 142316
rect 109558 142372 109614 142381
rect 109558 142307 109614 142316
rect 111238 142372 111294 142381
rect 111238 142307 111294 142316
rect 112918 142372 112974 142381
rect 112918 142307 112974 142316
rect 114598 142372 114654 142381
rect 114598 142307 114654 142316
rect 116278 142372 116334 142381
rect 116278 142307 116334 142316
rect 117958 142372 118014 142381
rect 117958 142307 118014 142316
rect 119638 142372 119694 142381
rect 119638 142307 119694 142316
rect 121318 142372 121374 142381
rect 121318 142307 121374 142316
rect 122998 142372 123054 142381
rect 122998 142307 123054 142316
rect 124678 142372 124734 142381
rect 124678 142307 124734 142316
rect 126358 142372 126414 142381
rect 126358 142307 126414 142316
rect 128038 142372 128094 142381
rect 128038 142307 128094 142316
rect 129718 142372 129774 142381
rect 129718 142307 129774 142316
rect 131398 142372 131454 142381
rect 131398 142307 131454 142316
rect 133078 142372 133134 142381
rect 133078 142307 133134 142316
rect 134758 142372 134814 142381
rect 134758 142307 134814 142316
rect 136438 142372 136494 142381
rect 136438 142307 136494 142316
rect 138118 142372 138174 142381
rect 138118 142307 138174 142316
rect 139798 142372 139854 142381
rect 139798 142307 139854 142316
rect 141478 142372 141534 142381
rect 141478 142307 141534 142316
rect 143158 142372 143214 142381
rect 143158 142307 143214 142316
rect 144838 142372 144894 142381
rect 144838 142307 144894 142316
rect 146518 142372 146574 142381
rect 146518 142307 146574 142316
rect 148198 142372 148254 142381
rect 148198 142307 148254 142316
rect 149878 142372 149934 142381
rect 149878 142307 149934 142316
rect 151558 142372 151614 142381
rect 151558 142307 151614 142316
rect 153238 142372 153294 142381
rect 153238 142307 153294 142316
rect 154918 142372 154974 142381
rect 154918 142307 154974 142316
rect 156598 142372 156654 142381
rect 156598 142307 156654 142316
rect 158278 142372 158334 142381
rect 158278 142307 158334 142316
rect 159958 142372 160014 142381
rect 159958 142307 160014 142316
rect 161638 142372 161694 142381
rect 161638 142307 161694 142316
rect 163318 142372 163374 142381
rect 163318 142307 163374 142316
rect 164998 142372 165054 142381
rect 164998 142307 165054 142316
rect 166678 142372 166734 142381
rect 166678 142307 166734 142316
rect 168358 142372 168414 142381
rect 168358 142307 168414 142316
rect 170038 142372 170094 142381
rect 170038 142307 170094 142316
rect 171718 142372 171774 142381
rect 171718 142307 171774 142316
rect 173398 142372 173454 142381
rect 173398 142307 173454 142316
rect 175078 142372 175134 142381
rect 175078 142307 175134 142316
rect 176758 142372 176814 142381
rect 176758 142307 176814 142316
rect 178438 142372 178494 142381
rect 178438 142307 178494 142316
rect 180118 142372 180174 142381
rect 180118 142307 180174 142316
rect 181798 142372 181854 142381
rect 181798 142307 181854 142316
rect 183478 142372 183534 142381
rect 183478 142307 183534 142316
rect 185158 142372 185214 142381
rect 185158 142307 185214 142316
rect 186838 142372 186894 142381
rect 186838 142307 186894 142316
rect 188518 142372 188574 142381
rect 188518 142307 188574 142316
rect 190198 142372 190254 142381
rect 190198 142307 190254 142316
rect 191878 142372 191934 142381
rect 191878 142307 191934 142316
rect 193558 142372 193614 142381
rect 193558 142307 193614 142316
rect 195238 142372 195294 142381
rect 195238 142307 195294 142316
rect 196918 142372 196974 142381
rect 196918 142307 196974 142316
rect 198598 142372 198654 142381
rect 198598 142307 198654 142316
rect 200278 142372 200334 142381
rect 200278 142307 200334 142316
rect 201958 142372 202014 142381
rect 201958 142307 202014 142316
rect 203638 142372 203694 142381
rect 203638 142307 203694 142316
rect 205318 142372 205374 142381
rect 205318 142307 205374 142316
rect 206998 142372 207054 142381
rect 206998 142307 207054 142316
rect 208678 142372 208734 142381
rect 208678 142307 208734 142316
rect 210358 142372 210414 142381
rect 210358 142307 210414 142316
rect 212038 142372 212094 142381
rect 212038 142307 212094 142316
rect 213718 142372 213774 142381
rect 213718 142307 213774 142316
rect 215398 142372 215454 142381
rect 215398 142307 215454 142316
rect 1618 141934 1704 141986
rect 1756 141934 1842 141986
rect 1618 141652 1842 141934
rect 216824 141986 217048 142456
rect 216824 141934 216910 141986
rect 216962 141934 217048 141986
rect 203400 141728 203456 141737
rect 203400 141663 203456 141672
rect 1618 141596 1702 141652
rect 1758 141596 1842 141652
rect 1618 141314 1842 141596
rect 198642 141472 198698 141481
rect 198642 141407 198698 141416
rect 199810 141472 199866 141481
rect 199810 141407 199866 141416
rect 200978 141472 201034 141481
rect 200978 141407 201034 141416
rect 1618 141262 1704 141314
rect 1756 141262 1842 141314
rect 1618 140978 1842 141262
rect 1618 140926 1704 140978
rect 1756 140926 1842 140978
rect 1618 140642 1842 140926
rect 1618 140590 1704 140642
rect 1756 140590 1842 140642
rect 1618 140306 1842 140590
rect 1618 140254 1704 140306
rect 1756 140254 1842 140306
rect 1618 139972 1842 140254
rect 1618 139916 1702 139972
rect 1758 139916 1842 139972
rect 1618 139634 1842 139916
rect 1618 139582 1704 139634
rect 1756 139582 1842 139634
rect 1618 139298 1842 139582
rect 1618 139246 1704 139298
rect 1756 139246 1842 139298
rect 1618 138962 1842 139246
rect 1618 138910 1704 138962
rect 1756 138910 1842 138962
rect 1618 138626 1842 138910
rect 1618 138574 1704 138626
rect 1756 138574 1842 138626
rect 1618 138292 1842 138574
rect 1618 138236 1702 138292
rect 1758 138236 1842 138292
rect 1618 137954 1842 138236
rect 1618 137902 1704 137954
rect 1756 137902 1842 137954
rect 1618 137618 1842 137902
rect 1618 137566 1704 137618
rect 1756 137566 1842 137618
rect 1618 137282 1842 137566
rect 1618 137230 1704 137282
rect 1756 137230 1842 137282
rect 1618 136946 1842 137230
rect 1618 136894 1704 136946
rect 1756 136894 1842 136946
rect 1618 136612 1842 136894
rect 1618 136556 1702 136612
rect 1758 136556 1842 136612
rect 1618 136274 1842 136556
rect 1618 136222 1704 136274
rect 1756 136222 1842 136274
rect 1618 135938 1842 136222
rect 1618 135886 1704 135938
rect 1756 135886 1842 135938
rect 1618 135602 1842 135886
rect 1618 135550 1704 135602
rect 1756 135550 1842 135602
rect 1618 135266 1842 135550
rect 1618 135214 1704 135266
rect 1756 135214 1842 135266
rect 1618 134932 1842 135214
rect 1618 134876 1702 134932
rect 1758 134876 1842 134932
rect 1618 134594 1842 134876
rect 1618 134542 1704 134594
rect 1756 134542 1842 134594
rect 1618 134258 1842 134542
rect 1618 134206 1704 134258
rect 1756 134206 1842 134258
rect 1618 133922 1842 134206
rect 1618 133870 1704 133922
rect 1756 133870 1842 133922
rect 1618 133586 1842 133870
rect 1618 133534 1704 133586
rect 1756 133534 1842 133586
rect 1618 133252 1842 133534
rect 1618 133196 1702 133252
rect 1758 133196 1842 133252
rect 1618 132914 1842 133196
rect 203414 134662 203442 141663
rect 216824 141652 217048 141934
rect 216824 141596 216908 141652
rect 216964 141596 217048 141652
rect 216824 141314 217048 141596
rect 216824 141262 216910 141314
rect 216962 141262 217048 141314
rect 216824 140978 217048 141262
rect 216824 140926 216910 140978
rect 216962 140926 217048 140978
rect 216824 140642 217048 140926
rect 216824 140590 216910 140642
rect 216962 140590 217048 140642
rect 216824 140306 217048 140590
rect 216824 140254 216910 140306
rect 216962 140254 217048 140306
rect 216824 139972 217048 140254
rect 216824 139916 216908 139972
rect 216964 139916 217048 139972
rect 216824 139634 217048 139916
rect 216824 139582 216910 139634
rect 216962 139582 217048 139634
rect 216824 139298 217048 139582
rect 216824 139246 216910 139298
rect 216962 139246 217048 139298
rect 216824 138962 217048 139246
rect 216824 138910 216910 138962
rect 216962 138910 217048 138962
rect 216824 138626 217048 138910
rect 216824 138574 216910 138626
rect 216962 138574 217048 138626
rect 216824 138292 217048 138574
rect 216824 138236 216908 138292
rect 216964 138236 217048 138292
rect 216824 137954 217048 138236
rect 216824 137902 216910 137954
rect 216962 137902 217048 137954
rect 216824 137618 217048 137902
rect 216824 137566 216910 137618
rect 216962 137566 217048 137618
rect 216824 137282 217048 137566
rect 216824 137230 216910 137282
rect 216962 137230 217048 137282
rect 216824 136946 217048 137230
rect 216824 136894 216910 136946
rect 216962 136894 217048 136946
rect 216824 136612 217048 136894
rect 216824 136556 216908 136612
rect 216964 136556 217048 136612
rect 216824 136274 217048 136556
rect 216824 136222 216910 136274
rect 216962 136222 217048 136274
rect 216824 135938 217048 136222
rect 216824 135886 216910 135938
rect 216962 135886 217048 135938
rect 216824 135602 217048 135886
rect 216824 135550 216910 135602
rect 216962 135550 217048 135602
rect 216824 135266 217048 135550
rect 216824 135214 216910 135266
rect 216962 135214 217048 135266
rect 216824 134932 217048 135214
rect 216824 134876 216908 134932
rect 216964 134876 217048 134932
rect 216284 134819 216340 134828
rect 216284 134754 216340 134763
rect 213183 134714 213239 134723
rect 203414 134634 203512 134662
rect 213183 134649 213239 134658
rect 29560 133094 29616 133103
rect 29560 133029 29616 133038
rect 34552 133094 34608 133103
rect 34552 133029 34608 133038
rect 39544 133094 39600 133103
rect 39544 133029 39600 133038
rect 44536 133094 44592 133103
rect 44536 133029 44592 133038
rect 49528 133094 49584 133103
rect 49528 133029 49584 133038
rect 54520 133094 54576 133103
rect 54520 133029 54576 133038
rect 59512 133094 59568 133103
rect 59512 133029 59568 133038
rect 64504 133094 64560 133103
rect 64504 133029 64560 133038
rect 69496 133094 69552 133103
rect 69496 133029 69552 133038
rect 74488 133094 74544 133103
rect 74488 133029 74544 133038
rect 79480 133094 79536 133103
rect 79480 133029 79536 133038
rect 84472 133094 84528 133103
rect 84472 133029 84528 133038
rect 89464 133094 89520 133103
rect 89464 133029 89520 133038
rect 94456 133094 94512 133103
rect 94456 133029 94512 133038
rect 99448 133094 99504 133103
rect 99448 133029 99504 133038
rect 104440 133094 104496 133103
rect 104440 133029 104496 133038
rect 109432 133094 109488 133103
rect 109432 133029 109488 133038
rect 114424 133094 114480 133103
rect 114424 133029 114480 133038
rect 119416 133094 119472 133103
rect 119416 133029 119472 133038
rect 124408 133094 124464 133103
rect 124408 133029 124464 133038
rect 129400 133094 129456 133103
rect 129400 133029 129456 133038
rect 134392 133094 134448 133103
rect 134392 133029 134448 133038
rect 139384 133094 139440 133103
rect 139384 133029 139440 133038
rect 144376 133094 144432 133103
rect 144376 133029 144432 133038
rect 149368 133094 149424 133103
rect 149368 133029 149424 133038
rect 154360 133094 154416 133103
rect 154360 133029 154416 133038
rect 159352 133094 159408 133103
rect 159352 133029 159408 133038
rect 164344 133094 164400 133103
rect 164344 133029 164400 133038
rect 169336 133094 169392 133103
rect 169336 133029 169392 133038
rect 174328 133094 174384 133103
rect 174328 133029 174384 133038
rect 179320 133094 179376 133103
rect 179320 133029 179376 133038
rect 184312 133094 184368 133103
rect 184312 133029 184368 133038
rect 1618 132862 1704 132914
rect 1756 132862 1842 132914
rect 1618 132578 1842 132862
rect 1618 132526 1704 132578
rect 1756 132526 1842 132578
rect 1618 132242 1842 132526
rect 1618 132190 1704 132242
rect 1756 132190 1842 132242
rect 1618 131906 1842 132190
rect 1618 131854 1704 131906
rect 1756 131854 1842 131906
rect 1618 131572 1842 131854
rect 1618 131516 1702 131572
rect 1758 131516 1842 131572
rect 1618 131234 1842 131516
rect 1618 131182 1704 131234
rect 1756 131182 1842 131234
rect 1618 130898 1842 131182
rect 1618 130846 1704 130898
rect 1756 130846 1842 130898
rect 1618 130562 1842 130846
rect 1618 130510 1704 130562
rect 1756 130510 1842 130562
rect 1618 130226 1842 130510
rect 190875 130434 190931 130443
rect 190875 130369 190931 130378
rect 1618 130174 1704 130226
rect 1756 130174 1842 130226
rect 1618 129892 1842 130174
rect 1618 129836 1702 129892
rect 1758 129836 1842 129892
rect 1618 129554 1842 129836
rect 1618 129502 1704 129554
rect 1756 129502 1842 129554
rect 1618 129218 1842 129502
rect 1618 129166 1704 129218
rect 1756 129166 1842 129218
rect 1618 128882 1842 129166
rect 1618 128830 1704 128882
rect 1756 128830 1842 128882
rect 1618 128546 1842 128830
rect 1618 128494 1704 128546
rect 1756 128494 1842 128546
rect 1618 128212 1842 128494
rect 1618 128156 1702 128212
rect 1758 128156 1842 128212
rect 1618 127874 1842 128156
rect 1618 127822 1704 127874
rect 1756 127822 1842 127874
rect 1618 127538 1842 127822
rect 1618 127486 1704 127538
rect 1756 127486 1842 127538
rect 1618 127202 1842 127486
rect 1618 127150 1704 127202
rect 1756 127150 1842 127202
rect 1618 126866 1842 127150
rect 1618 126814 1704 126866
rect 1756 126814 1842 126866
rect 1618 126532 1842 126814
rect 190889 126733 190917 130369
rect 190999 129020 191055 129029
rect 190999 128955 191055 128964
rect 191013 126733 191041 128955
rect 194858 127606 194914 127615
rect 194858 127541 194914 127550
rect 1618 126476 1702 126532
rect 1758 126476 1842 126532
rect 1618 126194 1842 126476
rect 194872 126256 194900 127541
rect 1618 126142 1704 126194
rect 1756 126142 1842 126194
rect 1618 125858 1842 126142
rect 1618 125806 1704 125858
rect 1756 125806 1842 125858
rect 1618 125522 1842 125806
rect 1618 125470 1704 125522
rect 1756 125470 1842 125522
rect 1618 125186 1842 125470
rect 1618 125134 1704 125186
rect 1756 125134 1842 125186
rect 1618 124852 1842 125134
rect 1618 124796 1702 124852
rect 1758 124796 1842 124852
rect 1618 124514 1842 124796
rect 1618 124462 1704 124514
rect 1756 124462 1842 124514
rect 1618 124178 1842 124462
rect 1618 124126 1704 124178
rect 1756 124126 1842 124178
rect 1618 123842 1842 124126
rect 1618 123790 1704 123842
rect 1756 123790 1842 123842
rect 1618 123506 1842 123790
rect 1618 123454 1704 123506
rect 1756 123454 1842 123506
rect 1618 123172 1842 123454
rect 1618 123116 1702 123172
rect 1758 123116 1842 123172
rect 1618 122834 1842 123116
rect 1618 122782 1704 122834
rect 1756 122782 1842 122834
rect 1618 122498 1842 122782
rect 1618 122446 1704 122498
rect 1756 122446 1842 122498
rect 1618 122162 1842 122446
rect 1618 122110 1704 122162
rect 1756 122110 1842 122162
rect 1618 121826 1842 122110
rect 1618 121774 1704 121826
rect 1756 121774 1842 121826
rect 1618 121492 1842 121774
rect 1618 121436 1702 121492
rect 1758 121436 1842 121492
rect 1618 121154 1842 121436
rect 1618 121102 1704 121154
rect 1756 121102 1842 121154
rect 1618 120818 1842 121102
rect 1618 120766 1704 120818
rect 1756 120766 1842 120818
rect 1618 120482 1842 120766
rect 1618 120430 1704 120482
rect 1756 120430 1842 120482
rect 1618 120146 1842 120430
rect 1618 120094 1704 120146
rect 1756 120094 1842 120146
rect 1618 119812 1842 120094
rect 1618 119756 1702 119812
rect 1758 119756 1842 119812
rect 1618 119474 1842 119756
rect 1618 119422 1704 119474
rect 1756 119422 1842 119474
rect 1618 119138 1842 119422
rect 1618 119086 1704 119138
rect 1756 119086 1842 119138
rect 1618 118802 1842 119086
rect 1618 118750 1704 118802
rect 1756 118750 1842 118802
rect 1618 118466 1842 118750
rect 1618 118414 1704 118466
rect 1756 118414 1842 118466
rect 1618 118132 1842 118414
rect 1618 118076 1702 118132
rect 1758 118076 1842 118132
rect 1618 117794 1842 118076
rect 1618 117742 1704 117794
rect 1756 117742 1842 117794
rect 1618 117458 1842 117742
rect 1618 117406 1704 117458
rect 1756 117406 1842 117458
rect 1618 117122 1842 117406
rect 1618 117070 1704 117122
rect 1756 117070 1842 117122
rect 1618 116786 1842 117070
rect 1618 116734 1704 116786
rect 1756 116734 1842 116786
rect 1618 116452 1842 116734
rect 1618 116396 1702 116452
rect 1758 116396 1842 116452
rect 1618 116114 1842 116396
rect 1618 116062 1704 116114
rect 1756 116062 1842 116114
rect 1618 115778 1842 116062
rect 1618 115726 1704 115778
rect 1756 115726 1842 115778
rect 1618 115442 1842 115726
rect 1618 115390 1704 115442
rect 1756 115390 1842 115442
rect 1618 115106 1842 115390
rect 1618 115054 1704 115106
rect 1756 115054 1842 115106
rect 1618 114772 1842 115054
rect 1618 114716 1702 114772
rect 1758 114716 1842 114772
rect 1618 114434 1842 114716
rect 1618 114382 1704 114434
rect 1756 114382 1842 114434
rect 1618 114098 1842 114382
rect 1618 114046 1704 114098
rect 1756 114046 1842 114098
rect 1618 113762 1842 114046
rect 1618 113710 1704 113762
rect 1756 113710 1842 113762
rect 1618 113426 1842 113710
rect 1618 113374 1704 113426
rect 1756 113374 1842 113426
rect 1618 113092 1842 113374
rect 1618 113036 1702 113092
rect 1758 113036 1842 113092
rect 1618 112754 1842 113036
rect 1618 112702 1704 112754
rect 1756 112702 1842 112754
rect 1618 112418 1842 112702
rect 1618 112366 1704 112418
rect 1756 112366 1842 112418
rect 1618 112082 1842 112366
rect 1618 112030 1704 112082
rect 1756 112030 1842 112082
rect 1618 111746 1842 112030
rect 1618 111694 1704 111746
rect 1756 111694 1842 111746
rect 1618 111412 1842 111694
rect 1618 111356 1702 111412
rect 1758 111356 1842 111412
rect 1618 111074 1842 111356
rect 1618 111022 1704 111074
rect 1756 111022 1842 111074
rect 1618 110738 1842 111022
rect 1618 110686 1704 110738
rect 1756 110686 1842 110738
rect 1618 110402 1842 110686
rect 1618 110350 1704 110402
rect 1756 110350 1842 110402
rect 1618 110066 1842 110350
rect 1618 110014 1704 110066
rect 1756 110014 1842 110066
rect 1618 109732 1842 110014
rect 1618 109676 1702 109732
rect 1758 109676 1842 109732
rect 1618 109394 1842 109676
rect 1618 109342 1704 109394
rect 1756 109342 1842 109394
rect 1618 109058 1842 109342
rect 1618 109006 1704 109058
rect 1756 109006 1842 109058
rect 1618 108722 1842 109006
rect 1618 108670 1704 108722
rect 1756 108670 1842 108722
rect 1618 108386 1842 108670
rect 1618 108334 1704 108386
rect 1756 108334 1842 108386
rect 1618 108052 1842 108334
rect 1618 107996 1702 108052
rect 1758 107996 1842 108052
rect 1618 107714 1842 107996
rect 1618 107662 1704 107714
rect 1756 107662 1842 107714
rect 1618 107378 1842 107662
rect 1618 107326 1704 107378
rect 1756 107326 1842 107378
rect 1618 107042 1842 107326
rect 1618 106990 1704 107042
rect 1756 106990 1842 107042
rect 1618 106706 1842 106990
rect 1618 106654 1704 106706
rect 1756 106654 1842 106706
rect 1618 106372 1842 106654
rect 1618 106316 1702 106372
rect 1758 106316 1842 106372
rect 1618 106034 1842 106316
rect 1618 105982 1704 106034
rect 1756 105982 1842 106034
rect 1618 105698 1842 105982
rect 1618 105646 1704 105698
rect 1756 105646 1842 105698
rect 1618 105362 1842 105646
rect 1618 105310 1704 105362
rect 1756 105310 1842 105362
rect 1618 105026 1842 105310
rect 1618 104974 1704 105026
rect 1756 104974 1842 105026
rect 1618 104692 1842 104974
rect 1618 104636 1702 104692
rect 1758 104636 1842 104692
rect 1618 104354 1842 104636
rect 1618 104302 1704 104354
rect 1756 104302 1842 104354
rect 1618 104018 1842 104302
rect 1618 103966 1704 104018
rect 1756 103966 1842 104018
rect 1618 103682 1842 103966
rect 1618 103630 1704 103682
rect 1756 103630 1842 103682
rect 1618 103346 1842 103630
rect 1618 103294 1704 103346
rect 1756 103294 1842 103346
rect 1618 103012 1842 103294
rect 1618 102956 1702 103012
rect 1758 102956 1842 103012
rect 1618 102674 1842 102956
rect 1618 102622 1704 102674
rect 1756 102622 1842 102674
rect 1618 102338 1842 102622
rect 1618 102286 1704 102338
rect 1756 102286 1842 102338
rect 1618 102002 1842 102286
rect 1618 101950 1704 102002
rect 1756 101950 1842 102002
rect 1618 101666 1842 101950
rect 1618 101614 1704 101666
rect 1756 101614 1842 101666
rect 1618 101332 1842 101614
rect 1618 101276 1702 101332
rect 1758 101276 1842 101332
rect 1618 100994 1842 101276
rect 1618 100942 1704 100994
rect 1756 100942 1842 100994
rect 1618 100658 1842 100942
rect 1618 100606 1704 100658
rect 1756 100606 1842 100658
rect 1618 100322 1842 100606
rect 1618 100270 1704 100322
rect 1756 100270 1842 100322
rect 1618 99986 1842 100270
rect 1618 99934 1704 99986
rect 1756 99934 1842 99986
rect 1618 99652 1842 99934
rect 1618 99596 1702 99652
rect 1758 99596 1842 99652
rect 1618 99314 1842 99596
rect 1618 99262 1704 99314
rect 1756 99262 1842 99314
rect 1618 98978 1842 99262
rect 1618 98926 1704 98978
rect 1756 98926 1842 98978
rect 1618 98642 1842 98926
rect 1618 98590 1704 98642
rect 1756 98590 1842 98642
rect 1618 98306 1842 98590
rect 1618 98254 1704 98306
rect 1756 98254 1842 98306
rect 1618 97972 1842 98254
rect 1618 97916 1702 97972
rect 1758 97916 1842 97972
rect 1618 97634 1842 97916
rect 1618 97582 1704 97634
rect 1756 97582 1842 97634
rect 1618 97298 1842 97582
rect 1618 97246 1704 97298
rect 1756 97246 1842 97298
rect 1618 96962 1842 97246
rect 1618 96910 1704 96962
rect 1756 96910 1842 96962
rect 1618 96626 1842 96910
rect 1618 96574 1704 96626
rect 1756 96574 1842 96626
rect 1618 96292 1842 96574
rect 1618 96236 1702 96292
rect 1758 96236 1842 96292
rect 1618 95954 1842 96236
rect 1618 95902 1704 95954
rect 1756 95902 1842 95954
rect 1618 95618 1842 95902
rect 1618 95566 1704 95618
rect 1756 95566 1842 95618
rect 1618 95282 1842 95566
rect 1618 95230 1704 95282
rect 1756 95230 1842 95282
rect 1618 94946 1842 95230
rect 1618 94894 1704 94946
rect 1756 94894 1842 94946
rect 1618 94612 1842 94894
rect 1618 94556 1702 94612
rect 1758 94556 1842 94612
rect 1618 94274 1842 94556
rect 1618 94222 1704 94274
rect 1756 94222 1842 94274
rect 1618 93938 1842 94222
rect 1618 93886 1704 93938
rect 1756 93886 1842 93938
rect 1618 93602 1842 93886
rect 1618 93550 1704 93602
rect 1756 93550 1842 93602
rect 1618 93266 1842 93550
rect 1618 93214 1704 93266
rect 1756 93214 1842 93266
rect 1618 92932 1842 93214
rect 1618 92876 1702 92932
rect 1758 92876 1842 92932
rect 1618 92594 1842 92876
rect 1618 92542 1704 92594
rect 1756 92542 1842 92594
rect 1618 92258 1842 92542
rect 1618 92206 1704 92258
rect 1756 92206 1842 92258
rect 1618 91922 1842 92206
rect 1618 91870 1704 91922
rect 1756 91870 1842 91922
rect 1618 91586 1842 91870
rect 1618 91534 1704 91586
rect 1756 91534 1842 91586
rect 1618 91252 1842 91534
rect 1618 91196 1702 91252
rect 1758 91196 1842 91252
rect 1618 90914 1842 91196
rect 1618 90862 1704 90914
rect 1756 90862 1842 90914
rect 1618 90578 1842 90862
rect 1618 90526 1704 90578
rect 1756 90526 1842 90578
rect 1618 90242 1842 90526
rect 1618 90190 1704 90242
rect 1756 90190 1842 90242
rect 1618 89906 1842 90190
rect 1618 89854 1704 89906
rect 1756 89854 1842 89906
rect 1618 89572 1842 89854
rect 1618 89516 1702 89572
rect 1758 89516 1842 89572
rect 1618 89234 1842 89516
rect 1618 89182 1704 89234
rect 1756 89182 1842 89234
rect 1618 88898 1842 89182
rect 1618 88846 1704 88898
rect 1756 88846 1842 88898
rect 1618 88562 1842 88846
rect 1618 88510 1704 88562
rect 1756 88510 1842 88562
rect 1618 88226 1842 88510
rect 1618 88174 1704 88226
rect 1756 88174 1842 88226
rect 1618 87892 1842 88174
rect 1618 87836 1702 87892
rect 1758 87836 1842 87892
rect 1618 87554 1842 87836
rect 1618 87502 1704 87554
rect 1756 87502 1842 87554
rect 1618 87218 1842 87502
rect 1618 87166 1704 87218
rect 1756 87166 1842 87218
rect 1618 86882 1842 87166
rect 1618 86830 1704 86882
rect 1756 86830 1842 86882
rect 1618 86546 1842 86830
rect 1618 86494 1704 86546
rect 1756 86494 1842 86546
rect 1618 86212 1842 86494
rect 1618 86156 1702 86212
rect 1758 86156 1842 86212
rect 1618 85874 1842 86156
rect 1618 85822 1704 85874
rect 1756 85822 1842 85874
rect 1618 85538 1842 85822
rect 1618 85486 1704 85538
rect 1756 85486 1842 85538
rect 1618 85202 1842 85486
rect 1618 85150 1704 85202
rect 1756 85150 1842 85202
rect 1618 84866 1842 85150
rect 1618 84814 1704 84866
rect 1756 84814 1842 84866
rect 1618 84532 1842 84814
rect 1618 84476 1702 84532
rect 1758 84476 1842 84532
rect 1618 84194 1842 84476
rect 1618 84142 1704 84194
rect 1756 84142 1842 84194
rect 1618 83858 1842 84142
rect 1618 83806 1704 83858
rect 1756 83806 1842 83858
rect 1618 83522 1842 83806
rect 1618 83470 1704 83522
rect 1756 83470 1842 83522
rect 1618 83186 1842 83470
rect 1618 83134 1704 83186
rect 1756 83134 1842 83186
rect 1618 82852 1842 83134
rect 1618 82796 1702 82852
rect 1758 82796 1842 82852
rect 1618 82514 1842 82796
rect 1618 82462 1704 82514
rect 1756 82462 1842 82514
rect 1618 82178 1842 82462
rect 1618 82126 1704 82178
rect 1756 82126 1842 82178
rect 1618 81842 1842 82126
rect 1618 81790 1704 81842
rect 1756 81790 1842 81842
rect 1618 81506 1842 81790
rect 1618 81454 1704 81506
rect 1756 81454 1842 81506
rect 1618 81172 1842 81454
rect 1618 81116 1702 81172
rect 1758 81116 1842 81172
rect 1618 80834 1842 81116
rect 1618 80782 1704 80834
rect 1756 80782 1842 80834
rect 1618 80498 1842 80782
rect 1618 80446 1704 80498
rect 1756 80446 1842 80498
rect 1618 80162 1842 80446
rect 1618 80110 1704 80162
rect 1756 80110 1842 80162
rect 1618 79826 1842 80110
rect 1618 79774 1704 79826
rect 1756 79774 1842 79826
rect 1618 79492 1842 79774
rect 1618 79436 1702 79492
rect 1758 79436 1842 79492
rect 1618 79154 1842 79436
rect 1618 79102 1704 79154
rect 1756 79102 1842 79154
rect 1618 78818 1842 79102
rect 1618 78766 1704 78818
rect 1756 78766 1842 78818
rect 1618 78482 1842 78766
rect 1618 78430 1704 78482
rect 1756 78430 1842 78482
rect 1618 78146 1842 78430
rect 1618 78094 1704 78146
rect 1756 78094 1842 78146
rect 1618 77812 1842 78094
rect 1618 77756 1702 77812
rect 1758 77756 1842 77812
rect 1618 77474 1842 77756
rect 1618 77422 1704 77474
rect 1756 77422 1842 77474
rect 1618 77138 1842 77422
rect 1618 77086 1704 77138
rect 1756 77086 1842 77138
rect 1618 76802 1842 77086
rect 1618 76750 1704 76802
rect 1756 76750 1842 76802
rect 1618 76466 1842 76750
rect 1618 76414 1704 76466
rect 1756 76414 1842 76466
rect 1618 76132 1842 76414
rect 1618 76076 1702 76132
rect 1758 76076 1842 76132
rect 1618 75794 1842 76076
rect 1618 75742 1704 75794
rect 1756 75742 1842 75794
rect 1618 75458 1842 75742
rect 1618 75406 1704 75458
rect 1756 75406 1842 75458
rect 1618 75122 1842 75406
rect 1618 75070 1704 75122
rect 1756 75070 1842 75122
rect 1618 74786 1842 75070
rect 1618 74734 1704 74786
rect 1756 74734 1842 74786
rect 1618 74452 1842 74734
rect 1618 74396 1702 74452
rect 1758 74396 1842 74452
rect 1618 74114 1842 74396
rect 1618 74062 1704 74114
rect 1756 74062 1842 74114
rect 1618 73778 1842 74062
rect 1618 73726 1704 73778
rect 1756 73726 1842 73778
rect 1618 73442 1842 73726
rect 1618 73390 1704 73442
rect 1756 73390 1842 73442
rect 1618 73106 1842 73390
rect 1618 73054 1704 73106
rect 1756 73054 1842 73106
rect 1618 72772 1842 73054
rect 1618 72716 1702 72772
rect 1758 72716 1842 72772
rect 1618 72434 1842 72716
rect 1618 72382 1704 72434
rect 1756 72382 1842 72434
rect 1618 72098 1842 72382
rect 1618 72046 1704 72098
rect 1756 72046 1842 72098
rect 1618 71762 1842 72046
rect 1618 71710 1704 71762
rect 1756 71710 1842 71762
rect 1618 71426 1842 71710
rect 1618 71374 1704 71426
rect 1756 71374 1842 71426
rect 1618 71092 1842 71374
rect 1618 71036 1702 71092
rect 1758 71036 1842 71092
rect 1618 70754 1842 71036
rect 1618 70702 1704 70754
rect 1756 70702 1842 70754
rect 1618 70418 1842 70702
rect 1618 70366 1704 70418
rect 1756 70366 1842 70418
rect 1618 70082 1842 70366
rect 1618 70030 1704 70082
rect 1756 70030 1842 70082
rect 1618 69746 1842 70030
rect 1618 69694 1704 69746
rect 1756 69694 1842 69746
rect 1618 69412 1842 69694
rect 1618 69356 1702 69412
rect 1758 69356 1842 69412
rect 1618 69074 1842 69356
rect 1618 69022 1704 69074
rect 1756 69022 1842 69074
rect 1618 68738 1842 69022
rect 1618 68686 1704 68738
rect 1756 68686 1842 68738
rect 1618 68402 1842 68686
rect 1618 68350 1704 68402
rect 1756 68350 1842 68402
rect 1618 68066 1842 68350
rect 1618 68014 1704 68066
rect 1756 68014 1842 68066
rect 1618 67732 1842 68014
rect 1618 67676 1702 67732
rect 1758 67676 1842 67732
rect 1618 67394 1842 67676
rect 1618 67342 1704 67394
rect 1756 67342 1842 67394
rect 1618 67058 1842 67342
rect 1618 67006 1704 67058
rect 1756 67006 1842 67058
rect 1618 66722 1842 67006
rect 1618 66670 1704 66722
rect 1756 66670 1842 66722
rect 1618 66386 1842 66670
rect 1618 66334 1704 66386
rect 1756 66334 1842 66386
rect 1618 66052 1842 66334
rect 1618 65996 1702 66052
rect 1758 65996 1842 66052
rect 1618 65714 1842 65996
rect 1618 65662 1704 65714
rect 1756 65662 1842 65714
rect 1618 65378 1842 65662
rect 1618 65326 1704 65378
rect 1756 65326 1842 65378
rect 1618 65042 1842 65326
rect 1618 64990 1704 65042
rect 1756 64990 1842 65042
rect 1618 64706 1842 64990
rect 1618 64654 1704 64706
rect 1756 64654 1842 64706
rect 1618 64372 1842 64654
rect 1618 64316 1702 64372
rect 1758 64316 1842 64372
rect 1618 64034 1842 64316
rect 1618 63982 1704 64034
rect 1756 63982 1842 64034
rect 1618 63698 1842 63982
rect 1618 63646 1704 63698
rect 1756 63646 1842 63698
rect 1618 63362 1842 63646
rect 1618 63310 1704 63362
rect 1756 63310 1842 63362
rect 1618 63026 1842 63310
rect 1618 62974 1704 63026
rect 1756 62974 1842 63026
rect 1618 62692 1842 62974
rect 1618 62636 1702 62692
rect 1758 62636 1842 62692
rect 1618 62354 1842 62636
rect 1618 62302 1704 62354
rect 1756 62302 1842 62354
rect 1618 62018 1842 62302
rect 1618 61966 1704 62018
rect 1756 61966 1842 62018
rect 1618 61682 1842 61966
rect 1618 61630 1704 61682
rect 1756 61630 1842 61682
rect 1618 61346 1842 61630
rect 1618 61294 1704 61346
rect 1756 61294 1842 61346
rect 1618 61012 1842 61294
rect 1618 60956 1702 61012
rect 1758 60956 1842 61012
rect 1618 60674 1842 60956
rect 1618 60622 1704 60674
rect 1756 60622 1842 60674
rect 1618 60338 1842 60622
rect 1618 60286 1704 60338
rect 1756 60286 1842 60338
rect 1618 60002 1842 60286
rect 1618 59950 1704 60002
rect 1756 59950 1842 60002
rect 1618 59666 1842 59950
rect 1618 59614 1704 59666
rect 1756 59614 1842 59666
rect 1618 59332 1842 59614
rect 1618 59276 1702 59332
rect 1758 59276 1842 59332
rect 1618 58994 1842 59276
rect 1618 58942 1704 58994
rect 1756 58942 1842 58994
rect 1618 58658 1842 58942
rect 1618 58606 1704 58658
rect 1756 58606 1842 58658
rect 1618 58322 1842 58606
rect 1618 58270 1704 58322
rect 1756 58270 1842 58322
rect 1618 57986 1842 58270
rect 1618 57934 1704 57986
rect 1756 57934 1842 57986
rect 1618 57652 1842 57934
rect 1618 57596 1702 57652
rect 1758 57596 1842 57652
rect 1618 57314 1842 57596
rect 1618 57262 1704 57314
rect 1756 57262 1842 57314
rect 1618 56978 1842 57262
rect 1618 56926 1704 56978
rect 1756 56926 1842 56978
rect 1618 56642 1842 56926
rect 1618 56590 1704 56642
rect 1756 56590 1842 56642
rect 1618 56306 1842 56590
rect 1618 56254 1704 56306
rect 1756 56254 1842 56306
rect 1618 55972 1842 56254
rect 1618 55916 1702 55972
rect 1758 55916 1842 55972
rect 1618 55634 1842 55916
rect 1618 55582 1704 55634
rect 1756 55582 1842 55634
rect 1618 55298 1842 55582
rect 1618 55246 1704 55298
rect 1756 55246 1842 55298
rect 1618 54962 1842 55246
rect 1618 54910 1704 54962
rect 1756 54910 1842 54962
rect 1618 54626 1842 54910
rect 1618 54574 1704 54626
rect 1756 54574 1842 54626
rect 1618 54292 1842 54574
rect 1618 54236 1702 54292
rect 1758 54236 1842 54292
rect 1618 53954 1842 54236
rect 1618 53902 1704 53954
rect 1756 53902 1842 53954
rect 1618 53618 1842 53902
rect 1618 53566 1704 53618
rect 1756 53566 1842 53618
rect 1618 53282 1842 53566
rect 1618 53230 1704 53282
rect 1756 53230 1842 53282
rect 1618 52946 1842 53230
rect 1618 52894 1704 52946
rect 1756 52894 1842 52946
rect 1618 52612 1842 52894
rect 1618 52556 1702 52612
rect 1758 52556 1842 52612
rect 1618 52274 1842 52556
rect 1618 52222 1704 52274
rect 1756 52222 1842 52274
rect 1618 51938 1842 52222
rect 1618 51886 1704 51938
rect 1756 51886 1842 51938
rect 1618 51602 1842 51886
rect 1618 51550 1704 51602
rect 1756 51550 1842 51602
rect 1618 51266 1842 51550
rect 1618 51214 1704 51266
rect 1756 51214 1842 51266
rect 1618 50932 1842 51214
rect 1618 50876 1702 50932
rect 1758 50876 1842 50932
rect 1618 50594 1842 50876
rect 1618 50542 1704 50594
rect 1756 50542 1842 50594
rect 1618 50258 1842 50542
rect 1618 50206 1704 50258
rect 1756 50206 1842 50258
rect 1618 49922 1842 50206
rect 1618 49870 1704 49922
rect 1756 49870 1842 49922
rect 1618 49586 1842 49870
rect 1618 49534 1704 49586
rect 1756 49534 1842 49586
rect 1618 49252 1842 49534
rect 1618 49196 1702 49252
rect 1758 49196 1842 49252
rect 1618 48914 1842 49196
rect 1618 48862 1704 48914
rect 1756 48862 1842 48914
rect 1618 48578 1842 48862
rect 1618 48526 1704 48578
rect 1756 48526 1842 48578
rect 1618 48242 1842 48526
rect 1618 48190 1704 48242
rect 1756 48190 1842 48242
rect 1618 47906 1842 48190
rect 1618 47854 1704 47906
rect 1756 47854 1842 47906
rect 1618 47572 1842 47854
rect 1618 47516 1702 47572
rect 1758 47516 1842 47572
rect 1618 47234 1842 47516
rect 1618 47182 1704 47234
rect 1756 47182 1842 47234
rect 1618 46898 1842 47182
rect 1618 46846 1704 46898
rect 1756 46846 1842 46898
rect 1618 46562 1842 46846
rect 1618 46510 1704 46562
rect 1756 46510 1842 46562
rect 1618 46226 1842 46510
rect 1618 46174 1704 46226
rect 1756 46174 1842 46226
rect 1618 45892 1842 46174
rect 1618 45836 1702 45892
rect 1758 45836 1842 45892
rect 1618 45554 1842 45836
rect 1618 45502 1704 45554
rect 1756 45502 1842 45554
rect 1618 45218 1842 45502
rect 1618 45166 1704 45218
rect 1756 45166 1842 45218
rect 1618 44882 1842 45166
rect 14212 45093 14268 45102
rect 14212 45028 14268 45037
rect 15157 45022 15213 45031
rect 15157 44957 15213 44966
rect 15971 45022 16027 45031
rect 15971 44957 16027 44966
rect 1618 44830 1704 44882
rect 1756 44830 1842 44882
rect 1618 44546 1842 44830
rect 1618 44494 1704 44546
rect 1756 44494 1842 44546
rect 1618 44212 1842 44494
rect 1618 44156 1702 44212
rect 1758 44156 1842 44212
rect 1618 43874 1842 44156
rect 1618 43822 1704 43874
rect 1756 43822 1842 43874
rect 1618 43538 1842 43822
rect 1618 43486 1704 43538
rect 1756 43486 1842 43538
rect 1618 43202 1842 43486
rect 15157 43464 15213 43473
rect 14212 43393 14268 43402
rect 15157 43399 15213 43408
rect 15891 43464 15947 43473
rect 15891 43399 15947 43408
rect 14212 43328 14268 43337
rect 1618 43150 1704 43202
rect 1756 43150 1842 43202
rect 1618 42866 1842 43150
rect 1618 42814 1704 42866
rect 1756 42814 1842 42866
rect 1618 42532 1842 42814
rect 1618 42476 1702 42532
rect 1758 42476 1842 42532
rect 1618 42194 1842 42476
rect 14212 42265 14268 42274
rect 14212 42200 14268 42209
rect 1618 42142 1704 42194
rect 1756 42142 1842 42194
rect 1618 41858 1842 42142
rect 15157 42194 15213 42203
rect 15157 42129 15213 42138
rect 15811 42194 15867 42203
rect 15811 42129 15867 42138
rect 1618 41806 1704 41858
rect 1756 41806 1842 41858
rect 1618 41522 1842 41806
rect 1618 41470 1704 41522
rect 1756 41470 1842 41522
rect 1618 41186 1842 41470
rect 1618 41134 1704 41186
rect 1756 41134 1842 41186
rect 1618 40852 1842 41134
rect 1618 40796 1702 40852
rect 1758 40796 1842 40852
rect 1618 40514 1842 40796
rect 15157 40636 15213 40645
rect 1618 40462 1704 40514
rect 1756 40462 1842 40514
rect 14212 40565 14268 40574
rect 15157 40571 15213 40580
rect 15731 40636 15787 40645
rect 15731 40571 15787 40580
rect 14212 40500 14268 40509
rect 1618 40178 1842 40462
rect 1618 40126 1704 40178
rect 1756 40126 1842 40178
rect 1618 39842 1842 40126
rect 1618 39790 1704 39842
rect 1756 39790 1842 39842
rect 1618 39506 1842 39790
rect 1618 39454 1704 39506
rect 1756 39454 1842 39506
rect 1618 39172 1842 39454
rect 14212 39437 14268 39446
rect 14212 39372 14268 39381
rect 15157 39366 15213 39375
rect 15157 39301 15213 39310
rect 15651 39366 15707 39375
rect 15651 39301 15707 39310
rect 1618 39116 1702 39172
rect 1758 39116 1842 39172
rect 1618 38834 1842 39116
rect 1618 38782 1704 38834
rect 1756 38782 1842 38834
rect 1618 38498 1842 38782
rect 1618 38446 1704 38498
rect 1756 38446 1842 38498
rect 1618 38162 1842 38446
rect 1618 38110 1704 38162
rect 1756 38110 1842 38162
rect 1618 37826 1842 38110
rect 1618 37774 1704 37826
rect 1756 37774 1842 37826
rect 1618 37492 1842 37774
rect 15157 37808 15213 37817
rect 14212 37737 14268 37746
rect 15157 37743 15213 37752
rect 15571 37808 15627 37817
rect 15571 37743 15627 37752
rect 14212 37672 14268 37681
rect 1618 37436 1702 37492
rect 1758 37436 1842 37492
rect 1618 37154 1842 37436
rect 1618 37102 1704 37154
rect 1756 37102 1842 37154
rect 1618 36818 1842 37102
rect 1618 36766 1704 36818
rect 1756 36766 1842 36818
rect 1618 36482 1842 36766
rect 14212 36609 14268 36618
rect 14212 36544 14268 36553
rect 1618 36430 1704 36482
rect 1756 36430 1842 36482
rect 15157 36538 15213 36547
rect 15157 36473 15213 36482
rect 15491 36538 15547 36547
rect 15491 36473 15547 36482
rect 1618 36146 1842 36430
rect 1618 36094 1704 36146
rect 1756 36094 1842 36146
rect 1618 35812 1842 36094
rect 1618 35756 1702 35812
rect 1758 35756 1842 35812
rect 1618 35474 1842 35756
rect 1618 35422 1704 35474
rect 1756 35422 1842 35474
rect 1618 35138 1842 35422
rect 1618 35086 1704 35138
rect 1756 35086 1842 35138
rect 1618 34802 1842 35086
rect 15157 34980 15213 34989
rect 14212 34909 14268 34918
rect 15157 34915 15213 34924
rect 15411 34980 15467 34989
rect 15411 34915 15467 34924
rect 14212 34844 14268 34853
rect 1618 34750 1704 34802
rect 1756 34750 1842 34802
rect 1618 34466 1842 34750
rect 15294 34653 15350 34662
rect 15294 34588 15350 34597
rect 1618 34414 1704 34466
rect 1756 34414 1842 34466
rect 1618 34132 1842 34414
rect 1618 34076 1702 34132
rect 1758 34076 1842 34132
rect 1618 33794 1842 34076
rect 1618 33742 1704 33794
rect 1756 33742 1842 33794
rect 1618 33458 1842 33742
rect 1618 33406 1704 33458
rect 1756 33406 1842 33458
rect 1618 33122 1842 33406
rect 1618 33070 1704 33122
rect 1756 33070 1842 33122
rect 1618 32786 1842 33070
rect 1618 32734 1704 32786
rect 1756 32734 1842 32786
rect 1618 32452 1842 32734
rect 1618 32396 1702 32452
rect 1758 32396 1842 32452
rect 1618 32114 1842 32396
rect 1618 32062 1704 32114
rect 1756 32062 1842 32114
rect 1618 31778 1842 32062
rect 1618 31726 1704 31778
rect 1756 31726 1842 31778
rect 1618 31442 1842 31726
rect 1618 31390 1704 31442
rect 1756 31390 1842 31442
rect 1618 31106 1842 31390
rect 1618 31054 1704 31106
rect 1756 31054 1842 31106
rect 1618 30772 1842 31054
rect 1618 30716 1702 30772
rect 1758 30716 1842 30772
rect 1618 30434 1842 30716
rect 1618 30382 1704 30434
rect 1756 30382 1842 30434
rect 1618 30098 1842 30382
rect 2113 30352 2169 30361
rect 2113 30287 2169 30296
rect 1618 30046 1704 30098
rect 1756 30046 1842 30098
rect 1618 29762 1842 30046
rect 1618 29710 1704 29762
rect 1756 29710 1842 29762
rect 1618 29426 1842 29710
rect 1618 29374 1704 29426
rect 1756 29374 1842 29426
rect 1618 29092 1842 29374
rect 1618 29036 1702 29092
rect 1758 29036 1842 29092
rect 1618 28754 1842 29036
rect 1618 28702 1704 28754
rect 1756 28702 1842 28754
rect 1618 28418 1842 28702
rect 1618 28366 1704 28418
rect 1756 28366 1842 28418
rect 1618 28082 1842 28366
rect 1618 28030 1704 28082
rect 1756 28030 1842 28082
rect 1618 27746 1842 28030
rect 1618 27694 1704 27746
rect 1756 27694 1842 27746
rect 1618 27412 1842 27694
rect 1618 27356 1702 27412
rect 1758 27356 1842 27412
rect 1618 27074 1842 27356
rect 1618 27022 1704 27074
rect 1756 27022 1842 27074
rect 1618 26738 1842 27022
rect 1618 26686 1704 26738
rect 1756 26686 1842 26738
rect 1618 26402 1842 26686
rect 1618 26350 1704 26402
rect 1756 26350 1842 26402
rect 1618 26066 1842 26350
rect 1618 26014 1704 26066
rect 1756 26014 1842 26066
rect 1618 25732 1842 26014
rect 1618 25676 1702 25732
rect 1758 25676 1842 25732
rect 1618 25394 1842 25676
rect 1618 25342 1704 25394
rect 1756 25342 1842 25394
rect 1618 25058 1842 25342
rect 1618 25006 1704 25058
rect 1756 25006 1842 25058
rect 1618 24722 1842 25006
rect 1618 24670 1704 24722
rect 1756 24670 1842 24722
rect 1618 24386 1842 24670
rect 1618 24334 1704 24386
rect 1756 24334 1842 24386
rect 1618 24052 1842 24334
rect 1618 23996 1702 24052
rect 1758 23996 1842 24052
rect 1618 23714 1842 23996
rect 1618 23662 1704 23714
rect 1756 23662 1842 23714
rect 1618 23378 1842 23662
rect 1618 23326 1704 23378
rect 1756 23326 1842 23378
rect 1618 23042 1842 23326
rect 15210 23244 15266 23253
rect 15210 23179 15266 23188
rect 1618 22990 1704 23042
rect 1756 22990 1842 23042
rect 1618 22706 1842 22990
rect 1618 22654 1704 22706
rect 1756 22654 1842 22706
rect 1618 22372 1842 22654
rect 1618 22316 1702 22372
rect 1758 22316 1842 22372
rect 1618 22034 1842 22316
rect 1618 21982 1704 22034
rect 1756 21982 1842 22034
rect 1618 21698 1842 21982
rect 1618 21646 1704 21698
rect 1756 21646 1842 21698
rect 1618 21362 1842 21646
rect 1618 21310 1704 21362
rect 1756 21310 1842 21362
rect 1618 21026 1842 21310
rect 1618 20974 1704 21026
rect 1756 20974 1842 21026
rect 1618 20692 1842 20974
rect 1618 20636 1702 20692
rect 1758 20636 1842 20692
rect 1618 20354 1842 20636
rect 1618 20302 1704 20354
rect 1756 20302 1842 20354
rect 15210 20416 15266 20425
rect 15210 20351 15266 20360
rect 1618 20018 1842 20302
rect 1618 19966 1704 20018
rect 1756 19966 1842 20018
rect 1618 19682 1842 19966
rect 1618 19630 1704 19682
rect 1756 19630 1842 19682
rect 1618 19346 1842 19630
rect 1618 19294 1704 19346
rect 1756 19294 1842 19346
rect 1618 19012 1842 19294
rect 1618 18956 1702 19012
rect 1758 18956 1842 19012
rect 1618 18674 1842 18956
rect 15210 19002 15266 19011
rect 15210 18937 15266 18946
rect 1618 18622 1704 18674
rect 1756 18622 1842 18674
rect 1618 18338 1842 18622
rect 1618 18286 1704 18338
rect 1756 18286 1842 18338
rect 1618 18002 1842 18286
rect 1618 17950 1704 18002
rect 1756 17950 1842 18002
rect 1618 17666 1842 17950
rect 1618 17614 1704 17666
rect 1756 17614 1842 17666
rect 1618 17332 1842 17614
rect 15210 17588 15266 17597
rect 15210 17523 15266 17532
rect 1618 17276 1702 17332
rect 1758 17276 1842 17332
rect 1618 16994 1842 17276
rect 1618 16942 1704 16994
rect 1756 16942 1842 16994
rect 1618 16658 1842 16942
rect 1618 16606 1704 16658
rect 1756 16606 1842 16658
rect 1618 16322 1842 16606
rect 1618 16270 1704 16322
rect 1756 16270 1842 16322
rect 1618 15986 1842 16270
rect 1618 15934 1704 15986
rect 1756 15934 1842 15986
rect 1618 15652 1842 15934
rect 1618 15596 1702 15652
rect 1758 15596 1842 15652
rect 1618 15314 1842 15596
rect 1618 15262 1704 15314
rect 1756 15262 1842 15314
rect 1618 14978 1842 15262
rect 1618 14926 1704 14978
rect 1756 14926 1842 14978
rect 1618 14642 1842 14926
rect 2326 14903 2382 14912
rect 2326 14838 2382 14847
rect 1618 14590 1704 14642
rect 1756 14590 1842 14642
rect 1618 14306 1842 14590
rect 1618 14254 1704 14306
rect 1756 14254 1842 14306
rect 1618 13972 1842 14254
rect 1618 13916 1702 13972
rect 1758 13916 1842 13972
rect 1618 13634 1842 13916
rect 1618 13582 1704 13634
rect 1756 13582 1842 13634
rect 1618 13298 1842 13582
rect 15308 13332 15336 34588
rect 203414 24566 203442 134634
rect 216824 134594 217048 134876
rect 216824 134542 216910 134594
rect 216962 134542 217048 134594
rect 216824 134258 217048 134542
rect 216824 134206 216910 134258
rect 216962 134206 217048 134258
rect 216824 133922 217048 134206
rect 216824 133870 216910 133922
rect 216962 133870 217048 133922
rect 216824 133586 217048 133870
rect 216824 133534 216910 133586
rect 216962 133534 217048 133586
rect 216824 133252 217048 133534
rect 216824 133196 216908 133252
rect 216964 133196 217048 133252
rect 216824 132914 217048 133196
rect 216824 132862 216910 132914
rect 216962 132862 217048 132914
rect 216824 132578 217048 132862
rect 216824 132526 216910 132578
rect 216962 132526 217048 132578
rect 216824 132242 217048 132526
rect 216824 132190 216910 132242
rect 216962 132190 217048 132242
rect 216824 131906 217048 132190
rect 216824 131854 216910 131906
rect 216962 131854 217048 131906
rect 216824 131572 217048 131854
rect 216824 131516 216908 131572
rect 216964 131516 217048 131572
rect 216824 131234 217048 131516
rect 216824 131182 216910 131234
rect 216962 131182 217048 131234
rect 216824 130898 217048 131182
rect 216824 130846 216910 130898
rect 216962 130846 217048 130898
rect 216824 130562 217048 130846
rect 216824 130510 216910 130562
rect 216962 130510 217048 130562
rect 203484 130434 203540 130443
rect 203484 130369 203540 130378
rect 216824 130226 217048 130510
rect 216824 130174 216910 130226
rect 216962 130174 217048 130226
rect 216824 129892 217048 130174
rect 216824 129836 216908 129892
rect 216964 129836 217048 129892
rect 216824 129554 217048 129836
rect 216824 129502 216910 129554
rect 216962 129502 217048 129554
rect 216824 129218 217048 129502
rect 216824 129166 216910 129218
rect 216962 129166 217048 129218
rect 203484 129020 203540 129029
rect 203484 128955 203540 128964
rect 216824 128882 217048 129166
rect 216824 128830 216910 128882
rect 216962 128830 217048 128882
rect 216824 128546 217048 128830
rect 216824 128494 216910 128546
rect 216962 128494 217048 128546
rect 216824 128212 217048 128494
rect 216824 128156 216908 128212
rect 216964 128156 217048 128212
rect 216824 127874 217048 128156
rect 216824 127822 216910 127874
rect 216962 127822 217048 127874
rect 203484 127606 203540 127615
rect 203484 127541 203540 127550
rect 216824 127538 217048 127822
rect 216824 127486 216910 127538
rect 216962 127486 217048 127538
rect 216824 127202 217048 127486
rect 216824 127150 216910 127202
rect 216962 127150 217048 127202
rect 216824 126866 217048 127150
rect 216824 126814 216910 126866
rect 216962 126814 217048 126866
rect 216824 126532 217048 126814
rect 216824 126476 216908 126532
rect 216964 126476 217048 126532
rect 216824 126194 217048 126476
rect 216824 126142 216910 126194
rect 216962 126142 217048 126194
rect 216824 125858 217048 126142
rect 216824 125806 216910 125858
rect 216962 125806 217048 125858
rect 216824 125522 217048 125806
rect 216824 125470 216910 125522
rect 216962 125470 217048 125522
rect 216824 125186 217048 125470
rect 216824 125134 216910 125186
rect 216962 125134 217048 125186
rect 216824 124852 217048 125134
rect 216824 124796 216908 124852
rect 216964 124796 217048 124852
rect 216824 124514 217048 124796
rect 216824 124462 216910 124514
rect 216962 124462 217048 124514
rect 216824 124178 217048 124462
rect 216824 124126 216910 124178
rect 216962 124126 217048 124178
rect 216824 123842 217048 124126
rect 216824 123790 216910 123842
rect 216962 123790 217048 123842
rect 216824 123506 217048 123790
rect 216824 123454 216910 123506
rect 216962 123454 217048 123506
rect 216824 123172 217048 123454
rect 216824 123116 216908 123172
rect 216964 123116 217048 123172
rect 216824 122834 217048 123116
rect 216824 122782 216910 122834
rect 216962 122782 217048 122834
rect 216824 122498 217048 122782
rect 216824 122446 216910 122498
rect 216962 122446 217048 122498
rect 216824 122162 217048 122446
rect 216824 122110 216910 122162
rect 216962 122110 217048 122162
rect 216824 121826 217048 122110
rect 216824 121774 216910 121826
rect 216962 121774 217048 121826
rect 216824 121492 217048 121774
rect 216824 121436 216908 121492
rect 216964 121436 217048 121492
rect 216824 121154 217048 121436
rect 216824 121102 216910 121154
rect 216962 121102 217048 121154
rect 216824 120818 217048 121102
rect 216824 120766 216910 120818
rect 216962 120766 217048 120818
rect 216824 120482 217048 120766
rect 216824 120430 216910 120482
rect 216962 120430 217048 120482
rect 216824 120146 217048 120430
rect 216824 120094 216910 120146
rect 216962 120094 217048 120146
rect 216824 119812 217048 120094
rect 216824 119756 216908 119812
rect 216964 119756 217048 119812
rect 216824 119474 217048 119756
rect 216824 119422 216910 119474
rect 216962 119422 217048 119474
rect 216824 119138 217048 119422
rect 216824 119086 216910 119138
rect 216962 119086 217048 119138
rect 216824 118802 217048 119086
rect 216824 118750 216910 118802
rect 216962 118750 217048 118802
rect 216824 118466 217048 118750
rect 216824 118414 216910 118466
rect 216962 118414 217048 118466
rect 216824 118132 217048 118414
rect 216824 118076 216908 118132
rect 216964 118076 217048 118132
rect 216824 117794 217048 118076
rect 216824 117742 216910 117794
rect 216962 117742 217048 117794
rect 216497 117670 216553 117679
rect 216497 117605 216553 117614
rect 216824 117458 217048 117742
rect 216824 117406 216910 117458
rect 216962 117406 217048 117458
rect 216824 117122 217048 117406
rect 216824 117070 216910 117122
rect 216962 117070 217048 117122
rect 216824 116786 217048 117070
rect 216824 116734 216910 116786
rect 216962 116734 217048 116786
rect 216824 116452 217048 116734
rect 216824 116396 216908 116452
rect 216964 116396 217048 116452
rect 216824 116114 217048 116396
rect 216824 116062 216910 116114
rect 216962 116062 217048 116114
rect 216824 115778 217048 116062
rect 216824 115726 216910 115778
rect 216962 115726 217048 115778
rect 216824 115442 217048 115726
rect 216824 115390 216910 115442
rect 216962 115390 217048 115442
rect 216824 115106 217048 115390
rect 216824 115054 216910 115106
rect 216962 115054 217048 115106
rect 216824 114772 217048 115054
rect 216824 114716 216908 114772
rect 216964 114716 217048 114772
rect 216824 114434 217048 114716
rect 216824 114382 216910 114434
rect 216962 114382 217048 114434
rect 216824 114098 217048 114382
rect 216824 114046 216910 114098
rect 216962 114046 217048 114098
rect 216824 113762 217048 114046
rect 216824 113710 216910 113762
rect 216962 113710 217048 113762
rect 216824 113426 217048 113710
rect 216824 113374 216910 113426
rect 216962 113374 217048 113426
rect 216824 113092 217048 113374
rect 216824 113036 216908 113092
rect 216964 113036 217048 113092
rect 216824 112754 217048 113036
rect 216824 112702 216910 112754
rect 216962 112702 217048 112754
rect 216824 112418 217048 112702
rect 216824 112366 216910 112418
rect 216962 112366 217048 112418
rect 216824 112082 217048 112366
rect 216824 112030 216910 112082
rect 216962 112030 217048 112082
rect 216824 111746 217048 112030
rect 216824 111694 216910 111746
rect 216962 111694 217048 111746
rect 216824 111412 217048 111694
rect 216824 111356 216908 111412
rect 216964 111356 217048 111412
rect 216824 111074 217048 111356
rect 216824 111022 216910 111074
rect 216962 111022 217048 111074
rect 216824 110738 217048 111022
rect 216824 110686 216910 110738
rect 216962 110686 217048 110738
rect 216824 110402 217048 110686
rect 216824 110350 216910 110402
rect 216962 110350 217048 110402
rect 216824 110066 217048 110350
rect 216824 110014 216910 110066
rect 216962 110014 217048 110066
rect 216824 109732 217048 110014
rect 216824 109676 216908 109732
rect 216964 109676 217048 109732
rect 216824 109394 217048 109676
rect 216824 109342 216910 109394
rect 216962 109342 217048 109394
rect 216824 109058 217048 109342
rect 216824 109006 216910 109058
rect 216962 109006 217048 109058
rect 216824 108722 217048 109006
rect 216824 108670 216910 108722
rect 216962 108670 217048 108722
rect 216824 108386 217048 108670
rect 216824 108334 216910 108386
rect 216962 108334 217048 108386
rect 216824 108052 217048 108334
rect 216824 107996 216908 108052
rect 216964 107996 217048 108052
rect 216824 107714 217048 107996
rect 216824 107662 216910 107714
rect 216962 107662 217048 107714
rect 216824 107378 217048 107662
rect 216824 107326 216910 107378
rect 216962 107326 217048 107378
rect 216824 107042 217048 107326
rect 216824 106990 216910 107042
rect 216962 106990 217048 107042
rect 216824 106706 217048 106990
rect 216824 106654 216910 106706
rect 216962 106654 217048 106706
rect 216824 106372 217048 106654
rect 216824 106316 216908 106372
rect 216964 106316 217048 106372
rect 216824 106034 217048 106316
rect 216824 105982 216910 106034
rect 216962 105982 217048 106034
rect 216824 105698 217048 105982
rect 216824 105646 216910 105698
rect 216962 105646 217048 105698
rect 216824 105362 217048 105646
rect 216824 105310 216910 105362
rect 216962 105310 217048 105362
rect 216824 105026 217048 105310
rect 216824 104974 216910 105026
rect 216962 104974 217048 105026
rect 216824 104692 217048 104974
rect 216824 104636 216908 104692
rect 216964 104636 217048 104692
rect 216824 104354 217048 104636
rect 216824 104302 216910 104354
rect 216962 104302 217048 104354
rect 216824 104018 217048 104302
rect 216824 103966 216910 104018
rect 216962 103966 217048 104018
rect 216824 103682 217048 103966
rect 216824 103630 216910 103682
rect 216962 103630 217048 103682
rect 216824 103346 217048 103630
rect 216824 103294 216910 103346
rect 216962 103294 217048 103346
rect 216824 103012 217048 103294
rect 216824 102956 216908 103012
rect 216964 102956 217048 103012
rect 216824 102674 217048 102956
rect 216824 102622 216910 102674
rect 216962 102622 217048 102674
rect 216824 102338 217048 102622
rect 216824 102286 216910 102338
rect 216962 102286 217048 102338
rect 216824 102002 217048 102286
rect 216824 101950 216910 102002
rect 216962 101950 217048 102002
rect 216824 101666 217048 101950
rect 216824 101614 216910 101666
rect 216962 101614 217048 101666
rect 216824 101332 217048 101614
rect 216824 101276 216908 101332
rect 216964 101276 217048 101332
rect 216824 100994 217048 101276
rect 216824 100942 216910 100994
rect 216962 100942 217048 100994
rect 216824 100658 217048 100942
rect 216824 100606 216910 100658
rect 216962 100606 217048 100658
rect 216824 100322 217048 100606
rect 216824 100270 216910 100322
rect 216962 100270 217048 100322
rect 216824 99986 217048 100270
rect 216824 99934 216910 99986
rect 216962 99934 217048 99986
rect 216824 99652 217048 99934
rect 216824 99596 216908 99652
rect 216964 99596 217048 99652
rect 216824 99314 217048 99596
rect 216824 99262 216910 99314
rect 216962 99262 217048 99314
rect 216824 98978 217048 99262
rect 216824 98926 216910 98978
rect 216962 98926 217048 98978
rect 216824 98642 217048 98926
rect 216824 98590 216910 98642
rect 216962 98590 217048 98642
rect 216824 98306 217048 98590
rect 216824 98254 216910 98306
rect 216962 98254 217048 98306
rect 216824 97972 217048 98254
rect 216824 97916 216908 97972
rect 216964 97916 217048 97972
rect 216824 97634 217048 97916
rect 216824 97582 216910 97634
rect 216962 97582 217048 97634
rect 216824 97298 217048 97582
rect 216824 97246 216910 97298
rect 216962 97246 217048 97298
rect 216824 96962 217048 97246
rect 216824 96910 216910 96962
rect 216962 96910 217048 96962
rect 216824 96626 217048 96910
rect 216824 96574 216910 96626
rect 216962 96574 217048 96626
rect 216824 96292 217048 96574
rect 216824 96236 216908 96292
rect 216964 96236 217048 96292
rect 216824 95954 217048 96236
rect 216824 95902 216910 95954
rect 216962 95902 217048 95954
rect 216824 95618 217048 95902
rect 216824 95566 216910 95618
rect 216962 95566 217048 95618
rect 216824 95282 217048 95566
rect 216824 95230 216910 95282
rect 216962 95230 217048 95282
rect 216824 94946 217048 95230
rect 216824 94894 216910 94946
rect 216962 94894 217048 94946
rect 216824 94612 217048 94894
rect 216824 94556 216908 94612
rect 216964 94556 217048 94612
rect 216824 94274 217048 94556
rect 216824 94222 216910 94274
rect 216962 94222 217048 94274
rect 216824 93938 217048 94222
rect 216824 93886 216910 93938
rect 216962 93886 217048 93938
rect 216824 93602 217048 93886
rect 216824 93550 216910 93602
rect 216962 93550 217048 93602
rect 216824 93266 217048 93550
rect 216824 93214 216910 93266
rect 216962 93214 217048 93266
rect 216824 92932 217048 93214
rect 216824 92876 216908 92932
rect 216964 92876 217048 92932
rect 216824 92594 217048 92876
rect 216824 92542 216910 92594
rect 216962 92542 217048 92594
rect 216824 92258 217048 92542
rect 216824 92206 216910 92258
rect 216962 92206 217048 92258
rect 216824 91922 217048 92206
rect 216824 91870 216910 91922
rect 216962 91870 217048 91922
rect 216824 91586 217048 91870
rect 216824 91534 216910 91586
rect 216962 91534 217048 91586
rect 216824 91252 217048 91534
rect 216824 91196 216908 91252
rect 216964 91196 217048 91252
rect 216824 90914 217048 91196
rect 216824 90862 216910 90914
rect 216962 90862 217048 90914
rect 216824 90578 217048 90862
rect 216824 90526 216910 90578
rect 216962 90526 217048 90578
rect 216824 90242 217048 90526
rect 216824 90190 216910 90242
rect 216962 90190 217048 90242
rect 216824 89906 217048 90190
rect 216824 89854 216910 89906
rect 216962 89854 217048 89906
rect 216824 89572 217048 89854
rect 216824 89516 216908 89572
rect 216964 89516 217048 89572
rect 216824 89234 217048 89516
rect 216824 89182 216910 89234
rect 216962 89182 217048 89234
rect 216824 88898 217048 89182
rect 216824 88846 216910 88898
rect 216962 88846 217048 88898
rect 216824 88562 217048 88846
rect 216824 88510 216910 88562
rect 216962 88510 217048 88562
rect 216824 88226 217048 88510
rect 216824 88174 216910 88226
rect 216962 88174 217048 88226
rect 216824 87892 217048 88174
rect 216824 87836 216908 87892
rect 216964 87836 217048 87892
rect 216824 87554 217048 87836
rect 216824 87502 216910 87554
rect 216962 87502 217048 87554
rect 216824 87218 217048 87502
rect 216824 87166 216910 87218
rect 216962 87166 217048 87218
rect 216824 86882 217048 87166
rect 216824 86830 216910 86882
rect 216962 86830 217048 86882
rect 216824 86546 217048 86830
rect 216824 86494 216910 86546
rect 216962 86494 217048 86546
rect 216824 86212 217048 86494
rect 216824 86156 216908 86212
rect 216964 86156 217048 86212
rect 216824 85874 217048 86156
rect 216824 85822 216910 85874
rect 216962 85822 217048 85874
rect 216824 85538 217048 85822
rect 216824 85486 216910 85538
rect 216962 85486 217048 85538
rect 216824 85202 217048 85486
rect 216824 85150 216910 85202
rect 216962 85150 217048 85202
rect 216824 84866 217048 85150
rect 216824 84814 216910 84866
rect 216962 84814 217048 84866
rect 216824 84532 217048 84814
rect 216824 84476 216908 84532
rect 216964 84476 217048 84532
rect 216824 84194 217048 84476
rect 216824 84142 216910 84194
rect 216962 84142 217048 84194
rect 216824 83858 217048 84142
rect 216824 83806 216910 83858
rect 216962 83806 217048 83858
rect 216824 83522 217048 83806
rect 216824 83470 216910 83522
rect 216962 83470 217048 83522
rect 216824 83186 217048 83470
rect 216824 83134 216910 83186
rect 216962 83134 217048 83186
rect 216824 82852 217048 83134
rect 216824 82796 216908 82852
rect 216964 82796 217048 82852
rect 216824 82514 217048 82796
rect 216824 82462 216910 82514
rect 216962 82462 217048 82514
rect 216824 82178 217048 82462
rect 216824 82126 216910 82178
rect 216962 82126 217048 82178
rect 216824 81842 217048 82126
rect 216824 81790 216910 81842
rect 216962 81790 217048 81842
rect 216824 81506 217048 81790
rect 216824 81454 216910 81506
rect 216962 81454 217048 81506
rect 216824 81172 217048 81454
rect 216824 81116 216908 81172
rect 216964 81116 217048 81172
rect 216824 80834 217048 81116
rect 216824 80782 216910 80834
rect 216962 80782 217048 80834
rect 216824 80498 217048 80782
rect 216824 80446 216910 80498
rect 216962 80446 217048 80498
rect 216824 80162 217048 80446
rect 216824 80110 216910 80162
rect 216962 80110 217048 80162
rect 216824 79826 217048 80110
rect 216824 79774 216910 79826
rect 216962 79774 217048 79826
rect 216824 79492 217048 79774
rect 216824 79436 216908 79492
rect 216964 79436 217048 79492
rect 216824 79154 217048 79436
rect 216824 79102 216910 79154
rect 216962 79102 217048 79154
rect 216824 78818 217048 79102
rect 216824 78766 216910 78818
rect 216962 78766 217048 78818
rect 216824 78482 217048 78766
rect 216824 78430 216910 78482
rect 216962 78430 217048 78482
rect 216824 78146 217048 78430
rect 216824 78094 216910 78146
rect 216962 78094 217048 78146
rect 216824 77812 217048 78094
rect 216824 77756 216908 77812
rect 216964 77756 217048 77812
rect 216824 77474 217048 77756
rect 216824 77422 216910 77474
rect 216962 77422 217048 77474
rect 216824 77138 217048 77422
rect 216824 77086 216910 77138
rect 216962 77086 217048 77138
rect 216824 76802 217048 77086
rect 216824 76750 216910 76802
rect 216962 76750 217048 76802
rect 216824 76466 217048 76750
rect 216824 76414 216910 76466
rect 216962 76414 217048 76466
rect 216824 76132 217048 76414
rect 216824 76076 216908 76132
rect 216964 76076 217048 76132
rect 216824 75794 217048 76076
rect 216824 75742 216910 75794
rect 216962 75742 217048 75794
rect 216824 75458 217048 75742
rect 216824 75406 216910 75458
rect 216962 75406 217048 75458
rect 216824 75122 217048 75406
rect 216824 75070 216910 75122
rect 216962 75070 217048 75122
rect 216824 74786 217048 75070
rect 216824 74734 216910 74786
rect 216962 74734 217048 74786
rect 216824 74452 217048 74734
rect 216824 74396 216908 74452
rect 216964 74396 217048 74452
rect 216824 74114 217048 74396
rect 216824 74062 216910 74114
rect 216962 74062 217048 74114
rect 216824 73778 217048 74062
rect 216824 73726 216910 73778
rect 216962 73726 217048 73778
rect 216824 73442 217048 73726
rect 216824 73390 216910 73442
rect 216962 73390 217048 73442
rect 216824 73106 217048 73390
rect 216824 73054 216910 73106
rect 216962 73054 217048 73106
rect 216824 72772 217048 73054
rect 216824 72716 216908 72772
rect 216964 72716 217048 72772
rect 216824 72434 217048 72716
rect 216824 72382 216910 72434
rect 216962 72382 217048 72434
rect 216824 72098 217048 72382
rect 216824 72046 216910 72098
rect 216962 72046 217048 72098
rect 216824 71762 217048 72046
rect 216824 71710 216910 71762
rect 216962 71710 217048 71762
rect 216824 71426 217048 71710
rect 216824 71374 216910 71426
rect 216962 71374 217048 71426
rect 216824 71092 217048 71374
rect 216824 71036 216908 71092
rect 216964 71036 217048 71092
rect 216824 70754 217048 71036
rect 216824 70702 216910 70754
rect 216962 70702 217048 70754
rect 216824 70418 217048 70702
rect 216824 70366 216910 70418
rect 216962 70366 217048 70418
rect 216824 70082 217048 70366
rect 216824 70030 216910 70082
rect 216962 70030 217048 70082
rect 216824 69746 217048 70030
rect 216824 69694 216910 69746
rect 216962 69694 217048 69746
rect 216824 69412 217048 69694
rect 216824 69356 216908 69412
rect 216964 69356 217048 69412
rect 216824 69074 217048 69356
rect 216824 69022 216910 69074
rect 216962 69022 217048 69074
rect 216824 68738 217048 69022
rect 216824 68686 216910 68738
rect 216962 68686 217048 68738
rect 216824 68402 217048 68686
rect 216824 68350 216910 68402
rect 216962 68350 217048 68402
rect 216824 68066 217048 68350
rect 216824 68014 216910 68066
rect 216962 68014 217048 68066
rect 216824 67732 217048 68014
rect 216824 67676 216908 67732
rect 216964 67676 217048 67732
rect 216824 67394 217048 67676
rect 216824 67342 216910 67394
rect 216962 67342 217048 67394
rect 216824 67058 217048 67342
rect 216824 67006 216910 67058
rect 216962 67006 217048 67058
rect 216824 66722 217048 67006
rect 216824 66670 216910 66722
rect 216962 66670 217048 66722
rect 216824 66386 217048 66670
rect 216824 66334 216910 66386
rect 216962 66334 217048 66386
rect 216824 66052 217048 66334
rect 216824 65996 216908 66052
rect 216964 65996 217048 66052
rect 216824 65714 217048 65996
rect 216824 65662 216910 65714
rect 216962 65662 217048 65714
rect 216824 65378 217048 65662
rect 216824 65326 216910 65378
rect 216962 65326 217048 65378
rect 216824 65042 217048 65326
rect 216824 64990 216910 65042
rect 216962 64990 217048 65042
rect 216824 64706 217048 64990
rect 216824 64654 216910 64706
rect 216962 64654 217048 64706
rect 216824 64372 217048 64654
rect 216824 64316 216908 64372
rect 216964 64316 217048 64372
rect 216824 64034 217048 64316
rect 216824 63982 216910 64034
rect 216962 63982 217048 64034
rect 216824 63698 217048 63982
rect 216824 63646 216910 63698
rect 216962 63646 217048 63698
rect 216824 63362 217048 63646
rect 216824 63310 216910 63362
rect 216962 63310 217048 63362
rect 216824 63026 217048 63310
rect 216824 62974 216910 63026
rect 216962 62974 217048 63026
rect 216824 62692 217048 62974
rect 216824 62636 216908 62692
rect 216964 62636 217048 62692
rect 216824 62354 217048 62636
rect 216824 62302 216910 62354
rect 216962 62302 217048 62354
rect 216824 62018 217048 62302
rect 216824 61966 216910 62018
rect 216962 61966 217048 62018
rect 216824 61682 217048 61966
rect 216824 61630 216910 61682
rect 216962 61630 217048 61682
rect 216824 61346 217048 61630
rect 216824 61294 216910 61346
rect 216962 61294 217048 61346
rect 216824 61012 217048 61294
rect 216824 60956 216908 61012
rect 216964 60956 217048 61012
rect 216824 60674 217048 60956
rect 216824 60622 216910 60674
rect 216962 60622 217048 60674
rect 216824 60338 217048 60622
rect 216824 60286 216910 60338
rect 216962 60286 217048 60338
rect 216824 60002 217048 60286
rect 216824 59950 216910 60002
rect 216962 59950 217048 60002
rect 216824 59666 217048 59950
rect 216824 59614 216910 59666
rect 216962 59614 217048 59666
rect 216824 59332 217048 59614
rect 216824 59276 216908 59332
rect 216964 59276 217048 59332
rect 216824 58994 217048 59276
rect 216824 58942 216910 58994
rect 216962 58942 217048 58994
rect 216824 58658 217048 58942
rect 216824 58606 216910 58658
rect 216962 58606 217048 58658
rect 216824 58322 217048 58606
rect 216824 58270 216910 58322
rect 216962 58270 217048 58322
rect 216824 57986 217048 58270
rect 216824 57934 216910 57986
rect 216962 57934 217048 57986
rect 216824 57652 217048 57934
rect 216824 57596 216908 57652
rect 216964 57596 217048 57652
rect 216824 57314 217048 57596
rect 216824 57262 216910 57314
rect 216962 57262 217048 57314
rect 216824 56978 217048 57262
rect 216824 56926 216910 56978
rect 216962 56926 217048 56978
rect 216824 56642 217048 56926
rect 216824 56590 216910 56642
rect 216962 56590 217048 56642
rect 216824 56306 217048 56590
rect 216824 56254 216910 56306
rect 216962 56254 217048 56306
rect 216824 55972 217048 56254
rect 216824 55916 216908 55972
rect 216964 55916 217048 55972
rect 216824 55634 217048 55916
rect 216824 55582 216910 55634
rect 216962 55582 217048 55634
rect 216824 55298 217048 55582
rect 216824 55246 216910 55298
rect 216962 55246 217048 55298
rect 216824 54962 217048 55246
rect 216824 54910 216910 54962
rect 216962 54910 217048 54962
rect 216824 54626 217048 54910
rect 216824 54574 216910 54626
rect 216962 54574 217048 54626
rect 216824 54292 217048 54574
rect 216824 54236 216908 54292
rect 216964 54236 217048 54292
rect 216824 53954 217048 54236
rect 216824 53902 216910 53954
rect 216962 53902 217048 53954
rect 216824 53618 217048 53902
rect 216824 53566 216910 53618
rect 216962 53566 217048 53618
rect 216824 53282 217048 53566
rect 216824 53230 216910 53282
rect 216962 53230 217048 53282
rect 216824 52946 217048 53230
rect 216824 52894 216910 52946
rect 216962 52894 217048 52946
rect 216824 52612 217048 52894
rect 216824 52556 216908 52612
rect 216964 52556 217048 52612
rect 216824 52274 217048 52556
rect 216824 52222 216910 52274
rect 216962 52222 217048 52274
rect 216824 51938 217048 52222
rect 216824 51886 216910 51938
rect 216962 51886 217048 51938
rect 216824 51602 217048 51886
rect 216824 51550 216910 51602
rect 216962 51550 217048 51602
rect 216824 51266 217048 51550
rect 216824 51214 216910 51266
rect 216962 51214 217048 51266
rect 216824 50932 217048 51214
rect 216824 50876 216908 50932
rect 216964 50876 217048 50932
rect 216824 50594 217048 50876
rect 216824 50542 216910 50594
rect 216962 50542 217048 50594
rect 216824 50258 217048 50542
rect 216824 50206 216910 50258
rect 216962 50206 217048 50258
rect 216824 49922 217048 50206
rect 216824 49870 216910 49922
rect 216962 49870 217048 49922
rect 216824 49586 217048 49870
rect 216824 49534 216910 49586
rect 216962 49534 217048 49586
rect 216824 49252 217048 49534
rect 216824 49196 216908 49252
rect 216964 49196 217048 49252
rect 216824 48914 217048 49196
rect 216824 48862 216910 48914
rect 216962 48862 217048 48914
rect 216824 48578 217048 48862
rect 216824 48526 216910 48578
rect 216962 48526 217048 48578
rect 216824 48242 217048 48526
rect 216824 48190 216910 48242
rect 216962 48190 217048 48242
rect 216824 47906 217048 48190
rect 216824 47854 216910 47906
rect 216962 47854 217048 47906
rect 216824 47572 217048 47854
rect 216824 47516 216908 47572
rect 216964 47516 217048 47572
rect 216824 47234 217048 47516
rect 216824 47182 216910 47234
rect 216962 47182 217048 47234
rect 216824 46898 217048 47182
rect 216824 46846 216910 46898
rect 216962 46846 217048 46898
rect 216824 46562 217048 46846
rect 216824 46510 216910 46562
rect 216962 46510 217048 46562
rect 216824 46226 217048 46510
rect 216824 46174 216910 46226
rect 216962 46174 217048 46226
rect 216824 45892 217048 46174
rect 216824 45836 216908 45892
rect 216964 45836 217048 45892
rect 216824 45554 217048 45836
rect 216824 45502 216910 45554
rect 216962 45502 217048 45554
rect 216824 45218 217048 45502
rect 216824 45166 216910 45218
rect 216962 45166 217048 45218
rect 216824 44882 217048 45166
rect 216824 44830 216910 44882
rect 216962 44830 217048 44882
rect 216824 44546 217048 44830
rect 216824 44494 216910 44546
rect 216962 44494 217048 44546
rect 216824 44212 217048 44494
rect 216824 44156 216908 44212
rect 216964 44156 217048 44212
rect 216824 43874 217048 44156
rect 216824 43822 216910 43874
rect 216962 43822 217048 43874
rect 216824 43538 217048 43822
rect 216824 43486 216910 43538
rect 216962 43486 217048 43538
rect 216824 43202 217048 43486
rect 216824 43150 216910 43202
rect 216962 43150 217048 43202
rect 216824 42866 217048 43150
rect 216824 42814 216910 42866
rect 216962 42814 217048 42866
rect 216824 42532 217048 42814
rect 216824 42476 216908 42532
rect 216964 42476 217048 42532
rect 216824 42194 217048 42476
rect 216824 42142 216910 42194
rect 216962 42142 217048 42194
rect 216824 41858 217048 42142
rect 216824 41806 216910 41858
rect 216962 41806 217048 41858
rect 216824 41522 217048 41806
rect 216824 41470 216910 41522
rect 216962 41470 217048 41522
rect 216824 41186 217048 41470
rect 216824 41134 216910 41186
rect 216962 41134 217048 41186
rect 216824 40852 217048 41134
rect 216824 40796 216908 40852
rect 216964 40796 217048 40852
rect 216824 40514 217048 40796
rect 216824 40462 216910 40514
rect 216962 40462 217048 40514
rect 216824 40178 217048 40462
rect 216824 40126 216910 40178
rect 216962 40126 217048 40178
rect 216824 39842 217048 40126
rect 216824 39790 216910 39842
rect 216962 39790 217048 39842
rect 216824 39506 217048 39790
rect 216824 39454 216910 39506
rect 216962 39454 217048 39506
rect 216824 39172 217048 39454
rect 216824 39116 216908 39172
rect 216964 39116 217048 39172
rect 216824 38834 217048 39116
rect 216824 38782 216910 38834
rect 216962 38782 217048 38834
rect 216824 38498 217048 38782
rect 216824 38446 216910 38498
rect 216962 38446 217048 38498
rect 216824 38162 217048 38446
rect 216824 38110 216910 38162
rect 216962 38110 217048 38162
rect 216824 37826 217048 38110
rect 216824 37774 216910 37826
rect 216962 37774 217048 37826
rect 216824 37492 217048 37774
rect 216824 37436 216908 37492
rect 216964 37436 217048 37492
rect 216824 37154 217048 37436
rect 216824 37102 216910 37154
rect 216962 37102 217048 37154
rect 216824 36818 217048 37102
rect 216824 36766 216910 36818
rect 216962 36766 217048 36818
rect 216824 36482 217048 36766
rect 216824 36430 216910 36482
rect 216962 36430 217048 36482
rect 216824 36146 217048 36430
rect 216824 36094 216910 36146
rect 216962 36094 217048 36146
rect 216824 35812 217048 36094
rect 216824 35756 216908 35812
rect 216964 35756 217048 35812
rect 216824 35474 217048 35756
rect 216824 35422 216910 35474
rect 216962 35422 217048 35474
rect 216824 35138 217048 35422
rect 216824 35086 216910 35138
rect 216962 35086 217048 35138
rect 216824 34802 217048 35086
rect 216824 34750 216910 34802
rect 216962 34750 217048 34802
rect 216824 34466 217048 34750
rect 216824 34414 216910 34466
rect 216962 34414 217048 34466
rect 216824 34132 217048 34414
rect 216824 34076 216908 34132
rect 216964 34076 217048 34132
rect 216824 33794 217048 34076
rect 216824 33742 216910 33794
rect 216962 33742 217048 33794
rect 216824 33458 217048 33742
rect 216824 33406 216910 33458
rect 216962 33406 217048 33458
rect 216824 33122 217048 33406
rect 216824 33070 216910 33122
rect 216962 33070 217048 33122
rect 216824 32786 217048 33070
rect 216824 32734 216910 32786
rect 216962 32734 217048 32786
rect 216824 32452 217048 32734
rect 216824 32396 216908 32452
rect 216964 32396 217048 32452
rect 216824 32114 217048 32396
rect 216824 32062 216910 32114
rect 216962 32062 217048 32114
rect 216824 31778 217048 32062
rect 216824 31726 216910 31778
rect 216962 31726 217048 31778
rect 216824 31442 217048 31726
rect 216824 31390 216910 31442
rect 216962 31390 217048 31442
rect 216824 31106 217048 31390
rect 216824 31054 216910 31106
rect 216962 31054 217048 31106
rect 216824 30772 217048 31054
rect 216824 30716 216908 30772
rect 216964 30716 217048 30772
rect 216824 30434 217048 30716
rect 216824 30382 216910 30434
rect 216962 30382 217048 30434
rect 216824 30098 217048 30382
rect 216824 30046 216910 30098
rect 216962 30046 217048 30098
rect 216824 29762 217048 30046
rect 216824 29710 216910 29762
rect 216962 29710 217048 29762
rect 216824 29426 217048 29710
rect 216824 29374 216910 29426
rect 216962 29374 217048 29426
rect 216824 29092 217048 29374
rect 216824 29036 216908 29092
rect 216964 29036 217048 29092
rect 216824 28754 217048 29036
rect 216824 28702 216910 28754
rect 216962 28702 217048 28754
rect 216824 28418 217048 28702
rect 216824 28366 216910 28418
rect 216962 28366 217048 28418
rect 216824 28082 217048 28366
rect 216824 28030 216910 28082
rect 216962 28030 217048 28082
rect 216824 27746 217048 28030
rect 216824 27694 216910 27746
rect 216962 27694 217048 27746
rect 216824 27412 217048 27694
rect 216824 27356 216908 27412
rect 216964 27356 217048 27412
rect 216824 27074 217048 27356
rect 216824 27022 216910 27074
rect 216962 27022 217048 27074
rect 216824 26738 217048 27022
rect 216824 26686 216910 26738
rect 216962 26686 217048 26738
rect 216824 26402 217048 26686
rect 216824 26350 216910 26402
rect 216962 26350 217048 26402
rect 216824 26066 217048 26350
rect 216824 26014 216910 26066
rect 216962 26014 217048 26066
rect 216824 25732 217048 26014
rect 216824 25676 216908 25732
rect 216964 25676 217048 25732
rect 216824 25394 217048 25676
rect 216824 25342 216910 25394
rect 216962 25342 217048 25394
rect 216824 25058 217048 25342
rect 216824 25006 216910 25058
rect 216962 25006 217048 25058
rect 216824 24722 217048 25006
rect 216824 24670 216910 24722
rect 216962 24670 217048 24722
rect 203400 24557 203456 24566
rect 23766 23253 23794 24538
rect 203400 24492 203456 24501
rect 216824 24386 217048 24670
rect 216824 24334 216910 24386
rect 216962 24334 217048 24386
rect 204482 24301 204538 24310
rect 203199 24230 203255 24239
rect 203199 24165 203255 24174
rect 203537 24230 203593 24239
rect 204482 24236 204538 24245
rect 203537 24165 203593 24174
rect 23752 23244 23808 23253
rect 23752 23179 23808 23188
rect 27467 20425 27495 24061
rect 27453 20416 27509 20425
rect 27453 20351 27509 20360
rect 27591 17597 27619 24061
rect 27715 19011 27743 24061
rect 216824 24052 217048 24334
rect 216824 23996 216908 24052
rect 216964 23996 217048 24052
rect 216824 23714 217048 23996
rect 216824 23662 216910 23714
rect 216962 23662 217048 23714
rect 216824 23378 217048 23662
rect 216824 23326 216910 23378
rect 216962 23326 217048 23378
rect 216824 23042 217048 23326
rect 216824 22990 216910 23042
rect 216962 22990 217048 23042
rect 216824 22706 217048 22990
rect 203119 22672 203175 22681
rect 203119 22607 203175 22616
rect 203537 22672 203593 22681
rect 203537 22607 203593 22616
rect 216824 22654 216910 22706
rect 216962 22654 217048 22706
rect 204482 22601 204538 22610
rect 204482 22536 204538 22545
rect 216824 22372 217048 22654
rect 216824 22316 216908 22372
rect 216964 22316 217048 22372
rect 216824 22034 217048 22316
rect 216824 21982 216910 22034
rect 216962 21982 217048 22034
rect 216824 21698 217048 21982
rect 216824 21646 216910 21698
rect 216962 21646 217048 21698
rect 204482 21473 204538 21482
rect 203039 21402 203095 21411
rect 203039 21337 203095 21346
rect 203537 21402 203593 21411
rect 204482 21408 204538 21417
rect 203537 21337 203593 21346
rect 216824 21362 217048 21646
rect 216824 21310 216910 21362
rect 216962 21310 217048 21362
rect 216824 21026 217048 21310
rect 216824 20974 216910 21026
rect 216962 20974 217048 21026
rect 216824 20692 217048 20974
rect 216824 20636 216908 20692
rect 216964 20636 217048 20692
rect 216824 20354 217048 20636
rect 216824 20302 216910 20354
rect 216962 20302 217048 20354
rect 216824 20018 217048 20302
rect 216824 19966 216910 20018
rect 216962 19966 217048 20018
rect 202959 19844 203015 19853
rect 202959 19779 203015 19788
rect 203537 19844 203593 19853
rect 203537 19779 203593 19788
rect 204482 19773 204538 19782
rect 204482 19708 204538 19717
rect 216824 19682 217048 19966
rect 216824 19630 216910 19682
rect 216962 19630 217048 19682
rect 216824 19346 217048 19630
rect 216824 19294 216910 19346
rect 216962 19294 217048 19346
rect 216824 19012 217048 19294
rect 27701 19002 27757 19011
rect 27701 18937 27757 18946
rect 216824 18956 216908 19012
rect 216964 18956 217048 19012
rect 216824 18674 217048 18956
rect 204482 18645 204538 18654
rect 202879 18574 202935 18583
rect 202879 18509 202935 18518
rect 203537 18574 203593 18583
rect 204482 18580 204538 18589
rect 216824 18622 216910 18674
rect 216962 18622 217048 18674
rect 203537 18509 203593 18518
rect 216824 18338 217048 18622
rect 216824 18286 216910 18338
rect 216962 18286 217048 18338
rect 216824 18002 217048 18286
rect 216824 17950 216910 18002
rect 216962 17950 217048 18002
rect 29560 17756 29616 17765
rect 29560 17691 29616 17700
rect 34552 17756 34608 17765
rect 34552 17691 34608 17700
rect 39544 17756 39600 17765
rect 39544 17691 39600 17700
rect 44536 17756 44592 17765
rect 44536 17691 44592 17700
rect 49528 17756 49584 17765
rect 49528 17691 49584 17700
rect 54520 17756 54576 17765
rect 54520 17691 54576 17700
rect 59512 17756 59568 17765
rect 59512 17691 59568 17700
rect 64504 17756 64560 17765
rect 64504 17691 64560 17700
rect 69496 17756 69552 17765
rect 69496 17691 69552 17700
rect 74488 17756 74544 17765
rect 74488 17691 74544 17700
rect 79480 17756 79536 17765
rect 79480 17691 79536 17700
rect 84472 17756 84528 17765
rect 84472 17691 84528 17700
rect 89464 17756 89520 17765
rect 89464 17691 89520 17700
rect 94456 17756 94512 17765
rect 94456 17691 94512 17700
rect 99448 17756 99504 17765
rect 99448 17691 99504 17700
rect 104440 17756 104496 17765
rect 104440 17691 104496 17700
rect 109432 17756 109488 17765
rect 109432 17691 109488 17700
rect 114424 17756 114480 17765
rect 114424 17691 114480 17700
rect 119416 17756 119472 17765
rect 119416 17691 119472 17700
rect 124408 17756 124464 17765
rect 124408 17691 124464 17700
rect 129400 17756 129456 17765
rect 129400 17691 129456 17700
rect 134392 17756 134448 17765
rect 134392 17691 134448 17700
rect 139384 17756 139440 17765
rect 139384 17691 139440 17700
rect 144376 17756 144432 17765
rect 144376 17691 144432 17700
rect 149368 17756 149424 17765
rect 149368 17691 149424 17700
rect 154360 17756 154416 17765
rect 154360 17691 154416 17700
rect 159352 17756 159408 17765
rect 159352 17691 159408 17700
rect 164344 17756 164400 17765
rect 164344 17691 164400 17700
rect 169336 17756 169392 17765
rect 169336 17691 169392 17700
rect 174328 17756 174384 17765
rect 174328 17691 174384 17700
rect 179320 17756 179376 17765
rect 179320 17691 179376 17700
rect 184312 17756 184368 17765
rect 184312 17691 184368 17700
rect 216824 17666 217048 17950
rect 216824 17614 216910 17666
rect 216962 17614 217048 17666
rect 27577 17588 27633 17597
rect 27577 17523 27633 17532
rect 216824 17332 217048 17614
rect 216824 17276 216908 17332
rect 216964 17276 217048 17332
rect 202799 17016 202855 17025
rect 202799 16951 202855 16960
rect 203537 17016 203593 17025
rect 203537 16951 203593 16960
rect 216824 16994 217048 17276
rect 204482 16945 204538 16954
rect 204482 16880 204538 16889
rect 216824 16942 216910 16994
rect 216962 16942 217048 16994
rect 216824 16658 217048 16942
rect 216824 16606 216910 16658
rect 216962 16606 217048 16658
rect 216824 16322 217048 16606
rect 216824 16270 216910 16322
rect 216962 16270 217048 16322
rect 216824 15986 217048 16270
rect 216824 15934 216910 15986
rect 216962 15934 217048 15986
rect 204482 15817 204538 15826
rect 202719 15746 202775 15755
rect 202719 15681 202775 15690
rect 203537 15746 203593 15755
rect 204482 15752 204538 15761
rect 203537 15681 203593 15690
rect 216824 15652 217048 15934
rect 216824 15596 216908 15652
rect 216964 15596 217048 15652
rect 216824 15314 217048 15596
rect 216824 15262 216910 15314
rect 216962 15262 217048 15314
rect 216824 14978 217048 15262
rect 216824 14926 216910 14978
rect 216962 14926 217048 14978
rect 216824 14642 217048 14926
rect 216824 14590 216910 14642
rect 216962 14590 217048 14642
rect 216824 14306 217048 14590
rect 216824 14254 216910 14306
rect 216962 14254 217048 14306
rect 202639 14188 202695 14197
rect 202639 14123 202695 14132
rect 203537 14188 203593 14197
rect 203537 14123 203593 14132
rect 204482 14117 204538 14126
rect 204482 14052 204538 14061
rect 1618 13246 1704 13298
rect 1756 13246 1842 13298
rect 1618 12962 1842 13246
rect 5511 13308 5567 13317
rect 15238 13304 15336 13332
rect 5511 13243 5567 13252
rect 2326 13203 2382 13212
rect 2326 13138 2382 13147
rect 1618 12910 1704 12962
rect 1756 12910 1842 12962
rect 1618 12626 1842 12910
rect 1618 12574 1704 12626
rect 1756 12574 1842 12626
rect 1618 12292 1842 12574
rect 1618 12236 1702 12292
rect 1758 12236 1842 12292
rect 1618 11954 1842 12236
rect 1618 11902 1704 11954
rect 1756 11902 1842 11954
rect 1618 11618 1842 11902
rect 1618 11566 1704 11618
rect 1756 11566 1842 11618
rect 1618 11282 1842 11566
rect 1618 11230 1704 11282
rect 1756 11230 1842 11282
rect 1618 10946 1842 11230
rect 1618 10894 1704 10946
rect 1756 10894 1842 10946
rect 1618 10612 1842 10894
rect 1618 10556 1702 10612
rect 1758 10556 1842 10612
rect 1618 10274 1842 10556
rect 1618 10222 1704 10274
rect 1756 10222 1842 10274
rect 1618 9938 1842 10222
rect 1618 9886 1704 9938
rect 1756 9886 1842 9938
rect 1618 9602 1842 9886
rect 1618 9550 1704 9602
rect 1756 9550 1842 9602
rect 1618 9266 1842 9550
rect 1618 9214 1704 9266
rect 1756 9214 1842 9266
rect 1618 8932 1842 9214
rect 1618 8876 1702 8932
rect 1758 8876 1842 8932
rect 1618 8594 1842 8876
rect 1618 8542 1704 8594
rect 1756 8542 1842 8594
rect 1618 8258 1842 8542
rect 1618 8206 1704 8258
rect 1756 8206 1842 8258
rect 1618 7922 1842 8206
rect 1618 7870 1704 7922
rect 1756 7870 1842 7922
rect 1618 7586 1842 7870
rect 1618 7534 1704 7586
rect 1756 7534 1842 7586
rect 1618 7252 1842 7534
rect 1618 7196 1702 7252
rect 1758 7196 1842 7252
rect 1618 6914 1842 7196
rect 1618 6862 1704 6914
rect 1756 6862 1842 6914
rect 1618 6578 1842 6862
rect 1618 6526 1704 6578
rect 1756 6526 1842 6578
rect 1618 6242 1842 6526
rect 1618 6190 1704 6242
rect 1756 6190 1842 6242
rect 1618 5906 1842 6190
rect 1618 5854 1704 5906
rect 1756 5854 1842 5906
rect 1618 5572 1842 5854
rect 1618 5516 1702 5572
rect 1758 5516 1842 5572
rect 1618 5234 1842 5516
rect 1618 5182 1704 5234
rect 1756 5182 1842 5234
rect 1618 4898 1842 5182
rect 1618 4846 1704 4898
rect 1756 4846 1842 4898
rect 1618 4562 1842 4846
rect 1618 4510 1704 4562
rect 1756 4510 1842 4562
rect 1618 4226 1842 4510
rect 1618 4174 1704 4226
rect 1756 4174 1842 4226
rect 1618 3892 1842 4174
rect 1618 3836 1702 3892
rect 1758 3836 1842 3892
rect 1618 3554 1842 3836
rect 1618 3502 1704 3554
rect 1756 3502 1842 3554
rect 1618 3218 1842 3502
rect 1618 3166 1704 3218
rect 1756 3166 1842 3218
rect 1618 2882 1842 3166
rect 1618 2830 1704 2882
rect 1756 2830 1842 2882
rect 1618 2546 1842 2830
rect 1618 2494 1704 2546
rect 1756 2494 1842 2546
rect 15308 2529 15336 13304
rect 216824 13972 217048 14254
rect 216824 13916 216908 13972
rect 216964 13916 217048 13972
rect 216824 13634 217048 13916
rect 216824 13582 216910 13634
rect 216962 13582 217048 13634
rect 216824 13298 217048 13582
rect 216824 13246 216910 13298
rect 216962 13246 217048 13298
rect 216824 12962 217048 13246
rect 216824 12910 216910 12962
rect 216962 12910 217048 12962
rect 216824 12626 217048 12910
rect 216824 12574 216910 12626
rect 216962 12574 217048 12626
rect 216824 12292 217048 12574
rect 216824 12236 216908 12292
rect 216964 12236 217048 12292
rect 216824 11954 217048 12236
rect 216824 11902 216910 11954
rect 216962 11902 217048 11954
rect 216824 11618 217048 11902
rect 216824 11566 216910 11618
rect 216962 11566 217048 11618
rect 216824 11282 217048 11566
rect 216824 11230 216910 11282
rect 216962 11230 217048 11282
rect 216824 10946 217048 11230
rect 216824 10894 216910 10946
rect 216962 10894 217048 10946
rect 216824 10612 217048 10894
rect 216824 10556 216908 10612
rect 216964 10556 217048 10612
rect 216824 10274 217048 10556
rect 216824 10222 216910 10274
rect 216962 10222 217048 10274
rect 216824 9938 217048 10222
rect 216824 9886 216910 9938
rect 216962 9886 217048 9938
rect 216824 9602 217048 9886
rect 216824 9550 216910 9602
rect 216962 9550 217048 9602
rect 216824 9266 217048 9550
rect 216824 9214 216910 9266
rect 216962 9214 217048 9266
rect 216824 8932 217048 9214
rect 216824 8876 216908 8932
rect 216964 8876 217048 8932
rect 216824 8594 217048 8876
rect 216824 8542 216910 8594
rect 216962 8542 217048 8594
rect 216824 8258 217048 8542
rect 216824 8206 216910 8258
rect 216962 8206 217048 8258
rect 216824 7922 217048 8206
rect 216824 7870 216910 7922
rect 216962 7870 217048 7922
rect 216824 7586 217048 7870
rect 216824 7534 216910 7586
rect 216962 7534 217048 7586
rect 216824 7252 217048 7534
rect 216824 7196 216908 7252
rect 216964 7196 217048 7252
rect 216824 6914 217048 7196
rect 216824 6862 216910 6914
rect 216962 6862 217048 6914
rect 216824 6578 217048 6862
rect 216824 6526 216910 6578
rect 216962 6526 217048 6578
rect 216824 6242 217048 6526
rect 216824 6190 216910 6242
rect 216962 6190 217048 6242
rect 216824 5906 217048 6190
rect 216824 5854 216910 5906
rect 216962 5854 217048 5906
rect 216824 5572 217048 5854
rect 216824 5516 216908 5572
rect 216964 5516 217048 5572
rect 216824 5234 217048 5516
rect 216824 5182 216910 5234
rect 216962 5182 217048 5234
rect 216824 4898 217048 5182
rect 216824 4846 216910 4898
rect 216962 4846 217048 4898
rect 216824 4562 217048 4846
rect 216824 4510 216910 4562
rect 216962 4510 217048 4562
rect 216824 4226 217048 4510
rect 216824 4174 216910 4226
rect 216962 4174 217048 4226
rect 216824 3892 217048 4174
rect 216824 3836 216908 3892
rect 216964 3836 217048 3892
rect 216824 3554 217048 3836
rect 216824 3502 216910 3554
rect 216962 3502 217048 3554
rect 216824 3218 217048 3502
rect 216824 3166 216910 3218
rect 216962 3166 217048 3218
rect 216824 2882 217048 3166
rect 216824 2830 216910 2882
rect 216962 2830 217048 2882
rect 16548 2776 16604 2785
rect 16548 2711 16604 2720
rect 17716 2776 17772 2785
rect 17716 2711 17772 2720
rect 18884 2776 18940 2785
rect 18884 2711 18940 2720
rect 20052 2776 20108 2785
rect 20052 2711 20108 2720
rect 21220 2776 21276 2785
rect 21220 2711 21276 2720
rect 22388 2776 22444 2785
rect 22388 2711 22444 2720
rect 23556 2776 23612 2785
rect 23556 2711 23612 2720
rect 24724 2776 24780 2785
rect 24724 2711 24780 2720
rect 25892 2776 25948 2785
rect 25892 2711 25948 2720
rect 27060 2776 27116 2785
rect 27060 2711 27116 2720
rect 28228 2776 28284 2785
rect 28228 2711 28284 2720
rect 29396 2776 29452 2785
rect 29396 2711 29452 2720
rect 30564 2776 30620 2785
rect 30564 2711 30620 2720
rect 31732 2776 31788 2785
rect 31732 2711 31788 2720
rect 32900 2776 32956 2785
rect 32900 2711 32956 2720
rect 34068 2776 34124 2785
rect 34068 2711 34124 2720
rect 35236 2776 35292 2785
rect 35236 2711 35292 2720
rect 36404 2776 36460 2785
rect 36404 2711 36460 2720
rect 37572 2776 37628 2785
rect 37572 2711 37628 2720
rect 38740 2776 38796 2785
rect 38740 2711 38796 2720
rect 39908 2776 39964 2785
rect 39908 2711 39964 2720
rect 41076 2776 41132 2785
rect 41076 2711 41132 2720
rect 42244 2776 42300 2785
rect 42244 2711 42300 2720
rect 43412 2776 43468 2785
rect 43412 2711 43468 2720
rect 44580 2776 44636 2785
rect 44580 2711 44636 2720
rect 45748 2776 45804 2785
rect 45748 2711 45804 2720
rect 46916 2776 46972 2785
rect 46916 2711 46972 2720
rect 48084 2776 48140 2785
rect 48084 2711 48140 2720
rect 49252 2776 49308 2785
rect 49252 2711 49308 2720
rect 50420 2776 50476 2785
rect 50420 2711 50476 2720
rect 51588 2776 51644 2785
rect 51588 2711 51644 2720
rect 52756 2776 52812 2785
rect 52756 2711 52812 2720
rect 53924 2776 53980 2785
rect 53924 2711 53980 2720
rect 55092 2776 55148 2785
rect 55092 2711 55148 2720
rect 56260 2776 56316 2785
rect 56260 2711 56316 2720
rect 57428 2776 57484 2785
rect 57428 2711 57484 2720
rect 58596 2776 58652 2785
rect 58596 2711 58652 2720
rect 59764 2776 59820 2785
rect 59764 2711 59820 2720
rect 60932 2776 60988 2785
rect 60932 2711 60988 2720
rect 216824 2546 217048 2830
rect 1618 2212 1842 2494
rect 15294 2520 15350 2529
rect 15294 2455 15350 2464
rect 216824 2494 216910 2546
rect 216962 2494 217048 2546
rect 1618 2156 1702 2212
rect 1758 2156 1842 2212
rect 1618 1736 1842 2156
rect 216824 2212 217048 2494
rect 216824 2156 216908 2212
rect 216964 2156 217048 2212
rect 2038 1876 2094 1885
rect 2038 1811 2094 1820
rect 3718 1876 3774 1885
rect 3718 1811 3774 1820
rect 5398 1876 5454 1885
rect 5398 1811 5454 1820
rect 7078 1876 7134 1885
rect 7078 1811 7134 1820
rect 8758 1876 8814 1885
rect 8758 1811 8814 1820
rect 10438 1876 10494 1885
rect 10438 1811 10494 1820
rect 12118 1876 12174 1885
rect 12118 1811 12174 1820
rect 13798 1876 13854 1885
rect 13798 1811 13854 1820
rect 15478 1876 15534 1885
rect 15478 1811 15534 1820
rect 17158 1876 17214 1885
rect 17158 1811 17214 1820
rect 18838 1876 18894 1885
rect 18838 1811 18894 1820
rect 20518 1876 20574 1885
rect 20518 1811 20574 1820
rect 22198 1876 22254 1885
rect 22198 1811 22254 1820
rect 23878 1876 23934 1885
rect 23878 1811 23934 1820
rect 25558 1876 25614 1885
rect 25558 1811 25614 1820
rect 27238 1876 27294 1885
rect 27238 1811 27294 1820
rect 28918 1876 28974 1885
rect 28918 1811 28974 1820
rect 30598 1876 30654 1885
rect 30598 1811 30654 1820
rect 32278 1876 32334 1885
rect 32278 1811 32334 1820
rect 33958 1876 34014 1885
rect 33958 1811 34014 1820
rect 35638 1876 35694 1885
rect 35638 1811 35694 1820
rect 37318 1876 37374 1885
rect 37318 1811 37374 1820
rect 38998 1876 39054 1885
rect 38998 1811 39054 1820
rect 40678 1876 40734 1885
rect 40678 1811 40734 1820
rect 42358 1876 42414 1885
rect 42358 1811 42414 1820
rect 44038 1876 44094 1885
rect 44038 1811 44094 1820
rect 45718 1876 45774 1885
rect 45718 1811 45774 1820
rect 47398 1876 47454 1885
rect 47398 1811 47454 1820
rect 49078 1876 49134 1885
rect 49078 1811 49134 1820
rect 50758 1876 50814 1885
rect 50758 1811 50814 1820
rect 52438 1876 52494 1885
rect 52438 1811 52494 1820
rect 54118 1876 54174 1885
rect 54118 1811 54174 1820
rect 55798 1876 55854 1885
rect 55798 1811 55854 1820
rect 57478 1876 57534 1885
rect 57478 1811 57534 1820
rect 59158 1876 59214 1885
rect 59158 1811 59214 1820
rect 60838 1876 60894 1885
rect 60838 1811 60894 1820
rect 62518 1876 62574 1885
rect 62518 1811 62574 1820
rect 64198 1876 64254 1885
rect 64198 1811 64254 1820
rect 65878 1876 65934 1885
rect 65878 1811 65934 1820
rect 67558 1876 67614 1885
rect 67558 1811 67614 1820
rect 69238 1876 69294 1885
rect 69238 1811 69294 1820
rect 70918 1876 70974 1885
rect 70918 1811 70974 1820
rect 72598 1876 72654 1885
rect 72598 1811 72654 1820
rect 74278 1876 74334 1885
rect 74278 1811 74334 1820
rect 75958 1876 76014 1885
rect 75958 1811 76014 1820
rect 77638 1876 77694 1885
rect 77638 1811 77694 1820
rect 79318 1876 79374 1885
rect 79318 1811 79374 1820
rect 80998 1876 81054 1885
rect 80998 1811 81054 1820
rect 82678 1876 82734 1885
rect 82678 1811 82734 1820
rect 84358 1876 84414 1885
rect 84358 1811 84414 1820
rect 86038 1876 86094 1885
rect 86038 1811 86094 1820
rect 87718 1876 87774 1885
rect 87718 1811 87774 1820
rect 89398 1876 89454 1885
rect 89398 1811 89454 1820
rect 91078 1876 91134 1885
rect 91078 1811 91134 1820
rect 92758 1876 92814 1885
rect 92758 1811 92814 1820
rect 94438 1876 94494 1885
rect 94438 1811 94494 1820
rect 96118 1876 96174 1885
rect 96118 1811 96174 1820
rect 97798 1876 97854 1885
rect 97798 1811 97854 1820
rect 99478 1876 99534 1885
rect 99478 1811 99534 1820
rect 101158 1876 101214 1885
rect 101158 1811 101214 1820
rect 102838 1876 102894 1885
rect 102838 1811 102894 1820
rect 104518 1876 104574 1885
rect 104518 1811 104574 1820
rect 106198 1876 106254 1885
rect 106198 1811 106254 1820
rect 107878 1876 107934 1885
rect 107878 1811 107934 1820
rect 109558 1876 109614 1885
rect 109558 1811 109614 1820
rect 111238 1876 111294 1885
rect 111238 1811 111294 1820
rect 112918 1876 112974 1885
rect 112918 1811 112974 1820
rect 114598 1876 114654 1885
rect 114598 1811 114654 1820
rect 116278 1876 116334 1885
rect 116278 1811 116334 1820
rect 117958 1876 118014 1885
rect 117958 1811 118014 1820
rect 119638 1876 119694 1885
rect 119638 1811 119694 1820
rect 121318 1876 121374 1885
rect 121318 1811 121374 1820
rect 122998 1876 123054 1885
rect 122998 1811 123054 1820
rect 124678 1876 124734 1885
rect 124678 1811 124734 1820
rect 126358 1876 126414 1885
rect 126358 1811 126414 1820
rect 128038 1876 128094 1885
rect 128038 1811 128094 1820
rect 129718 1876 129774 1885
rect 129718 1811 129774 1820
rect 131398 1876 131454 1885
rect 131398 1811 131454 1820
rect 133078 1876 133134 1885
rect 133078 1811 133134 1820
rect 134758 1876 134814 1885
rect 134758 1811 134814 1820
rect 136438 1876 136494 1885
rect 136438 1811 136494 1820
rect 138118 1876 138174 1885
rect 138118 1811 138174 1820
rect 139798 1876 139854 1885
rect 139798 1811 139854 1820
rect 141478 1876 141534 1885
rect 141478 1811 141534 1820
rect 143158 1876 143214 1885
rect 143158 1811 143214 1820
rect 144838 1876 144894 1885
rect 144838 1811 144894 1820
rect 146518 1876 146574 1885
rect 146518 1811 146574 1820
rect 148198 1876 148254 1885
rect 148198 1811 148254 1820
rect 149878 1876 149934 1885
rect 149878 1811 149934 1820
rect 151558 1876 151614 1885
rect 151558 1811 151614 1820
rect 153238 1876 153294 1885
rect 153238 1811 153294 1820
rect 154918 1876 154974 1885
rect 154918 1811 154974 1820
rect 156598 1876 156654 1885
rect 156598 1811 156654 1820
rect 158278 1876 158334 1885
rect 158278 1811 158334 1820
rect 159958 1876 160014 1885
rect 159958 1811 160014 1820
rect 161638 1876 161694 1885
rect 161638 1811 161694 1820
rect 163318 1876 163374 1885
rect 163318 1811 163374 1820
rect 164998 1876 165054 1885
rect 164998 1811 165054 1820
rect 166678 1876 166734 1885
rect 166678 1811 166734 1820
rect 168358 1876 168414 1885
rect 168358 1811 168414 1820
rect 170038 1876 170094 1885
rect 170038 1811 170094 1820
rect 171718 1876 171774 1885
rect 171718 1811 171774 1820
rect 173398 1876 173454 1885
rect 173398 1811 173454 1820
rect 175078 1876 175134 1885
rect 175078 1811 175134 1820
rect 176758 1876 176814 1885
rect 176758 1811 176814 1820
rect 178438 1876 178494 1885
rect 178438 1811 178494 1820
rect 180118 1876 180174 1885
rect 180118 1811 180174 1820
rect 181798 1876 181854 1885
rect 181798 1811 181854 1820
rect 183478 1876 183534 1885
rect 183478 1811 183534 1820
rect 185158 1876 185214 1885
rect 185158 1811 185214 1820
rect 186838 1876 186894 1885
rect 186838 1811 186894 1820
rect 188518 1876 188574 1885
rect 188518 1811 188574 1820
rect 190198 1876 190254 1885
rect 190198 1811 190254 1820
rect 191878 1876 191934 1885
rect 191878 1811 191934 1820
rect 193558 1876 193614 1885
rect 193558 1811 193614 1820
rect 195238 1876 195294 1885
rect 195238 1811 195294 1820
rect 196918 1876 196974 1885
rect 196918 1811 196974 1820
rect 198598 1876 198654 1885
rect 198598 1811 198654 1820
rect 200278 1876 200334 1885
rect 200278 1811 200334 1820
rect 201958 1876 202014 1885
rect 201958 1811 202014 1820
rect 203638 1876 203694 1885
rect 203638 1811 203694 1820
rect 205318 1876 205374 1885
rect 205318 1811 205374 1820
rect 206998 1876 207054 1885
rect 206998 1811 207054 1820
rect 208678 1876 208734 1885
rect 208678 1811 208734 1820
rect 210358 1876 210414 1885
rect 210358 1811 210414 1820
rect 212038 1876 212094 1885
rect 212038 1811 212094 1820
rect 213718 1876 213774 1885
rect 213718 1811 213774 1820
rect 215398 1876 215454 1885
rect 215398 1811 215454 1820
rect 216824 1736 217048 2156
<< via2 >>
rect 2038 142370 2094 142372
rect 2038 142318 2040 142370
rect 2040 142318 2092 142370
rect 2092 142318 2094 142370
rect 2038 142316 2094 142318
rect 3718 142370 3774 142372
rect 3718 142318 3720 142370
rect 3720 142318 3772 142370
rect 3772 142318 3774 142370
rect 3718 142316 3774 142318
rect 5398 142370 5454 142372
rect 5398 142318 5400 142370
rect 5400 142318 5452 142370
rect 5452 142318 5454 142370
rect 5398 142316 5454 142318
rect 7078 142370 7134 142372
rect 7078 142318 7080 142370
rect 7080 142318 7132 142370
rect 7132 142318 7134 142370
rect 7078 142316 7134 142318
rect 8758 142370 8814 142372
rect 8758 142318 8760 142370
rect 8760 142318 8812 142370
rect 8812 142318 8814 142370
rect 8758 142316 8814 142318
rect 10438 142370 10494 142372
rect 10438 142318 10440 142370
rect 10440 142318 10492 142370
rect 10492 142318 10494 142370
rect 10438 142316 10494 142318
rect 12118 142370 12174 142372
rect 12118 142318 12120 142370
rect 12120 142318 12172 142370
rect 12172 142318 12174 142370
rect 12118 142316 12174 142318
rect 13798 142370 13854 142372
rect 13798 142318 13800 142370
rect 13800 142318 13852 142370
rect 13852 142318 13854 142370
rect 13798 142316 13854 142318
rect 15478 142370 15534 142372
rect 15478 142318 15480 142370
rect 15480 142318 15532 142370
rect 15532 142318 15534 142370
rect 15478 142316 15534 142318
rect 17158 142370 17214 142372
rect 17158 142318 17160 142370
rect 17160 142318 17212 142370
rect 17212 142318 17214 142370
rect 17158 142316 17214 142318
rect 18838 142370 18894 142372
rect 18838 142318 18840 142370
rect 18840 142318 18892 142370
rect 18892 142318 18894 142370
rect 18838 142316 18894 142318
rect 20518 142370 20574 142372
rect 20518 142318 20520 142370
rect 20520 142318 20572 142370
rect 20572 142318 20574 142370
rect 20518 142316 20574 142318
rect 22198 142370 22254 142372
rect 22198 142318 22200 142370
rect 22200 142318 22252 142370
rect 22252 142318 22254 142370
rect 22198 142316 22254 142318
rect 23878 142370 23934 142372
rect 23878 142318 23880 142370
rect 23880 142318 23932 142370
rect 23932 142318 23934 142370
rect 23878 142316 23934 142318
rect 25558 142370 25614 142372
rect 25558 142318 25560 142370
rect 25560 142318 25612 142370
rect 25612 142318 25614 142370
rect 25558 142316 25614 142318
rect 27238 142370 27294 142372
rect 27238 142318 27240 142370
rect 27240 142318 27292 142370
rect 27292 142318 27294 142370
rect 27238 142316 27294 142318
rect 28918 142370 28974 142372
rect 28918 142318 28920 142370
rect 28920 142318 28972 142370
rect 28972 142318 28974 142370
rect 28918 142316 28974 142318
rect 30598 142370 30654 142372
rect 30598 142318 30600 142370
rect 30600 142318 30652 142370
rect 30652 142318 30654 142370
rect 30598 142316 30654 142318
rect 32278 142370 32334 142372
rect 32278 142318 32280 142370
rect 32280 142318 32332 142370
rect 32332 142318 32334 142370
rect 32278 142316 32334 142318
rect 33958 142370 34014 142372
rect 33958 142318 33960 142370
rect 33960 142318 34012 142370
rect 34012 142318 34014 142370
rect 33958 142316 34014 142318
rect 35638 142370 35694 142372
rect 35638 142318 35640 142370
rect 35640 142318 35692 142370
rect 35692 142318 35694 142370
rect 35638 142316 35694 142318
rect 37318 142370 37374 142372
rect 37318 142318 37320 142370
rect 37320 142318 37372 142370
rect 37372 142318 37374 142370
rect 37318 142316 37374 142318
rect 38998 142370 39054 142372
rect 38998 142318 39000 142370
rect 39000 142318 39052 142370
rect 39052 142318 39054 142370
rect 38998 142316 39054 142318
rect 40678 142370 40734 142372
rect 40678 142318 40680 142370
rect 40680 142318 40732 142370
rect 40732 142318 40734 142370
rect 40678 142316 40734 142318
rect 42358 142370 42414 142372
rect 42358 142318 42360 142370
rect 42360 142318 42412 142370
rect 42412 142318 42414 142370
rect 42358 142316 42414 142318
rect 44038 142370 44094 142372
rect 44038 142318 44040 142370
rect 44040 142318 44092 142370
rect 44092 142318 44094 142370
rect 44038 142316 44094 142318
rect 45718 142370 45774 142372
rect 45718 142318 45720 142370
rect 45720 142318 45772 142370
rect 45772 142318 45774 142370
rect 45718 142316 45774 142318
rect 47398 142370 47454 142372
rect 47398 142318 47400 142370
rect 47400 142318 47452 142370
rect 47452 142318 47454 142370
rect 47398 142316 47454 142318
rect 49078 142370 49134 142372
rect 49078 142318 49080 142370
rect 49080 142318 49132 142370
rect 49132 142318 49134 142370
rect 49078 142316 49134 142318
rect 50758 142370 50814 142372
rect 50758 142318 50760 142370
rect 50760 142318 50812 142370
rect 50812 142318 50814 142370
rect 50758 142316 50814 142318
rect 52438 142370 52494 142372
rect 52438 142318 52440 142370
rect 52440 142318 52492 142370
rect 52492 142318 52494 142370
rect 52438 142316 52494 142318
rect 54118 142370 54174 142372
rect 54118 142318 54120 142370
rect 54120 142318 54172 142370
rect 54172 142318 54174 142370
rect 54118 142316 54174 142318
rect 55798 142370 55854 142372
rect 55798 142318 55800 142370
rect 55800 142318 55852 142370
rect 55852 142318 55854 142370
rect 55798 142316 55854 142318
rect 57478 142370 57534 142372
rect 57478 142318 57480 142370
rect 57480 142318 57532 142370
rect 57532 142318 57534 142370
rect 57478 142316 57534 142318
rect 59158 142370 59214 142372
rect 59158 142318 59160 142370
rect 59160 142318 59212 142370
rect 59212 142318 59214 142370
rect 59158 142316 59214 142318
rect 60838 142370 60894 142372
rect 60838 142318 60840 142370
rect 60840 142318 60892 142370
rect 60892 142318 60894 142370
rect 60838 142316 60894 142318
rect 62518 142370 62574 142372
rect 62518 142318 62520 142370
rect 62520 142318 62572 142370
rect 62572 142318 62574 142370
rect 62518 142316 62574 142318
rect 64198 142370 64254 142372
rect 64198 142318 64200 142370
rect 64200 142318 64252 142370
rect 64252 142318 64254 142370
rect 64198 142316 64254 142318
rect 65878 142370 65934 142372
rect 65878 142318 65880 142370
rect 65880 142318 65932 142370
rect 65932 142318 65934 142370
rect 65878 142316 65934 142318
rect 67558 142370 67614 142372
rect 67558 142318 67560 142370
rect 67560 142318 67612 142370
rect 67612 142318 67614 142370
rect 67558 142316 67614 142318
rect 69238 142370 69294 142372
rect 69238 142318 69240 142370
rect 69240 142318 69292 142370
rect 69292 142318 69294 142370
rect 69238 142316 69294 142318
rect 70918 142370 70974 142372
rect 70918 142318 70920 142370
rect 70920 142318 70972 142370
rect 70972 142318 70974 142370
rect 70918 142316 70974 142318
rect 72598 142370 72654 142372
rect 72598 142318 72600 142370
rect 72600 142318 72652 142370
rect 72652 142318 72654 142370
rect 72598 142316 72654 142318
rect 74278 142370 74334 142372
rect 74278 142318 74280 142370
rect 74280 142318 74332 142370
rect 74332 142318 74334 142370
rect 74278 142316 74334 142318
rect 75958 142370 76014 142372
rect 75958 142318 75960 142370
rect 75960 142318 76012 142370
rect 76012 142318 76014 142370
rect 75958 142316 76014 142318
rect 77638 142370 77694 142372
rect 77638 142318 77640 142370
rect 77640 142318 77692 142370
rect 77692 142318 77694 142370
rect 77638 142316 77694 142318
rect 79318 142370 79374 142372
rect 79318 142318 79320 142370
rect 79320 142318 79372 142370
rect 79372 142318 79374 142370
rect 79318 142316 79374 142318
rect 80998 142370 81054 142372
rect 80998 142318 81000 142370
rect 81000 142318 81052 142370
rect 81052 142318 81054 142370
rect 80998 142316 81054 142318
rect 82678 142370 82734 142372
rect 82678 142318 82680 142370
rect 82680 142318 82732 142370
rect 82732 142318 82734 142370
rect 82678 142316 82734 142318
rect 84358 142370 84414 142372
rect 84358 142318 84360 142370
rect 84360 142318 84412 142370
rect 84412 142318 84414 142370
rect 84358 142316 84414 142318
rect 86038 142370 86094 142372
rect 86038 142318 86040 142370
rect 86040 142318 86092 142370
rect 86092 142318 86094 142370
rect 86038 142316 86094 142318
rect 87718 142370 87774 142372
rect 87718 142318 87720 142370
rect 87720 142318 87772 142370
rect 87772 142318 87774 142370
rect 87718 142316 87774 142318
rect 89398 142370 89454 142372
rect 89398 142318 89400 142370
rect 89400 142318 89452 142370
rect 89452 142318 89454 142370
rect 89398 142316 89454 142318
rect 91078 142370 91134 142372
rect 91078 142318 91080 142370
rect 91080 142318 91132 142370
rect 91132 142318 91134 142370
rect 91078 142316 91134 142318
rect 92758 142370 92814 142372
rect 92758 142318 92760 142370
rect 92760 142318 92812 142370
rect 92812 142318 92814 142370
rect 92758 142316 92814 142318
rect 94438 142370 94494 142372
rect 94438 142318 94440 142370
rect 94440 142318 94492 142370
rect 94492 142318 94494 142370
rect 94438 142316 94494 142318
rect 96118 142370 96174 142372
rect 96118 142318 96120 142370
rect 96120 142318 96172 142370
rect 96172 142318 96174 142370
rect 96118 142316 96174 142318
rect 97798 142370 97854 142372
rect 97798 142318 97800 142370
rect 97800 142318 97852 142370
rect 97852 142318 97854 142370
rect 97798 142316 97854 142318
rect 99478 142370 99534 142372
rect 99478 142318 99480 142370
rect 99480 142318 99532 142370
rect 99532 142318 99534 142370
rect 99478 142316 99534 142318
rect 101158 142370 101214 142372
rect 101158 142318 101160 142370
rect 101160 142318 101212 142370
rect 101212 142318 101214 142370
rect 101158 142316 101214 142318
rect 102838 142370 102894 142372
rect 102838 142318 102840 142370
rect 102840 142318 102892 142370
rect 102892 142318 102894 142370
rect 102838 142316 102894 142318
rect 104518 142370 104574 142372
rect 104518 142318 104520 142370
rect 104520 142318 104572 142370
rect 104572 142318 104574 142370
rect 104518 142316 104574 142318
rect 106198 142370 106254 142372
rect 106198 142318 106200 142370
rect 106200 142318 106252 142370
rect 106252 142318 106254 142370
rect 106198 142316 106254 142318
rect 107878 142370 107934 142372
rect 107878 142318 107880 142370
rect 107880 142318 107932 142370
rect 107932 142318 107934 142370
rect 107878 142316 107934 142318
rect 109558 142370 109614 142372
rect 109558 142318 109560 142370
rect 109560 142318 109612 142370
rect 109612 142318 109614 142370
rect 109558 142316 109614 142318
rect 111238 142370 111294 142372
rect 111238 142318 111240 142370
rect 111240 142318 111292 142370
rect 111292 142318 111294 142370
rect 111238 142316 111294 142318
rect 112918 142370 112974 142372
rect 112918 142318 112920 142370
rect 112920 142318 112972 142370
rect 112972 142318 112974 142370
rect 112918 142316 112974 142318
rect 114598 142370 114654 142372
rect 114598 142318 114600 142370
rect 114600 142318 114652 142370
rect 114652 142318 114654 142370
rect 114598 142316 114654 142318
rect 116278 142370 116334 142372
rect 116278 142318 116280 142370
rect 116280 142318 116332 142370
rect 116332 142318 116334 142370
rect 116278 142316 116334 142318
rect 117958 142370 118014 142372
rect 117958 142318 117960 142370
rect 117960 142318 118012 142370
rect 118012 142318 118014 142370
rect 117958 142316 118014 142318
rect 119638 142370 119694 142372
rect 119638 142318 119640 142370
rect 119640 142318 119692 142370
rect 119692 142318 119694 142370
rect 119638 142316 119694 142318
rect 121318 142370 121374 142372
rect 121318 142318 121320 142370
rect 121320 142318 121372 142370
rect 121372 142318 121374 142370
rect 121318 142316 121374 142318
rect 122998 142370 123054 142372
rect 122998 142318 123000 142370
rect 123000 142318 123052 142370
rect 123052 142318 123054 142370
rect 122998 142316 123054 142318
rect 124678 142370 124734 142372
rect 124678 142318 124680 142370
rect 124680 142318 124732 142370
rect 124732 142318 124734 142370
rect 124678 142316 124734 142318
rect 126358 142370 126414 142372
rect 126358 142318 126360 142370
rect 126360 142318 126412 142370
rect 126412 142318 126414 142370
rect 126358 142316 126414 142318
rect 128038 142370 128094 142372
rect 128038 142318 128040 142370
rect 128040 142318 128092 142370
rect 128092 142318 128094 142370
rect 128038 142316 128094 142318
rect 129718 142370 129774 142372
rect 129718 142318 129720 142370
rect 129720 142318 129772 142370
rect 129772 142318 129774 142370
rect 129718 142316 129774 142318
rect 131398 142370 131454 142372
rect 131398 142318 131400 142370
rect 131400 142318 131452 142370
rect 131452 142318 131454 142370
rect 131398 142316 131454 142318
rect 133078 142370 133134 142372
rect 133078 142318 133080 142370
rect 133080 142318 133132 142370
rect 133132 142318 133134 142370
rect 133078 142316 133134 142318
rect 134758 142370 134814 142372
rect 134758 142318 134760 142370
rect 134760 142318 134812 142370
rect 134812 142318 134814 142370
rect 134758 142316 134814 142318
rect 136438 142370 136494 142372
rect 136438 142318 136440 142370
rect 136440 142318 136492 142370
rect 136492 142318 136494 142370
rect 136438 142316 136494 142318
rect 138118 142370 138174 142372
rect 138118 142318 138120 142370
rect 138120 142318 138172 142370
rect 138172 142318 138174 142370
rect 138118 142316 138174 142318
rect 139798 142370 139854 142372
rect 139798 142318 139800 142370
rect 139800 142318 139852 142370
rect 139852 142318 139854 142370
rect 139798 142316 139854 142318
rect 141478 142370 141534 142372
rect 141478 142318 141480 142370
rect 141480 142318 141532 142370
rect 141532 142318 141534 142370
rect 141478 142316 141534 142318
rect 143158 142370 143214 142372
rect 143158 142318 143160 142370
rect 143160 142318 143212 142370
rect 143212 142318 143214 142370
rect 143158 142316 143214 142318
rect 144838 142370 144894 142372
rect 144838 142318 144840 142370
rect 144840 142318 144892 142370
rect 144892 142318 144894 142370
rect 144838 142316 144894 142318
rect 146518 142370 146574 142372
rect 146518 142318 146520 142370
rect 146520 142318 146572 142370
rect 146572 142318 146574 142370
rect 146518 142316 146574 142318
rect 148198 142370 148254 142372
rect 148198 142318 148200 142370
rect 148200 142318 148252 142370
rect 148252 142318 148254 142370
rect 148198 142316 148254 142318
rect 149878 142370 149934 142372
rect 149878 142318 149880 142370
rect 149880 142318 149932 142370
rect 149932 142318 149934 142370
rect 149878 142316 149934 142318
rect 151558 142370 151614 142372
rect 151558 142318 151560 142370
rect 151560 142318 151612 142370
rect 151612 142318 151614 142370
rect 151558 142316 151614 142318
rect 153238 142370 153294 142372
rect 153238 142318 153240 142370
rect 153240 142318 153292 142370
rect 153292 142318 153294 142370
rect 153238 142316 153294 142318
rect 154918 142370 154974 142372
rect 154918 142318 154920 142370
rect 154920 142318 154972 142370
rect 154972 142318 154974 142370
rect 154918 142316 154974 142318
rect 156598 142370 156654 142372
rect 156598 142318 156600 142370
rect 156600 142318 156652 142370
rect 156652 142318 156654 142370
rect 156598 142316 156654 142318
rect 158278 142370 158334 142372
rect 158278 142318 158280 142370
rect 158280 142318 158332 142370
rect 158332 142318 158334 142370
rect 158278 142316 158334 142318
rect 159958 142370 160014 142372
rect 159958 142318 159960 142370
rect 159960 142318 160012 142370
rect 160012 142318 160014 142370
rect 159958 142316 160014 142318
rect 161638 142370 161694 142372
rect 161638 142318 161640 142370
rect 161640 142318 161692 142370
rect 161692 142318 161694 142370
rect 161638 142316 161694 142318
rect 163318 142370 163374 142372
rect 163318 142318 163320 142370
rect 163320 142318 163372 142370
rect 163372 142318 163374 142370
rect 163318 142316 163374 142318
rect 164998 142370 165054 142372
rect 164998 142318 165000 142370
rect 165000 142318 165052 142370
rect 165052 142318 165054 142370
rect 164998 142316 165054 142318
rect 166678 142370 166734 142372
rect 166678 142318 166680 142370
rect 166680 142318 166732 142370
rect 166732 142318 166734 142370
rect 166678 142316 166734 142318
rect 168358 142370 168414 142372
rect 168358 142318 168360 142370
rect 168360 142318 168412 142370
rect 168412 142318 168414 142370
rect 168358 142316 168414 142318
rect 170038 142370 170094 142372
rect 170038 142318 170040 142370
rect 170040 142318 170092 142370
rect 170092 142318 170094 142370
rect 170038 142316 170094 142318
rect 171718 142370 171774 142372
rect 171718 142318 171720 142370
rect 171720 142318 171772 142370
rect 171772 142318 171774 142370
rect 171718 142316 171774 142318
rect 173398 142370 173454 142372
rect 173398 142318 173400 142370
rect 173400 142318 173452 142370
rect 173452 142318 173454 142370
rect 173398 142316 173454 142318
rect 175078 142370 175134 142372
rect 175078 142318 175080 142370
rect 175080 142318 175132 142370
rect 175132 142318 175134 142370
rect 175078 142316 175134 142318
rect 176758 142370 176814 142372
rect 176758 142318 176760 142370
rect 176760 142318 176812 142370
rect 176812 142318 176814 142370
rect 176758 142316 176814 142318
rect 178438 142370 178494 142372
rect 178438 142318 178440 142370
rect 178440 142318 178492 142370
rect 178492 142318 178494 142370
rect 178438 142316 178494 142318
rect 180118 142370 180174 142372
rect 180118 142318 180120 142370
rect 180120 142318 180172 142370
rect 180172 142318 180174 142370
rect 180118 142316 180174 142318
rect 181798 142370 181854 142372
rect 181798 142318 181800 142370
rect 181800 142318 181852 142370
rect 181852 142318 181854 142370
rect 181798 142316 181854 142318
rect 183478 142370 183534 142372
rect 183478 142318 183480 142370
rect 183480 142318 183532 142370
rect 183532 142318 183534 142370
rect 183478 142316 183534 142318
rect 185158 142370 185214 142372
rect 185158 142318 185160 142370
rect 185160 142318 185212 142370
rect 185212 142318 185214 142370
rect 185158 142316 185214 142318
rect 186838 142370 186894 142372
rect 186838 142318 186840 142370
rect 186840 142318 186892 142370
rect 186892 142318 186894 142370
rect 186838 142316 186894 142318
rect 188518 142370 188574 142372
rect 188518 142318 188520 142370
rect 188520 142318 188572 142370
rect 188572 142318 188574 142370
rect 188518 142316 188574 142318
rect 190198 142370 190254 142372
rect 190198 142318 190200 142370
rect 190200 142318 190252 142370
rect 190252 142318 190254 142370
rect 190198 142316 190254 142318
rect 191878 142370 191934 142372
rect 191878 142318 191880 142370
rect 191880 142318 191932 142370
rect 191932 142318 191934 142370
rect 191878 142316 191934 142318
rect 193558 142370 193614 142372
rect 193558 142318 193560 142370
rect 193560 142318 193612 142370
rect 193612 142318 193614 142370
rect 193558 142316 193614 142318
rect 195238 142370 195294 142372
rect 195238 142318 195240 142370
rect 195240 142318 195292 142370
rect 195292 142318 195294 142370
rect 195238 142316 195294 142318
rect 196918 142370 196974 142372
rect 196918 142318 196920 142370
rect 196920 142318 196972 142370
rect 196972 142318 196974 142370
rect 196918 142316 196974 142318
rect 198598 142370 198654 142372
rect 198598 142318 198600 142370
rect 198600 142318 198652 142370
rect 198652 142318 198654 142370
rect 198598 142316 198654 142318
rect 200278 142370 200334 142372
rect 200278 142318 200280 142370
rect 200280 142318 200332 142370
rect 200332 142318 200334 142370
rect 200278 142316 200334 142318
rect 201958 142370 202014 142372
rect 201958 142318 201960 142370
rect 201960 142318 202012 142370
rect 202012 142318 202014 142370
rect 201958 142316 202014 142318
rect 203638 142370 203694 142372
rect 203638 142318 203640 142370
rect 203640 142318 203692 142370
rect 203692 142318 203694 142370
rect 203638 142316 203694 142318
rect 205318 142370 205374 142372
rect 205318 142318 205320 142370
rect 205320 142318 205372 142370
rect 205372 142318 205374 142370
rect 205318 142316 205374 142318
rect 206998 142370 207054 142372
rect 206998 142318 207000 142370
rect 207000 142318 207052 142370
rect 207052 142318 207054 142370
rect 206998 142316 207054 142318
rect 208678 142370 208734 142372
rect 208678 142318 208680 142370
rect 208680 142318 208732 142370
rect 208732 142318 208734 142370
rect 208678 142316 208734 142318
rect 210358 142370 210414 142372
rect 210358 142318 210360 142370
rect 210360 142318 210412 142370
rect 210412 142318 210414 142370
rect 210358 142316 210414 142318
rect 212038 142370 212094 142372
rect 212038 142318 212040 142370
rect 212040 142318 212092 142370
rect 212092 142318 212094 142370
rect 212038 142316 212094 142318
rect 213718 142370 213774 142372
rect 213718 142318 213720 142370
rect 213720 142318 213772 142370
rect 213772 142318 213774 142370
rect 213718 142316 213774 142318
rect 215398 142370 215454 142372
rect 215398 142318 215400 142370
rect 215400 142318 215452 142370
rect 215452 142318 215454 142370
rect 215398 142316 215454 142318
rect 203400 141672 203456 141728
rect 1702 141650 1758 141652
rect 1702 141598 1704 141650
rect 1704 141598 1756 141650
rect 1756 141598 1758 141650
rect 1702 141596 1758 141598
rect 198642 141416 198698 141472
rect 199810 141416 199866 141472
rect 200978 141416 201034 141472
rect 1702 139970 1758 139972
rect 1702 139918 1704 139970
rect 1704 139918 1756 139970
rect 1756 139918 1758 139970
rect 1702 139916 1758 139918
rect 1702 138290 1758 138292
rect 1702 138238 1704 138290
rect 1704 138238 1756 138290
rect 1756 138238 1758 138290
rect 1702 138236 1758 138238
rect 1702 136610 1758 136612
rect 1702 136558 1704 136610
rect 1704 136558 1756 136610
rect 1756 136558 1758 136610
rect 1702 136556 1758 136558
rect 1702 134930 1758 134932
rect 1702 134878 1704 134930
rect 1704 134878 1756 134930
rect 1756 134878 1758 134930
rect 1702 134876 1758 134878
rect 1702 133250 1758 133252
rect 1702 133198 1704 133250
rect 1704 133198 1756 133250
rect 1756 133198 1758 133250
rect 1702 133196 1758 133198
rect 216908 141650 216964 141652
rect 216908 141598 216910 141650
rect 216910 141598 216962 141650
rect 216962 141598 216964 141650
rect 216908 141596 216964 141598
rect 216908 139970 216964 139972
rect 216908 139918 216910 139970
rect 216910 139918 216962 139970
rect 216962 139918 216964 139970
rect 216908 139916 216964 139918
rect 216908 138290 216964 138292
rect 216908 138238 216910 138290
rect 216910 138238 216962 138290
rect 216962 138238 216964 138290
rect 216908 138236 216964 138238
rect 216908 136610 216964 136612
rect 216908 136558 216910 136610
rect 216910 136558 216962 136610
rect 216962 136558 216964 136610
rect 216908 136556 216964 136558
rect 216908 134930 216964 134932
rect 216908 134878 216910 134930
rect 216910 134878 216962 134930
rect 216962 134878 216964 134930
rect 216908 134876 216964 134878
rect 216284 134763 216340 134819
rect 213183 134658 213239 134714
rect 29560 133092 29616 133094
rect 29560 133040 29562 133092
rect 29562 133040 29614 133092
rect 29614 133040 29616 133092
rect 29560 133038 29616 133040
rect 34552 133092 34608 133094
rect 34552 133040 34554 133092
rect 34554 133040 34606 133092
rect 34606 133040 34608 133092
rect 34552 133038 34608 133040
rect 39544 133092 39600 133094
rect 39544 133040 39546 133092
rect 39546 133040 39598 133092
rect 39598 133040 39600 133092
rect 39544 133038 39600 133040
rect 44536 133092 44592 133094
rect 44536 133040 44538 133092
rect 44538 133040 44590 133092
rect 44590 133040 44592 133092
rect 44536 133038 44592 133040
rect 49528 133092 49584 133094
rect 49528 133040 49530 133092
rect 49530 133040 49582 133092
rect 49582 133040 49584 133092
rect 49528 133038 49584 133040
rect 54520 133092 54576 133094
rect 54520 133040 54522 133092
rect 54522 133040 54574 133092
rect 54574 133040 54576 133092
rect 54520 133038 54576 133040
rect 59512 133092 59568 133094
rect 59512 133040 59514 133092
rect 59514 133040 59566 133092
rect 59566 133040 59568 133092
rect 59512 133038 59568 133040
rect 64504 133092 64560 133094
rect 64504 133040 64506 133092
rect 64506 133040 64558 133092
rect 64558 133040 64560 133092
rect 64504 133038 64560 133040
rect 69496 133092 69552 133094
rect 69496 133040 69498 133092
rect 69498 133040 69550 133092
rect 69550 133040 69552 133092
rect 69496 133038 69552 133040
rect 74488 133092 74544 133094
rect 74488 133040 74490 133092
rect 74490 133040 74542 133092
rect 74542 133040 74544 133092
rect 74488 133038 74544 133040
rect 79480 133092 79536 133094
rect 79480 133040 79482 133092
rect 79482 133040 79534 133092
rect 79534 133040 79536 133092
rect 79480 133038 79536 133040
rect 84472 133092 84528 133094
rect 84472 133040 84474 133092
rect 84474 133040 84526 133092
rect 84526 133040 84528 133092
rect 84472 133038 84528 133040
rect 89464 133092 89520 133094
rect 89464 133040 89466 133092
rect 89466 133040 89518 133092
rect 89518 133040 89520 133092
rect 89464 133038 89520 133040
rect 94456 133092 94512 133094
rect 94456 133040 94458 133092
rect 94458 133040 94510 133092
rect 94510 133040 94512 133092
rect 94456 133038 94512 133040
rect 99448 133092 99504 133094
rect 99448 133040 99450 133092
rect 99450 133040 99502 133092
rect 99502 133040 99504 133092
rect 99448 133038 99504 133040
rect 104440 133092 104496 133094
rect 104440 133040 104442 133092
rect 104442 133040 104494 133092
rect 104494 133040 104496 133092
rect 104440 133038 104496 133040
rect 109432 133092 109488 133094
rect 109432 133040 109434 133092
rect 109434 133040 109486 133092
rect 109486 133040 109488 133092
rect 109432 133038 109488 133040
rect 114424 133092 114480 133094
rect 114424 133040 114426 133092
rect 114426 133040 114478 133092
rect 114478 133040 114480 133092
rect 114424 133038 114480 133040
rect 119416 133092 119472 133094
rect 119416 133040 119418 133092
rect 119418 133040 119470 133092
rect 119470 133040 119472 133092
rect 119416 133038 119472 133040
rect 124408 133092 124464 133094
rect 124408 133040 124410 133092
rect 124410 133040 124462 133092
rect 124462 133040 124464 133092
rect 124408 133038 124464 133040
rect 129400 133092 129456 133094
rect 129400 133040 129402 133092
rect 129402 133040 129454 133092
rect 129454 133040 129456 133092
rect 129400 133038 129456 133040
rect 134392 133092 134448 133094
rect 134392 133040 134394 133092
rect 134394 133040 134446 133092
rect 134446 133040 134448 133092
rect 134392 133038 134448 133040
rect 139384 133092 139440 133094
rect 139384 133040 139386 133092
rect 139386 133040 139438 133092
rect 139438 133040 139440 133092
rect 139384 133038 139440 133040
rect 144376 133092 144432 133094
rect 144376 133040 144378 133092
rect 144378 133040 144430 133092
rect 144430 133040 144432 133092
rect 144376 133038 144432 133040
rect 149368 133092 149424 133094
rect 149368 133040 149370 133092
rect 149370 133040 149422 133092
rect 149422 133040 149424 133092
rect 149368 133038 149424 133040
rect 154360 133092 154416 133094
rect 154360 133040 154362 133092
rect 154362 133040 154414 133092
rect 154414 133040 154416 133092
rect 154360 133038 154416 133040
rect 159352 133092 159408 133094
rect 159352 133040 159354 133092
rect 159354 133040 159406 133092
rect 159406 133040 159408 133092
rect 159352 133038 159408 133040
rect 164344 133092 164400 133094
rect 164344 133040 164346 133092
rect 164346 133040 164398 133092
rect 164398 133040 164400 133092
rect 164344 133038 164400 133040
rect 169336 133092 169392 133094
rect 169336 133040 169338 133092
rect 169338 133040 169390 133092
rect 169390 133040 169392 133092
rect 169336 133038 169392 133040
rect 174328 133092 174384 133094
rect 174328 133040 174330 133092
rect 174330 133040 174382 133092
rect 174382 133040 174384 133092
rect 174328 133038 174384 133040
rect 179320 133092 179376 133094
rect 179320 133040 179322 133092
rect 179322 133040 179374 133092
rect 179374 133040 179376 133092
rect 179320 133038 179376 133040
rect 184312 133092 184368 133094
rect 184312 133040 184314 133092
rect 184314 133040 184366 133092
rect 184366 133040 184368 133092
rect 184312 133038 184368 133040
rect 1702 131570 1758 131572
rect 1702 131518 1704 131570
rect 1704 131518 1756 131570
rect 1756 131518 1758 131570
rect 1702 131516 1758 131518
rect 190875 130378 190931 130434
rect 1702 129890 1758 129892
rect 1702 129838 1704 129890
rect 1704 129838 1756 129890
rect 1756 129838 1758 129890
rect 1702 129836 1758 129838
rect 1702 128210 1758 128212
rect 1702 128158 1704 128210
rect 1704 128158 1756 128210
rect 1756 128158 1758 128210
rect 1702 128156 1758 128158
rect 190999 128964 191055 129020
rect 194858 127550 194914 127606
rect 1702 126530 1758 126532
rect 1702 126478 1704 126530
rect 1704 126478 1756 126530
rect 1756 126478 1758 126530
rect 1702 126476 1758 126478
rect 1702 124850 1758 124852
rect 1702 124798 1704 124850
rect 1704 124798 1756 124850
rect 1756 124798 1758 124850
rect 1702 124796 1758 124798
rect 1702 123170 1758 123172
rect 1702 123118 1704 123170
rect 1704 123118 1756 123170
rect 1756 123118 1758 123170
rect 1702 123116 1758 123118
rect 1702 121490 1758 121492
rect 1702 121438 1704 121490
rect 1704 121438 1756 121490
rect 1756 121438 1758 121490
rect 1702 121436 1758 121438
rect 1702 119810 1758 119812
rect 1702 119758 1704 119810
rect 1704 119758 1756 119810
rect 1756 119758 1758 119810
rect 1702 119756 1758 119758
rect 1702 118130 1758 118132
rect 1702 118078 1704 118130
rect 1704 118078 1756 118130
rect 1756 118078 1758 118130
rect 1702 118076 1758 118078
rect 1702 116450 1758 116452
rect 1702 116398 1704 116450
rect 1704 116398 1756 116450
rect 1756 116398 1758 116450
rect 1702 116396 1758 116398
rect 1702 114770 1758 114772
rect 1702 114718 1704 114770
rect 1704 114718 1756 114770
rect 1756 114718 1758 114770
rect 1702 114716 1758 114718
rect 1702 113090 1758 113092
rect 1702 113038 1704 113090
rect 1704 113038 1756 113090
rect 1756 113038 1758 113090
rect 1702 113036 1758 113038
rect 1702 111410 1758 111412
rect 1702 111358 1704 111410
rect 1704 111358 1756 111410
rect 1756 111358 1758 111410
rect 1702 111356 1758 111358
rect 1702 109730 1758 109732
rect 1702 109678 1704 109730
rect 1704 109678 1756 109730
rect 1756 109678 1758 109730
rect 1702 109676 1758 109678
rect 1702 108050 1758 108052
rect 1702 107998 1704 108050
rect 1704 107998 1756 108050
rect 1756 107998 1758 108050
rect 1702 107996 1758 107998
rect 1702 106370 1758 106372
rect 1702 106318 1704 106370
rect 1704 106318 1756 106370
rect 1756 106318 1758 106370
rect 1702 106316 1758 106318
rect 1702 104690 1758 104692
rect 1702 104638 1704 104690
rect 1704 104638 1756 104690
rect 1756 104638 1758 104690
rect 1702 104636 1758 104638
rect 1702 103010 1758 103012
rect 1702 102958 1704 103010
rect 1704 102958 1756 103010
rect 1756 102958 1758 103010
rect 1702 102956 1758 102958
rect 1702 101330 1758 101332
rect 1702 101278 1704 101330
rect 1704 101278 1756 101330
rect 1756 101278 1758 101330
rect 1702 101276 1758 101278
rect 1702 99650 1758 99652
rect 1702 99598 1704 99650
rect 1704 99598 1756 99650
rect 1756 99598 1758 99650
rect 1702 99596 1758 99598
rect 1702 97970 1758 97972
rect 1702 97918 1704 97970
rect 1704 97918 1756 97970
rect 1756 97918 1758 97970
rect 1702 97916 1758 97918
rect 1702 96290 1758 96292
rect 1702 96238 1704 96290
rect 1704 96238 1756 96290
rect 1756 96238 1758 96290
rect 1702 96236 1758 96238
rect 1702 94610 1758 94612
rect 1702 94558 1704 94610
rect 1704 94558 1756 94610
rect 1756 94558 1758 94610
rect 1702 94556 1758 94558
rect 1702 92930 1758 92932
rect 1702 92878 1704 92930
rect 1704 92878 1756 92930
rect 1756 92878 1758 92930
rect 1702 92876 1758 92878
rect 1702 91250 1758 91252
rect 1702 91198 1704 91250
rect 1704 91198 1756 91250
rect 1756 91198 1758 91250
rect 1702 91196 1758 91198
rect 1702 89570 1758 89572
rect 1702 89518 1704 89570
rect 1704 89518 1756 89570
rect 1756 89518 1758 89570
rect 1702 89516 1758 89518
rect 1702 87890 1758 87892
rect 1702 87838 1704 87890
rect 1704 87838 1756 87890
rect 1756 87838 1758 87890
rect 1702 87836 1758 87838
rect 1702 86210 1758 86212
rect 1702 86158 1704 86210
rect 1704 86158 1756 86210
rect 1756 86158 1758 86210
rect 1702 86156 1758 86158
rect 1702 84530 1758 84532
rect 1702 84478 1704 84530
rect 1704 84478 1756 84530
rect 1756 84478 1758 84530
rect 1702 84476 1758 84478
rect 1702 82850 1758 82852
rect 1702 82798 1704 82850
rect 1704 82798 1756 82850
rect 1756 82798 1758 82850
rect 1702 82796 1758 82798
rect 1702 81170 1758 81172
rect 1702 81118 1704 81170
rect 1704 81118 1756 81170
rect 1756 81118 1758 81170
rect 1702 81116 1758 81118
rect 1702 79490 1758 79492
rect 1702 79438 1704 79490
rect 1704 79438 1756 79490
rect 1756 79438 1758 79490
rect 1702 79436 1758 79438
rect 1702 77810 1758 77812
rect 1702 77758 1704 77810
rect 1704 77758 1756 77810
rect 1756 77758 1758 77810
rect 1702 77756 1758 77758
rect 1702 76130 1758 76132
rect 1702 76078 1704 76130
rect 1704 76078 1756 76130
rect 1756 76078 1758 76130
rect 1702 76076 1758 76078
rect 1702 74450 1758 74452
rect 1702 74398 1704 74450
rect 1704 74398 1756 74450
rect 1756 74398 1758 74450
rect 1702 74396 1758 74398
rect 1702 72770 1758 72772
rect 1702 72718 1704 72770
rect 1704 72718 1756 72770
rect 1756 72718 1758 72770
rect 1702 72716 1758 72718
rect 1702 71090 1758 71092
rect 1702 71038 1704 71090
rect 1704 71038 1756 71090
rect 1756 71038 1758 71090
rect 1702 71036 1758 71038
rect 1702 69410 1758 69412
rect 1702 69358 1704 69410
rect 1704 69358 1756 69410
rect 1756 69358 1758 69410
rect 1702 69356 1758 69358
rect 1702 67730 1758 67732
rect 1702 67678 1704 67730
rect 1704 67678 1756 67730
rect 1756 67678 1758 67730
rect 1702 67676 1758 67678
rect 1702 66050 1758 66052
rect 1702 65998 1704 66050
rect 1704 65998 1756 66050
rect 1756 65998 1758 66050
rect 1702 65996 1758 65998
rect 1702 64370 1758 64372
rect 1702 64318 1704 64370
rect 1704 64318 1756 64370
rect 1756 64318 1758 64370
rect 1702 64316 1758 64318
rect 1702 62690 1758 62692
rect 1702 62638 1704 62690
rect 1704 62638 1756 62690
rect 1756 62638 1758 62690
rect 1702 62636 1758 62638
rect 1702 61010 1758 61012
rect 1702 60958 1704 61010
rect 1704 60958 1756 61010
rect 1756 60958 1758 61010
rect 1702 60956 1758 60958
rect 1702 59330 1758 59332
rect 1702 59278 1704 59330
rect 1704 59278 1756 59330
rect 1756 59278 1758 59330
rect 1702 59276 1758 59278
rect 1702 57650 1758 57652
rect 1702 57598 1704 57650
rect 1704 57598 1756 57650
rect 1756 57598 1758 57650
rect 1702 57596 1758 57598
rect 1702 55970 1758 55972
rect 1702 55918 1704 55970
rect 1704 55918 1756 55970
rect 1756 55918 1758 55970
rect 1702 55916 1758 55918
rect 1702 54290 1758 54292
rect 1702 54238 1704 54290
rect 1704 54238 1756 54290
rect 1756 54238 1758 54290
rect 1702 54236 1758 54238
rect 1702 52610 1758 52612
rect 1702 52558 1704 52610
rect 1704 52558 1756 52610
rect 1756 52558 1758 52610
rect 1702 52556 1758 52558
rect 1702 50930 1758 50932
rect 1702 50878 1704 50930
rect 1704 50878 1756 50930
rect 1756 50878 1758 50930
rect 1702 50876 1758 50878
rect 1702 49250 1758 49252
rect 1702 49198 1704 49250
rect 1704 49198 1756 49250
rect 1756 49198 1758 49250
rect 1702 49196 1758 49198
rect 1702 47570 1758 47572
rect 1702 47518 1704 47570
rect 1704 47518 1756 47570
rect 1756 47518 1758 47570
rect 1702 47516 1758 47518
rect 1702 45890 1758 45892
rect 1702 45838 1704 45890
rect 1704 45838 1756 45890
rect 1756 45838 1758 45890
rect 1702 45836 1758 45838
rect 14212 45037 14268 45093
rect 15157 44966 15213 45022
rect 15971 45020 16027 45022
rect 15971 44968 15973 45020
rect 15973 44968 16025 45020
rect 16025 44968 16027 45020
rect 15971 44966 16027 44968
rect 1702 44210 1758 44212
rect 1702 44158 1704 44210
rect 1704 44158 1756 44210
rect 1756 44158 1758 44210
rect 1702 44156 1758 44158
rect 15157 43408 15213 43464
rect 15891 43462 15947 43464
rect 15891 43410 15893 43462
rect 15893 43410 15945 43462
rect 15945 43410 15947 43462
rect 15891 43408 15947 43410
rect 14212 43337 14268 43393
rect 1702 42530 1758 42532
rect 1702 42478 1704 42530
rect 1704 42478 1756 42530
rect 1756 42478 1758 42530
rect 1702 42476 1758 42478
rect 14212 42209 14268 42265
rect 15157 42138 15213 42194
rect 15811 42192 15867 42194
rect 15811 42140 15813 42192
rect 15813 42140 15865 42192
rect 15865 42140 15867 42192
rect 15811 42138 15867 42140
rect 1702 40850 1758 40852
rect 1702 40798 1704 40850
rect 1704 40798 1756 40850
rect 1756 40798 1758 40850
rect 1702 40796 1758 40798
rect 15157 40580 15213 40636
rect 15731 40634 15787 40636
rect 15731 40582 15733 40634
rect 15733 40582 15785 40634
rect 15785 40582 15787 40634
rect 15731 40580 15787 40582
rect 14212 40509 14268 40565
rect 14212 39381 14268 39437
rect 15157 39310 15213 39366
rect 15651 39364 15707 39366
rect 15651 39312 15653 39364
rect 15653 39312 15705 39364
rect 15705 39312 15707 39364
rect 15651 39310 15707 39312
rect 1702 39170 1758 39172
rect 1702 39118 1704 39170
rect 1704 39118 1756 39170
rect 1756 39118 1758 39170
rect 1702 39116 1758 39118
rect 15157 37752 15213 37808
rect 15571 37806 15627 37808
rect 15571 37754 15573 37806
rect 15573 37754 15625 37806
rect 15625 37754 15627 37806
rect 15571 37752 15627 37754
rect 14212 37681 14268 37737
rect 1702 37490 1758 37492
rect 1702 37438 1704 37490
rect 1704 37438 1756 37490
rect 1756 37438 1758 37490
rect 1702 37436 1758 37438
rect 14212 36553 14268 36609
rect 15157 36482 15213 36538
rect 15491 36536 15547 36538
rect 15491 36484 15493 36536
rect 15493 36484 15545 36536
rect 15545 36484 15547 36536
rect 15491 36482 15547 36484
rect 1702 35810 1758 35812
rect 1702 35758 1704 35810
rect 1704 35758 1756 35810
rect 1756 35758 1758 35810
rect 1702 35756 1758 35758
rect 15157 34924 15213 34980
rect 15411 34978 15467 34980
rect 15411 34926 15413 34978
rect 15413 34926 15465 34978
rect 15465 34926 15467 34978
rect 15411 34924 15467 34926
rect 14212 34853 14268 34909
rect 15294 34597 15350 34653
rect 1702 34130 1758 34132
rect 1702 34078 1704 34130
rect 1704 34078 1756 34130
rect 1756 34078 1758 34130
rect 1702 34076 1758 34078
rect 1702 32450 1758 32452
rect 1702 32398 1704 32450
rect 1704 32398 1756 32450
rect 1756 32398 1758 32450
rect 1702 32396 1758 32398
rect 1702 30770 1758 30772
rect 1702 30718 1704 30770
rect 1704 30718 1756 30770
rect 1756 30718 1758 30770
rect 1702 30716 1758 30718
rect 2113 30296 2169 30352
rect 1702 29090 1758 29092
rect 1702 29038 1704 29090
rect 1704 29038 1756 29090
rect 1756 29038 1758 29090
rect 1702 29036 1758 29038
rect 1702 27410 1758 27412
rect 1702 27358 1704 27410
rect 1704 27358 1756 27410
rect 1756 27358 1758 27410
rect 1702 27356 1758 27358
rect 1702 25730 1758 25732
rect 1702 25678 1704 25730
rect 1704 25678 1756 25730
rect 1756 25678 1758 25730
rect 1702 25676 1758 25678
rect 1702 24050 1758 24052
rect 1702 23998 1704 24050
rect 1704 23998 1756 24050
rect 1756 23998 1758 24050
rect 1702 23996 1758 23998
rect 15210 23188 15266 23244
rect 1702 22370 1758 22372
rect 1702 22318 1704 22370
rect 1704 22318 1756 22370
rect 1756 22318 1758 22370
rect 1702 22316 1758 22318
rect 1702 20690 1758 20692
rect 1702 20638 1704 20690
rect 1704 20638 1756 20690
rect 1756 20638 1758 20690
rect 1702 20636 1758 20638
rect 15210 20360 15266 20416
rect 1702 19010 1758 19012
rect 1702 18958 1704 19010
rect 1704 18958 1756 19010
rect 1756 18958 1758 19010
rect 1702 18956 1758 18958
rect 15210 18946 15266 19002
rect 15210 17532 15266 17588
rect 1702 17330 1758 17332
rect 1702 17278 1704 17330
rect 1704 17278 1756 17330
rect 1756 17278 1758 17330
rect 1702 17276 1758 17278
rect 1702 15650 1758 15652
rect 1702 15598 1704 15650
rect 1704 15598 1756 15650
rect 1756 15598 1758 15650
rect 1702 15596 1758 15598
rect 2326 14847 2382 14903
rect 1702 13970 1758 13972
rect 1702 13918 1704 13970
rect 1704 13918 1756 13970
rect 1756 13918 1758 13970
rect 1702 13916 1758 13918
rect 216908 133250 216964 133252
rect 216908 133198 216910 133250
rect 216910 133198 216962 133250
rect 216962 133198 216964 133250
rect 216908 133196 216964 133198
rect 216908 131570 216964 131572
rect 216908 131518 216910 131570
rect 216910 131518 216962 131570
rect 216962 131518 216964 131570
rect 216908 131516 216964 131518
rect 203484 130378 203540 130434
rect 216908 129890 216964 129892
rect 216908 129838 216910 129890
rect 216910 129838 216962 129890
rect 216962 129838 216964 129890
rect 216908 129836 216964 129838
rect 203484 128964 203540 129020
rect 216908 128210 216964 128212
rect 216908 128158 216910 128210
rect 216910 128158 216962 128210
rect 216962 128158 216964 128210
rect 216908 128156 216964 128158
rect 203484 127550 203540 127606
rect 216908 126530 216964 126532
rect 216908 126478 216910 126530
rect 216910 126478 216962 126530
rect 216962 126478 216964 126530
rect 216908 126476 216964 126478
rect 216908 124850 216964 124852
rect 216908 124798 216910 124850
rect 216910 124798 216962 124850
rect 216962 124798 216964 124850
rect 216908 124796 216964 124798
rect 216908 123170 216964 123172
rect 216908 123118 216910 123170
rect 216910 123118 216962 123170
rect 216962 123118 216964 123170
rect 216908 123116 216964 123118
rect 216908 121490 216964 121492
rect 216908 121438 216910 121490
rect 216910 121438 216962 121490
rect 216962 121438 216964 121490
rect 216908 121436 216964 121438
rect 216908 119810 216964 119812
rect 216908 119758 216910 119810
rect 216910 119758 216962 119810
rect 216962 119758 216964 119810
rect 216908 119756 216964 119758
rect 216908 118130 216964 118132
rect 216908 118078 216910 118130
rect 216910 118078 216962 118130
rect 216962 118078 216964 118130
rect 216908 118076 216964 118078
rect 216497 117614 216553 117670
rect 216908 116450 216964 116452
rect 216908 116398 216910 116450
rect 216910 116398 216962 116450
rect 216962 116398 216964 116450
rect 216908 116396 216964 116398
rect 216908 114770 216964 114772
rect 216908 114718 216910 114770
rect 216910 114718 216962 114770
rect 216962 114718 216964 114770
rect 216908 114716 216964 114718
rect 216908 113090 216964 113092
rect 216908 113038 216910 113090
rect 216910 113038 216962 113090
rect 216962 113038 216964 113090
rect 216908 113036 216964 113038
rect 216908 111410 216964 111412
rect 216908 111358 216910 111410
rect 216910 111358 216962 111410
rect 216962 111358 216964 111410
rect 216908 111356 216964 111358
rect 216908 109730 216964 109732
rect 216908 109678 216910 109730
rect 216910 109678 216962 109730
rect 216962 109678 216964 109730
rect 216908 109676 216964 109678
rect 216908 108050 216964 108052
rect 216908 107998 216910 108050
rect 216910 107998 216962 108050
rect 216962 107998 216964 108050
rect 216908 107996 216964 107998
rect 216908 106370 216964 106372
rect 216908 106318 216910 106370
rect 216910 106318 216962 106370
rect 216962 106318 216964 106370
rect 216908 106316 216964 106318
rect 216908 104690 216964 104692
rect 216908 104638 216910 104690
rect 216910 104638 216962 104690
rect 216962 104638 216964 104690
rect 216908 104636 216964 104638
rect 216908 103010 216964 103012
rect 216908 102958 216910 103010
rect 216910 102958 216962 103010
rect 216962 102958 216964 103010
rect 216908 102956 216964 102958
rect 216908 101330 216964 101332
rect 216908 101278 216910 101330
rect 216910 101278 216962 101330
rect 216962 101278 216964 101330
rect 216908 101276 216964 101278
rect 216908 99650 216964 99652
rect 216908 99598 216910 99650
rect 216910 99598 216962 99650
rect 216962 99598 216964 99650
rect 216908 99596 216964 99598
rect 216908 97970 216964 97972
rect 216908 97918 216910 97970
rect 216910 97918 216962 97970
rect 216962 97918 216964 97970
rect 216908 97916 216964 97918
rect 216908 96290 216964 96292
rect 216908 96238 216910 96290
rect 216910 96238 216962 96290
rect 216962 96238 216964 96290
rect 216908 96236 216964 96238
rect 216908 94610 216964 94612
rect 216908 94558 216910 94610
rect 216910 94558 216962 94610
rect 216962 94558 216964 94610
rect 216908 94556 216964 94558
rect 216908 92930 216964 92932
rect 216908 92878 216910 92930
rect 216910 92878 216962 92930
rect 216962 92878 216964 92930
rect 216908 92876 216964 92878
rect 216908 91250 216964 91252
rect 216908 91198 216910 91250
rect 216910 91198 216962 91250
rect 216962 91198 216964 91250
rect 216908 91196 216964 91198
rect 216908 89570 216964 89572
rect 216908 89518 216910 89570
rect 216910 89518 216962 89570
rect 216962 89518 216964 89570
rect 216908 89516 216964 89518
rect 216908 87890 216964 87892
rect 216908 87838 216910 87890
rect 216910 87838 216962 87890
rect 216962 87838 216964 87890
rect 216908 87836 216964 87838
rect 216908 86210 216964 86212
rect 216908 86158 216910 86210
rect 216910 86158 216962 86210
rect 216962 86158 216964 86210
rect 216908 86156 216964 86158
rect 216908 84530 216964 84532
rect 216908 84478 216910 84530
rect 216910 84478 216962 84530
rect 216962 84478 216964 84530
rect 216908 84476 216964 84478
rect 216908 82850 216964 82852
rect 216908 82798 216910 82850
rect 216910 82798 216962 82850
rect 216962 82798 216964 82850
rect 216908 82796 216964 82798
rect 216908 81170 216964 81172
rect 216908 81118 216910 81170
rect 216910 81118 216962 81170
rect 216962 81118 216964 81170
rect 216908 81116 216964 81118
rect 216908 79490 216964 79492
rect 216908 79438 216910 79490
rect 216910 79438 216962 79490
rect 216962 79438 216964 79490
rect 216908 79436 216964 79438
rect 216908 77810 216964 77812
rect 216908 77758 216910 77810
rect 216910 77758 216962 77810
rect 216962 77758 216964 77810
rect 216908 77756 216964 77758
rect 216908 76130 216964 76132
rect 216908 76078 216910 76130
rect 216910 76078 216962 76130
rect 216962 76078 216964 76130
rect 216908 76076 216964 76078
rect 216908 74450 216964 74452
rect 216908 74398 216910 74450
rect 216910 74398 216962 74450
rect 216962 74398 216964 74450
rect 216908 74396 216964 74398
rect 216908 72770 216964 72772
rect 216908 72718 216910 72770
rect 216910 72718 216962 72770
rect 216962 72718 216964 72770
rect 216908 72716 216964 72718
rect 216908 71090 216964 71092
rect 216908 71038 216910 71090
rect 216910 71038 216962 71090
rect 216962 71038 216964 71090
rect 216908 71036 216964 71038
rect 216908 69410 216964 69412
rect 216908 69358 216910 69410
rect 216910 69358 216962 69410
rect 216962 69358 216964 69410
rect 216908 69356 216964 69358
rect 216908 67730 216964 67732
rect 216908 67678 216910 67730
rect 216910 67678 216962 67730
rect 216962 67678 216964 67730
rect 216908 67676 216964 67678
rect 216908 66050 216964 66052
rect 216908 65998 216910 66050
rect 216910 65998 216962 66050
rect 216962 65998 216964 66050
rect 216908 65996 216964 65998
rect 216908 64370 216964 64372
rect 216908 64318 216910 64370
rect 216910 64318 216962 64370
rect 216962 64318 216964 64370
rect 216908 64316 216964 64318
rect 216908 62690 216964 62692
rect 216908 62638 216910 62690
rect 216910 62638 216962 62690
rect 216962 62638 216964 62690
rect 216908 62636 216964 62638
rect 216908 61010 216964 61012
rect 216908 60958 216910 61010
rect 216910 60958 216962 61010
rect 216962 60958 216964 61010
rect 216908 60956 216964 60958
rect 216908 59330 216964 59332
rect 216908 59278 216910 59330
rect 216910 59278 216962 59330
rect 216962 59278 216964 59330
rect 216908 59276 216964 59278
rect 216908 57650 216964 57652
rect 216908 57598 216910 57650
rect 216910 57598 216962 57650
rect 216962 57598 216964 57650
rect 216908 57596 216964 57598
rect 216908 55970 216964 55972
rect 216908 55918 216910 55970
rect 216910 55918 216962 55970
rect 216962 55918 216964 55970
rect 216908 55916 216964 55918
rect 216908 54290 216964 54292
rect 216908 54238 216910 54290
rect 216910 54238 216962 54290
rect 216962 54238 216964 54290
rect 216908 54236 216964 54238
rect 216908 52610 216964 52612
rect 216908 52558 216910 52610
rect 216910 52558 216962 52610
rect 216962 52558 216964 52610
rect 216908 52556 216964 52558
rect 216908 50930 216964 50932
rect 216908 50878 216910 50930
rect 216910 50878 216962 50930
rect 216962 50878 216964 50930
rect 216908 50876 216964 50878
rect 216908 49250 216964 49252
rect 216908 49198 216910 49250
rect 216910 49198 216962 49250
rect 216962 49198 216964 49250
rect 216908 49196 216964 49198
rect 216908 47570 216964 47572
rect 216908 47518 216910 47570
rect 216910 47518 216962 47570
rect 216962 47518 216964 47570
rect 216908 47516 216964 47518
rect 216908 45890 216964 45892
rect 216908 45838 216910 45890
rect 216910 45838 216962 45890
rect 216962 45838 216964 45890
rect 216908 45836 216964 45838
rect 216908 44210 216964 44212
rect 216908 44158 216910 44210
rect 216910 44158 216962 44210
rect 216962 44158 216964 44210
rect 216908 44156 216964 44158
rect 216908 42530 216964 42532
rect 216908 42478 216910 42530
rect 216910 42478 216962 42530
rect 216962 42478 216964 42530
rect 216908 42476 216964 42478
rect 216908 40850 216964 40852
rect 216908 40798 216910 40850
rect 216910 40798 216962 40850
rect 216962 40798 216964 40850
rect 216908 40796 216964 40798
rect 216908 39170 216964 39172
rect 216908 39118 216910 39170
rect 216910 39118 216962 39170
rect 216962 39118 216964 39170
rect 216908 39116 216964 39118
rect 216908 37490 216964 37492
rect 216908 37438 216910 37490
rect 216910 37438 216962 37490
rect 216962 37438 216964 37490
rect 216908 37436 216964 37438
rect 216908 35810 216964 35812
rect 216908 35758 216910 35810
rect 216910 35758 216962 35810
rect 216962 35758 216964 35810
rect 216908 35756 216964 35758
rect 216908 34130 216964 34132
rect 216908 34078 216910 34130
rect 216910 34078 216962 34130
rect 216962 34078 216964 34130
rect 216908 34076 216964 34078
rect 216908 32450 216964 32452
rect 216908 32398 216910 32450
rect 216910 32398 216962 32450
rect 216962 32398 216964 32450
rect 216908 32396 216964 32398
rect 216908 30770 216964 30772
rect 216908 30718 216910 30770
rect 216910 30718 216962 30770
rect 216962 30718 216964 30770
rect 216908 30716 216964 30718
rect 216908 29090 216964 29092
rect 216908 29038 216910 29090
rect 216910 29038 216962 29090
rect 216962 29038 216964 29090
rect 216908 29036 216964 29038
rect 216908 27410 216964 27412
rect 216908 27358 216910 27410
rect 216910 27358 216962 27410
rect 216962 27358 216964 27410
rect 216908 27356 216964 27358
rect 216908 25730 216964 25732
rect 216908 25678 216910 25730
rect 216910 25678 216962 25730
rect 216962 25678 216964 25730
rect 216908 25676 216964 25678
rect 203400 24501 203456 24557
rect 204482 24245 204538 24301
rect 203199 24228 203255 24230
rect 203199 24176 203201 24228
rect 203201 24176 203253 24228
rect 203253 24176 203255 24228
rect 203199 24174 203255 24176
rect 203537 24174 203593 24230
rect 23752 23188 23808 23244
rect 27453 20360 27509 20416
rect 216908 24050 216964 24052
rect 216908 23998 216910 24050
rect 216910 23998 216962 24050
rect 216962 23998 216964 24050
rect 216908 23996 216964 23998
rect 203119 22670 203175 22672
rect 203119 22618 203121 22670
rect 203121 22618 203173 22670
rect 203173 22618 203175 22670
rect 203119 22616 203175 22618
rect 203537 22616 203593 22672
rect 204482 22545 204538 22601
rect 216908 22370 216964 22372
rect 216908 22318 216910 22370
rect 216910 22318 216962 22370
rect 216962 22318 216964 22370
rect 216908 22316 216964 22318
rect 204482 21417 204538 21473
rect 203039 21400 203095 21402
rect 203039 21348 203041 21400
rect 203041 21348 203093 21400
rect 203093 21348 203095 21400
rect 203039 21346 203095 21348
rect 203537 21346 203593 21402
rect 216908 20690 216964 20692
rect 216908 20638 216910 20690
rect 216910 20638 216962 20690
rect 216962 20638 216964 20690
rect 216908 20636 216964 20638
rect 202959 19842 203015 19844
rect 202959 19790 202961 19842
rect 202961 19790 203013 19842
rect 203013 19790 203015 19842
rect 202959 19788 203015 19790
rect 203537 19788 203593 19844
rect 204482 19717 204538 19773
rect 27701 18946 27757 19002
rect 216908 19010 216964 19012
rect 216908 18958 216910 19010
rect 216910 18958 216962 19010
rect 216962 18958 216964 19010
rect 216908 18956 216964 18958
rect 204482 18589 204538 18645
rect 202879 18572 202935 18574
rect 202879 18520 202881 18572
rect 202881 18520 202933 18572
rect 202933 18520 202935 18572
rect 202879 18518 202935 18520
rect 203537 18518 203593 18574
rect 29560 17754 29616 17756
rect 29560 17702 29562 17754
rect 29562 17702 29614 17754
rect 29614 17702 29616 17754
rect 29560 17700 29616 17702
rect 34552 17754 34608 17756
rect 34552 17702 34554 17754
rect 34554 17702 34606 17754
rect 34606 17702 34608 17754
rect 34552 17700 34608 17702
rect 39544 17754 39600 17756
rect 39544 17702 39546 17754
rect 39546 17702 39598 17754
rect 39598 17702 39600 17754
rect 39544 17700 39600 17702
rect 44536 17754 44592 17756
rect 44536 17702 44538 17754
rect 44538 17702 44590 17754
rect 44590 17702 44592 17754
rect 44536 17700 44592 17702
rect 49528 17754 49584 17756
rect 49528 17702 49530 17754
rect 49530 17702 49582 17754
rect 49582 17702 49584 17754
rect 49528 17700 49584 17702
rect 54520 17754 54576 17756
rect 54520 17702 54522 17754
rect 54522 17702 54574 17754
rect 54574 17702 54576 17754
rect 54520 17700 54576 17702
rect 59512 17754 59568 17756
rect 59512 17702 59514 17754
rect 59514 17702 59566 17754
rect 59566 17702 59568 17754
rect 59512 17700 59568 17702
rect 64504 17754 64560 17756
rect 64504 17702 64506 17754
rect 64506 17702 64558 17754
rect 64558 17702 64560 17754
rect 64504 17700 64560 17702
rect 69496 17754 69552 17756
rect 69496 17702 69498 17754
rect 69498 17702 69550 17754
rect 69550 17702 69552 17754
rect 69496 17700 69552 17702
rect 74488 17754 74544 17756
rect 74488 17702 74490 17754
rect 74490 17702 74542 17754
rect 74542 17702 74544 17754
rect 74488 17700 74544 17702
rect 79480 17754 79536 17756
rect 79480 17702 79482 17754
rect 79482 17702 79534 17754
rect 79534 17702 79536 17754
rect 79480 17700 79536 17702
rect 84472 17754 84528 17756
rect 84472 17702 84474 17754
rect 84474 17702 84526 17754
rect 84526 17702 84528 17754
rect 84472 17700 84528 17702
rect 89464 17754 89520 17756
rect 89464 17702 89466 17754
rect 89466 17702 89518 17754
rect 89518 17702 89520 17754
rect 89464 17700 89520 17702
rect 94456 17754 94512 17756
rect 94456 17702 94458 17754
rect 94458 17702 94510 17754
rect 94510 17702 94512 17754
rect 94456 17700 94512 17702
rect 99448 17754 99504 17756
rect 99448 17702 99450 17754
rect 99450 17702 99502 17754
rect 99502 17702 99504 17754
rect 99448 17700 99504 17702
rect 104440 17754 104496 17756
rect 104440 17702 104442 17754
rect 104442 17702 104494 17754
rect 104494 17702 104496 17754
rect 104440 17700 104496 17702
rect 109432 17754 109488 17756
rect 109432 17702 109434 17754
rect 109434 17702 109486 17754
rect 109486 17702 109488 17754
rect 109432 17700 109488 17702
rect 114424 17754 114480 17756
rect 114424 17702 114426 17754
rect 114426 17702 114478 17754
rect 114478 17702 114480 17754
rect 114424 17700 114480 17702
rect 119416 17754 119472 17756
rect 119416 17702 119418 17754
rect 119418 17702 119470 17754
rect 119470 17702 119472 17754
rect 119416 17700 119472 17702
rect 124408 17754 124464 17756
rect 124408 17702 124410 17754
rect 124410 17702 124462 17754
rect 124462 17702 124464 17754
rect 124408 17700 124464 17702
rect 129400 17754 129456 17756
rect 129400 17702 129402 17754
rect 129402 17702 129454 17754
rect 129454 17702 129456 17754
rect 129400 17700 129456 17702
rect 134392 17754 134448 17756
rect 134392 17702 134394 17754
rect 134394 17702 134446 17754
rect 134446 17702 134448 17754
rect 134392 17700 134448 17702
rect 139384 17754 139440 17756
rect 139384 17702 139386 17754
rect 139386 17702 139438 17754
rect 139438 17702 139440 17754
rect 139384 17700 139440 17702
rect 144376 17754 144432 17756
rect 144376 17702 144378 17754
rect 144378 17702 144430 17754
rect 144430 17702 144432 17754
rect 144376 17700 144432 17702
rect 149368 17754 149424 17756
rect 149368 17702 149370 17754
rect 149370 17702 149422 17754
rect 149422 17702 149424 17754
rect 149368 17700 149424 17702
rect 154360 17754 154416 17756
rect 154360 17702 154362 17754
rect 154362 17702 154414 17754
rect 154414 17702 154416 17754
rect 154360 17700 154416 17702
rect 159352 17754 159408 17756
rect 159352 17702 159354 17754
rect 159354 17702 159406 17754
rect 159406 17702 159408 17754
rect 159352 17700 159408 17702
rect 164344 17754 164400 17756
rect 164344 17702 164346 17754
rect 164346 17702 164398 17754
rect 164398 17702 164400 17754
rect 164344 17700 164400 17702
rect 169336 17754 169392 17756
rect 169336 17702 169338 17754
rect 169338 17702 169390 17754
rect 169390 17702 169392 17754
rect 169336 17700 169392 17702
rect 174328 17754 174384 17756
rect 174328 17702 174330 17754
rect 174330 17702 174382 17754
rect 174382 17702 174384 17754
rect 174328 17700 174384 17702
rect 179320 17754 179376 17756
rect 179320 17702 179322 17754
rect 179322 17702 179374 17754
rect 179374 17702 179376 17754
rect 179320 17700 179376 17702
rect 184312 17754 184368 17756
rect 184312 17702 184314 17754
rect 184314 17702 184366 17754
rect 184366 17702 184368 17754
rect 184312 17700 184368 17702
rect 27577 17532 27633 17588
rect 216908 17330 216964 17332
rect 216908 17278 216910 17330
rect 216910 17278 216962 17330
rect 216962 17278 216964 17330
rect 216908 17276 216964 17278
rect 202799 17014 202855 17016
rect 202799 16962 202801 17014
rect 202801 16962 202853 17014
rect 202853 16962 202855 17014
rect 202799 16960 202855 16962
rect 203537 16960 203593 17016
rect 204482 16889 204538 16945
rect 204482 15761 204538 15817
rect 202719 15744 202775 15746
rect 202719 15692 202721 15744
rect 202721 15692 202773 15744
rect 202773 15692 202775 15744
rect 202719 15690 202775 15692
rect 203537 15690 203593 15746
rect 216908 15650 216964 15652
rect 216908 15598 216910 15650
rect 216910 15598 216962 15650
rect 216962 15598 216964 15650
rect 216908 15596 216964 15598
rect 202639 14186 202695 14188
rect 202639 14134 202641 14186
rect 202641 14134 202693 14186
rect 202693 14134 202695 14186
rect 202639 14132 202695 14134
rect 203537 14132 203593 14188
rect 204482 14061 204538 14117
rect 5511 13252 5567 13308
rect 2326 13147 2382 13203
rect 1702 12290 1758 12292
rect 1702 12238 1704 12290
rect 1704 12238 1756 12290
rect 1756 12238 1758 12290
rect 1702 12236 1758 12238
rect 1702 10610 1758 10612
rect 1702 10558 1704 10610
rect 1704 10558 1756 10610
rect 1756 10558 1758 10610
rect 1702 10556 1758 10558
rect 1702 8930 1758 8932
rect 1702 8878 1704 8930
rect 1704 8878 1756 8930
rect 1756 8878 1758 8930
rect 1702 8876 1758 8878
rect 1702 7250 1758 7252
rect 1702 7198 1704 7250
rect 1704 7198 1756 7250
rect 1756 7198 1758 7250
rect 1702 7196 1758 7198
rect 1702 5570 1758 5572
rect 1702 5518 1704 5570
rect 1704 5518 1756 5570
rect 1756 5518 1758 5570
rect 1702 5516 1758 5518
rect 1702 3890 1758 3892
rect 1702 3838 1704 3890
rect 1704 3838 1756 3890
rect 1756 3838 1758 3890
rect 1702 3836 1758 3838
rect 216908 13970 216964 13972
rect 216908 13918 216910 13970
rect 216910 13918 216962 13970
rect 216962 13918 216964 13970
rect 216908 13916 216964 13918
rect 216908 12290 216964 12292
rect 216908 12238 216910 12290
rect 216910 12238 216962 12290
rect 216962 12238 216964 12290
rect 216908 12236 216964 12238
rect 216908 10610 216964 10612
rect 216908 10558 216910 10610
rect 216910 10558 216962 10610
rect 216962 10558 216964 10610
rect 216908 10556 216964 10558
rect 216908 8930 216964 8932
rect 216908 8878 216910 8930
rect 216910 8878 216962 8930
rect 216962 8878 216964 8930
rect 216908 8876 216964 8878
rect 216908 7250 216964 7252
rect 216908 7198 216910 7250
rect 216910 7198 216962 7250
rect 216962 7198 216964 7250
rect 216908 7196 216964 7198
rect 216908 5570 216964 5572
rect 216908 5518 216910 5570
rect 216910 5518 216962 5570
rect 216962 5518 216964 5570
rect 216908 5516 216964 5518
rect 216908 3890 216964 3892
rect 216908 3838 216910 3890
rect 216910 3838 216962 3890
rect 216962 3838 216964 3890
rect 216908 3836 216964 3838
rect 16548 2720 16604 2776
rect 17716 2720 17772 2776
rect 18884 2720 18940 2776
rect 20052 2720 20108 2776
rect 21220 2720 21276 2776
rect 22388 2720 22444 2776
rect 23556 2720 23612 2776
rect 24724 2720 24780 2776
rect 25892 2720 25948 2776
rect 27060 2720 27116 2776
rect 28228 2720 28284 2776
rect 29396 2720 29452 2776
rect 30564 2720 30620 2776
rect 31732 2720 31788 2776
rect 32900 2720 32956 2776
rect 34068 2720 34124 2776
rect 35236 2720 35292 2776
rect 36404 2720 36460 2776
rect 37572 2720 37628 2776
rect 38740 2720 38796 2776
rect 39908 2720 39964 2776
rect 41076 2720 41132 2776
rect 42244 2720 42300 2776
rect 43412 2720 43468 2776
rect 44580 2720 44636 2776
rect 45748 2720 45804 2776
rect 46916 2720 46972 2776
rect 48084 2720 48140 2776
rect 49252 2720 49308 2776
rect 50420 2720 50476 2776
rect 51588 2720 51644 2776
rect 52756 2720 52812 2776
rect 53924 2720 53980 2776
rect 55092 2720 55148 2776
rect 56260 2720 56316 2776
rect 57428 2720 57484 2776
rect 58596 2720 58652 2776
rect 59764 2720 59820 2776
rect 60932 2720 60988 2776
rect 15294 2464 15350 2520
rect 1702 2210 1758 2212
rect 1702 2158 1704 2210
rect 1704 2158 1756 2210
rect 1756 2158 1758 2210
rect 1702 2156 1758 2158
rect 216908 2210 216964 2212
rect 216908 2158 216910 2210
rect 216910 2158 216962 2210
rect 216962 2158 216964 2210
rect 216908 2156 216964 2158
rect 2038 1874 2094 1876
rect 2038 1822 2040 1874
rect 2040 1822 2092 1874
rect 2092 1822 2094 1874
rect 2038 1820 2094 1822
rect 3718 1874 3774 1876
rect 3718 1822 3720 1874
rect 3720 1822 3772 1874
rect 3772 1822 3774 1874
rect 3718 1820 3774 1822
rect 5398 1874 5454 1876
rect 5398 1822 5400 1874
rect 5400 1822 5452 1874
rect 5452 1822 5454 1874
rect 5398 1820 5454 1822
rect 7078 1874 7134 1876
rect 7078 1822 7080 1874
rect 7080 1822 7132 1874
rect 7132 1822 7134 1874
rect 7078 1820 7134 1822
rect 8758 1874 8814 1876
rect 8758 1822 8760 1874
rect 8760 1822 8812 1874
rect 8812 1822 8814 1874
rect 8758 1820 8814 1822
rect 10438 1874 10494 1876
rect 10438 1822 10440 1874
rect 10440 1822 10492 1874
rect 10492 1822 10494 1874
rect 10438 1820 10494 1822
rect 12118 1874 12174 1876
rect 12118 1822 12120 1874
rect 12120 1822 12172 1874
rect 12172 1822 12174 1874
rect 12118 1820 12174 1822
rect 13798 1874 13854 1876
rect 13798 1822 13800 1874
rect 13800 1822 13852 1874
rect 13852 1822 13854 1874
rect 13798 1820 13854 1822
rect 15478 1874 15534 1876
rect 15478 1822 15480 1874
rect 15480 1822 15532 1874
rect 15532 1822 15534 1874
rect 15478 1820 15534 1822
rect 17158 1874 17214 1876
rect 17158 1822 17160 1874
rect 17160 1822 17212 1874
rect 17212 1822 17214 1874
rect 17158 1820 17214 1822
rect 18838 1874 18894 1876
rect 18838 1822 18840 1874
rect 18840 1822 18892 1874
rect 18892 1822 18894 1874
rect 18838 1820 18894 1822
rect 20518 1874 20574 1876
rect 20518 1822 20520 1874
rect 20520 1822 20572 1874
rect 20572 1822 20574 1874
rect 20518 1820 20574 1822
rect 22198 1874 22254 1876
rect 22198 1822 22200 1874
rect 22200 1822 22252 1874
rect 22252 1822 22254 1874
rect 22198 1820 22254 1822
rect 23878 1874 23934 1876
rect 23878 1822 23880 1874
rect 23880 1822 23932 1874
rect 23932 1822 23934 1874
rect 23878 1820 23934 1822
rect 25558 1874 25614 1876
rect 25558 1822 25560 1874
rect 25560 1822 25612 1874
rect 25612 1822 25614 1874
rect 25558 1820 25614 1822
rect 27238 1874 27294 1876
rect 27238 1822 27240 1874
rect 27240 1822 27292 1874
rect 27292 1822 27294 1874
rect 27238 1820 27294 1822
rect 28918 1874 28974 1876
rect 28918 1822 28920 1874
rect 28920 1822 28972 1874
rect 28972 1822 28974 1874
rect 28918 1820 28974 1822
rect 30598 1874 30654 1876
rect 30598 1822 30600 1874
rect 30600 1822 30652 1874
rect 30652 1822 30654 1874
rect 30598 1820 30654 1822
rect 32278 1874 32334 1876
rect 32278 1822 32280 1874
rect 32280 1822 32332 1874
rect 32332 1822 32334 1874
rect 32278 1820 32334 1822
rect 33958 1874 34014 1876
rect 33958 1822 33960 1874
rect 33960 1822 34012 1874
rect 34012 1822 34014 1874
rect 33958 1820 34014 1822
rect 35638 1874 35694 1876
rect 35638 1822 35640 1874
rect 35640 1822 35692 1874
rect 35692 1822 35694 1874
rect 35638 1820 35694 1822
rect 37318 1874 37374 1876
rect 37318 1822 37320 1874
rect 37320 1822 37372 1874
rect 37372 1822 37374 1874
rect 37318 1820 37374 1822
rect 38998 1874 39054 1876
rect 38998 1822 39000 1874
rect 39000 1822 39052 1874
rect 39052 1822 39054 1874
rect 38998 1820 39054 1822
rect 40678 1874 40734 1876
rect 40678 1822 40680 1874
rect 40680 1822 40732 1874
rect 40732 1822 40734 1874
rect 40678 1820 40734 1822
rect 42358 1874 42414 1876
rect 42358 1822 42360 1874
rect 42360 1822 42412 1874
rect 42412 1822 42414 1874
rect 42358 1820 42414 1822
rect 44038 1874 44094 1876
rect 44038 1822 44040 1874
rect 44040 1822 44092 1874
rect 44092 1822 44094 1874
rect 44038 1820 44094 1822
rect 45718 1874 45774 1876
rect 45718 1822 45720 1874
rect 45720 1822 45772 1874
rect 45772 1822 45774 1874
rect 45718 1820 45774 1822
rect 47398 1874 47454 1876
rect 47398 1822 47400 1874
rect 47400 1822 47452 1874
rect 47452 1822 47454 1874
rect 47398 1820 47454 1822
rect 49078 1874 49134 1876
rect 49078 1822 49080 1874
rect 49080 1822 49132 1874
rect 49132 1822 49134 1874
rect 49078 1820 49134 1822
rect 50758 1874 50814 1876
rect 50758 1822 50760 1874
rect 50760 1822 50812 1874
rect 50812 1822 50814 1874
rect 50758 1820 50814 1822
rect 52438 1874 52494 1876
rect 52438 1822 52440 1874
rect 52440 1822 52492 1874
rect 52492 1822 52494 1874
rect 52438 1820 52494 1822
rect 54118 1874 54174 1876
rect 54118 1822 54120 1874
rect 54120 1822 54172 1874
rect 54172 1822 54174 1874
rect 54118 1820 54174 1822
rect 55798 1874 55854 1876
rect 55798 1822 55800 1874
rect 55800 1822 55852 1874
rect 55852 1822 55854 1874
rect 55798 1820 55854 1822
rect 57478 1874 57534 1876
rect 57478 1822 57480 1874
rect 57480 1822 57532 1874
rect 57532 1822 57534 1874
rect 57478 1820 57534 1822
rect 59158 1874 59214 1876
rect 59158 1822 59160 1874
rect 59160 1822 59212 1874
rect 59212 1822 59214 1874
rect 59158 1820 59214 1822
rect 60838 1874 60894 1876
rect 60838 1822 60840 1874
rect 60840 1822 60892 1874
rect 60892 1822 60894 1874
rect 60838 1820 60894 1822
rect 62518 1874 62574 1876
rect 62518 1822 62520 1874
rect 62520 1822 62572 1874
rect 62572 1822 62574 1874
rect 62518 1820 62574 1822
rect 64198 1874 64254 1876
rect 64198 1822 64200 1874
rect 64200 1822 64252 1874
rect 64252 1822 64254 1874
rect 64198 1820 64254 1822
rect 65878 1874 65934 1876
rect 65878 1822 65880 1874
rect 65880 1822 65932 1874
rect 65932 1822 65934 1874
rect 65878 1820 65934 1822
rect 67558 1874 67614 1876
rect 67558 1822 67560 1874
rect 67560 1822 67612 1874
rect 67612 1822 67614 1874
rect 67558 1820 67614 1822
rect 69238 1874 69294 1876
rect 69238 1822 69240 1874
rect 69240 1822 69292 1874
rect 69292 1822 69294 1874
rect 69238 1820 69294 1822
rect 70918 1874 70974 1876
rect 70918 1822 70920 1874
rect 70920 1822 70972 1874
rect 70972 1822 70974 1874
rect 70918 1820 70974 1822
rect 72598 1874 72654 1876
rect 72598 1822 72600 1874
rect 72600 1822 72652 1874
rect 72652 1822 72654 1874
rect 72598 1820 72654 1822
rect 74278 1874 74334 1876
rect 74278 1822 74280 1874
rect 74280 1822 74332 1874
rect 74332 1822 74334 1874
rect 74278 1820 74334 1822
rect 75958 1874 76014 1876
rect 75958 1822 75960 1874
rect 75960 1822 76012 1874
rect 76012 1822 76014 1874
rect 75958 1820 76014 1822
rect 77638 1874 77694 1876
rect 77638 1822 77640 1874
rect 77640 1822 77692 1874
rect 77692 1822 77694 1874
rect 77638 1820 77694 1822
rect 79318 1874 79374 1876
rect 79318 1822 79320 1874
rect 79320 1822 79372 1874
rect 79372 1822 79374 1874
rect 79318 1820 79374 1822
rect 80998 1874 81054 1876
rect 80998 1822 81000 1874
rect 81000 1822 81052 1874
rect 81052 1822 81054 1874
rect 80998 1820 81054 1822
rect 82678 1874 82734 1876
rect 82678 1822 82680 1874
rect 82680 1822 82732 1874
rect 82732 1822 82734 1874
rect 82678 1820 82734 1822
rect 84358 1874 84414 1876
rect 84358 1822 84360 1874
rect 84360 1822 84412 1874
rect 84412 1822 84414 1874
rect 84358 1820 84414 1822
rect 86038 1874 86094 1876
rect 86038 1822 86040 1874
rect 86040 1822 86092 1874
rect 86092 1822 86094 1874
rect 86038 1820 86094 1822
rect 87718 1874 87774 1876
rect 87718 1822 87720 1874
rect 87720 1822 87772 1874
rect 87772 1822 87774 1874
rect 87718 1820 87774 1822
rect 89398 1874 89454 1876
rect 89398 1822 89400 1874
rect 89400 1822 89452 1874
rect 89452 1822 89454 1874
rect 89398 1820 89454 1822
rect 91078 1874 91134 1876
rect 91078 1822 91080 1874
rect 91080 1822 91132 1874
rect 91132 1822 91134 1874
rect 91078 1820 91134 1822
rect 92758 1874 92814 1876
rect 92758 1822 92760 1874
rect 92760 1822 92812 1874
rect 92812 1822 92814 1874
rect 92758 1820 92814 1822
rect 94438 1874 94494 1876
rect 94438 1822 94440 1874
rect 94440 1822 94492 1874
rect 94492 1822 94494 1874
rect 94438 1820 94494 1822
rect 96118 1874 96174 1876
rect 96118 1822 96120 1874
rect 96120 1822 96172 1874
rect 96172 1822 96174 1874
rect 96118 1820 96174 1822
rect 97798 1874 97854 1876
rect 97798 1822 97800 1874
rect 97800 1822 97852 1874
rect 97852 1822 97854 1874
rect 97798 1820 97854 1822
rect 99478 1874 99534 1876
rect 99478 1822 99480 1874
rect 99480 1822 99532 1874
rect 99532 1822 99534 1874
rect 99478 1820 99534 1822
rect 101158 1874 101214 1876
rect 101158 1822 101160 1874
rect 101160 1822 101212 1874
rect 101212 1822 101214 1874
rect 101158 1820 101214 1822
rect 102838 1874 102894 1876
rect 102838 1822 102840 1874
rect 102840 1822 102892 1874
rect 102892 1822 102894 1874
rect 102838 1820 102894 1822
rect 104518 1874 104574 1876
rect 104518 1822 104520 1874
rect 104520 1822 104572 1874
rect 104572 1822 104574 1874
rect 104518 1820 104574 1822
rect 106198 1874 106254 1876
rect 106198 1822 106200 1874
rect 106200 1822 106252 1874
rect 106252 1822 106254 1874
rect 106198 1820 106254 1822
rect 107878 1874 107934 1876
rect 107878 1822 107880 1874
rect 107880 1822 107932 1874
rect 107932 1822 107934 1874
rect 107878 1820 107934 1822
rect 109558 1874 109614 1876
rect 109558 1822 109560 1874
rect 109560 1822 109612 1874
rect 109612 1822 109614 1874
rect 109558 1820 109614 1822
rect 111238 1874 111294 1876
rect 111238 1822 111240 1874
rect 111240 1822 111292 1874
rect 111292 1822 111294 1874
rect 111238 1820 111294 1822
rect 112918 1874 112974 1876
rect 112918 1822 112920 1874
rect 112920 1822 112972 1874
rect 112972 1822 112974 1874
rect 112918 1820 112974 1822
rect 114598 1874 114654 1876
rect 114598 1822 114600 1874
rect 114600 1822 114652 1874
rect 114652 1822 114654 1874
rect 114598 1820 114654 1822
rect 116278 1874 116334 1876
rect 116278 1822 116280 1874
rect 116280 1822 116332 1874
rect 116332 1822 116334 1874
rect 116278 1820 116334 1822
rect 117958 1874 118014 1876
rect 117958 1822 117960 1874
rect 117960 1822 118012 1874
rect 118012 1822 118014 1874
rect 117958 1820 118014 1822
rect 119638 1874 119694 1876
rect 119638 1822 119640 1874
rect 119640 1822 119692 1874
rect 119692 1822 119694 1874
rect 119638 1820 119694 1822
rect 121318 1874 121374 1876
rect 121318 1822 121320 1874
rect 121320 1822 121372 1874
rect 121372 1822 121374 1874
rect 121318 1820 121374 1822
rect 122998 1874 123054 1876
rect 122998 1822 123000 1874
rect 123000 1822 123052 1874
rect 123052 1822 123054 1874
rect 122998 1820 123054 1822
rect 124678 1874 124734 1876
rect 124678 1822 124680 1874
rect 124680 1822 124732 1874
rect 124732 1822 124734 1874
rect 124678 1820 124734 1822
rect 126358 1874 126414 1876
rect 126358 1822 126360 1874
rect 126360 1822 126412 1874
rect 126412 1822 126414 1874
rect 126358 1820 126414 1822
rect 128038 1874 128094 1876
rect 128038 1822 128040 1874
rect 128040 1822 128092 1874
rect 128092 1822 128094 1874
rect 128038 1820 128094 1822
rect 129718 1874 129774 1876
rect 129718 1822 129720 1874
rect 129720 1822 129772 1874
rect 129772 1822 129774 1874
rect 129718 1820 129774 1822
rect 131398 1874 131454 1876
rect 131398 1822 131400 1874
rect 131400 1822 131452 1874
rect 131452 1822 131454 1874
rect 131398 1820 131454 1822
rect 133078 1874 133134 1876
rect 133078 1822 133080 1874
rect 133080 1822 133132 1874
rect 133132 1822 133134 1874
rect 133078 1820 133134 1822
rect 134758 1874 134814 1876
rect 134758 1822 134760 1874
rect 134760 1822 134812 1874
rect 134812 1822 134814 1874
rect 134758 1820 134814 1822
rect 136438 1874 136494 1876
rect 136438 1822 136440 1874
rect 136440 1822 136492 1874
rect 136492 1822 136494 1874
rect 136438 1820 136494 1822
rect 138118 1874 138174 1876
rect 138118 1822 138120 1874
rect 138120 1822 138172 1874
rect 138172 1822 138174 1874
rect 138118 1820 138174 1822
rect 139798 1874 139854 1876
rect 139798 1822 139800 1874
rect 139800 1822 139852 1874
rect 139852 1822 139854 1874
rect 139798 1820 139854 1822
rect 141478 1874 141534 1876
rect 141478 1822 141480 1874
rect 141480 1822 141532 1874
rect 141532 1822 141534 1874
rect 141478 1820 141534 1822
rect 143158 1874 143214 1876
rect 143158 1822 143160 1874
rect 143160 1822 143212 1874
rect 143212 1822 143214 1874
rect 143158 1820 143214 1822
rect 144838 1874 144894 1876
rect 144838 1822 144840 1874
rect 144840 1822 144892 1874
rect 144892 1822 144894 1874
rect 144838 1820 144894 1822
rect 146518 1874 146574 1876
rect 146518 1822 146520 1874
rect 146520 1822 146572 1874
rect 146572 1822 146574 1874
rect 146518 1820 146574 1822
rect 148198 1874 148254 1876
rect 148198 1822 148200 1874
rect 148200 1822 148252 1874
rect 148252 1822 148254 1874
rect 148198 1820 148254 1822
rect 149878 1874 149934 1876
rect 149878 1822 149880 1874
rect 149880 1822 149932 1874
rect 149932 1822 149934 1874
rect 149878 1820 149934 1822
rect 151558 1874 151614 1876
rect 151558 1822 151560 1874
rect 151560 1822 151612 1874
rect 151612 1822 151614 1874
rect 151558 1820 151614 1822
rect 153238 1874 153294 1876
rect 153238 1822 153240 1874
rect 153240 1822 153292 1874
rect 153292 1822 153294 1874
rect 153238 1820 153294 1822
rect 154918 1874 154974 1876
rect 154918 1822 154920 1874
rect 154920 1822 154972 1874
rect 154972 1822 154974 1874
rect 154918 1820 154974 1822
rect 156598 1874 156654 1876
rect 156598 1822 156600 1874
rect 156600 1822 156652 1874
rect 156652 1822 156654 1874
rect 156598 1820 156654 1822
rect 158278 1874 158334 1876
rect 158278 1822 158280 1874
rect 158280 1822 158332 1874
rect 158332 1822 158334 1874
rect 158278 1820 158334 1822
rect 159958 1874 160014 1876
rect 159958 1822 159960 1874
rect 159960 1822 160012 1874
rect 160012 1822 160014 1874
rect 159958 1820 160014 1822
rect 161638 1874 161694 1876
rect 161638 1822 161640 1874
rect 161640 1822 161692 1874
rect 161692 1822 161694 1874
rect 161638 1820 161694 1822
rect 163318 1874 163374 1876
rect 163318 1822 163320 1874
rect 163320 1822 163372 1874
rect 163372 1822 163374 1874
rect 163318 1820 163374 1822
rect 164998 1874 165054 1876
rect 164998 1822 165000 1874
rect 165000 1822 165052 1874
rect 165052 1822 165054 1874
rect 164998 1820 165054 1822
rect 166678 1874 166734 1876
rect 166678 1822 166680 1874
rect 166680 1822 166732 1874
rect 166732 1822 166734 1874
rect 166678 1820 166734 1822
rect 168358 1874 168414 1876
rect 168358 1822 168360 1874
rect 168360 1822 168412 1874
rect 168412 1822 168414 1874
rect 168358 1820 168414 1822
rect 170038 1874 170094 1876
rect 170038 1822 170040 1874
rect 170040 1822 170092 1874
rect 170092 1822 170094 1874
rect 170038 1820 170094 1822
rect 171718 1874 171774 1876
rect 171718 1822 171720 1874
rect 171720 1822 171772 1874
rect 171772 1822 171774 1874
rect 171718 1820 171774 1822
rect 173398 1874 173454 1876
rect 173398 1822 173400 1874
rect 173400 1822 173452 1874
rect 173452 1822 173454 1874
rect 173398 1820 173454 1822
rect 175078 1874 175134 1876
rect 175078 1822 175080 1874
rect 175080 1822 175132 1874
rect 175132 1822 175134 1874
rect 175078 1820 175134 1822
rect 176758 1874 176814 1876
rect 176758 1822 176760 1874
rect 176760 1822 176812 1874
rect 176812 1822 176814 1874
rect 176758 1820 176814 1822
rect 178438 1874 178494 1876
rect 178438 1822 178440 1874
rect 178440 1822 178492 1874
rect 178492 1822 178494 1874
rect 178438 1820 178494 1822
rect 180118 1874 180174 1876
rect 180118 1822 180120 1874
rect 180120 1822 180172 1874
rect 180172 1822 180174 1874
rect 180118 1820 180174 1822
rect 181798 1874 181854 1876
rect 181798 1822 181800 1874
rect 181800 1822 181852 1874
rect 181852 1822 181854 1874
rect 181798 1820 181854 1822
rect 183478 1874 183534 1876
rect 183478 1822 183480 1874
rect 183480 1822 183532 1874
rect 183532 1822 183534 1874
rect 183478 1820 183534 1822
rect 185158 1874 185214 1876
rect 185158 1822 185160 1874
rect 185160 1822 185212 1874
rect 185212 1822 185214 1874
rect 185158 1820 185214 1822
rect 186838 1874 186894 1876
rect 186838 1822 186840 1874
rect 186840 1822 186892 1874
rect 186892 1822 186894 1874
rect 186838 1820 186894 1822
rect 188518 1874 188574 1876
rect 188518 1822 188520 1874
rect 188520 1822 188572 1874
rect 188572 1822 188574 1874
rect 188518 1820 188574 1822
rect 190198 1874 190254 1876
rect 190198 1822 190200 1874
rect 190200 1822 190252 1874
rect 190252 1822 190254 1874
rect 190198 1820 190254 1822
rect 191878 1874 191934 1876
rect 191878 1822 191880 1874
rect 191880 1822 191932 1874
rect 191932 1822 191934 1874
rect 191878 1820 191934 1822
rect 193558 1874 193614 1876
rect 193558 1822 193560 1874
rect 193560 1822 193612 1874
rect 193612 1822 193614 1874
rect 193558 1820 193614 1822
rect 195238 1874 195294 1876
rect 195238 1822 195240 1874
rect 195240 1822 195292 1874
rect 195292 1822 195294 1874
rect 195238 1820 195294 1822
rect 196918 1874 196974 1876
rect 196918 1822 196920 1874
rect 196920 1822 196972 1874
rect 196972 1822 196974 1874
rect 196918 1820 196974 1822
rect 198598 1874 198654 1876
rect 198598 1822 198600 1874
rect 198600 1822 198652 1874
rect 198652 1822 198654 1874
rect 198598 1820 198654 1822
rect 200278 1874 200334 1876
rect 200278 1822 200280 1874
rect 200280 1822 200332 1874
rect 200332 1822 200334 1874
rect 200278 1820 200334 1822
rect 201958 1874 202014 1876
rect 201958 1822 201960 1874
rect 201960 1822 202012 1874
rect 202012 1822 202014 1874
rect 201958 1820 202014 1822
rect 203638 1874 203694 1876
rect 203638 1822 203640 1874
rect 203640 1822 203692 1874
rect 203692 1822 203694 1874
rect 203638 1820 203694 1822
rect 205318 1874 205374 1876
rect 205318 1822 205320 1874
rect 205320 1822 205372 1874
rect 205372 1822 205374 1874
rect 205318 1820 205374 1822
rect 206998 1874 207054 1876
rect 206998 1822 207000 1874
rect 207000 1822 207052 1874
rect 207052 1822 207054 1874
rect 206998 1820 207054 1822
rect 208678 1874 208734 1876
rect 208678 1822 208680 1874
rect 208680 1822 208732 1874
rect 208732 1822 208734 1874
rect 208678 1820 208734 1822
rect 210358 1874 210414 1876
rect 210358 1822 210360 1874
rect 210360 1822 210412 1874
rect 210412 1822 210414 1874
rect 210358 1820 210414 1822
rect 212038 1874 212094 1876
rect 212038 1822 212040 1874
rect 212040 1822 212092 1874
rect 212092 1822 212094 1874
rect 212038 1820 212094 1822
rect 213718 1874 213774 1876
rect 213718 1822 213720 1874
rect 213720 1822 213772 1874
rect 213772 1822 213774 1874
rect 213718 1820 213774 1822
rect 215398 1874 215454 1876
rect 215398 1822 215400 1874
rect 215400 1822 215452 1874
rect 215452 1822 215454 1874
rect 215398 1820 215454 1822
<< metal3 >>
rect 272 143822 218492 143828
rect 272 143758 278 143822
rect 342 143758 414 143822
rect 478 143758 550 143822
rect 614 143758 218150 143822
rect 218214 143758 218286 143822
rect 218350 143758 218422 143822
rect 218486 143758 218492 143822
rect 272 143686 218492 143758
rect 272 143622 278 143686
rect 342 143622 414 143686
rect 478 143622 550 143686
rect 614 143622 218150 143686
rect 218214 143622 218286 143686
rect 218350 143622 218422 143686
rect 218486 143622 218492 143686
rect 272 143550 218492 143622
rect 272 143486 278 143550
rect 342 143486 414 143550
rect 478 143486 550 143550
rect 614 143486 198158 143550
rect 198222 143486 218150 143550
rect 218214 143486 218286 143550
rect 218350 143486 218422 143550
rect 218486 143486 218492 143550
rect 272 143480 218492 143486
rect 952 143142 217812 143148
rect 952 143078 958 143142
rect 1022 143078 1094 143142
rect 1158 143078 1230 143142
rect 1294 143078 217470 143142
rect 217534 143078 217606 143142
rect 217670 143078 217742 143142
rect 217806 143078 217812 143142
rect 952 143006 217812 143078
rect 952 142942 958 143006
rect 1022 142942 1094 143006
rect 1158 142942 1230 143006
rect 1294 142942 217470 143006
rect 217534 142942 217606 143006
rect 217670 142942 217742 143006
rect 217806 142942 217812 143006
rect 952 142870 217812 142942
rect 952 142806 958 142870
rect 1022 142806 1094 142870
rect 1158 142806 1230 142870
rect 1294 142806 1910 142870
rect 1974 142806 3678 142870
rect 3742 142806 5446 142870
rect 5510 142806 7214 142870
rect 7278 142806 8710 142870
rect 8774 142806 10478 142870
rect 10542 142806 12246 142870
rect 12310 142806 13742 142870
rect 13806 142806 15374 142870
rect 15438 142806 17142 142870
rect 17206 142806 18910 142870
rect 18974 142806 20406 142870
rect 20470 142806 22174 142870
rect 22238 142806 23942 142870
rect 24006 142806 25438 142870
rect 25502 142806 27206 142870
rect 27270 142806 28974 142870
rect 29038 142806 30470 142870
rect 30534 142806 32238 142870
rect 32302 142806 33870 142870
rect 33934 142806 35502 142870
rect 35566 142806 37406 142870
rect 37470 142806 38902 142870
rect 38966 142806 40670 142870
rect 40734 142806 42438 142870
rect 42502 142806 43934 142870
rect 43998 142806 45702 142870
rect 45766 142806 47470 142870
rect 47534 142806 48966 142870
rect 49030 142806 50734 142870
rect 50798 142806 52366 142870
rect 52430 142806 53998 142870
rect 54062 142806 55902 142870
rect 55966 142806 57398 142870
rect 57462 142806 59166 142870
rect 59230 142806 60934 142870
rect 60998 142806 62430 142870
rect 62494 142806 64062 142870
rect 64126 142806 65966 142870
rect 66030 142806 67462 142870
rect 67526 142806 69366 142870
rect 69430 142806 70862 142870
rect 70926 142806 72494 142870
rect 72558 142806 74262 142870
rect 74326 142806 75894 142870
rect 75958 142806 77662 142870
rect 77726 142806 79430 142870
rect 79494 142806 80926 142870
rect 80990 142806 82694 142870
rect 82758 142806 84598 142870
rect 84662 142806 85958 142870
rect 86022 142806 87726 142870
rect 87790 142806 89494 142870
rect 89558 142806 90990 142870
rect 91054 142806 92894 142870
rect 92958 142806 94390 142870
rect 94454 142806 96158 142870
rect 96222 142806 97790 142870
rect 97854 142806 99558 142870
rect 99622 142806 101190 142870
rect 101254 142806 102958 142870
rect 103022 142806 104454 142870
rect 104518 142806 106222 142870
rect 106286 142806 107854 142870
rect 107918 142806 109622 142870
rect 109686 142806 111118 142870
rect 111182 142806 112886 142870
rect 112950 142806 114654 142870
rect 114718 142806 116150 142870
rect 116214 142806 117918 142870
rect 117982 142806 119686 142870
rect 119750 142806 121318 142870
rect 121382 142806 122950 142870
rect 123014 142806 124718 142870
rect 124782 142806 126214 142870
rect 126278 142806 127982 142870
rect 128046 142806 129614 142870
rect 129678 142806 131382 142870
rect 131446 142806 133150 142870
rect 133214 142806 134646 142870
rect 134710 142806 136414 142870
rect 136478 142806 138182 142870
rect 138246 142806 139678 142870
rect 139742 142806 141446 142870
rect 141510 142806 143214 142870
rect 143278 142806 144710 142870
rect 144774 142806 146478 142870
rect 146542 142806 148110 142870
rect 148174 142806 149742 142870
rect 149806 142806 151646 142870
rect 151710 142806 153142 142870
rect 153206 142806 154774 142870
rect 154838 142806 156678 142870
rect 156742 142806 158174 142870
rect 158238 142806 159942 142870
rect 160006 142806 161710 142870
rect 161774 142806 163206 142870
rect 163270 142806 164974 142870
rect 165038 142806 166606 142870
rect 166670 142806 168238 142870
rect 168302 142806 170142 142870
rect 170206 142806 171638 142870
rect 171702 142806 173406 142870
rect 173470 142806 175174 142870
rect 175238 142806 176670 142870
rect 176734 142806 178438 142870
rect 178502 142806 180206 142870
rect 180270 142806 181702 142870
rect 181766 142806 183334 142870
rect 183398 142806 185102 142870
rect 185166 142806 186734 142870
rect 186798 142806 188638 142870
rect 188702 142806 190134 142870
rect 190198 142806 191902 142870
rect 191966 142806 193670 142870
rect 193734 142806 195166 142870
rect 195230 142806 196934 142870
rect 196998 142806 198838 142870
rect 198902 142806 200198 142870
rect 200262 142806 201966 142870
rect 202030 142806 203598 142870
rect 203662 142806 205230 142870
rect 205294 142806 206862 142870
rect 206926 142806 208630 142870
rect 208694 142806 210398 142870
rect 210462 142806 212030 142870
rect 212094 142806 213662 142870
rect 213726 142806 215430 142870
rect 215494 142806 217470 142870
rect 217534 142806 217606 142870
rect 217670 142806 217742 142870
rect 217806 142806 217812 142870
rect 952 142800 217812 142806
rect 1904 142462 2116 142468
rect 1904 142398 1910 142462
rect 1974 142398 2116 142462
rect 1904 142372 2116 142398
rect 1904 142316 2038 142372
rect 2094 142316 2116 142372
rect 1904 142256 2116 142316
rect 3672 142462 3884 142468
rect 3672 142398 3678 142462
rect 3742 142398 3884 142462
rect 3672 142372 3884 142398
rect 3672 142316 3718 142372
rect 3774 142316 3884 142372
rect 3672 142256 3884 142316
rect 5304 142462 5516 142468
rect 5304 142398 5446 142462
rect 5510 142398 5516 142462
rect 5304 142372 5516 142398
rect 5304 142316 5398 142372
rect 5454 142316 5516 142372
rect 5304 142256 5516 142316
rect 6936 142462 7284 142468
rect 6936 142398 7214 142462
rect 7278 142398 7284 142462
rect 6936 142372 7284 142398
rect 6936 142316 7078 142372
rect 7134 142316 7284 142372
rect 6936 142256 7284 142316
rect 8704 142462 8916 142468
rect 8704 142398 8710 142462
rect 8774 142398 8916 142462
rect 8704 142372 8916 142398
rect 8704 142316 8758 142372
rect 8814 142316 8916 142372
rect 8704 142256 8916 142316
rect 10336 142462 10548 142468
rect 10336 142398 10478 142462
rect 10542 142398 10548 142462
rect 10336 142372 10548 142398
rect 10336 142316 10438 142372
rect 10494 142316 10548 142372
rect 10336 142256 10548 142316
rect 11968 142462 12316 142468
rect 11968 142398 12246 142462
rect 12310 142398 12316 142462
rect 11968 142372 12316 142398
rect 11968 142316 12118 142372
rect 12174 142316 12316 142372
rect 11968 142256 12316 142316
rect 13736 142462 13948 142468
rect 13736 142398 13742 142462
rect 13806 142398 13948 142462
rect 13736 142372 13948 142398
rect 13736 142316 13798 142372
rect 13854 142316 13948 142372
rect 13736 142256 13948 142316
rect 15368 142462 15580 142468
rect 15368 142398 15374 142462
rect 15438 142398 15580 142462
rect 15368 142372 15580 142398
rect 15368 142316 15478 142372
rect 15534 142316 15580 142372
rect 15368 142256 15580 142316
rect 17136 142462 17348 142468
rect 17136 142398 17142 142462
rect 17206 142398 17348 142462
rect 17136 142372 17348 142398
rect 17136 142316 17158 142372
rect 17214 142316 17348 142372
rect 17136 142256 17348 142316
rect 18768 142462 18980 142468
rect 18768 142398 18910 142462
rect 18974 142398 18980 142462
rect 18768 142372 18980 142398
rect 18768 142316 18838 142372
rect 18894 142316 18980 142372
rect 18768 142256 18980 142316
rect 20400 142462 20612 142468
rect 20400 142398 20406 142462
rect 20470 142398 20612 142462
rect 20400 142372 20612 142398
rect 20400 142316 20518 142372
rect 20574 142316 20612 142372
rect 20400 142256 20612 142316
rect 22168 142462 22380 142468
rect 22168 142398 22174 142462
rect 22238 142398 22380 142462
rect 22168 142372 22380 142398
rect 22168 142316 22198 142372
rect 22254 142316 22380 142372
rect 22168 142256 22380 142316
rect 23800 142462 24012 142468
rect 23800 142398 23942 142462
rect 24006 142398 24012 142462
rect 23800 142372 24012 142398
rect 23800 142316 23878 142372
rect 23934 142316 24012 142372
rect 23800 142256 24012 142316
rect 25432 142462 25644 142468
rect 25432 142398 25438 142462
rect 25502 142398 25644 142462
rect 25432 142372 25644 142398
rect 25432 142316 25558 142372
rect 25614 142316 25644 142372
rect 25432 142256 25644 142316
rect 27200 142462 27412 142468
rect 27200 142398 27206 142462
rect 27270 142398 27412 142462
rect 27200 142372 27412 142398
rect 27200 142316 27238 142372
rect 27294 142316 27412 142372
rect 27200 142256 27412 142316
rect 28832 142462 29044 142468
rect 28832 142398 28974 142462
rect 29038 142398 29044 142462
rect 28832 142372 29044 142398
rect 28832 142316 28918 142372
rect 28974 142316 29044 142372
rect 28832 142256 29044 142316
rect 30464 142462 30676 142468
rect 30464 142398 30470 142462
rect 30534 142398 30676 142462
rect 30464 142372 30676 142398
rect 30464 142316 30598 142372
rect 30654 142316 30676 142372
rect 30464 142256 30676 142316
rect 32232 142462 32444 142468
rect 32232 142398 32238 142462
rect 32302 142398 32444 142462
rect 32232 142372 32444 142398
rect 32232 142316 32278 142372
rect 32334 142316 32444 142372
rect 32232 142256 32444 142316
rect 33864 142462 34076 142468
rect 33864 142398 33870 142462
rect 33934 142398 34076 142462
rect 33864 142372 34076 142398
rect 33864 142316 33958 142372
rect 34014 142316 34076 142372
rect 33864 142256 34076 142316
rect 35496 142462 35844 142468
rect 35496 142398 35502 142462
rect 35566 142398 35844 142462
rect 35496 142372 35844 142398
rect 35496 142316 35638 142372
rect 35694 142316 35844 142372
rect 35496 142256 35844 142316
rect 37264 142462 37476 142468
rect 37264 142398 37406 142462
rect 37470 142398 37476 142462
rect 37264 142372 37476 142398
rect 37264 142316 37318 142372
rect 37374 142316 37476 142372
rect 37264 142256 37476 142316
rect 38896 142462 39108 142468
rect 38896 142398 38902 142462
rect 38966 142398 39108 142462
rect 38896 142372 39108 142398
rect 38896 142316 38998 142372
rect 39054 142316 39108 142372
rect 38896 142256 39108 142316
rect 40528 142462 40876 142468
rect 40528 142398 40670 142462
rect 40734 142398 40876 142462
rect 40528 142372 40876 142398
rect 40528 142316 40678 142372
rect 40734 142316 40876 142372
rect 40528 142256 40876 142316
rect 42296 142462 42508 142468
rect 42296 142398 42438 142462
rect 42502 142398 42508 142462
rect 42296 142372 42508 142398
rect 42296 142316 42358 142372
rect 42414 142316 42508 142372
rect 42296 142256 42508 142316
rect 43928 142462 44140 142468
rect 43928 142398 43934 142462
rect 43998 142398 44140 142462
rect 43928 142372 44140 142398
rect 43928 142316 44038 142372
rect 44094 142316 44140 142372
rect 43928 142256 44140 142316
rect 45696 142462 45908 142468
rect 45696 142398 45702 142462
rect 45766 142398 45908 142462
rect 45696 142372 45908 142398
rect 45696 142316 45718 142372
rect 45774 142316 45908 142372
rect 45696 142256 45908 142316
rect 47328 142462 47540 142468
rect 47328 142398 47470 142462
rect 47534 142398 47540 142462
rect 47328 142372 47540 142398
rect 47328 142316 47398 142372
rect 47454 142316 47540 142372
rect 47328 142256 47540 142316
rect 48960 142462 49172 142468
rect 48960 142398 48966 142462
rect 49030 142398 49172 142462
rect 48960 142372 49172 142398
rect 48960 142316 49078 142372
rect 49134 142316 49172 142372
rect 48960 142256 49172 142316
rect 50728 142462 50940 142468
rect 50728 142398 50734 142462
rect 50798 142398 50940 142462
rect 50728 142372 50940 142398
rect 50728 142316 50758 142372
rect 50814 142316 50940 142372
rect 50728 142256 50940 142316
rect 52360 142462 52572 142468
rect 52360 142398 52366 142462
rect 52430 142398 52572 142462
rect 52360 142372 52572 142398
rect 52360 142316 52438 142372
rect 52494 142316 52572 142372
rect 52360 142256 52572 142316
rect 53992 142462 54204 142468
rect 53992 142398 53998 142462
rect 54062 142398 54204 142462
rect 53992 142372 54204 142398
rect 53992 142316 54118 142372
rect 54174 142316 54204 142372
rect 53992 142256 54204 142316
rect 55760 142462 55972 142468
rect 55760 142398 55902 142462
rect 55966 142398 55972 142462
rect 55760 142372 55972 142398
rect 55760 142316 55798 142372
rect 55854 142316 55972 142372
rect 55760 142256 55972 142316
rect 57392 142462 57604 142468
rect 57392 142398 57398 142462
rect 57462 142398 57604 142462
rect 57392 142372 57604 142398
rect 57392 142316 57478 142372
rect 57534 142316 57604 142372
rect 57392 142256 57604 142316
rect 59024 142462 59236 142468
rect 59024 142398 59166 142462
rect 59230 142398 59236 142462
rect 59024 142372 59236 142398
rect 59024 142316 59158 142372
rect 59214 142316 59236 142372
rect 59024 142256 59236 142316
rect 60792 142462 61004 142468
rect 60792 142398 60934 142462
rect 60998 142398 61004 142462
rect 60792 142372 61004 142398
rect 60792 142316 60838 142372
rect 60894 142316 61004 142372
rect 60792 142256 61004 142316
rect 62424 142462 62636 142468
rect 62424 142398 62430 142462
rect 62494 142398 62636 142462
rect 62424 142372 62636 142398
rect 62424 142316 62518 142372
rect 62574 142316 62636 142372
rect 62424 142256 62636 142316
rect 64056 142462 64404 142468
rect 64056 142398 64062 142462
rect 64126 142398 64404 142462
rect 64056 142372 64404 142398
rect 64056 142316 64198 142372
rect 64254 142316 64404 142372
rect 64056 142256 64404 142316
rect 65824 142462 66036 142468
rect 65824 142398 65966 142462
rect 66030 142398 66036 142462
rect 65824 142372 66036 142398
rect 65824 142316 65878 142372
rect 65934 142316 66036 142372
rect 65824 142256 66036 142316
rect 67456 142462 67668 142468
rect 67456 142398 67462 142462
rect 67526 142398 67668 142462
rect 67456 142372 67668 142398
rect 67456 142316 67558 142372
rect 67614 142316 67668 142372
rect 67456 142256 67668 142316
rect 69088 142462 69436 142468
rect 69088 142398 69366 142462
rect 69430 142398 69436 142462
rect 69088 142372 69436 142398
rect 69088 142316 69238 142372
rect 69294 142316 69436 142372
rect 69088 142256 69436 142316
rect 70856 142462 71068 142468
rect 70856 142398 70862 142462
rect 70926 142398 71068 142462
rect 70856 142372 71068 142398
rect 70856 142316 70918 142372
rect 70974 142316 71068 142372
rect 70856 142256 71068 142316
rect 72488 142462 72700 142468
rect 72488 142398 72494 142462
rect 72558 142398 72700 142462
rect 72488 142372 72700 142398
rect 72488 142316 72598 142372
rect 72654 142316 72700 142372
rect 72488 142256 72700 142316
rect 74256 142462 74468 142468
rect 74256 142398 74262 142462
rect 74326 142398 74468 142462
rect 74256 142372 74468 142398
rect 74256 142316 74278 142372
rect 74334 142316 74468 142372
rect 74256 142256 74468 142316
rect 75888 142462 76100 142468
rect 75888 142398 75894 142462
rect 75958 142398 76100 142462
rect 75888 142372 76100 142398
rect 75888 142316 75958 142372
rect 76014 142316 76100 142372
rect 75888 142256 76100 142316
rect 77520 142462 77732 142468
rect 77520 142398 77662 142462
rect 77726 142398 77732 142462
rect 77520 142372 77732 142398
rect 77520 142316 77638 142372
rect 77694 142316 77732 142372
rect 77520 142256 77732 142316
rect 79288 142462 79500 142468
rect 79288 142398 79430 142462
rect 79494 142398 79500 142462
rect 79288 142372 79500 142398
rect 79288 142316 79318 142372
rect 79374 142316 79500 142372
rect 79288 142256 79500 142316
rect 80920 142462 81132 142468
rect 80920 142398 80926 142462
rect 80990 142398 81132 142462
rect 80920 142372 81132 142398
rect 80920 142316 80998 142372
rect 81054 142316 81132 142372
rect 80920 142256 81132 142316
rect 82552 142462 82764 142468
rect 82552 142398 82694 142462
rect 82758 142398 82764 142462
rect 82552 142372 82764 142398
rect 82552 142316 82678 142372
rect 82734 142316 82764 142372
rect 82552 142256 82764 142316
rect 84320 142462 84668 142468
rect 84320 142398 84598 142462
rect 84662 142398 84668 142462
rect 84320 142392 84668 142398
rect 85952 142462 86164 142468
rect 85952 142398 85958 142462
rect 86022 142398 86164 142462
rect 84320 142372 84532 142392
rect 84320 142316 84358 142372
rect 84414 142316 84532 142372
rect 84320 142256 84532 142316
rect 85952 142372 86164 142398
rect 85952 142316 86038 142372
rect 86094 142316 86164 142372
rect 85952 142256 86164 142316
rect 87584 142462 87796 142468
rect 87584 142398 87726 142462
rect 87790 142398 87796 142462
rect 87584 142372 87796 142398
rect 87584 142316 87718 142372
rect 87774 142316 87796 142372
rect 87584 142256 87796 142316
rect 89352 142462 89564 142468
rect 89352 142398 89494 142462
rect 89558 142398 89564 142462
rect 89352 142372 89564 142398
rect 89352 142316 89398 142372
rect 89454 142316 89564 142372
rect 89352 142256 89564 142316
rect 90984 142462 91196 142468
rect 90984 142398 90990 142462
rect 91054 142398 91196 142462
rect 90984 142372 91196 142398
rect 90984 142316 91078 142372
rect 91134 142316 91196 142372
rect 90984 142256 91196 142316
rect 92616 142462 92964 142468
rect 92616 142398 92894 142462
rect 92958 142398 92964 142462
rect 92616 142372 92964 142398
rect 92616 142316 92758 142372
rect 92814 142316 92964 142372
rect 92616 142256 92964 142316
rect 94384 142462 94596 142468
rect 94384 142398 94390 142462
rect 94454 142398 94596 142462
rect 94384 142372 94596 142398
rect 94384 142316 94438 142372
rect 94494 142316 94596 142372
rect 94384 142256 94596 142316
rect 96016 142462 96228 142468
rect 96016 142398 96158 142462
rect 96222 142398 96228 142462
rect 96016 142372 96228 142398
rect 96016 142316 96118 142372
rect 96174 142316 96228 142372
rect 96016 142256 96228 142316
rect 97648 142462 97996 142468
rect 97648 142398 97790 142462
rect 97854 142398 97996 142462
rect 97648 142372 97996 142398
rect 97648 142316 97798 142372
rect 97854 142316 97996 142372
rect 97648 142256 97996 142316
rect 99416 142462 99628 142468
rect 99416 142398 99558 142462
rect 99622 142398 99628 142462
rect 99416 142372 99628 142398
rect 99416 142316 99478 142372
rect 99534 142316 99628 142372
rect 99416 142256 99628 142316
rect 101048 142462 101260 142468
rect 101048 142398 101190 142462
rect 101254 142398 101260 142462
rect 101048 142372 101260 142398
rect 101048 142316 101158 142372
rect 101214 142316 101260 142372
rect 101048 142256 101260 142316
rect 102816 142462 103028 142468
rect 102816 142398 102958 142462
rect 103022 142398 103028 142462
rect 102816 142372 103028 142398
rect 102816 142316 102838 142372
rect 102894 142316 103028 142372
rect 102816 142256 103028 142316
rect 104448 142462 104660 142468
rect 104448 142398 104454 142462
rect 104518 142398 104660 142462
rect 104448 142372 104660 142398
rect 104448 142316 104518 142372
rect 104574 142316 104660 142372
rect 104448 142256 104660 142316
rect 106080 142462 106292 142468
rect 106080 142398 106222 142462
rect 106286 142398 106292 142462
rect 106080 142372 106292 142398
rect 106080 142316 106198 142372
rect 106254 142316 106292 142372
rect 106080 142256 106292 142316
rect 107848 142462 108060 142468
rect 107848 142398 107854 142462
rect 107918 142398 108060 142462
rect 107848 142372 108060 142398
rect 107848 142316 107878 142372
rect 107934 142316 108060 142372
rect 107848 142256 108060 142316
rect 109480 142462 109692 142468
rect 109480 142398 109622 142462
rect 109686 142398 109692 142462
rect 109480 142372 109692 142398
rect 109480 142316 109558 142372
rect 109614 142316 109692 142372
rect 109480 142256 109692 142316
rect 111112 142462 111324 142468
rect 111112 142398 111118 142462
rect 111182 142398 111324 142462
rect 111112 142372 111324 142398
rect 111112 142316 111238 142372
rect 111294 142316 111324 142372
rect 111112 142256 111324 142316
rect 112880 142462 113092 142468
rect 112880 142398 112886 142462
rect 112950 142398 113092 142462
rect 112880 142372 113092 142398
rect 112880 142316 112918 142372
rect 112974 142316 113092 142372
rect 112880 142256 113092 142316
rect 114512 142462 114724 142468
rect 114512 142398 114654 142462
rect 114718 142398 114724 142462
rect 114512 142372 114724 142398
rect 114512 142316 114598 142372
rect 114654 142316 114724 142372
rect 114512 142256 114724 142316
rect 116144 142462 116356 142468
rect 116144 142398 116150 142462
rect 116214 142398 116356 142462
rect 116144 142372 116356 142398
rect 116144 142316 116278 142372
rect 116334 142316 116356 142372
rect 116144 142256 116356 142316
rect 117912 142462 118124 142468
rect 117912 142398 117918 142462
rect 117982 142398 118124 142462
rect 117912 142372 118124 142398
rect 117912 142316 117958 142372
rect 118014 142316 118124 142372
rect 117912 142256 118124 142316
rect 119544 142462 119756 142468
rect 119544 142398 119686 142462
rect 119750 142398 119756 142462
rect 119544 142372 119756 142398
rect 119544 142316 119638 142372
rect 119694 142316 119756 142372
rect 119544 142256 119756 142316
rect 121176 142462 121524 142468
rect 121176 142398 121318 142462
rect 121382 142398 121524 142462
rect 121176 142372 121524 142398
rect 121176 142316 121318 142372
rect 121374 142316 121524 142372
rect 121176 142256 121524 142316
rect 122944 142462 123156 142468
rect 122944 142398 122950 142462
rect 123014 142398 123156 142462
rect 122944 142372 123156 142398
rect 122944 142316 122998 142372
rect 123054 142316 123156 142372
rect 122944 142256 123156 142316
rect 124576 142462 124788 142468
rect 124576 142398 124718 142462
rect 124782 142398 124788 142462
rect 124576 142372 124788 142398
rect 124576 142316 124678 142372
rect 124734 142316 124788 142372
rect 124576 142256 124788 142316
rect 126208 142462 126556 142468
rect 126208 142398 126214 142462
rect 126278 142398 126556 142462
rect 126208 142372 126556 142398
rect 126208 142316 126358 142372
rect 126414 142316 126556 142372
rect 126208 142256 126556 142316
rect 127976 142462 128188 142468
rect 127976 142398 127982 142462
rect 128046 142398 128188 142462
rect 127976 142372 128188 142398
rect 127976 142316 128038 142372
rect 128094 142316 128188 142372
rect 127976 142256 128188 142316
rect 129608 142462 129820 142468
rect 129608 142398 129614 142462
rect 129678 142398 129820 142462
rect 129608 142372 129820 142398
rect 129608 142316 129718 142372
rect 129774 142316 129820 142372
rect 129608 142256 129820 142316
rect 131376 142462 131588 142468
rect 131376 142398 131382 142462
rect 131446 142398 131588 142462
rect 131376 142372 131588 142398
rect 131376 142316 131398 142372
rect 131454 142316 131588 142372
rect 131376 142256 131588 142316
rect 133008 142462 133220 142468
rect 133008 142398 133150 142462
rect 133214 142398 133220 142462
rect 133008 142372 133220 142398
rect 133008 142316 133078 142372
rect 133134 142316 133220 142372
rect 133008 142256 133220 142316
rect 134640 142462 134852 142468
rect 134640 142398 134646 142462
rect 134710 142398 134852 142462
rect 134640 142372 134852 142398
rect 134640 142316 134758 142372
rect 134814 142316 134852 142372
rect 134640 142256 134852 142316
rect 136408 142462 136620 142468
rect 136408 142398 136414 142462
rect 136478 142398 136620 142462
rect 136408 142372 136620 142398
rect 136408 142316 136438 142372
rect 136494 142316 136620 142372
rect 136408 142256 136620 142316
rect 138040 142462 138252 142468
rect 138040 142398 138182 142462
rect 138246 142398 138252 142462
rect 138040 142372 138252 142398
rect 138040 142316 138118 142372
rect 138174 142316 138252 142372
rect 138040 142256 138252 142316
rect 139672 142462 139884 142468
rect 139672 142398 139678 142462
rect 139742 142398 139884 142462
rect 139672 142372 139884 142398
rect 139672 142316 139798 142372
rect 139854 142316 139884 142372
rect 139672 142256 139884 142316
rect 141440 142462 141652 142468
rect 141440 142398 141446 142462
rect 141510 142398 141652 142462
rect 141440 142372 141652 142398
rect 141440 142316 141478 142372
rect 141534 142316 141652 142372
rect 141440 142256 141652 142316
rect 143072 142462 143284 142468
rect 143072 142398 143214 142462
rect 143278 142398 143284 142462
rect 143072 142372 143284 142398
rect 143072 142316 143158 142372
rect 143214 142316 143284 142372
rect 143072 142256 143284 142316
rect 144704 142462 144916 142468
rect 144704 142398 144710 142462
rect 144774 142398 144916 142462
rect 144704 142372 144916 142398
rect 144704 142316 144838 142372
rect 144894 142316 144916 142372
rect 144704 142256 144916 142316
rect 146472 142462 146684 142468
rect 146472 142398 146478 142462
rect 146542 142398 146684 142462
rect 146472 142372 146684 142398
rect 146472 142316 146518 142372
rect 146574 142316 146684 142372
rect 146472 142256 146684 142316
rect 148104 142462 148316 142468
rect 148104 142398 148110 142462
rect 148174 142398 148316 142462
rect 148104 142372 148316 142398
rect 148104 142316 148198 142372
rect 148254 142316 148316 142372
rect 148104 142256 148316 142316
rect 149736 142462 150084 142468
rect 149736 142398 149742 142462
rect 149806 142398 150084 142462
rect 149736 142372 150084 142398
rect 149736 142316 149878 142372
rect 149934 142316 150084 142372
rect 149736 142256 150084 142316
rect 151504 142462 151716 142468
rect 151504 142398 151646 142462
rect 151710 142398 151716 142462
rect 151504 142372 151716 142398
rect 151504 142316 151558 142372
rect 151614 142316 151716 142372
rect 151504 142256 151716 142316
rect 153136 142462 153348 142468
rect 153136 142398 153142 142462
rect 153206 142398 153348 142462
rect 153136 142372 153348 142398
rect 153136 142316 153238 142372
rect 153294 142316 153348 142372
rect 153136 142256 153348 142316
rect 154768 142462 155116 142468
rect 154768 142398 154774 142462
rect 154838 142398 155116 142462
rect 154768 142372 155116 142398
rect 154768 142316 154918 142372
rect 154974 142316 155116 142372
rect 154768 142256 155116 142316
rect 156536 142462 156748 142468
rect 156536 142398 156678 142462
rect 156742 142398 156748 142462
rect 156536 142372 156748 142398
rect 156536 142316 156598 142372
rect 156654 142316 156748 142372
rect 156536 142256 156748 142316
rect 158168 142462 158380 142468
rect 158168 142398 158174 142462
rect 158238 142398 158380 142462
rect 158168 142372 158380 142398
rect 158168 142316 158278 142372
rect 158334 142316 158380 142372
rect 158168 142256 158380 142316
rect 159936 142462 160148 142468
rect 159936 142398 159942 142462
rect 160006 142398 160148 142462
rect 159936 142372 160148 142398
rect 159936 142316 159958 142372
rect 160014 142316 160148 142372
rect 159936 142256 160148 142316
rect 161568 142462 161780 142468
rect 161568 142398 161710 142462
rect 161774 142398 161780 142462
rect 161568 142372 161780 142398
rect 161568 142316 161638 142372
rect 161694 142316 161780 142372
rect 161568 142256 161780 142316
rect 163200 142462 163412 142468
rect 163200 142398 163206 142462
rect 163270 142398 163412 142462
rect 163200 142372 163412 142398
rect 163200 142316 163318 142372
rect 163374 142316 163412 142372
rect 163200 142256 163412 142316
rect 164968 142462 165180 142468
rect 164968 142398 164974 142462
rect 165038 142398 165180 142462
rect 164968 142372 165180 142398
rect 164968 142316 164998 142372
rect 165054 142316 165180 142372
rect 164968 142256 165180 142316
rect 166600 142462 166812 142468
rect 166600 142398 166606 142462
rect 166670 142398 166812 142462
rect 166600 142372 166812 142398
rect 166600 142316 166678 142372
rect 166734 142316 166812 142372
rect 166600 142256 166812 142316
rect 168232 142462 168444 142468
rect 168232 142398 168238 142462
rect 168302 142398 168444 142462
rect 168232 142372 168444 142398
rect 168232 142316 168358 142372
rect 168414 142316 168444 142372
rect 168232 142256 168444 142316
rect 170000 142462 170212 142468
rect 170000 142398 170142 142462
rect 170206 142398 170212 142462
rect 170000 142372 170212 142398
rect 170000 142316 170038 142372
rect 170094 142316 170212 142372
rect 170000 142256 170212 142316
rect 171632 142462 171844 142468
rect 171632 142398 171638 142462
rect 171702 142398 171844 142462
rect 171632 142372 171844 142398
rect 171632 142316 171718 142372
rect 171774 142316 171844 142372
rect 171632 142256 171844 142316
rect 173264 142462 173476 142468
rect 173264 142398 173406 142462
rect 173470 142398 173476 142462
rect 173264 142372 173476 142398
rect 173264 142316 173398 142372
rect 173454 142316 173476 142372
rect 173264 142256 173476 142316
rect 175032 142462 175244 142468
rect 175032 142398 175174 142462
rect 175238 142398 175244 142462
rect 175032 142372 175244 142398
rect 175032 142316 175078 142372
rect 175134 142316 175244 142372
rect 175032 142256 175244 142316
rect 176664 142462 176876 142468
rect 176664 142398 176670 142462
rect 176734 142398 176876 142462
rect 176664 142372 176876 142398
rect 176664 142316 176758 142372
rect 176814 142316 176876 142372
rect 176664 142256 176876 142316
rect 178296 142462 178644 142468
rect 178296 142398 178438 142462
rect 178502 142398 178644 142462
rect 178296 142372 178644 142398
rect 178296 142316 178438 142372
rect 178494 142316 178644 142372
rect 178296 142256 178644 142316
rect 180064 142462 180276 142468
rect 180064 142398 180206 142462
rect 180270 142398 180276 142462
rect 180064 142372 180276 142398
rect 180064 142316 180118 142372
rect 180174 142316 180276 142372
rect 180064 142256 180276 142316
rect 181696 142462 181908 142468
rect 181696 142398 181702 142462
rect 181766 142398 181908 142462
rect 181696 142372 181908 142398
rect 181696 142316 181798 142372
rect 181854 142316 181908 142372
rect 181696 142256 181908 142316
rect 183328 142462 183676 142468
rect 183328 142398 183334 142462
rect 183398 142398 183676 142462
rect 183328 142372 183676 142398
rect 183328 142316 183478 142372
rect 183534 142316 183676 142372
rect 183328 142256 183676 142316
rect 185096 142462 185308 142468
rect 185096 142398 185102 142462
rect 185166 142398 185308 142462
rect 185096 142372 185308 142398
rect 185096 142316 185158 142372
rect 185214 142316 185308 142372
rect 185096 142256 185308 142316
rect 186728 142462 186940 142468
rect 186728 142398 186734 142462
rect 186798 142398 186940 142462
rect 186728 142372 186940 142398
rect 186728 142316 186838 142372
rect 186894 142316 186940 142372
rect 186728 142256 186940 142316
rect 188496 142462 188708 142468
rect 188496 142398 188638 142462
rect 188702 142398 188708 142462
rect 188496 142372 188708 142398
rect 188496 142316 188518 142372
rect 188574 142316 188708 142372
rect 188496 142256 188708 142316
rect 190128 142462 190340 142468
rect 190128 142398 190134 142462
rect 190198 142398 190340 142462
rect 190128 142372 190340 142398
rect 190128 142316 190198 142372
rect 190254 142316 190340 142372
rect 190128 142256 190340 142316
rect 191760 142462 191972 142468
rect 191760 142398 191902 142462
rect 191966 142398 191972 142462
rect 191760 142372 191972 142398
rect 191760 142316 191878 142372
rect 191934 142316 191972 142372
rect 191760 142256 191972 142316
rect 193528 142462 193740 142468
rect 193528 142398 193670 142462
rect 193734 142398 193740 142462
rect 193528 142372 193740 142398
rect 193528 142316 193558 142372
rect 193614 142316 193740 142372
rect 193528 142256 193740 142316
rect 195160 142462 195372 142468
rect 195160 142398 195166 142462
rect 195230 142398 195372 142462
rect 195160 142372 195372 142398
rect 195160 142316 195238 142372
rect 195294 142316 195372 142372
rect 195160 142256 195372 142316
rect 196792 142462 197004 142468
rect 196792 142398 196934 142462
rect 196998 142398 197004 142462
rect 196792 142372 197004 142398
rect 196792 142316 196918 142372
rect 196974 142316 197004 142372
rect 196792 142256 197004 142316
rect 198560 142462 198908 142468
rect 198560 142398 198838 142462
rect 198902 142398 198908 142462
rect 198560 142392 198908 142398
rect 200192 142462 200404 142468
rect 200192 142398 200198 142462
rect 200262 142398 200404 142462
rect 198560 142372 198772 142392
rect 198560 142316 198598 142372
rect 198654 142332 198772 142372
rect 200192 142372 200404 142398
rect 198654 142326 199316 142332
rect 198654 142316 199246 142326
rect 198560 142262 199246 142316
rect 199310 142262 199316 142326
rect 198560 142256 199316 142262
rect 200192 142316 200278 142372
rect 200334 142332 200404 142372
rect 201824 142462 202036 142468
rect 201824 142398 201966 142462
rect 202030 142398 202036 142462
rect 201824 142372 202036 142398
rect 200334 142326 200540 142332
rect 200334 142316 200470 142326
rect 200192 142262 200470 142316
rect 200534 142262 200540 142326
rect 200192 142256 200540 142262
rect 201824 142316 201958 142372
rect 202014 142316 202036 142372
rect 201824 142256 202036 142316
rect 203592 142462 203804 142468
rect 203592 142398 203598 142462
rect 203662 142398 203804 142462
rect 203592 142372 203804 142398
rect 203592 142316 203638 142372
rect 203694 142316 203804 142372
rect 203592 142256 203804 142316
rect 205224 142462 205436 142468
rect 205224 142398 205230 142462
rect 205294 142398 205436 142462
rect 205224 142372 205436 142398
rect 205224 142316 205318 142372
rect 205374 142316 205436 142372
rect 205224 142256 205436 142316
rect 206856 142462 207204 142468
rect 206856 142398 206862 142462
rect 206926 142398 207204 142462
rect 206856 142372 207204 142398
rect 206856 142316 206998 142372
rect 207054 142316 207204 142372
rect 206856 142256 207204 142316
rect 208624 142462 208836 142468
rect 208624 142398 208630 142462
rect 208694 142398 208836 142462
rect 208624 142372 208836 142398
rect 208624 142316 208678 142372
rect 208734 142316 208836 142372
rect 208624 142256 208836 142316
rect 210256 142462 210468 142468
rect 210256 142398 210398 142462
rect 210462 142398 210468 142462
rect 210256 142372 210468 142398
rect 210256 142316 210358 142372
rect 210414 142316 210468 142372
rect 210256 142256 210468 142316
rect 211888 142462 212236 142468
rect 211888 142398 212030 142462
rect 212094 142398 212236 142462
rect 211888 142372 212236 142398
rect 211888 142316 212038 142372
rect 212094 142316 212236 142372
rect 211888 142256 212236 142316
rect 213656 142462 213868 142468
rect 213656 142398 213662 142462
rect 213726 142398 213868 142462
rect 213656 142372 213868 142398
rect 213656 142316 213718 142372
rect 213774 142316 213868 142372
rect 213656 142256 213868 142316
rect 215288 142462 215500 142468
rect 215288 142398 215430 142462
rect 215494 142398 215500 142462
rect 215288 142372 215500 142398
rect 215288 142316 215398 142372
rect 215454 142316 215500 142372
rect 215288 142256 215500 142316
rect 198560 142060 198636 142256
rect 198152 141984 198636 142060
rect 199240 142054 199588 142060
rect 199240 141990 199246 142054
rect 199310 141990 199588 142054
rect 198152 141918 198364 141984
rect 198152 141854 198294 141918
rect 198358 141854 198364 141918
rect 198152 141848 198364 141854
rect 199240 141848 199588 141990
rect 200464 142054 200676 142060
rect 200464 141990 200470 142054
rect 200534 141990 200676 142054
rect 200464 141848 200676 141990
rect 1224 141782 1844 141788
rect 1224 141718 1230 141782
rect 1294 141718 1844 141782
rect 216784 141782 217540 141788
rect 203395 141730 203461 141733
rect 1224 141712 1844 141718
rect 1632 141652 1844 141712
rect 199424 141728 203461 141730
rect 199424 141672 203400 141728
rect 203456 141672 203461 141728
rect 199424 141670 203461 141672
rect 203395 141667 203461 141670
rect 216784 141718 217470 141782
rect 217534 141718 217540 141782
rect 216784 141712 217540 141718
rect 1632 141596 1702 141652
rect 1758 141596 1844 141652
rect 1632 141440 1844 141596
rect 216784 141652 216996 141712
rect 216784 141596 216908 141652
rect 216964 141596 216996 141652
rect 198560 141510 198772 141516
rect 198560 141446 198566 141510
rect 198630 141472 198772 141510
rect 198630 141446 198642 141472
rect 198560 141416 198642 141446
rect 198698 141416 198772 141472
rect 198560 141304 198772 141416
rect 199784 141510 199996 141516
rect 199784 141472 199926 141510
rect 199784 141416 199810 141472
rect 199866 141446 199926 141472
rect 199990 141446 199996 141510
rect 199866 141416 199996 141446
rect 199784 141304 199996 141416
rect 200872 141510 201084 141516
rect 200872 141472 201014 141510
rect 200872 141416 200978 141472
rect 201078 141446 201084 141510
rect 201034 141416 201084 141446
rect 216784 141440 216996 141596
rect 200872 141304 201084 141416
rect 198152 140694 198364 140700
rect 198152 140630 198158 140694
rect 198222 140630 198364 140694
rect 198152 140564 198364 140630
rect 199240 140564 199588 140700
rect 200464 140564 200676 140700
rect 198152 140558 200676 140564
rect 198152 140494 198158 140558
rect 198222 140494 200676 140558
rect 198152 140488 200676 140494
rect 1632 139972 1844 140020
rect 1632 139916 1702 139972
rect 1758 139916 1844 139972
rect 1632 139884 1844 139916
rect 216784 140014 217540 140020
rect 216784 139972 217470 140014
rect 216784 139916 216908 139972
rect 216964 139950 217470 139972
rect 217534 139950 217540 140014
rect 216964 139944 217540 139950
rect 216964 139916 216996 139944
rect 1224 139878 1844 139884
rect 1224 139814 1230 139878
rect 1294 139814 1844 139878
rect 1224 139808 1844 139814
rect 196520 139878 198364 139884
rect 196520 139814 198294 139878
rect 198358 139814 198364 139878
rect 196520 139808 198364 139814
rect 216784 139808 216996 139916
rect 196520 139672 196732 139808
rect 197880 139742 198092 139808
rect 197880 139678 197886 139742
rect 197950 139678 198092 139742
rect 197880 139672 198092 139678
rect 196520 138388 196732 138524
rect 197880 138518 198228 138524
rect 197880 138454 198158 138518
rect 198222 138454 198228 138518
rect 197880 138448 198228 138454
rect 197880 138388 198092 138448
rect 1632 138292 1844 138388
rect 196520 138382 198092 138388
rect 196520 138318 196662 138382
rect 196726 138318 198092 138382
rect 196520 138312 198092 138318
rect 216784 138382 217540 138388
rect 216784 138318 217470 138382
rect 217534 138318 217540 138382
rect 216784 138312 217540 138318
rect 1632 138252 1702 138292
rect 1224 138246 1702 138252
rect 1224 138182 1230 138246
rect 1294 138236 1702 138246
rect 1758 138236 1844 138292
rect 1294 138182 1844 138236
rect 1224 138176 1844 138182
rect 216784 138292 216996 138312
rect 216784 138236 216908 138292
rect 216964 138236 216996 138292
rect 216784 138176 216996 138236
rect 196520 137028 196732 137164
rect 197880 137158 198092 137164
rect 197880 137094 197886 137158
rect 197950 137094 198092 137158
rect 197880 137028 198092 137094
rect 196520 136952 198092 137028
rect 196520 136816 196732 136952
rect 197880 136886 198092 136952
rect 197880 136822 197886 136886
rect 197950 136822 198092 136886
rect 197880 136816 198092 136822
rect 1224 136750 1844 136756
rect 1224 136686 1230 136750
rect 1294 136686 1844 136750
rect 1224 136680 1844 136686
rect 1632 136612 1844 136680
rect 1632 136556 1702 136612
rect 1758 136556 1844 136612
rect 1632 136408 1844 136556
rect 216784 136620 216996 136756
rect 216784 136614 217540 136620
rect 216784 136612 217470 136614
rect 216784 136556 216908 136612
rect 216964 136556 217470 136612
rect 216784 136550 217470 136556
rect 217534 136550 217540 136614
rect 216784 136544 217540 136550
rect 216784 136408 216996 136544
rect 196520 135662 196732 135668
rect 196520 135598 196662 135662
rect 196726 135598 196732 135662
rect 196520 135532 196732 135598
rect 197880 135532 198092 135668
rect 196520 135526 198092 135532
rect 196520 135462 198022 135526
rect 198086 135462 198092 135526
rect 196520 135456 198092 135462
rect 203456 135260 203668 135532
rect 203358 135254 203668 135260
rect 203320 135190 203326 135254
rect 203390 135190 203668 135254
rect 203358 135184 203668 135190
rect 216376 135260 216588 135532
rect 216376 135254 216860 135260
rect 216376 135190 216790 135254
rect 216854 135190 216860 135254
rect 216376 135184 216860 135190
rect 1224 134982 1844 134988
rect 1224 134918 1230 134982
rect 1294 134932 1844 134982
rect 1294 134918 1702 134932
rect 1224 134912 1702 134918
rect 1632 134876 1702 134912
rect 1758 134876 1844 134932
rect 1632 134776 1844 134876
rect 216784 134982 216996 134988
rect 216784 134918 216790 134982
rect 216854 134932 216996 134982
rect 216854 134918 216908 134932
rect 216784 134876 216908 134918
rect 216964 134876 216996 134932
rect 216784 134852 216996 134876
rect 213112 134716 213324 134852
rect 216240 134819 216452 134852
rect 216240 134763 216284 134819
rect 216340 134763 216452 134819
rect 216784 134846 217540 134852
rect 216784 134782 217470 134846
rect 217534 134782 217540 134846
rect 216784 134776 217540 134782
rect 216240 134716 216452 134763
rect 213112 134714 216180 134716
rect 213112 134658 213183 134714
rect 213239 134658 216180 134714
rect 213112 134640 216180 134658
rect 216240 134640 218764 134716
rect 213112 134504 213324 134640
rect 216104 134580 216180 134640
rect 216104 134504 218764 134580
rect 196520 134172 196732 134308
rect 197880 134302 198092 134308
rect 197880 134238 197886 134302
rect 197950 134238 198092 134302
rect 197880 134172 198092 134238
rect 196520 134166 198092 134172
rect 196520 134102 196662 134166
rect 196726 134102 198092 134166
rect 196520 134096 198092 134102
rect 203456 133894 203668 134036
rect 203456 133830 203462 133894
rect 203526 133830 203598 133894
rect 203662 133830 203668 133894
rect 203456 133824 203668 133830
rect 216376 133900 216588 134036
rect 216376 133894 218220 133900
rect 216376 133830 218150 133894
rect 218214 133830 218220 133894
rect 216376 133824 218220 133830
rect 1632 133252 1844 133356
rect 1632 133220 1702 133252
rect 1224 133214 1702 133220
rect 1224 133150 1230 133214
rect 1294 133196 1702 133214
rect 1758 133196 1844 133252
rect 216784 133350 217540 133356
rect 216784 133286 217470 133350
rect 217534 133286 217540 133350
rect 216784 133280 217540 133286
rect 216784 133252 216996 133280
rect 1294 133150 1844 133196
rect 1224 133144 1844 133150
rect 29512 133214 29724 133220
rect 29512 133150 29518 133214
rect 29582 133150 29724 133214
rect 29512 133094 29724 133150
rect 29920 133134 29996 133220
rect 29512 133038 29560 133094
rect 29616 133038 29724 133094
rect 29512 133008 29724 133038
rect 29793 133078 29996 133134
rect 29793 133036 29926 133078
rect 29920 133014 29926 133036
rect 29990 133014 29996 133078
rect 29920 133008 29996 133014
rect 34408 133214 34620 133220
rect 34408 133150 34414 133214
rect 34478 133150 34620 133214
rect 34408 133115 34620 133150
rect 34816 133134 34892 133220
rect 34408 133094 34629 133115
rect 34408 133038 34552 133094
rect 34608 133038 34629 133094
rect 34408 133017 34629 133038
rect 34785 133078 34892 133134
rect 34785 133036 34822 133078
rect 34408 133008 34620 133017
rect 34816 133014 34822 133036
rect 34886 133014 34892 133078
rect 34816 133008 34892 133014
rect 39440 133214 39652 133220
rect 39440 133150 39446 133214
rect 39510 133150 39652 133214
rect 39440 133094 39652 133150
rect 39440 133038 39544 133094
rect 39600 133038 39652 133094
rect 39440 133008 39652 133038
rect 39712 133078 39924 133220
rect 39712 133014 39854 133078
rect 39918 133014 39924 133078
rect 39712 133008 39924 133014
rect 44472 133214 44684 133220
rect 44472 133150 44478 133214
rect 44542 133150 44684 133214
rect 44472 133094 44684 133150
rect 44880 133134 44956 133220
rect 44472 133038 44536 133094
rect 44592 133038 44684 133094
rect 44472 133008 44684 133038
rect 44769 133078 44956 133134
rect 44769 133036 44886 133078
rect 44880 133014 44886 133036
rect 44950 133014 44956 133078
rect 44880 133008 44956 133014
rect 49504 133214 49580 133220
rect 49504 133150 49510 133214
rect 49574 133150 49580 133214
rect 49504 133115 49580 133150
rect 49776 133134 49988 133220
rect 49504 133094 49605 133115
rect 49504 133038 49528 133094
rect 49584 133038 49605 133094
rect 49504 133017 49605 133038
rect 49761 133078 49988 133134
rect 49761 133036 49918 133078
rect 49504 133008 49580 133017
rect 49776 133014 49918 133036
rect 49982 133014 49988 133078
rect 49776 133008 49988 133014
rect 54400 133214 54612 133220
rect 54400 133150 54542 133214
rect 54606 133150 54612 133214
rect 54400 133094 54612 133150
rect 54808 133134 54884 133220
rect 54400 133038 54520 133094
rect 54576 133038 54612 133094
rect 54400 133008 54612 133038
rect 54753 133078 54884 133134
rect 54753 133036 54814 133078
rect 54808 133014 54814 133036
rect 54878 133014 54884 133078
rect 54808 133008 54884 133014
rect 59432 133214 59644 133220
rect 59432 133150 59438 133214
rect 59502 133150 59644 133214
rect 59432 133094 59644 133150
rect 59840 133134 59916 133220
rect 59432 133038 59512 133094
rect 59568 133038 59644 133094
rect 59432 133008 59644 133038
rect 59745 133078 59916 133134
rect 59745 133036 59846 133078
rect 59840 133014 59846 133036
rect 59910 133014 59916 133078
rect 59840 133008 59916 133014
rect 64464 133214 64676 133220
rect 64464 133150 64470 133214
rect 64534 133150 64676 133214
rect 64464 133094 64676 133150
rect 64464 133038 64504 133094
rect 64560 133038 64676 133094
rect 64464 133008 64676 133038
rect 64736 133078 64948 133220
rect 64736 133014 64742 133078
rect 64806 133014 64948 133078
rect 64736 133008 64948 133014
rect 69360 133214 69572 133220
rect 69360 133150 69502 133214
rect 69566 133150 69572 133214
rect 69360 133115 69572 133150
rect 69768 133134 69844 133220
rect 69360 133094 69573 133115
rect 69360 133038 69496 133094
rect 69552 133038 69573 133094
rect 69360 133017 69573 133038
rect 69729 133084 69844 133134
rect 74392 133214 74604 133220
rect 74392 133150 74534 133214
rect 74598 133150 74604 133214
rect 74392 133094 74604 133150
rect 74800 133134 74876 133220
rect 69729 133078 69980 133084
rect 69729 133036 69910 133078
rect 69360 133008 69572 133017
rect 69768 133014 69910 133036
rect 69974 133014 69980 133078
rect 69768 133008 69980 133014
rect 74392 133038 74488 133094
rect 74544 133038 74604 133094
rect 74392 133008 74604 133038
rect 74721 133078 74876 133134
rect 74721 133036 74806 133078
rect 74800 133014 74806 133036
rect 74870 133014 74876 133078
rect 74800 133008 74876 133014
rect 79424 133214 79636 133220
rect 79424 133150 79566 133214
rect 79630 133150 79636 133214
rect 79424 133094 79636 133150
rect 79832 133134 79908 133220
rect 79424 133038 79480 133094
rect 79536 133038 79636 133094
rect 79424 133008 79636 133038
rect 79713 133078 79908 133134
rect 79713 133036 79838 133078
rect 79832 133014 79838 133036
rect 79902 133014 79908 133078
rect 79832 133008 79908 133014
rect 84320 133214 84532 133220
rect 84320 133150 84326 133214
rect 84390 133150 84532 133214
rect 84320 133115 84532 133150
rect 84728 133134 84804 133220
rect 84320 133094 84549 133115
rect 84320 133038 84472 133094
rect 84528 133038 84549 133094
rect 84320 133017 84549 133038
rect 84705 133084 84804 133134
rect 89352 133214 89564 133220
rect 89352 133150 89358 133214
rect 89422 133150 89564 133214
rect 89352 133094 89564 133150
rect 89760 133134 89836 133220
rect 84705 133078 84940 133084
rect 84705 133036 84870 133078
rect 84320 133008 84532 133017
rect 84728 133014 84870 133036
rect 84934 133014 84940 133078
rect 84728 133008 84940 133014
rect 89352 133038 89464 133094
rect 89520 133038 89564 133094
rect 89352 133008 89564 133038
rect 89697 133084 89836 133134
rect 94384 133214 94596 133220
rect 94384 133150 94526 133214
rect 94590 133150 94596 133214
rect 94384 133094 94596 133150
rect 94792 133134 94868 133220
rect 89697 133078 89972 133084
rect 89697 133036 89902 133078
rect 89760 133014 89902 133036
rect 89966 133014 89972 133078
rect 89760 133008 89972 133014
rect 94384 133038 94456 133094
rect 94512 133038 94596 133094
rect 94384 133008 94596 133038
rect 94689 133084 94868 133134
rect 99416 133214 99492 133220
rect 99416 133150 99422 133214
rect 99486 133150 99492 133214
rect 99416 133115 99492 133150
rect 99688 133134 99900 133220
rect 99416 133094 99525 133115
rect 94689 133078 95004 133084
rect 94689 133036 94934 133078
rect 94792 133014 94934 133036
rect 94998 133014 95004 133078
rect 94792 133008 95004 133014
rect 99416 133038 99448 133094
rect 99504 133038 99525 133094
rect 99416 133017 99525 133038
rect 99681 133078 99900 133134
rect 99681 133036 99830 133078
rect 99416 133008 99492 133017
rect 99688 133014 99830 133036
rect 99894 133014 99900 133078
rect 99688 133008 99900 133014
rect 104312 133214 104524 133220
rect 104312 133150 104318 133214
rect 104382 133150 104524 133214
rect 104312 133094 104524 133150
rect 104720 133134 104796 133220
rect 104312 133038 104440 133094
rect 104496 133038 104524 133094
rect 104312 133008 104524 133038
rect 104673 133078 104796 133134
rect 104673 133036 104726 133078
rect 104720 133014 104726 133036
rect 104790 133014 104796 133078
rect 104720 133008 104796 133014
rect 109344 133214 109556 133220
rect 109344 133150 109350 133214
rect 109414 133150 109556 133214
rect 109344 133094 109556 133150
rect 109752 133134 109828 133220
rect 109344 133038 109432 133094
rect 109488 133038 109556 133094
rect 109344 133008 109556 133038
rect 109665 133084 109828 133134
rect 114376 133214 114588 133220
rect 114376 133150 114382 133214
rect 114446 133150 114588 133214
rect 114376 133094 114588 133150
rect 114784 133134 114860 133220
rect 109665 133078 109964 133084
rect 109665 133036 109894 133078
rect 109752 133014 109894 133036
rect 109958 133014 109964 133078
rect 109752 133008 109964 133014
rect 114376 133038 114424 133094
rect 114480 133038 114588 133094
rect 114376 133008 114588 133038
rect 114657 133078 114860 133134
rect 114657 133036 114790 133078
rect 114784 133014 114790 133036
rect 114854 133014 114860 133078
rect 114784 133008 114860 133014
rect 119272 133214 119484 133220
rect 119272 133150 119278 133214
rect 119342 133150 119484 133214
rect 119272 133115 119484 133150
rect 119680 133134 119756 133220
rect 119272 133094 119493 133115
rect 119272 133038 119416 133094
rect 119472 133038 119493 133094
rect 119272 133017 119493 133038
rect 119649 133078 119756 133134
rect 119649 133036 119686 133078
rect 119272 133008 119484 133017
rect 119680 133014 119686 133036
rect 119750 133014 119756 133078
rect 119680 133008 119756 133014
rect 124304 133214 124516 133220
rect 124304 133150 124310 133214
rect 124374 133150 124516 133214
rect 124304 133094 124516 133150
rect 124712 133134 124788 133220
rect 124304 133038 124408 133094
rect 124464 133038 124516 133094
rect 124304 133008 124516 133038
rect 124641 133078 124788 133134
rect 124641 133036 124718 133078
rect 124712 133014 124718 133036
rect 124782 133014 124788 133078
rect 124712 133008 124788 133014
rect 129336 133214 129548 133220
rect 129336 133150 129342 133214
rect 129406 133150 129548 133214
rect 129336 133094 129548 133150
rect 129744 133134 129820 133220
rect 129336 133038 129400 133094
rect 129456 133038 129548 133094
rect 129336 133008 129548 133038
rect 129633 133078 129820 133134
rect 129633 133036 129750 133078
rect 129744 133014 129750 133036
rect 129814 133014 129820 133078
rect 129744 133008 129820 133014
rect 134368 133214 134444 133220
rect 134368 133150 134374 133214
rect 134438 133150 134444 133214
rect 134368 133115 134444 133150
rect 134640 133134 134852 133220
rect 134368 133094 134469 133115
rect 134368 133038 134392 133094
rect 134448 133038 134469 133094
rect 134368 133017 134469 133038
rect 134625 133078 134852 133134
rect 134625 133036 134782 133078
rect 134368 133008 134444 133017
rect 134640 133014 134782 133036
rect 134846 133014 134852 133078
rect 134640 133008 134852 133014
rect 139264 133214 139476 133220
rect 139264 133150 139406 133214
rect 139470 133150 139476 133214
rect 139264 133094 139476 133150
rect 139672 133134 139748 133220
rect 139264 133038 139384 133094
rect 139440 133038 139476 133094
rect 139264 133008 139476 133038
rect 139617 133078 139748 133134
rect 139617 133036 139678 133078
rect 139672 133014 139678 133036
rect 139742 133014 139748 133078
rect 139672 133008 139748 133014
rect 144296 133214 144508 133220
rect 144296 133150 144302 133214
rect 144366 133150 144508 133214
rect 144296 133094 144508 133150
rect 144704 133134 144780 133220
rect 144296 133038 144376 133094
rect 144432 133038 144508 133094
rect 144296 133008 144508 133038
rect 144609 133078 144780 133134
rect 144609 133036 144710 133078
rect 144704 133014 144710 133036
rect 144774 133014 144780 133078
rect 144704 133008 144780 133014
rect 149328 133214 149540 133220
rect 149328 133150 149334 133214
rect 149398 133150 149540 133214
rect 149328 133094 149540 133150
rect 149736 133134 149812 133220
rect 149328 133038 149368 133094
rect 149424 133038 149540 133094
rect 149328 133008 149540 133038
rect 149601 133078 149812 133134
rect 149601 133036 149742 133078
rect 149736 133014 149742 133036
rect 149806 133014 149812 133078
rect 149736 133008 149812 133014
rect 154224 133214 154436 133220
rect 154224 133150 154366 133214
rect 154430 133150 154436 133214
rect 154224 133115 154436 133150
rect 154632 133134 154708 133220
rect 154224 133094 154437 133115
rect 154224 133038 154360 133094
rect 154416 133038 154437 133094
rect 154224 133017 154437 133038
rect 154593 133084 154708 133134
rect 159256 133214 159468 133220
rect 159256 133150 159398 133214
rect 159462 133150 159468 133214
rect 159256 133094 159468 133150
rect 159664 133134 159740 133220
rect 154593 133078 154844 133084
rect 154593 133036 154774 133078
rect 154224 133008 154436 133017
rect 154632 133014 154774 133036
rect 154838 133014 154844 133078
rect 154632 133008 154844 133014
rect 159256 133038 159352 133094
rect 159408 133038 159468 133094
rect 159256 133008 159468 133038
rect 159585 133084 159740 133134
rect 164288 133214 164500 133220
rect 164288 133150 164430 133214
rect 164494 133150 164500 133214
rect 164288 133094 164500 133150
rect 159585 133078 159876 133084
rect 159585 133036 159806 133078
rect 159664 133014 159806 133036
rect 159870 133014 159876 133078
rect 159664 133008 159876 133014
rect 164288 133038 164344 133094
rect 164400 133038 164500 133094
rect 164288 133008 164500 133038
rect 164560 133078 164772 133220
rect 164560 133014 164702 133078
rect 164766 133014 164772 133078
rect 164560 133008 164772 133014
rect 169184 133214 169396 133220
rect 169184 133150 169190 133214
rect 169254 133150 169396 133214
rect 169184 133115 169396 133150
rect 169592 133134 169668 133220
rect 169184 133094 169413 133115
rect 169184 133038 169336 133094
rect 169392 133038 169413 133094
rect 169184 133017 169413 133038
rect 169569 133084 169668 133134
rect 174216 133214 174428 133220
rect 174216 133150 174222 133214
rect 174286 133150 174428 133214
rect 174216 133094 174428 133150
rect 174624 133134 174700 133220
rect 169569 133078 169804 133084
rect 169569 133036 169734 133078
rect 169184 133008 169396 133017
rect 169592 133014 169734 133036
rect 169798 133014 169804 133078
rect 169592 133008 169804 133014
rect 174216 133038 174328 133094
rect 174384 133038 174428 133094
rect 174216 133008 174428 133038
rect 174561 133084 174700 133134
rect 179248 133214 179460 133220
rect 179248 133150 179390 133214
rect 179454 133150 179460 133214
rect 179248 133094 179460 133150
rect 179656 133134 179732 133220
rect 174561 133078 174836 133084
rect 174561 133036 174766 133078
rect 174624 133014 174766 133036
rect 174830 133014 174836 133078
rect 174624 133008 174836 133014
rect 179248 133038 179320 133094
rect 179376 133038 179460 133094
rect 179248 133008 179460 133038
rect 179553 133084 179732 133134
rect 184280 133214 184356 133220
rect 184280 133150 184286 133214
rect 184350 133150 184356 133214
rect 184280 133115 184356 133150
rect 184552 133134 184764 133220
rect 216784 133196 216908 133252
rect 216964 133196 216996 133252
rect 216784 133144 216996 133196
rect 184280 133094 184389 133115
rect 179553 133078 179868 133084
rect 179553 133036 179798 133078
rect 179656 133014 179798 133036
rect 179862 133014 179868 133078
rect 179656 133008 179868 133014
rect 184280 133038 184312 133094
rect 184368 133038 184389 133094
rect 184280 133017 184389 133038
rect 184545 133078 184764 133134
rect 184545 133036 184558 133078
rect 184280 133008 184356 133017
rect 184552 133014 184558 133036
rect 184622 133014 184764 133078
rect 184552 133008 184764 133014
rect 29784 132670 29996 132948
rect 29784 132606 29790 132670
rect 29854 132606 29996 132670
rect 29784 132600 29996 132606
rect 34680 132670 34892 132948
rect 34680 132606 34686 132670
rect 34750 132606 34892 132670
rect 34680 132600 34892 132606
rect 39712 132670 39924 132948
rect 39712 132606 39718 132670
rect 39782 132606 39924 132670
rect 39712 132600 39924 132606
rect 44744 132670 44956 132948
rect 49640 132872 49988 132948
rect 49761 132676 49859 132872
rect 44744 132606 44750 132670
rect 44814 132606 44956 132670
rect 44744 132600 44956 132606
rect 49640 132670 49988 132676
rect 49640 132606 49646 132670
rect 49710 132606 49988 132670
rect 49640 132600 49988 132606
rect 54672 132670 54884 132948
rect 54672 132606 54678 132670
rect 54742 132606 54884 132670
rect 54672 132600 54884 132606
rect 59704 132670 59916 132948
rect 59704 132606 59710 132670
rect 59774 132606 59916 132670
rect 59704 132600 59916 132606
rect 64736 132872 64948 132948
rect 64736 132676 64835 132872
rect 64736 132670 64948 132676
rect 64736 132606 64878 132670
rect 64942 132606 64948 132670
rect 64736 132600 64948 132606
rect 69632 132670 69844 132948
rect 69632 132606 69774 132670
rect 69838 132606 69844 132670
rect 69632 132600 69844 132606
rect 74664 132670 74876 132948
rect 74664 132606 74670 132670
rect 74734 132606 74876 132670
rect 74664 132600 74876 132606
rect 79696 132670 79908 132948
rect 84592 132872 84804 132948
rect 84705 132676 84804 132872
rect 79696 132606 79702 132670
rect 79766 132606 79908 132670
rect 79696 132600 79908 132606
rect 84592 132670 84804 132676
rect 84592 132606 84734 132670
rect 84798 132606 84804 132670
rect 84592 132600 84804 132606
rect 89624 132670 89836 132948
rect 89624 132606 89766 132670
rect 89830 132606 89836 132670
rect 89624 132600 89836 132606
rect 94656 132670 94868 132948
rect 99552 132872 99900 132948
rect 99681 132676 99779 132872
rect 94656 132606 94798 132670
rect 94862 132606 94868 132670
rect 94656 132600 94868 132606
rect 99552 132670 99900 132676
rect 99552 132606 99694 132670
rect 99758 132606 99900 132670
rect 99552 132600 99900 132606
rect 104584 132670 104796 132948
rect 104584 132606 104590 132670
rect 104654 132606 104796 132670
rect 104584 132600 104796 132606
rect 109616 132670 109828 132948
rect 109616 132606 109758 132670
rect 109822 132606 109828 132670
rect 109616 132600 109828 132606
rect 114648 132670 114860 132948
rect 114648 132606 114790 132670
rect 114854 132606 114860 132670
rect 114648 132600 114860 132606
rect 119544 132670 119756 132948
rect 119544 132606 119550 132670
rect 119614 132606 119756 132670
rect 119544 132600 119756 132606
rect 124576 132670 124788 132948
rect 124576 132606 124582 132670
rect 124646 132606 124788 132670
rect 124576 132600 124788 132606
rect 129608 132670 129820 132948
rect 134504 132872 134852 132948
rect 134625 132676 134723 132872
rect 129608 132606 129614 132670
rect 129678 132606 129820 132670
rect 129608 132600 129820 132606
rect 134504 132670 134852 132676
rect 134504 132606 134646 132670
rect 134710 132606 134852 132670
rect 134504 132600 134852 132606
rect 139536 132670 139748 132948
rect 139536 132606 139542 132670
rect 139606 132606 139748 132670
rect 139536 132600 139748 132606
rect 144568 132670 144780 132948
rect 144568 132606 144574 132670
rect 144638 132606 144780 132670
rect 144568 132600 144780 132606
rect 149600 132872 149812 132948
rect 149600 132676 149699 132872
rect 149600 132670 149812 132676
rect 149600 132606 149606 132670
rect 149670 132606 149812 132670
rect 149600 132600 149812 132606
rect 154496 132670 154708 132948
rect 154496 132606 154638 132670
rect 154702 132606 154708 132670
rect 154496 132600 154708 132606
rect 159528 132670 159740 132948
rect 159528 132606 159670 132670
rect 159734 132606 159740 132670
rect 159528 132600 159740 132606
rect 164560 132670 164772 132948
rect 169456 132872 169668 132948
rect 169569 132676 169668 132872
rect 164560 132606 164566 132670
rect 164630 132606 164772 132670
rect 164560 132600 164772 132606
rect 169456 132670 169668 132676
rect 169456 132606 169598 132670
rect 169662 132606 169668 132670
rect 169456 132600 169668 132606
rect 174488 132670 174700 132948
rect 174488 132606 174630 132670
rect 174694 132606 174700 132670
rect 174488 132600 174700 132606
rect 179520 132670 179732 132948
rect 184416 132872 184764 132948
rect 184545 132676 184643 132872
rect 196520 132676 196732 132812
rect 197880 132806 203532 132812
rect 197880 132742 198022 132806
rect 198086 132742 203462 132806
rect 203526 132742 203532 132806
rect 197880 132736 203532 132742
rect 197880 132676 198092 132736
rect 179520 132606 179662 132670
rect 179726 132606 179732 132670
rect 179520 132600 179732 132606
rect 184416 132670 184764 132676
rect 184416 132606 184422 132670
rect 184486 132606 184764 132670
rect 184416 132600 184764 132606
rect 196520 132670 198092 132676
rect 196520 132606 196526 132670
rect 196590 132606 198092 132670
rect 196520 132600 198092 132606
rect 203320 132670 203668 132676
rect 203320 132606 203326 132670
rect 203390 132606 203668 132670
rect 203320 132600 203668 132606
rect 203456 132540 203668 132600
rect 203320 132534 203668 132540
rect 203320 132470 203326 132534
rect 203390 132470 203462 132534
rect 203526 132470 203668 132534
rect 203320 132464 203668 132470
rect 29648 131990 29996 131996
rect 29648 131926 29790 131990
rect 29854 131926 29996 131990
rect 29648 131854 29996 131926
rect 29648 131790 29654 131854
rect 29718 131790 29996 131854
rect 29648 131784 29996 131790
rect 34680 131990 34892 131996
rect 34680 131926 34686 131990
rect 34750 131926 34892 131990
rect 34680 131860 34892 131926
rect 39712 131990 39924 131996
rect 39712 131926 39718 131990
rect 39782 131926 39924 131990
rect 34680 131854 35844 131860
rect 34680 131790 35774 131854
rect 35838 131790 35844 131854
rect 34680 131784 35844 131790
rect 39712 131854 39924 131926
rect 44744 131990 44956 131996
rect 44744 131926 44750 131990
rect 44814 131926 44956 131990
rect 44744 131860 44956 131926
rect 44374 131854 44956 131860
rect 39712 131790 39718 131854
rect 39782 131790 39924 131854
rect 44336 131790 44342 131854
rect 44406 131790 44956 131854
rect 39712 131784 39924 131790
rect 44374 131784 44956 131790
rect 49640 131990 49852 131996
rect 49640 131926 49646 131990
rect 49710 131926 49852 131990
rect 49640 131860 49852 131926
rect 54672 131990 54884 131996
rect 54672 131926 54678 131990
rect 54742 131926 54884 131990
rect 49640 131854 50804 131860
rect 49640 131790 50734 131854
rect 50798 131790 50804 131854
rect 49640 131784 50804 131790
rect 54672 131854 54884 131926
rect 54672 131790 54678 131854
rect 54742 131790 54884 131854
rect 54672 131784 54884 131790
rect 59704 131990 59916 131996
rect 59704 131926 59710 131990
rect 59774 131926 59916 131990
rect 59704 131860 59916 131926
rect 64600 131990 64948 131996
rect 64600 131926 64878 131990
rect 64942 131926 64948 131990
rect 59704 131854 60868 131860
rect 59704 131790 60798 131854
rect 60862 131790 60868 131854
rect 59704 131784 60868 131790
rect 64600 131854 64948 131926
rect 69632 131990 69844 131996
rect 69632 131926 69774 131990
rect 69838 131926 69844 131990
rect 69632 131860 69844 131926
rect 69262 131854 69844 131860
rect 64600 131790 64606 131854
rect 64670 131790 64948 131854
rect 69224 131790 69230 131854
rect 69294 131790 69844 131854
rect 64600 131784 64948 131790
rect 69262 131784 69844 131790
rect 74664 131990 74876 131996
rect 74664 131926 74670 131990
rect 74734 131926 74876 131990
rect 74664 131854 74876 131926
rect 79696 131990 79908 131996
rect 79696 131926 79702 131990
rect 79766 131926 79908 131990
rect 79696 131860 79908 131926
rect 84592 131990 84804 131996
rect 84592 131926 84734 131990
rect 84798 131926 84804 131990
rect 84592 131860 84804 131926
rect 79326 131854 79908 131860
rect 84222 131854 84804 131860
rect 74664 131790 74670 131854
rect 74734 131790 74876 131854
rect 79288 131790 79294 131854
rect 79358 131790 79908 131854
rect 84184 131790 84190 131854
rect 84254 131790 84804 131854
rect 74664 131784 74876 131790
rect 79326 131784 79908 131790
rect 84222 131784 84804 131790
rect 89624 131990 89836 131996
rect 89624 131926 89766 131990
rect 89830 131926 89836 131990
rect 89624 131854 89836 131926
rect 89624 131790 89630 131854
rect 89694 131790 89836 131854
rect 89624 131784 89836 131790
rect 94656 131990 94868 131996
rect 94656 131926 94798 131990
rect 94862 131926 94868 131990
rect 94656 131854 94868 131926
rect 94656 131790 94662 131854
rect 94726 131790 94868 131854
rect 94656 131784 94868 131790
rect 99552 131990 99900 131996
rect 99552 131926 99694 131990
rect 99758 131926 99900 131990
rect 99552 131854 99900 131926
rect 104584 131990 104796 131996
rect 104584 131926 104590 131990
rect 104654 131926 104796 131990
rect 104584 131860 104796 131926
rect 104350 131854 104796 131860
rect 99552 131790 99558 131854
rect 99622 131790 99900 131854
rect 104312 131790 104318 131854
rect 104382 131790 104796 131854
rect 99552 131784 99900 131790
rect 104350 131784 104796 131790
rect 109616 131990 109828 131996
rect 109616 131926 109758 131990
rect 109822 131926 109828 131990
rect 109616 131854 109828 131926
rect 114512 131990 114860 131996
rect 114512 131926 114790 131990
rect 114854 131926 114860 131990
rect 114512 131860 114860 131926
rect 114278 131854 114860 131860
rect 109616 131790 109622 131854
rect 109686 131790 109828 131854
rect 114240 131790 114246 131854
rect 114310 131790 114860 131854
rect 109616 131784 109828 131790
rect 114278 131784 114860 131790
rect 119544 131990 119756 131996
rect 119544 131926 119550 131990
rect 119614 131926 119756 131990
rect 119544 131860 119756 131926
rect 124576 131990 124788 131996
rect 124576 131926 124582 131990
rect 124646 131926 124788 131990
rect 119544 131854 120300 131860
rect 119544 131790 120230 131854
rect 120294 131790 120300 131854
rect 119544 131784 120300 131790
rect 124576 131854 124788 131926
rect 129608 131990 129820 131996
rect 129608 131926 129614 131990
rect 129678 131926 129820 131990
rect 129608 131860 129820 131926
rect 129238 131854 129820 131860
rect 124576 131790 124582 131854
rect 124646 131790 124788 131854
rect 129200 131790 129206 131854
rect 129270 131790 129820 131854
rect 124576 131784 124788 131790
rect 129238 131784 129820 131790
rect 134504 131990 134716 131996
rect 134504 131926 134646 131990
rect 134710 131926 134716 131990
rect 134504 131860 134716 131926
rect 139536 131990 139748 131996
rect 139536 131926 139542 131990
rect 139606 131926 139748 131990
rect 134504 131854 135668 131860
rect 134504 131790 135598 131854
rect 135662 131790 135668 131854
rect 134504 131784 135668 131790
rect 139536 131854 139748 131926
rect 139536 131790 139542 131854
rect 139606 131790 139748 131854
rect 139536 131784 139748 131790
rect 144568 131990 144780 131996
rect 144568 131926 144574 131990
rect 144638 131926 144780 131990
rect 144568 131860 144780 131926
rect 149464 131990 149812 131996
rect 149464 131926 149606 131990
rect 149670 131926 149812 131990
rect 144568 131854 145324 131860
rect 144568 131790 145254 131854
rect 145318 131790 145324 131854
rect 144568 131784 145324 131790
rect 149464 131854 149812 131926
rect 154496 131990 154708 131996
rect 154496 131926 154638 131990
rect 154702 131926 154708 131990
rect 154496 131860 154708 131926
rect 154126 131854 154708 131860
rect 149464 131790 149470 131854
rect 149534 131790 149812 131854
rect 154088 131790 154094 131854
rect 154158 131790 154708 131854
rect 149464 131784 149812 131790
rect 154126 131784 154708 131790
rect 159528 131990 159740 131996
rect 159528 131926 159670 131990
rect 159734 131926 159740 131990
rect 159528 131860 159740 131926
rect 164560 131990 164772 131996
rect 164560 131926 164566 131990
rect 164630 131926 164772 131990
rect 164560 131860 164772 131926
rect 169456 131990 169668 131996
rect 169456 131926 169598 131990
rect 169662 131926 169668 131990
rect 169456 131860 169668 131926
rect 174488 131990 174700 131996
rect 174488 131926 174630 131990
rect 174694 131926 174700 131990
rect 159528 131854 160284 131860
rect 159528 131790 160214 131854
rect 160278 131790 160284 131854
rect 159528 131784 160284 131790
rect 164560 131854 165588 131860
rect 164560 131790 165518 131854
rect 165582 131790 165588 131854
rect 164560 131784 165588 131790
rect 169456 131854 170212 131860
rect 169456 131790 170142 131854
rect 170206 131790 170212 131854
rect 169456 131784 170212 131790
rect 174488 131854 174700 131926
rect 174488 131790 174494 131854
rect 174558 131790 174700 131854
rect 174488 131784 174700 131790
rect 179520 131990 179732 131996
rect 179520 131926 179662 131990
rect 179726 131926 179732 131990
rect 179520 131854 179732 131926
rect 179520 131790 179526 131854
rect 179590 131790 179732 131854
rect 179520 131784 179732 131790
rect 184416 131990 184764 131996
rect 184416 131926 184422 131990
rect 184486 131926 184764 131990
rect 184416 131854 184764 131926
rect 184416 131790 184422 131854
rect 184486 131790 184764 131854
rect 184416 131784 184764 131790
rect 1632 131588 1844 131724
rect 1224 131582 1844 131588
rect 1224 131518 1230 131582
rect 1294 131572 1844 131582
rect 1294 131518 1702 131572
rect 1224 131516 1702 131518
rect 1758 131516 1844 131572
rect 1224 131512 1844 131516
rect 1632 131376 1844 131512
rect 216784 131588 216996 131724
rect 216784 131582 217540 131588
rect 216784 131572 217470 131582
rect 216784 131516 216908 131572
rect 216964 131518 217470 131572
rect 217534 131518 217540 131582
rect 216964 131516 217540 131518
rect 216784 131512 217540 131516
rect 196520 131446 196732 131452
rect 196520 131382 196662 131446
rect 196726 131382 196732 131446
rect 196520 131316 196732 131382
rect 197880 131446 203532 131452
rect 197880 131382 203462 131446
rect 203526 131382 203532 131446
rect 197880 131376 203532 131382
rect 216784 131376 216996 131512
rect 197880 131316 198092 131376
rect 29784 131310 29996 131316
rect 29784 131246 29926 131310
rect 29990 131246 29996 131310
rect 29784 131174 29996 131246
rect 29784 131110 29926 131174
rect 29990 131110 29996 131174
rect 29784 131104 29996 131110
rect 34816 131310 35028 131316
rect 34816 131246 34822 131310
rect 34886 131246 35028 131310
rect 34816 131174 35028 131246
rect 34816 131110 34958 131174
rect 35022 131110 35028 131174
rect 34816 131104 35028 131110
rect 39712 131310 40060 131316
rect 39712 131246 39854 131310
rect 39918 131246 40060 131310
rect 39712 131174 40060 131246
rect 39712 131110 39990 131174
rect 40054 131110 40060 131174
rect 39712 131104 40060 131110
rect 44744 131310 44956 131316
rect 44744 131246 44886 131310
rect 44950 131246 44956 131310
rect 44744 131174 44956 131246
rect 44744 131110 44886 131174
rect 44950 131110 44956 131174
rect 44744 131104 44956 131110
rect 49776 131310 49988 131316
rect 49776 131246 49918 131310
rect 49982 131246 49988 131310
rect 49776 131174 49988 131246
rect 49776 131110 49918 131174
rect 49982 131110 49988 131174
rect 49776 131104 49988 131110
rect 54808 131310 55020 131316
rect 54808 131246 54814 131310
rect 54878 131246 55020 131310
rect 54808 131174 55020 131246
rect 54808 131110 54814 131174
rect 54878 131110 55020 131174
rect 54808 131104 55020 131110
rect 59704 131310 59916 131316
rect 59704 131246 59846 131310
rect 59910 131246 59916 131310
rect 59704 131180 59916 131246
rect 64736 131310 64948 131316
rect 64736 131246 64742 131310
rect 64806 131246 64948 131310
rect 59704 131174 60052 131180
rect 59704 131110 59982 131174
rect 60046 131110 60052 131174
rect 59704 131104 60052 131110
rect 64736 131174 64948 131246
rect 64736 131110 64878 131174
rect 64942 131110 64948 131174
rect 64736 131104 64948 131110
rect 69768 131310 69980 131316
rect 69768 131246 69910 131310
rect 69974 131246 69980 131310
rect 69768 131174 69980 131246
rect 69768 131110 69910 131174
rect 69974 131110 69980 131174
rect 69768 131104 69980 131110
rect 74664 131310 75012 131316
rect 74664 131246 74806 131310
rect 74870 131246 75012 131310
rect 74664 131174 75012 131246
rect 74664 131110 74942 131174
rect 75006 131110 75012 131174
rect 74664 131104 75012 131110
rect 79696 131310 79908 131316
rect 79696 131246 79838 131310
rect 79902 131246 79908 131310
rect 79696 131174 79908 131246
rect 79696 131110 79838 131174
rect 79902 131110 79908 131174
rect 79696 131104 79908 131110
rect 84728 131310 84940 131316
rect 84728 131246 84870 131310
rect 84934 131246 84940 131310
rect 84728 131174 84940 131246
rect 84728 131110 84870 131174
rect 84934 131110 84940 131174
rect 84728 131104 84940 131110
rect 89760 131310 89972 131316
rect 89760 131246 89902 131310
rect 89966 131246 89972 131310
rect 89760 131174 89972 131246
rect 89760 131110 89902 131174
rect 89966 131110 89972 131174
rect 89760 131104 89972 131110
rect 94656 131310 94966 131316
rect 99688 131310 99900 131316
rect 94656 131246 94934 131310
rect 94998 131246 95004 131310
rect 99688 131246 99830 131310
rect 99894 131246 99900 131310
rect 94656 131240 94966 131246
rect 94656 131180 94868 131240
rect 94656 131174 95004 131180
rect 94656 131110 94934 131174
rect 94998 131110 95004 131174
rect 94656 131104 95004 131110
rect 99688 131174 99900 131246
rect 99688 131110 99830 131174
rect 99894 131110 99900 131174
rect 99688 131104 99900 131110
rect 104720 131310 104932 131316
rect 104720 131246 104726 131310
rect 104790 131246 104932 131310
rect 104720 131174 104932 131246
rect 104720 131110 104862 131174
rect 104926 131110 104932 131174
rect 104720 131104 104932 131110
rect 109616 131310 109964 131316
rect 109616 131246 109894 131310
rect 109958 131246 109964 131310
rect 109616 131174 109964 131246
rect 109616 131110 109894 131174
rect 109958 131110 109964 131174
rect 109616 131104 109964 131110
rect 114648 131310 114860 131316
rect 114648 131246 114654 131310
rect 114718 131246 114860 131310
rect 114648 131174 114860 131246
rect 114648 131110 114654 131174
rect 114718 131110 114860 131174
rect 114648 131104 114860 131110
rect 119680 131310 119892 131316
rect 119680 131246 119686 131310
rect 119750 131246 119892 131310
rect 119680 131174 119892 131246
rect 119680 131110 119822 131174
rect 119886 131110 119892 131174
rect 119680 131104 119892 131110
rect 124576 131310 124924 131316
rect 124576 131246 124718 131310
rect 124782 131246 124924 131310
rect 124576 131174 124924 131246
rect 124576 131110 124854 131174
rect 124918 131110 124924 131174
rect 124576 131104 124924 131110
rect 129608 131310 129820 131316
rect 129608 131246 129750 131310
rect 129814 131246 129820 131310
rect 129608 131174 129820 131246
rect 129608 131110 129750 131174
rect 129814 131110 129820 131174
rect 129608 131104 129820 131110
rect 134640 131310 134852 131316
rect 134640 131246 134782 131310
rect 134846 131246 134852 131310
rect 134640 131174 134852 131246
rect 134640 131110 134782 131174
rect 134846 131110 134852 131174
rect 134640 131104 134852 131110
rect 139672 131310 139884 131316
rect 139672 131246 139678 131310
rect 139742 131246 139884 131310
rect 139672 131174 139884 131246
rect 139672 131110 139814 131174
rect 139878 131110 139884 131174
rect 139672 131104 139884 131110
rect 144568 131310 144780 131316
rect 144568 131246 144710 131310
rect 144774 131246 144780 131310
rect 144568 131180 144780 131246
rect 149600 131310 149812 131316
rect 149600 131246 149742 131310
rect 149806 131246 149812 131310
rect 144568 131174 144916 131180
rect 144568 131110 144846 131174
rect 144910 131110 144916 131174
rect 144568 131104 144916 131110
rect 149600 131174 149812 131246
rect 149600 131110 149606 131174
rect 149670 131110 149812 131174
rect 149600 131104 149812 131110
rect 154632 131310 154844 131316
rect 154632 131246 154774 131310
rect 154838 131246 154844 131310
rect 154632 131174 154844 131246
rect 154632 131110 154774 131174
rect 154838 131110 154844 131174
rect 154632 131104 154844 131110
rect 159528 131310 159876 131316
rect 159528 131246 159806 131310
rect 159870 131246 159876 131310
rect 159528 131174 159876 131246
rect 159528 131110 159806 131174
rect 159870 131110 159876 131174
rect 159528 131104 159876 131110
rect 164560 131310 164772 131316
rect 164560 131246 164702 131310
rect 164766 131246 164772 131310
rect 164560 131174 164772 131246
rect 164560 131110 164702 131174
rect 164766 131110 164772 131174
rect 164560 131104 164772 131110
rect 169592 131310 169804 131316
rect 169592 131246 169734 131310
rect 169798 131246 169804 131310
rect 169592 131174 169804 131246
rect 169592 131110 169734 131174
rect 169798 131110 169804 131174
rect 169592 131104 169804 131110
rect 174624 131310 174836 131316
rect 174624 131246 174766 131310
rect 174830 131246 174836 131310
rect 174624 131174 174836 131246
rect 174624 131110 174630 131174
rect 174694 131110 174836 131174
rect 174624 131104 174836 131110
rect 179520 131310 179830 131316
rect 184552 131310 184764 131316
rect 179520 131246 179798 131310
rect 179862 131246 179868 131310
rect 184552 131246 184558 131310
rect 184622 131246 184764 131310
rect 179520 131240 179830 131246
rect 179520 131180 179732 131240
rect 179520 131174 179868 131180
rect 179520 131110 179798 131174
rect 179862 131110 179868 131174
rect 179520 131104 179868 131110
rect 184552 131174 184764 131246
rect 196520 131310 198092 131316
rect 196520 131246 197886 131310
rect 197950 131246 198092 131310
rect 196520 131240 198092 131246
rect 184552 131110 184694 131174
rect 184758 131110 184764 131174
rect 184552 131104 184764 131110
rect 203456 131174 203668 131180
rect 203456 131110 203598 131174
rect 203662 131110 203668 131174
rect 29863 131102 29961 131104
rect 34855 131102 34953 131104
rect 39847 131102 39945 131104
rect 44839 131102 44937 131104
rect 49831 131102 49929 131104
rect 54823 131102 54921 131104
rect 59815 131102 59913 131104
rect 64807 131102 64905 131104
rect 69799 131102 69897 131104
rect 74791 131102 74889 131104
rect 79783 131102 79881 131104
rect 84775 131102 84873 131104
rect 89767 131102 89865 131104
rect 94759 131102 94857 131104
rect 99751 131102 99849 131104
rect 104743 131102 104841 131104
rect 109735 131102 109833 131104
rect 114727 131102 114825 131104
rect 119719 131102 119817 131104
rect 124711 131102 124809 131104
rect 129703 131102 129801 131104
rect 134695 131102 134793 131104
rect 139687 131102 139785 131104
rect 144679 131102 144777 131104
rect 149671 131102 149769 131104
rect 154663 131102 154761 131104
rect 159655 131102 159753 131104
rect 164647 131102 164745 131104
rect 169639 131102 169737 131104
rect 174631 131102 174729 131104
rect 179623 131102 179721 131104
rect 184615 131102 184713 131104
rect 203456 131038 203668 131110
rect 203456 130974 203598 131038
rect 203662 130974 203668 131038
rect 203456 130968 203668 130974
rect 190870 130436 190936 130439
rect 203479 130436 203545 130439
rect 190870 130434 203545 130436
rect 190870 130378 190875 130434
rect 190931 130378 203484 130434
rect 203540 130378 203545 130434
rect 190870 130376 203545 130378
rect 190870 130373 190936 130376
rect 203479 130373 203545 130376
rect 196520 130086 198092 130092
rect 196520 130022 196526 130086
rect 196590 130022 198092 130086
rect 196520 130016 198092 130022
rect 1632 129892 1844 129956
rect 1632 129836 1702 129892
rect 1758 129836 1844 129892
rect 1632 129820 1844 129836
rect 1224 129814 1844 129820
rect 1224 129750 1230 129814
rect 1294 129750 1844 129814
rect 1224 129744 1844 129750
rect 196520 129814 196732 130016
rect 196520 129750 196526 129814
rect 196590 129750 196732 129814
rect 196520 129744 196732 129750
rect 197880 129744 198092 130016
rect 216784 129950 217540 129956
rect 216784 129892 217470 129950
rect 216784 129836 216908 129892
rect 216964 129886 217470 129892
rect 217534 129886 217540 129950
rect 216964 129880 217540 129886
rect 216964 129836 216996 129880
rect 203358 129814 203668 129820
rect 203320 129750 203326 129814
rect 203390 129750 203668 129814
rect 203358 129744 203668 129750
rect 203456 129678 203668 129744
rect 203456 129614 203462 129678
rect 203526 129614 203668 129678
rect 203456 129608 203668 129614
rect 215016 129684 215228 129820
rect 215696 129684 215908 129820
rect 216784 129744 216996 129836
rect 215016 129678 218220 129684
rect 215016 129614 218150 129678
rect 218214 129614 218220 129678
rect 215016 129608 218220 129614
rect 190994 129022 191060 129025
rect 203479 129022 203545 129025
rect 190994 129020 203545 129022
rect 190994 128964 190999 129020
rect 191055 128964 203484 129020
rect 203540 128964 203545 129020
rect 190994 128962 203545 128964
rect 190994 128959 191060 128962
rect 203479 128959 203545 128962
rect 29920 128726 31492 128732
rect 29920 128662 29926 128726
rect 29990 128662 31492 128726
rect 29920 128656 31492 128662
rect 29920 128596 30268 128656
rect 28870 128590 30268 128596
rect 28832 128526 28838 128590
rect 28902 128526 30268 128590
rect 28870 128520 30268 128526
rect 31280 128596 31492 128656
rect 32504 128726 35164 128732
rect 32504 128662 34958 128726
rect 35022 128662 35164 128726
rect 32504 128656 35164 128662
rect 32504 128596 32716 128656
rect 31280 128520 32716 128596
rect 33728 128520 33940 128656
rect 34952 128596 35164 128656
rect 36176 128596 36388 128732
rect 37400 128596 37748 128732
rect 38760 128596 38972 128732
rect 39984 128726 40196 128732
rect 39984 128662 39990 128726
rect 40054 128662 40196 128726
rect 39984 128596 40196 128662
rect 41208 128656 43868 128732
rect 41208 128596 41420 128656
rect 34952 128520 41420 128596
rect 42432 128520 42644 128656
rect 43656 128596 43868 128656
rect 44880 128726 48900 128732
rect 44880 128662 44886 128726
rect 44950 128662 48900 128726
rect 44880 128656 48900 128662
rect 44880 128596 45228 128656
rect 43656 128520 45228 128596
rect 46240 128520 46452 128656
rect 47464 128520 47676 128656
rect 48688 128596 48900 128656
rect 49912 128726 52708 128732
rect 49912 128662 49918 128726
rect 49982 128662 52708 128726
rect 49912 128656 52708 128662
rect 49912 128596 50124 128656
rect 48688 128520 50124 128596
rect 51136 128520 51484 128656
rect 52496 128596 52708 128656
rect 53720 128726 54884 128732
rect 53720 128662 54814 128726
rect 54878 128662 54884 128726
rect 53720 128656 54884 128662
rect 54944 128656 56380 128732
rect 53720 128596 53932 128656
rect 54944 128596 55156 128656
rect 52496 128520 55156 128596
rect 56168 128596 56380 128656
rect 57392 128596 57604 128732
rect 58616 128726 60188 128732
rect 58616 128662 59982 128726
rect 60046 128662 60188 128726
rect 58616 128656 60188 128662
rect 58616 128596 58964 128656
rect 56168 128520 58964 128596
rect 59976 128596 60188 128656
rect 61200 128596 61412 128732
rect 62424 128726 70116 128732
rect 62424 128662 64878 128726
rect 64942 128662 69910 128726
rect 69974 128662 70116 128726
rect 62424 128656 70116 128662
rect 62424 128596 62636 128656
rect 59976 128520 62636 128596
rect 63648 128520 63860 128656
rect 64872 128520 65084 128656
rect 66096 128520 66444 128656
rect 67456 128520 67668 128656
rect 68680 128520 68892 128656
rect 69904 128596 70116 128656
rect 71128 128656 73924 128732
rect 71128 128596 71340 128656
rect 69904 128520 71340 128596
rect 72352 128520 72700 128656
rect 73712 128596 73924 128656
rect 74936 128726 77596 128732
rect 74936 128662 74942 128726
rect 75006 128662 77596 128726
rect 74936 128656 77596 128662
rect 74936 128596 75148 128656
rect 73712 128520 75148 128596
rect 76160 128520 76372 128656
rect 77384 128596 77596 128656
rect 78608 128596 78820 128732
rect 79832 128726 80180 128732
rect 79832 128662 79838 128726
rect 79902 128662 80180 128726
rect 79832 128596 80180 128662
rect 81192 128596 81404 128732
rect 82416 128596 82628 128732
rect 83640 128726 86300 128732
rect 83640 128662 84870 128726
rect 84934 128662 86300 128726
rect 83640 128656 86300 128662
rect 83640 128596 83852 128656
rect 77384 128520 83852 128596
rect 84864 128520 85076 128656
rect 86088 128596 86300 128656
rect 87312 128726 90108 128732
rect 87312 128662 89902 128726
rect 89966 128662 90108 128726
rect 87312 128656 90108 128662
rect 87312 128596 87660 128656
rect 86088 128520 87660 128596
rect 88672 128520 88884 128656
rect 89896 128596 90108 128656
rect 91120 128596 91332 128732
rect 92344 128656 93916 128732
rect 92344 128596 92556 128656
rect 89896 128520 92556 128596
rect 93568 128596 93916 128656
rect 94928 128726 95140 128732
rect 94928 128662 94934 128726
rect 94998 128662 95140 128726
rect 94928 128596 95140 128662
rect 96152 128656 98812 128732
rect 96152 128596 96364 128656
rect 93568 128520 96364 128596
rect 97376 128520 97588 128656
rect 98600 128596 98812 128656
rect 99824 128726 100036 128732
rect 99824 128662 99830 128726
rect 99894 128662 100036 128726
rect 99824 128596 100036 128662
rect 101048 128596 101396 128732
rect 102408 128596 102620 128732
rect 103632 128596 103844 128732
rect 104856 128726 111324 128732
rect 104856 128662 104862 128726
rect 104926 128662 109894 128726
rect 109958 128662 111324 128726
rect 104856 128656 111324 128662
rect 104856 128596 105068 128656
rect 98600 128520 105068 128596
rect 106080 128520 106292 128656
rect 107304 128520 107516 128656
rect 108528 128520 108876 128656
rect 109888 128520 110100 128656
rect 111112 128596 111324 128656
rect 112336 128596 112548 128732
rect 113560 128726 114724 128732
rect 113560 128662 114654 128726
rect 114718 128662 114724 128726
rect 113560 128656 114724 128662
rect 114784 128656 116356 128732
rect 113560 128596 113772 128656
rect 114784 128596 115132 128656
rect 111112 128520 115132 128596
rect 116144 128596 116356 128656
rect 117368 128726 121252 128732
rect 117368 128662 119822 128726
rect 119886 128662 121252 128726
rect 117368 128656 121252 128662
rect 117368 128596 117580 128656
rect 116144 128520 117580 128596
rect 118592 128520 118804 128656
rect 119816 128520 120028 128656
rect 121040 128596 121252 128656
rect 122264 128656 123836 128732
rect 122264 128596 122612 128656
rect 121040 128520 122612 128596
rect 123624 128596 123836 128656
rect 124848 128726 125060 128732
rect 124848 128662 124854 128726
rect 124918 128662 125060 128726
rect 124848 128596 125060 128662
rect 126072 128656 128732 128732
rect 126072 128596 126284 128656
rect 123624 128520 126284 128596
rect 127296 128520 127508 128656
rect 128520 128596 128732 128656
rect 129744 128726 130092 128732
rect 129744 128662 129750 128726
rect 129814 128662 130092 128726
rect 129744 128596 130092 128662
rect 131104 128656 132540 128732
rect 131104 128596 131316 128656
rect 128520 128520 131316 128596
rect 132328 128596 132540 128656
rect 133552 128596 133764 128732
rect 134776 128726 137572 128732
rect 134776 128662 134782 128726
rect 134846 128662 137572 128726
rect 134776 128656 137572 128662
rect 134776 128596 134988 128656
rect 132328 128520 134988 128596
rect 136000 128520 136348 128656
rect 137360 128596 137572 128656
rect 138584 128726 141244 128732
rect 138584 128662 139814 128726
rect 139878 128662 141244 128726
rect 138584 128656 141244 128662
rect 138584 128596 138796 128656
rect 137360 128520 138796 128596
rect 139808 128520 140020 128656
rect 141032 128596 141244 128656
rect 142256 128596 142468 128732
rect 143480 128596 143828 128732
rect 144840 128726 146276 128732
rect 144840 128662 144846 128726
rect 144910 128662 146276 128726
rect 144840 128656 146276 128662
rect 144840 128596 145052 128656
rect 141032 128520 145052 128596
rect 146064 128596 146276 128656
rect 147288 128726 149676 128732
rect 147288 128662 149606 128726
rect 149670 128662 149676 128726
rect 147288 128656 149676 128662
rect 147288 128596 147500 128656
rect 146064 128520 147500 128596
rect 148512 128596 148724 128656
rect 149736 128596 149948 128732
rect 150960 128656 153756 128732
rect 150960 128596 151308 128656
rect 148512 128520 151308 128596
rect 152320 128520 152532 128656
rect 153544 128596 153756 128656
rect 154768 128726 154980 128732
rect 154768 128662 154774 128726
rect 154838 128662 154980 128726
rect 154768 128596 154980 128662
rect 155992 128656 157564 128732
rect 155992 128596 156204 128656
rect 153544 128520 156204 128596
rect 157216 128596 157564 128656
rect 158576 128596 158788 128732
rect 159800 128726 163684 128732
rect 159800 128662 159806 128726
rect 159870 128662 163684 128726
rect 159800 128656 163684 128662
rect 159800 128596 160012 128656
rect 157216 128520 160012 128596
rect 161024 128520 161236 128656
rect 162248 128520 162460 128656
rect 163472 128596 163684 128656
rect 164696 128726 165044 128732
rect 164696 128662 164702 128726
rect 164766 128662 165044 128726
rect 164696 128596 165044 128662
rect 166056 128596 166268 128732
rect 167280 128596 167492 128732
rect 168504 128726 171164 128732
rect 168504 128662 169734 128726
rect 169798 128662 171164 128726
rect 168504 128656 171164 128662
rect 168504 128596 168716 128656
rect 163472 128520 168716 128596
rect 169728 128520 169940 128656
rect 170952 128596 171164 128656
rect 172176 128726 174700 128732
rect 172176 128662 174630 128726
rect 174694 128662 174700 128726
rect 172176 128656 174700 128662
rect 172176 128596 172524 128656
rect 170952 128520 172524 128596
rect 173536 128596 173748 128656
rect 174760 128596 174972 128732
rect 175984 128596 176196 128732
rect 177208 128726 180004 128732
rect 177208 128662 179798 128726
rect 179862 128662 180004 128726
rect 177208 128656 180004 128662
rect 177208 128596 177420 128656
rect 173536 128520 177420 128596
rect 178432 128520 178780 128656
rect 179792 128596 180004 128656
rect 181016 128656 183676 128732
rect 181016 128596 181228 128656
rect 179792 128520 181228 128596
rect 182240 128520 182452 128656
rect 183464 128596 183676 128656
rect 184688 128726 184900 128732
rect 184688 128662 184694 128726
rect 184758 128662 184900 128726
rect 184688 128596 184900 128662
rect 185912 128596 186260 128732
rect 187272 128656 188708 128732
rect 187272 128596 187484 128656
rect 183464 128520 187484 128596
rect 188496 128596 188708 128656
rect 188496 128590 190476 128596
rect 188496 128526 190406 128590
rect 190470 128526 190476 128590
rect 188496 128520 190476 128526
rect 196520 128460 196732 128596
rect 197880 128590 198092 128596
rect 197880 128526 197886 128590
rect 197950 128526 198092 128590
rect 197880 128460 198092 128526
rect 196520 128454 198092 128460
rect 196520 128390 196662 128454
rect 196726 128390 198092 128454
rect 196520 128384 198092 128390
rect 203456 128454 203668 128460
rect 203456 128390 203598 128454
rect 203662 128390 203668 128454
rect 1632 128212 1844 128324
rect 1632 128188 1702 128212
rect 1224 128182 1702 128188
rect 1224 128118 1230 128182
rect 1294 128156 1702 128182
rect 1758 128156 1844 128212
rect 1294 128118 1844 128156
rect 1224 128112 1844 128118
rect 203456 128112 203668 128390
rect 215016 128384 215908 128460
rect 215016 128112 215228 128384
rect 215696 128188 215908 128384
rect 216784 128318 217540 128324
rect 216784 128254 217470 128318
rect 217534 128254 217540 128318
rect 216784 128248 217540 128254
rect 216784 128212 216996 128248
rect 216784 128188 216908 128212
rect 215696 128156 216908 128188
rect 216964 128156 216996 128212
rect 215696 128112 216996 128156
rect 216487 127907 216493 127909
rect 196284 127847 196344 127907
rect 203344 127847 216493 127907
rect 216487 127845 216493 127847
rect 216557 127845 216563 127909
rect 194853 127608 194919 127611
rect 203479 127608 203545 127611
rect 194853 127606 203545 127608
rect 194853 127550 194858 127606
rect 194914 127550 203484 127606
rect 203540 127550 203545 127606
rect 194853 127548 203545 127550
rect 194853 127545 194919 127548
rect 203479 127545 203545 127548
rect 29512 127230 29724 127236
rect 29512 127166 29654 127230
rect 29718 127166 29724 127230
rect 29512 127094 29724 127166
rect 29512 127030 29654 127094
rect 29718 127030 29724 127094
rect 29512 127024 29724 127030
rect 30464 127160 31084 127236
rect 30464 127024 30676 127160
rect 30736 127094 31084 127160
rect 30736 127030 30878 127094
rect 30942 127030 31084 127094
rect 30736 127024 31084 127030
rect 31688 127100 31900 127236
rect 32096 127100 32308 127236
rect 31688 127094 32308 127100
rect 31688 127030 31694 127094
rect 31758 127030 32308 127094
rect 31688 127024 32308 127030
rect 32912 127160 33532 127236
rect 32912 127094 33124 127160
rect 32912 127030 32918 127094
rect 32982 127030 33124 127094
rect 32912 127024 33124 127030
rect 33320 127094 33532 127160
rect 33320 127030 33462 127094
rect 33526 127030 33532 127094
rect 33320 127024 33532 127030
rect 34136 127100 34348 127236
rect 34544 127100 34756 127236
rect 34136 127094 34756 127100
rect 34136 127030 34142 127094
rect 34206 127030 34686 127094
rect 34750 127030 34756 127094
rect 34136 127024 34756 127030
rect 35360 127230 35980 127236
rect 35360 127166 35774 127230
rect 35838 127166 35980 127230
rect 35360 127160 35980 127166
rect 35360 127024 35572 127160
rect 35768 127094 35980 127160
rect 35768 127030 35910 127094
rect 35974 127030 35980 127094
rect 35768 127024 35980 127030
rect 36584 127100 36932 127236
rect 36992 127100 37204 127236
rect 36584 127094 37204 127100
rect 36584 127030 36590 127094
rect 36654 127030 37134 127094
rect 37198 127030 37204 127094
rect 36584 127024 37204 127030
rect 37944 127100 38156 127236
rect 38216 127100 38564 127236
rect 37944 127094 38564 127100
rect 37944 127030 38086 127094
rect 38150 127030 38564 127094
rect 37944 127024 38564 127030
rect 39168 127230 39788 127236
rect 39168 127166 39718 127230
rect 39782 127166 39788 127230
rect 39168 127160 39788 127166
rect 39168 127100 39380 127160
rect 39168 127094 39516 127100
rect 39168 127030 39446 127094
rect 39510 127030 39516 127094
rect 39168 127024 39516 127030
rect 39576 127024 39788 127160
rect 40392 127100 40604 127236
rect 40800 127100 41012 127236
rect 40392 127094 41012 127100
rect 40392 127030 40398 127094
rect 40462 127030 41012 127094
rect 40392 127024 41012 127030
rect 41616 127160 42236 127236
rect 41616 127094 41828 127160
rect 41616 127030 41622 127094
rect 41686 127030 41828 127094
rect 41616 127024 41828 127030
rect 42024 127094 42236 127160
rect 42024 127030 42166 127094
rect 42230 127030 42236 127094
rect 42024 127024 42236 127030
rect 42840 127094 43052 127236
rect 42840 127030 42982 127094
rect 43046 127030 43052 127094
rect 42840 127024 43052 127030
rect 43248 127094 43460 127236
rect 43248 127030 43254 127094
rect 43318 127030 43460 127094
rect 43248 127024 43460 127030
rect 44064 127230 44684 127236
rect 44064 127166 44342 127230
rect 44406 127166 44684 127230
rect 44064 127160 44684 127166
rect 44064 127024 44412 127160
rect 44472 127094 44684 127160
rect 44472 127030 44614 127094
rect 44678 127030 44684 127094
rect 44472 127024 44684 127030
rect 45424 127160 46044 127236
rect 45424 127094 45636 127160
rect 45424 127030 45430 127094
rect 45494 127030 45636 127094
rect 45424 127024 45636 127030
rect 45696 127094 46044 127160
rect 45696 127030 45974 127094
rect 46038 127030 46044 127094
rect 45696 127024 46044 127030
rect 46648 127100 46860 127236
rect 47056 127160 48492 127236
rect 47056 127100 47268 127160
rect 46648 127094 47268 127100
rect 46648 127030 46654 127094
rect 46718 127030 46790 127094
rect 46854 127030 47268 127094
rect 46648 127024 47268 127030
rect 47872 127024 48084 127160
rect 48280 127094 48492 127160
rect 48280 127030 48422 127094
rect 48486 127030 48492 127094
rect 48280 127024 48492 127030
rect 49096 127100 49308 127236
rect 49504 127100 49716 127236
rect 49096 127094 49716 127100
rect 49096 127030 49102 127094
rect 49166 127030 49716 127094
rect 49096 127024 49716 127030
rect 50320 127230 50940 127236
rect 50320 127166 50734 127230
rect 50798 127166 50940 127230
rect 50320 127160 50940 127166
rect 50320 127094 50668 127160
rect 50320 127030 50326 127094
rect 50390 127030 50668 127094
rect 50320 127024 50668 127030
rect 50728 127094 50940 127160
rect 50728 127030 50870 127094
rect 50934 127030 50940 127094
rect 50728 127024 50940 127030
rect 51680 127160 52300 127236
rect 51680 127024 51892 127160
rect 51952 127100 52300 127160
rect 52904 127100 53116 127236
rect 53312 127100 53524 127236
rect 51952 127094 52844 127100
rect 51952 127030 52230 127094
rect 52294 127030 52774 127094
rect 52838 127030 52844 127094
rect 51952 127024 52844 127030
rect 52904 127094 53524 127100
rect 52904 127030 53318 127094
rect 53382 127030 53524 127094
rect 52904 127024 53524 127030
rect 54128 127230 54748 127236
rect 54128 127166 54678 127230
rect 54742 127166 54748 127230
rect 54128 127160 54748 127166
rect 54128 127094 54340 127160
rect 54128 127030 54134 127094
rect 54198 127030 54340 127094
rect 54128 127024 54340 127030
rect 54536 127094 54748 127160
rect 54536 127030 54678 127094
rect 54742 127030 54748 127094
rect 54536 127024 54748 127030
rect 55352 127100 55564 127236
rect 55760 127160 57196 127236
rect 55760 127100 55972 127160
rect 55352 127094 55972 127100
rect 55352 127030 55358 127094
rect 55422 127030 55902 127094
rect 55966 127030 55972 127094
rect 55352 127024 55972 127030
rect 56576 127024 56788 127160
rect 56984 127094 57196 127160
rect 56984 127030 57126 127094
rect 57190 127030 57196 127094
rect 56984 127024 57196 127030
rect 57800 127100 58148 127236
rect 58208 127100 58420 127236
rect 57800 127094 58420 127100
rect 57800 127030 57806 127094
rect 57870 127030 58420 127094
rect 57800 127024 58420 127030
rect 59160 127100 59372 127236
rect 59432 127100 59780 127236
rect 59160 127094 59780 127100
rect 59160 127030 59574 127094
rect 59638 127030 59780 127094
rect 59160 127024 59780 127030
rect 60384 127230 61004 127236
rect 60384 127166 60798 127230
rect 60862 127166 61004 127230
rect 60384 127160 61004 127166
rect 60384 127024 60596 127160
rect 60792 127100 61004 127160
rect 61608 127100 61820 127236
rect 62016 127100 62228 127236
rect 60792 127094 61548 127100
rect 60792 127030 60934 127094
rect 60998 127030 61478 127094
rect 61542 127030 61548 127094
rect 60792 127024 61548 127030
rect 61608 127094 62228 127100
rect 61608 127030 61614 127094
rect 61678 127030 62158 127094
rect 62222 127030 62228 127094
rect 61608 127024 62228 127030
rect 62832 127160 63452 127236
rect 62832 127094 63044 127160
rect 62832 127030 62838 127094
rect 62902 127030 63044 127094
rect 62832 127024 63044 127030
rect 63240 127094 63452 127160
rect 63240 127030 63382 127094
rect 63446 127030 63452 127094
rect 63240 127024 63452 127030
rect 64056 127100 64268 127236
rect 64464 127230 64676 127236
rect 64464 127166 64606 127230
rect 64670 127166 64676 127230
rect 64464 127100 64676 127166
rect 64056 127094 64676 127100
rect 64056 127030 64062 127094
rect 64126 127030 64676 127094
rect 64056 127024 64676 127030
rect 65280 127160 65900 127236
rect 65280 127024 65628 127160
rect 65688 127094 65900 127160
rect 65688 127030 65694 127094
rect 65758 127030 65900 127094
rect 65688 127024 65900 127030
rect 66640 127160 67260 127236
rect 66640 127094 66852 127160
rect 66640 127030 66646 127094
rect 66710 127030 66852 127094
rect 66640 127024 66852 127030
rect 66912 127094 67260 127160
rect 67864 127100 68076 127236
rect 68272 127100 68484 127236
rect 67358 127094 68484 127100
rect 66912 127030 67190 127094
rect 67254 127030 67260 127094
rect 67320 127030 67326 127094
rect 67390 127030 68414 127094
rect 68478 127030 68484 127094
rect 66912 127024 67260 127030
rect 67358 127024 68484 127030
rect 69088 127230 69708 127236
rect 69088 127166 69230 127230
rect 69294 127166 69708 127230
rect 69088 127160 69708 127166
rect 69088 127094 69300 127160
rect 69088 127030 69094 127094
rect 69158 127030 69300 127094
rect 69088 127024 69300 127030
rect 69496 127094 69708 127160
rect 69496 127030 69638 127094
rect 69702 127030 69708 127094
rect 69496 127024 69708 127030
rect 70312 127100 70524 127236
rect 70720 127100 70932 127236
rect 70312 127094 70932 127100
rect 70312 127030 70318 127094
rect 70382 127030 70862 127094
rect 70926 127030 70932 127094
rect 70312 127024 70932 127030
rect 71536 127160 72156 127236
rect 71536 127024 71884 127160
rect 71944 127094 72156 127160
rect 71944 127030 71950 127094
rect 72014 127030 72156 127094
rect 71944 127024 72156 127030
rect 72896 127160 73516 127236
rect 72896 127094 73108 127160
rect 72896 127030 72902 127094
rect 72966 127030 73108 127094
rect 72896 127024 73108 127030
rect 73168 127024 73516 127160
rect 74120 127100 74332 127236
rect 74528 127230 74740 127236
rect 74528 127166 74670 127230
rect 74734 127166 74740 127230
rect 74528 127100 74740 127166
rect 75344 127160 75964 127236
rect 74120 127094 75284 127100
rect 74120 127030 74126 127094
rect 74190 127030 75214 127094
rect 75278 127030 75284 127094
rect 74120 127024 75284 127030
rect 75344 127094 75556 127160
rect 75344 127030 75350 127094
rect 75414 127030 75556 127094
rect 75344 127024 75556 127030
rect 75752 127094 75964 127160
rect 75752 127030 75894 127094
rect 75958 127030 75964 127094
rect 75752 127024 75964 127030
rect 76568 127100 76780 127236
rect 76976 127100 77188 127236
rect 76568 127094 77188 127100
rect 76568 127030 76574 127094
rect 76638 127030 77118 127094
rect 77182 127030 77188 127094
rect 76568 127024 77188 127030
rect 77792 127160 78412 127236
rect 77792 127094 78004 127160
rect 77792 127030 77798 127094
rect 77862 127030 78004 127094
rect 77792 127024 78004 127030
rect 78200 127094 78412 127160
rect 78200 127030 78342 127094
rect 78406 127030 78412 127094
rect 78200 127024 78412 127030
rect 79016 127230 79636 127236
rect 79016 127166 79294 127230
rect 79358 127166 79636 127230
rect 79016 127160 79636 127166
rect 79016 127024 79364 127160
rect 79424 127094 79636 127160
rect 79424 127030 79566 127094
rect 79630 127030 79636 127094
rect 79424 127024 79636 127030
rect 80376 127100 80588 127236
rect 80648 127100 80996 127236
rect 81600 127160 82220 127236
rect 80376 127094 81540 127100
rect 80376 127030 80926 127094
rect 80990 127030 81470 127094
rect 81534 127030 81540 127094
rect 80376 127024 81540 127030
rect 81600 127094 81812 127160
rect 81600 127030 81606 127094
rect 81670 127030 81812 127094
rect 81600 127024 81812 127030
rect 82008 127094 82220 127160
rect 82008 127030 82014 127094
rect 82078 127030 82220 127094
rect 82008 127024 82220 127030
rect 82824 127100 83036 127236
rect 83232 127100 83444 127236
rect 82824 127094 83444 127100
rect 82824 127030 82830 127094
rect 82894 127030 83444 127094
rect 82824 127024 83444 127030
rect 84048 127230 84668 127236
rect 84048 127166 84190 127230
rect 84254 127166 84668 127230
rect 84048 127160 84668 127166
rect 84048 127094 84260 127160
rect 84048 127030 84054 127094
rect 84118 127030 84260 127094
rect 84048 127024 84260 127030
rect 84456 127094 84668 127160
rect 84456 127030 84598 127094
rect 84662 127030 84668 127094
rect 84456 127024 84668 127030
rect 85272 127100 85484 127236
rect 85680 127100 85892 127236
rect 85272 127094 85892 127100
rect 85272 127030 85278 127094
rect 85342 127030 85822 127094
rect 85886 127030 85892 127094
rect 85272 127024 85892 127030
rect 86496 127160 87116 127236
rect 86496 127094 86844 127160
rect 86496 127030 86502 127094
rect 86566 127030 86844 127094
rect 86496 127024 86844 127030
rect 86904 127094 87116 127160
rect 86904 127030 87046 127094
rect 87110 127030 87116 127094
rect 86904 127024 87116 127030
rect 87856 127160 88476 127236
rect 87856 127024 88068 127160
rect 88128 127094 88476 127160
rect 88128 127030 88406 127094
rect 88470 127030 88476 127094
rect 88128 127024 88476 127030
rect 89080 127100 89292 127236
rect 89488 127230 89700 127236
rect 89488 127166 89630 127230
rect 89694 127166 89700 127230
rect 89488 127100 89700 127166
rect 89080 127094 89700 127100
rect 89080 127030 89222 127094
rect 89286 127030 89700 127094
rect 89080 127024 89700 127030
rect 90304 127160 90924 127236
rect 90304 127094 90516 127160
rect 90304 127030 90310 127094
rect 90374 127030 90516 127094
rect 90304 127024 90516 127030
rect 90712 127094 90924 127160
rect 90712 127030 90854 127094
rect 90918 127030 90924 127094
rect 90712 127024 90924 127030
rect 91528 127100 91740 127236
rect 91936 127100 92148 127236
rect 91528 127094 92148 127100
rect 91528 127030 91534 127094
rect 91598 127030 92148 127094
rect 91528 127024 92148 127030
rect 92752 127160 93372 127236
rect 92752 127094 93100 127160
rect 92752 127030 92758 127094
rect 92822 127030 93100 127094
rect 92752 127024 93100 127030
rect 93160 127094 93372 127160
rect 93160 127030 93302 127094
rect 93366 127030 93372 127094
rect 93160 127024 93372 127030
rect 94112 127230 94732 127236
rect 94112 127166 94662 127230
rect 94726 127166 94732 127230
rect 94112 127160 94732 127166
rect 94112 127024 94324 127160
rect 94384 127094 94732 127160
rect 94384 127030 94662 127094
rect 94726 127030 94732 127094
rect 94384 127024 94732 127030
rect 95336 127100 95548 127236
rect 95744 127100 95956 127236
rect 95336 127094 95956 127100
rect 95336 127030 95342 127094
rect 95406 127030 95750 127094
rect 95814 127030 95956 127094
rect 95336 127024 95956 127030
rect 96560 127160 97180 127236
rect 96560 127094 96772 127160
rect 96560 127030 96566 127094
rect 96630 127030 96772 127094
rect 96560 127024 96772 127030
rect 96968 127094 97180 127160
rect 96968 127030 97110 127094
rect 97174 127030 97180 127094
rect 96968 127024 97180 127030
rect 97784 127100 97996 127236
rect 98192 127100 98404 127236
rect 97784 127094 98404 127100
rect 97784 127030 97926 127094
rect 97990 127030 98404 127094
rect 97784 127024 98404 127030
rect 99008 127230 99628 127236
rect 99008 127166 99558 127230
rect 99622 127166 99628 127230
rect 99008 127160 99628 127166
rect 99008 127024 99220 127160
rect 99416 127094 99628 127160
rect 99416 127030 99558 127094
rect 99622 127030 99628 127094
rect 99416 127024 99628 127030
rect 100232 127100 100580 127236
rect 100640 127100 100852 127236
rect 100232 127094 100852 127100
rect 100232 127030 100238 127094
rect 100302 127030 100510 127094
rect 100574 127030 100852 127094
rect 100232 127024 100852 127030
rect 101592 127100 101804 127236
rect 101864 127100 102212 127236
rect 101592 127094 102212 127100
rect 101592 127030 102006 127094
rect 102070 127030 102212 127094
rect 101592 127024 102212 127030
rect 102816 127160 103436 127236
rect 102816 127024 103028 127160
rect 103224 127094 103436 127160
rect 103224 127030 103366 127094
rect 103430 127030 103436 127094
rect 103224 127024 103436 127030
rect 104040 127230 104388 127236
rect 104040 127166 104318 127230
rect 104382 127166 104388 127230
rect 104040 127160 104388 127166
rect 104040 127100 104252 127160
rect 104448 127100 104660 127236
rect 104040 127094 104660 127100
rect 104040 127030 104046 127094
rect 104110 127030 104590 127094
rect 104654 127030 104660 127094
rect 104040 127024 104660 127030
rect 105264 127160 105884 127236
rect 105264 127094 105476 127160
rect 105264 127030 105270 127094
rect 105334 127030 105476 127094
rect 105264 127024 105476 127030
rect 105672 127094 105884 127160
rect 105672 127030 105814 127094
rect 105878 127030 105884 127094
rect 105672 127024 105884 127030
rect 106488 127100 106700 127236
rect 106896 127100 107108 127236
rect 106488 127094 107108 127100
rect 106488 127030 106494 127094
rect 106558 127030 107108 127094
rect 106488 127024 107108 127030
rect 107712 127160 108332 127236
rect 107712 127024 108060 127160
rect 108120 127094 108332 127160
rect 108120 127030 108126 127094
rect 108190 127030 108332 127094
rect 108120 127024 108332 127030
rect 109072 127230 109692 127236
rect 109072 127166 109622 127230
rect 109686 127166 109692 127230
rect 109072 127160 109692 127166
rect 109072 127094 109284 127160
rect 109072 127030 109214 127094
rect 109278 127030 109284 127094
rect 109072 127024 109284 127030
rect 109344 127024 109692 127160
rect 110296 127100 110508 127236
rect 110704 127100 110916 127236
rect 110296 127094 110916 127100
rect 110296 127030 110302 127094
rect 110366 127030 110846 127094
rect 110910 127030 110916 127094
rect 110296 127024 110916 127030
rect 111520 127160 112140 127236
rect 111520 127094 111732 127160
rect 111520 127030 111526 127094
rect 111590 127030 111732 127094
rect 111520 127024 111732 127030
rect 111928 127094 112140 127160
rect 111928 127030 112070 127094
rect 112134 127030 112140 127094
rect 111928 127024 112140 127030
rect 112744 127100 112956 127236
rect 113152 127100 113364 127236
rect 112744 127094 113364 127100
rect 112744 127030 112750 127094
rect 112814 127030 113294 127094
rect 113358 127030 113364 127094
rect 112744 127024 113364 127030
rect 113968 127230 114588 127236
rect 113968 127166 114246 127230
rect 114310 127166 114588 127230
rect 113968 127160 114588 127166
rect 113968 127024 114316 127160
rect 114376 127094 114588 127160
rect 114376 127030 114518 127094
rect 114582 127030 114588 127094
rect 114376 127024 114588 127030
rect 115328 127160 115948 127236
rect 115328 127024 115540 127160
rect 115600 127094 115948 127160
rect 115600 127030 115742 127094
rect 115806 127030 115948 127094
rect 115600 127024 115948 127030
rect 116552 127100 116764 127236
rect 116960 127100 117172 127236
rect 117776 127160 118396 127236
rect 116552 127094 117716 127100
rect 116552 127030 116558 127094
rect 116622 127030 117646 127094
rect 117710 127030 117716 127094
rect 116552 127024 117716 127030
rect 117776 127094 117988 127160
rect 117776 127030 117782 127094
rect 117846 127030 117988 127094
rect 117776 127024 117988 127030
rect 118184 127094 118396 127160
rect 118184 127030 118326 127094
rect 118390 127030 118396 127094
rect 118184 127024 118396 127030
rect 119000 127100 119212 127236
rect 119408 127100 119620 127236
rect 119000 127094 119620 127100
rect 119000 127030 119006 127094
rect 119070 127030 119550 127094
rect 119614 127030 119620 127094
rect 119000 127024 119620 127030
rect 120224 127230 120844 127236
rect 120224 127166 120230 127230
rect 120294 127166 120844 127230
rect 120224 127160 120844 127166
rect 120224 127024 120436 127160
rect 120632 127094 120844 127160
rect 120632 127030 120774 127094
rect 120838 127030 120844 127094
rect 120632 127024 120844 127030
rect 121448 127100 121796 127236
rect 121856 127100 122068 127236
rect 121448 127094 122068 127100
rect 121448 127030 121454 127094
rect 121518 127030 121998 127094
rect 122062 127030 122068 127094
rect 121448 127024 122068 127030
rect 122808 127100 123020 127236
rect 123080 127100 123428 127236
rect 124032 127230 124652 127236
rect 124032 127166 124582 127230
rect 124646 127166 124652 127230
rect 124032 127160 124652 127166
rect 124032 127100 124244 127160
rect 122808 127094 123972 127100
rect 122808 127030 122950 127094
rect 123014 127030 123902 127094
rect 123966 127030 123972 127094
rect 122808 127024 123972 127030
rect 124032 127094 124380 127100
rect 124032 127030 124310 127094
rect 124374 127030 124380 127094
rect 124032 127024 124380 127030
rect 124440 127024 124652 127160
rect 125256 127100 125468 127236
rect 125664 127100 125876 127236
rect 125256 127094 125876 127100
rect 125256 127030 125262 127094
rect 125326 127030 125806 127094
rect 125870 127030 125876 127094
rect 125256 127024 125876 127030
rect 126480 127160 127100 127236
rect 126480 127094 126692 127160
rect 126480 127030 126486 127094
rect 126550 127030 126692 127094
rect 126480 127024 126692 127030
rect 126888 127094 127100 127160
rect 126888 127030 127030 127094
rect 127094 127030 127100 127094
rect 126888 127024 127100 127030
rect 127704 127100 127916 127236
rect 128112 127100 128324 127236
rect 127704 127094 128324 127100
rect 127704 127030 128254 127094
rect 128318 127030 128324 127094
rect 127704 127024 128324 127030
rect 128928 127230 129276 127236
rect 128928 127166 129206 127230
rect 129270 127166 129276 127230
rect 128928 127100 129276 127166
rect 129336 127100 129548 127236
rect 128928 127094 129548 127100
rect 128928 127030 128934 127094
rect 128998 127030 129478 127094
rect 129542 127030 129548 127094
rect 128928 127024 129548 127030
rect 130288 127160 130908 127236
rect 130288 127094 130500 127160
rect 130288 127030 130294 127094
rect 130358 127030 130500 127094
rect 130288 127024 130500 127030
rect 130560 127094 130908 127160
rect 130560 127030 130838 127094
rect 130902 127030 130908 127094
rect 130560 127024 130908 127030
rect 131512 127100 131724 127236
rect 131920 127160 133356 127236
rect 131920 127100 132132 127160
rect 131512 127094 132132 127100
rect 131512 127030 132062 127094
rect 132126 127030 132132 127094
rect 131512 127024 132132 127030
rect 132736 127024 132948 127160
rect 133144 127094 133356 127160
rect 133144 127030 133286 127094
rect 133350 127030 133356 127094
rect 133144 127024 133356 127030
rect 133960 127100 134172 127236
rect 134368 127100 134580 127236
rect 133960 127094 134580 127100
rect 133960 127030 133966 127094
rect 134030 127030 134510 127094
rect 134574 127030 134580 127094
rect 133960 127024 134580 127030
rect 135184 127230 135804 127236
rect 135184 127166 135598 127230
rect 135662 127166 135804 127230
rect 135184 127160 135804 127166
rect 135184 127094 135532 127160
rect 135184 127030 135190 127094
rect 135254 127030 135462 127094
rect 135526 127030 135532 127094
rect 135184 127024 135532 127030
rect 135592 127024 135804 127160
rect 136544 127160 137164 127236
rect 136544 127024 136756 127160
rect 136816 127094 137164 127160
rect 136816 127030 137094 127094
rect 137158 127030 137164 127094
rect 136816 127024 137164 127030
rect 137768 127100 137980 127236
rect 138176 127100 138388 127236
rect 137768 127094 138388 127100
rect 137768 127030 138182 127094
rect 138246 127030 138388 127094
rect 137768 127024 138388 127030
rect 138992 127230 139612 127236
rect 138992 127166 139542 127230
rect 139606 127166 139612 127230
rect 138992 127160 139612 127166
rect 138992 127024 139204 127160
rect 139400 127094 139612 127160
rect 139400 127030 139542 127094
rect 139606 127030 139612 127094
rect 139400 127024 139612 127030
rect 140216 127100 140428 127236
rect 140624 127100 140836 127236
rect 140216 127094 140836 127100
rect 140216 127030 140358 127094
rect 140422 127030 140836 127094
rect 140216 127024 140836 127030
rect 141440 127160 142060 127236
rect 141440 127094 141652 127160
rect 141440 127030 141446 127094
rect 141510 127030 141652 127094
rect 141440 127024 141652 127030
rect 141848 127094 142060 127160
rect 141848 127030 141990 127094
rect 142054 127030 142060 127094
rect 141848 127024 142060 127030
rect 142664 127160 143284 127236
rect 142664 127094 143012 127160
rect 142664 127030 142670 127094
rect 142734 127030 143012 127094
rect 142664 127024 143012 127030
rect 143072 127024 143284 127160
rect 144024 127100 144236 127236
rect 144296 127100 144644 127236
rect 144024 127094 144644 127100
rect 144024 127030 144438 127094
rect 144502 127030 144644 127094
rect 144024 127024 144644 127030
rect 145248 127230 145868 127236
rect 145248 127166 145254 127230
rect 145318 127166 145868 127230
rect 145248 127160 145868 127166
rect 145248 127094 145460 127160
rect 145248 127030 145254 127094
rect 145318 127030 145460 127094
rect 145248 127024 145460 127030
rect 145656 127024 145868 127160
rect 146472 127100 146684 127236
rect 146880 127100 147092 127236
rect 146472 127094 147092 127100
rect 146472 127030 146478 127094
rect 146542 127030 147022 127094
rect 147086 127030 147092 127094
rect 146472 127024 147092 127030
rect 147696 127160 148316 127236
rect 147696 127094 147908 127160
rect 147696 127030 147702 127094
rect 147766 127030 147908 127094
rect 147696 127024 147908 127030
rect 148104 127094 148316 127160
rect 148104 127030 148246 127094
rect 148310 127030 148316 127094
rect 148104 127024 148316 127030
rect 148920 127100 149132 127236
rect 149328 127230 149540 127236
rect 149328 127166 149470 127230
rect 149534 127166 149540 127230
rect 149328 127100 149540 127166
rect 148920 127024 149540 127100
rect 150144 127100 150492 127236
rect 150552 127100 150764 127236
rect 150144 127094 150764 127100
rect 150144 127030 150150 127094
rect 150214 127030 150764 127094
rect 150144 127024 150764 127030
rect 151504 127160 152124 127236
rect 151504 127094 151716 127160
rect 151504 127030 151510 127094
rect 151574 127030 151716 127094
rect 151504 127024 151716 127030
rect 151776 127094 152124 127160
rect 151776 127030 151918 127094
rect 151982 127030 152124 127094
rect 151776 127024 152124 127030
rect 152728 127100 152940 127236
rect 153136 127100 153348 127236
rect 152728 127094 153348 127100
rect 152728 127030 153278 127094
rect 153342 127030 153348 127094
rect 152728 127024 153348 127030
rect 153952 127230 154572 127236
rect 153952 127166 154094 127230
rect 154158 127166 154572 127230
rect 153952 127160 154572 127166
rect 153952 127094 154164 127160
rect 153952 127030 153958 127094
rect 154022 127030 154164 127094
rect 153952 127024 154164 127030
rect 154360 127094 154572 127160
rect 154360 127030 154502 127094
rect 154566 127030 154572 127094
rect 154360 127024 154572 127030
rect 155176 127100 155388 127236
rect 155584 127100 155796 127236
rect 155176 127094 155796 127100
rect 155176 127030 155182 127094
rect 155246 127030 155726 127094
rect 155790 127030 155796 127094
rect 155176 127024 155796 127030
rect 156400 127100 156748 127236
rect 156808 127100 157020 127236
rect 156400 127094 157020 127100
rect 156400 127030 156678 127094
rect 156742 127030 157020 127094
rect 156400 127024 157020 127030
rect 157760 127160 158380 127236
rect 157760 127094 157972 127160
rect 157760 127030 157902 127094
rect 157966 127030 157972 127094
rect 157760 127024 157972 127030
rect 158032 127024 158380 127160
rect 158984 127100 159196 127236
rect 159392 127100 159604 127236
rect 158984 127094 159604 127100
rect 158984 127030 158990 127094
rect 159054 127030 159604 127094
rect 158984 127024 159604 127030
rect 160208 127230 160828 127236
rect 160208 127166 160214 127230
rect 160278 127166 160828 127230
rect 160208 127160 160828 127166
rect 160208 127094 160420 127160
rect 160208 127030 160214 127094
rect 160278 127030 160420 127094
rect 160208 127024 160420 127030
rect 160616 127094 160828 127160
rect 160616 127030 160758 127094
rect 160822 127030 160828 127094
rect 160616 127024 160828 127030
rect 161432 127100 161644 127236
rect 161840 127100 162052 127236
rect 161432 127094 162052 127100
rect 161432 127030 161982 127094
rect 162046 127030 162052 127094
rect 161432 127024 162052 127030
rect 162656 127160 163276 127236
rect 162656 127024 162868 127160
rect 163064 127094 163276 127160
rect 163064 127030 163206 127094
rect 163270 127030 163276 127094
rect 163064 127024 163276 127030
rect 163880 127100 164228 127236
rect 164288 127100 164500 127236
rect 163880 127094 164500 127100
rect 163880 127030 163886 127094
rect 163950 127030 164430 127094
rect 164494 127030 164500 127094
rect 163880 127024 164500 127030
rect 165240 127100 165452 127236
rect 165512 127230 165860 127236
rect 165512 127166 165518 127230
rect 165582 127166 165860 127230
rect 165512 127100 165860 127166
rect 166464 127160 167084 127236
rect 165240 127094 166404 127100
rect 165240 127030 165382 127094
rect 165446 127030 166334 127094
rect 166398 127030 166404 127094
rect 165240 127024 166404 127030
rect 166464 127094 166676 127160
rect 166464 127030 166470 127094
rect 166534 127030 166676 127094
rect 166464 127024 166676 127030
rect 166872 127024 167084 127160
rect 167688 127100 167900 127236
rect 168096 127100 168308 127236
rect 167688 127094 168308 127100
rect 167688 127030 168238 127094
rect 168302 127030 168308 127094
rect 167688 127024 168308 127030
rect 168912 127160 169532 127236
rect 168912 127094 169124 127160
rect 168912 127030 168918 127094
rect 168982 127030 169124 127094
rect 168912 127024 169124 127030
rect 169320 127094 169532 127160
rect 169320 127030 169462 127094
rect 169526 127030 169532 127094
rect 169320 127024 169532 127030
rect 170136 127230 170348 127236
rect 170136 127166 170142 127230
rect 170206 127166 170348 127230
rect 170136 127100 170348 127166
rect 170544 127100 170756 127236
rect 170136 127094 170756 127100
rect 170136 127030 170686 127094
rect 170750 127030 170756 127094
rect 170136 127024 170756 127030
rect 171360 127160 171980 127236
rect 171360 127094 171708 127160
rect 171360 127030 171366 127094
rect 171430 127030 171708 127094
rect 171360 127024 171708 127030
rect 171768 127094 171980 127160
rect 171768 127030 171910 127094
rect 171974 127030 171980 127094
rect 171768 127024 171980 127030
rect 172720 127160 173340 127236
rect 172720 127024 172932 127160
rect 172992 127094 173340 127160
rect 172992 127030 173134 127094
rect 173198 127030 173340 127094
rect 172992 127024 173340 127030
rect 173944 127100 174156 127236
rect 174352 127230 174564 127236
rect 174352 127166 174494 127230
rect 174558 127166 174564 127230
rect 174352 127100 174564 127166
rect 173944 127094 174564 127100
rect 173944 127030 174494 127094
rect 174558 127030 174564 127094
rect 173944 127024 174564 127030
rect 175168 127160 175788 127236
rect 175168 127094 175380 127160
rect 175168 127030 175174 127094
rect 175238 127030 175380 127094
rect 175168 127024 175380 127030
rect 175576 127094 175788 127160
rect 175576 127030 175718 127094
rect 175782 127030 175788 127094
rect 175576 127024 175788 127030
rect 176392 127100 176604 127236
rect 176800 127100 177012 127236
rect 176392 127094 177012 127100
rect 176392 127030 176942 127094
rect 177006 127030 177012 127094
rect 176392 127024 177012 127030
rect 177616 127100 177964 127236
rect 178024 127100 178236 127236
rect 177616 127094 178236 127100
rect 177616 127030 178166 127094
rect 178230 127030 178236 127094
rect 177616 127024 178236 127030
rect 178976 127230 179596 127236
rect 178976 127166 179526 127230
rect 179590 127166 179596 127230
rect 178976 127160 179596 127166
rect 178976 127094 179188 127160
rect 178976 127030 178982 127094
rect 179046 127030 179188 127094
rect 178976 127024 179188 127030
rect 179248 127024 179596 127160
rect 180200 127100 180412 127236
rect 180608 127100 180820 127236
rect 180200 127094 180820 127100
rect 180200 127030 180206 127094
rect 180270 127030 180614 127094
rect 180678 127030 180820 127094
rect 180200 127024 180820 127030
rect 181424 127160 182044 127236
rect 181424 127094 181636 127160
rect 181424 127030 181430 127094
rect 181494 127030 181636 127094
rect 181424 127024 181636 127030
rect 181832 127094 182044 127160
rect 181832 127030 181974 127094
rect 182038 127030 182044 127094
rect 181832 127024 182044 127030
rect 182648 127100 182860 127236
rect 183056 127100 183268 127236
rect 182648 127094 183268 127100
rect 182648 127030 183198 127094
rect 183262 127030 183268 127094
rect 182648 127024 183268 127030
rect 183872 127094 184084 127236
rect 183872 127030 184014 127094
rect 184078 127030 184084 127094
rect 183872 127024 184084 127030
rect 184280 127230 184492 127236
rect 184280 127166 184422 127230
rect 184486 127166 184492 127230
rect 184280 127094 184492 127166
rect 185096 127100 185444 127236
rect 185504 127100 185716 127236
rect 184998 127094 185716 127100
rect 184280 127030 184286 127094
rect 184350 127030 184492 127094
rect 184960 127030 184966 127094
rect 185030 127030 185238 127094
rect 185302 127030 185374 127094
rect 185438 127030 185716 127094
rect 184280 127024 184492 127030
rect 184998 127024 185716 127030
rect 186456 127100 186668 127236
rect 186728 127100 187076 127236
rect 186456 127094 187076 127100
rect 186456 127030 187006 127094
rect 187070 127030 187076 127094
rect 186456 127024 187076 127030
rect 187680 127160 188300 127236
rect 187680 127024 187892 127160
rect 188088 127094 188300 127160
rect 188088 127030 188230 127094
rect 188294 127030 188300 127094
rect 188088 127024 188300 127030
rect 188904 127100 189116 127236
rect 189312 127100 189524 127236
rect 188904 127094 189524 127100
rect 188904 127030 188910 127094
rect 188974 127030 189454 127094
rect 189518 127030 189524 127094
rect 188904 127024 189524 127030
rect 149056 126964 149132 127024
rect 149056 126958 149540 126964
rect 149056 126894 149470 126958
rect 149534 126894 149540 126958
rect 149056 126888 149540 126894
rect 203456 126958 203668 126964
rect 203456 126894 203462 126958
rect 203526 126894 203668 126958
rect 203456 126752 203668 126894
rect 215016 126828 215228 126964
rect 215696 126958 218220 126964
rect 215696 126894 218150 126958
rect 218214 126894 218220 126958
rect 215696 126888 218220 126894
rect 215696 126828 215908 126888
rect 215016 126752 215908 126828
rect 1224 126550 1844 126556
rect 1224 126486 1230 126550
rect 1294 126532 1844 126550
rect 1294 126486 1702 126532
rect 1224 126480 1702 126486
rect 1632 126476 1702 126480
rect 1758 126476 1844 126532
rect 1632 126344 1844 126476
rect 28968 126420 29316 126692
rect 29648 126686 29860 126692
rect 29648 126622 29654 126686
rect 29718 126622 29860 126686
rect 29648 126420 29860 126622
rect 30328 126420 30540 126692
rect 30872 126686 31084 126692
rect 30872 126622 30878 126686
rect 30942 126622 31084 126686
rect 30872 126556 31084 126622
rect 31552 126686 32444 126692
rect 31552 126622 31694 126686
rect 31758 126622 32444 126686
rect 31552 126616 32444 126622
rect 31552 126556 31764 126616
rect 30872 126480 31764 126556
rect 30872 126420 31084 126480
rect 28016 126414 28908 126420
rect 28016 126350 28838 126414
rect 28902 126350 28908 126414
rect 28016 126344 28908 126350
rect 28968 126344 31084 126420
rect 31552 126344 31764 126480
rect 32096 126556 32444 126616
rect 32776 126686 32988 126692
rect 32776 126622 32918 126686
rect 32982 126622 32988 126686
rect 32776 126556 32988 126622
rect 32096 126480 32988 126556
rect 32096 126344 32444 126480
rect 32776 126344 32988 126480
rect 33456 126686 33668 126692
rect 33456 126622 33462 126686
rect 33526 126622 33668 126686
rect 33456 126420 33668 126622
rect 34000 126686 34212 126692
rect 34000 126622 34142 126686
rect 34206 126622 34212 126686
rect 34000 126420 34212 126622
rect 33456 126344 34212 126420
rect 34680 126686 34892 126692
rect 34680 126622 34686 126686
rect 34750 126622 34892 126686
rect 34680 126420 34892 126622
rect 35224 126420 35572 126692
rect 35904 126686 36796 126692
rect 35904 126622 35910 126686
rect 35974 126622 36590 126686
rect 36654 126622 36796 126686
rect 35904 126616 36796 126622
rect 35904 126420 36116 126616
rect 34680 126344 36116 126420
rect 36584 126344 36796 126616
rect 37128 126686 38020 126692
rect 38118 126686 38564 126692
rect 37128 126622 37134 126686
rect 37198 126622 38020 126686
rect 38080 126622 38086 126686
rect 38150 126622 38564 126686
rect 37128 126616 38020 126622
rect 38118 126616 38564 126622
rect 37128 126344 37340 126616
rect 37808 126420 38020 126616
rect 38352 126420 38564 126616
rect 39032 126420 39244 126692
rect 39478 126686 39924 126692
rect 39440 126622 39446 126686
rect 39510 126622 39924 126686
rect 39478 126616 39924 126622
rect 39576 126420 39924 126616
rect 40256 126686 41148 126692
rect 40256 126622 40398 126686
rect 40462 126622 41148 126686
rect 40256 126616 41148 126622
rect 40256 126420 40468 126616
rect 37808 126344 40468 126420
rect 40936 126556 41148 126616
rect 41480 126686 41692 126692
rect 41480 126622 41622 126686
rect 41686 126622 41692 126686
rect 41480 126556 41692 126622
rect 40936 126480 41692 126556
rect 40936 126344 41148 126480
rect 41480 126344 41692 126480
rect 42160 126686 42372 126692
rect 42160 126622 42166 126686
rect 42230 126622 42372 126686
rect 42160 126420 42372 126622
rect 42704 126686 43324 126692
rect 42704 126622 42982 126686
rect 43046 126622 43254 126686
rect 43318 126622 43324 126686
rect 42704 126616 43324 126622
rect 42704 126556 43052 126616
rect 43384 126556 43596 126692
rect 42704 126480 43596 126556
rect 42704 126420 43052 126480
rect 42160 126344 43052 126420
rect 43384 126420 43596 126480
rect 44064 126420 44276 126692
rect 44608 126686 45500 126692
rect 44608 126622 44614 126686
rect 44678 126622 45430 126686
rect 45494 126622 45500 126686
rect 44608 126616 45500 126622
rect 44608 126420 44820 126616
rect 43384 126344 44820 126420
rect 45288 126344 45500 126616
rect 45832 126686 46724 126692
rect 46822 126686 47948 126692
rect 45832 126622 45974 126686
rect 46038 126622 46654 126686
rect 46718 126622 46724 126686
rect 46784 126622 46790 126686
rect 46854 126622 47948 126686
rect 45832 126616 46724 126622
rect 46822 126616 47948 126622
rect 45832 126344 46180 126616
rect 46512 126344 46724 126616
rect 47192 126344 47404 126616
rect 47736 126344 47948 126616
rect 48416 126686 48628 126692
rect 48416 126622 48422 126686
rect 48486 126622 48628 126686
rect 48416 126420 48628 126622
rect 48960 126686 49852 126692
rect 48960 126622 49102 126686
rect 49166 126622 49852 126686
rect 48960 126616 49852 126622
rect 48960 126420 49172 126616
rect 48416 126344 49172 126420
rect 49640 126556 49852 126616
rect 50184 126686 50532 126692
rect 50184 126622 50326 126686
rect 50390 126622 50532 126686
rect 50184 126556 50532 126622
rect 49640 126480 50532 126556
rect 49640 126344 49852 126480
rect 50184 126344 50532 126480
rect 50864 126686 51076 126692
rect 50864 126622 50870 126686
rect 50934 126622 51076 126686
rect 50864 126420 51076 126622
rect 51544 126686 52300 126692
rect 51544 126622 52230 126686
rect 52294 126622 52300 126686
rect 51544 126616 52300 126622
rect 51544 126420 51756 126616
rect 50864 126344 51756 126420
rect 52088 126344 52300 126616
rect 52768 126686 52980 126692
rect 52768 126622 52774 126686
rect 52838 126622 52980 126686
rect 52768 126420 52980 126622
rect 53312 126686 54204 126692
rect 53312 126622 53318 126686
rect 53382 126622 54134 126686
rect 54198 126622 54204 126686
rect 53312 126616 54204 126622
rect 53312 126420 53660 126616
rect 52768 126344 53660 126420
rect 53992 126344 54204 126616
rect 54672 126686 55428 126692
rect 54672 126622 54678 126686
rect 54742 126622 55358 126686
rect 55422 126622 55428 126686
rect 54672 126616 55428 126622
rect 54672 126344 54884 126616
rect 55216 126344 55428 126616
rect 55896 126686 56788 126692
rect 55896 126622 55902 126686
rect 55966 126622 56788 126686
rect 55896 126616 56788 126622
rect 55896 126344 56108 126616
rect 56440 126344 56788 126616
rect 57120 126686 57332 126692
rect 57120 126622 57126 126686
rect 57190 126622 57332 126686
rect 57120 126420 57332 126622
rect 57800 126686 58556 126692
rect 57800 126622 57806 126686
rect 57870 126622 58556 126686
rect 57800 126616 58556 126622
rect 57800 126420 58012 126616
rect 57120 126344 58012 126420
rect 58344 126556 58556 126616
rect 59024 126686 59780 126692
rect 59024 126622 59574 126686
rect 59638 126622 59780 126686
rect 59024 126616 59780 126622
rect 59024 126556 59236 126616
rect 58344 126480 59236 126556
rect 58344 126344 58556 126480
rect 59024 126344 59236 126480
rect 59568 126420 59780 126616
rect 60248 126686 61140 126692
rect 60248 126622 60934 126686
rect 60998 126622 61140 126686
rect 60248 126616 61140 126622
rect 60248 126420 60460 126616
rect 59568 126344 60460 126420
rect 60792 126344 61140 126616
rect 61472 126686 61684 126692
rect 61472 126622 61478 126686
rect 61542 126622 61614 126686
rect 61678 126622 61684 126686
rect 61472 126344 61684 126622
rect 62152 126686 62908 126692
rect 62152 126622 62158 126686
rect 62222 126622 62838 126686
rect 62902 126622 62908 126686
rect 62152 126616 62908 126622
rect 62152 126344 62364 126616
rect 62696 126344 62908 126616
rect 63376 126686 64268 126692
rect 63376 126622 63382 126686
rect 63446 126622 64062 126686
rect 64126 126622 64268 126686
rect 63376 126616 64268 126622
rect 63376 126344 63588 126616
rect 63920 126556 64268 126616
rect 64600 126686 65764 126692
rect 64600 126622 65694 126686
rect 65758 126622 65764 126686
rect 64600 126616 65764 126622
rect 64600 126556 64812 126616
rect 63920 126480 64812 126556
rect 63920 126344 64268 126480
rect 64600 126344 64812 126480
rect 65280 126556 65492 126616
rect 65824 126556 66036 126692
rect 65280 126480 66036 126556
rect 65280 126344 65492 126480
rect 65824 126420 66036 126480
rect 66504 126686 66716 126692
rect 66504 126622 66646 126686
rect 66710 126622 66716 126686
rect 66504 126420 66716 126622
rect 65824 126344 66716 126420
rect 67048 126686 67940 126692
rect 67048 126622 67190 126686
rect 67254 126622 67326 126686
rect 67390 126622 67940 126686
rect 67048 126616 67940 126622
rect 67048 126344 67396 126616
rect 67728 126344 67940 126616
rect 68408 126686 68620 126692
rect 68408 126622 68414 126686
rect 68478 126622 68620 126686
rect 68408 126556 68620 126622
rect 68952 126686 69164 126692
rect 68952 126622 69094 126686
rect 69158 126622 69164 126686
rect 68952 126556 69164 126622
rect 68408 126480 69164 126556
rect 68408 126344 68620 126480
rect 68952 126344 69164 126480
rect 69632 126686 69844 126692
rect 69632 126622 69638 126686
rect 69702 126622 69844 126686
rect 69632 126556 69844 126622
rect 70176 126686 70388 126692
rect 70176 126622 70318 126686
rect 70382 126622 70388 126686
rect 70176 126556 70388 126622
rect 69632 126480 70388 126556
rect 69632 126344 69844 126480
rect 70176 126344 70388 126480
rect 70856 126686 72020 126692
rect 70856 126622 70862 126686
rect 70926 126622 71950 126686
rect 72014 126622 72020 126686
rect 70856 126616 72020 126622
rect 72080 126686 72972 126692
rect 72080 126622 72902 126686
rect 72966 126622 72972 126686
rect 72080 126616 72972 126622
rect 70856 126344 71068 126616
rect 71400 126420 71748 126616
rect 72080 126420 72292 126616
rect 71400 126344 72292 126420
rect 72760 126556 72972 126616
rect 73304 126686 74196 126692
rect 73304 126622 74126 126686
rect 74190 126622 74196 126686
rect 73304 126616 74196 126622
rect 73304 126556 73516 126616
rect 72760 126480 73516 126556
rect 72760 126344 72972 126480
rect 73304 126344 73516 126480
rect 73984 126556 74196 126616
rect 74528 126556 74876 126692
rect 73984 126480 74876 126556
rect 73984 126344 74196 126480
rect 74528 126344 74876 126480
rect 75208 126686 75420 126692
rect 75208 126622 75214 126686
rect 75278 126622 75350 126686
rect 75414 126622 75420 126686
rect 75208 126344 75420 126622
rect 75888 126686 76644 126692
rect 75888 126622 75894 126686
rect 75958 126622 76574 126686
rect 76638 126622 76644 126686
rect 75888 126616 76644 126622
rect 75888 126344 76100 126616
rect 76432 126344 76644 126616
rect 77112 126686 77324 126692
rect 77112 126622 77118 126686
rect 77182 126622 77324 126686
rect 77112 126556 77324 126622
rect 77656 126686 78004 126692
rect 77656 126622 77798 126686
rect 77862 126622 78004 126686
rect 77656 126556 78004 126622
rect 77112 126480 78004 126556
rect 77112 126344 77324 126480
rect 77656 126344 78004 126480
rect 78336 126686 78548 126692
rect 78336 126622 78342 126686
rect 78406 126622 78548 126686
rect 78336 126556 78548 126622
rect 79016 126686 80996 126692
rect 79016 126622 79566 126686
rect 79630 126622 80926 126686
rect 80990 126622 80996 126686
rect 79016 126616 80996 126622
rect 79016 126556 79228 126616
rect 78336 126480 79228 126556
rect 78336 126344 78548 126480
rect 79016 126344 79228 126480
rect 79560 126344 79772 126616
rect 80240 126344 80452 126616
rect 80784 126344 80996 126616
rect 81464 126686 81676 126692
rect 81464 126622 81470 126686
rect 81534 126622 81606 126686
rect 81670 126622 81676 126686
rect 81464 126344 81676 126622
rect 82008 126686 82900 126692
rect 82008 126622 82014 126686
rect 82078 126622 82830 126686
rect 82894 126622 82900 126686
rect 82008 126616 82900 126622
rect 82008 126344 82356 126616
rect 82688 126556 82900 126616
rect 83368 126686 84124 126692
rect 83368 126622 84054 126686
rect 84118 126622 84124 126686
rect 83368 126616 84124 126622
rect 83368 126556 83580 126616
rect 82688 126480 83580 126556
rect 82688 126344 82900 126480
rect 83368 126344 83580 126480
rect 83912 126344 84124 126616
rect 84592 126686 85484 126692
rect 84592 126622 84598 126686
rect 84662 126622 85278 126686
rect 85342 126622 85484 126686
rect 84592 126616 85484 126622
rect 84592 126344 84804 126616
rect 85136 126344 85484 126616
rect 85816 126686 86028 126692
rect 85816 126622 85822 126686
rect 85886 126622 86028 126686
rect 85816 126556 86028 126622
rect 86496 126686 86708 126692
rect 86496 126622 86502 126686
rect 86566 126622 86708 126686
rect 86496 126556 86708 126622
rect 85816 126480 86708 126556
rect 85816 126344 86028 126480
rect 86496 126344 86708 126480
rect 87040 126686 87252 126692
rect 87040 126622 87046 126686
rect 87110 126622 87252 126686
rect 87040 126556 87252 126622
rect 87720 126686 88612 126692
rect 87720 126622 88406 126686
rect 88470 126622 88612 126686
rect 87720 126616 88612 126622
rect 87720 126556 87932 126616
rect 87040 126480 87932 126556
rect 87040 126344 87252 126480
rect 87720 126344 87932 126480
rect 88264 126556 88612 126616
rect 88944 126686 90380 126692
rect 88944 126622 90310 126686
rect 90374 126622 90380 126686
rect 88944 126616 90380 126622
rect 88944 126556 89156 126616
rect 89624 126556 89836 126616
rect 88264 126480 89156 126556
rect 89254 126550 89836 126556
rect 89216 126486 89222 126550
rect 89286 126486 89836 126550
rect 89254 126480 89836 126486
rect 88264 126344 88612 126480
rect 88944 126344 89156 126480
rect 89624 126344 89836 126480
rect 90168 126344 90380 126616
rect 90848 126686 91604 126692
rect 90848 126622 90854 126686
rect 90918 126622 91534 126686
rect 91598 126622 91604 126686
rect 90848 126616 91604 126622
rect 90848 126344 91060 126616
rect 91392 126556 91604 126616
rect 92072 126686 92964 126692
rect 92072 126622 92758 126686
rect 92822 126622 92964 126686
rect 92072 126616 92964 126622
rect 92072 126556 92284 126616
rect 91392 126480 92284 126556
rect 91392 126344 91604 126480
rect 92072 126344 92284 126480
rect 92616 126344 92964 126616
rect 93296 126686 94732 126692
rect 93296 126622 93302 126686
rect 93366 126622 94662 126686
rect 94726 126622 94732 126686
rect 93296 126616 94732 126622
rect 93296 126344 93508 126616
rect 93976 126344 94188 126616
rect 94520 126556 94732 126616
rect 95200 126686 95412 126692
rect 95200 126622 95342 126686
rect 95406 126622 95412 126686
rect 95200 126556 95412 126622
rect 94520 126480 95412 126556
rect 94520 126344 94732 126480
rect 95200 126344 95412 126480
rect 95744 126686 96092 126692
rect 95744 126622 95750 126686
rect 95814 126622 96092 126686
rect 95744 126420 96092 126622
rect 96424 126686 96636 126692
rect 96424 126622 96566 126686
rect 96630 126622 96636 126686
rect 96424 126420 96636 126622
rect 95744 126344 96636 126420
rect 97104 126686 97316 126692
rect 97104 126622 97110 126686
rect 97174 126622 97316 126686
rect 97104 126556 97316 126622
rect 97648 126616 99220 126692
rect 97648 126556 97860 126616
rect 98328 126556 98540 126616
rect 97104 126480 97860 126556
rect 97958 126550 98540 126556
rect 97920 126486 97926 126550
rect 97990 126486 98540 126550
rect 97958 126480 98540 126486
rect 97104 126344 97316 126480
rect 97648 126344 97860 126480
rect 98328 126344 98540 126480
rect 98872 126420 99220 126616
rect 99552 126686 100444 126692
rect 100542 126686 101668 126692
rect 99552 126622 99558 126686
rect 99622 126622 100238 126686
rect 100302 126622 100444 126686
rect 100504 126622 100510 126686
rect 100574 126622 101668 126686
rect 99552 126616 100444 126622
rect 100542 126616 101668 126622
rect 99552 126420 99764 126616
rect 98872 126344 99764 126420
rect 100232 126344 100444 126616
rect 100776 126344 100988 126616
rect 101456 126556 101668 126616
rect 102000 126686 103572 126692
rect 102000 126622 102006 126686
rect 102070 126622 103366 126686
rect 103430 126622 103572 126686
rect 102000 126616 103572 126622
rect 102000 126556 102212 126616
rect 101456 126480 102212 126556
rect 101456 126344 101668 126480
rect 102000 126344 102212 126480
rect 102680 126344 102892 126616
rect 103224 126420 103572 126616
rect 103904 126686 104116 126692
rect 103904 126622 104046 126686
rect 104110 126622 104116 126686
rect 103904 126420 104116 126622
rect 103224 126344 104116 126420
rect 104584 126686 104796 126692
rect 104584 126622 104590 126686
rect 104654 126622 104796 126686
rect 104584 126420 104796 126622
rect 105128 126686 105340 126692
rect 105128 126622 105270 126686
rect 105334 126622 105340 126686
rect 105128 126420 105340 126622
rect 104584 126344 105340 126420
rect 105808 126686 106020 126692
rect 105808 126622 105814 126686
rect 105878 126622 106020 126686
rect 105808 126556 106020 126622
rect 106352 126686 108196 126692
rect 106352 126622 106494 126686
rect 106558 126622 108126 126686
rect 108190 126622 108196 126686
rect 106352 126616 108196 126622
rect 108256 126616 109148 126692
rect 109246 126686 109828 126692
rect 109208 126622 109214 126686
rect 109278 126622 109828 126686
rect 109246 126616 109828 126622
rect 106352 126556 106700 126616
rect 105808 126480 106700 126556
rect 105808 126344 106020 126480
rect 106352 126344 106700 126480
rect 107032 126344 107244 126616
rect 107712 126420 107924 126616
rect 108256 126420 108468 126616
rect 107712 126344 108468 126420
rect 108936 126420 109148 126616
rect 109480 126556 109828 126616
rect 110160 126686 110372 126692
rect 110160 126622 110302 126686
rect 110366 126622 110372 126686
rect 110160 126556 110372 126622
rect 109480 126480 110372 126556
rect 109480 126420 109828 126480
rect 108936 126344 109828 126420
rect 110160 126344 110372 126480
rect 110840 126686 111596 126692
rect 110840 126622 110846 126686
rect 110910 126622 111526 126686
rect 111590 126622 111596 126686
rect 110840 126616 111596 126622
rect 110840 126344 111052 126616
rect 111384 126344 111596 126616
rect 112064 126686 112276 126692
rect 112064 126622 112070 126686
rect 112134 126622 112276 126686
rect 112064 126420 112276 126622
rect 112608 126686 112820 126692
rect 112608 126622 112750 126686
rect 112814 126622 112820 126686
rect 112608 126420 112820 126622
rect 112064 126344 112820 126420
rect 113288 126686 113500 126692
rect 113288 126622 113294 126686
rect 113358 126622 113500 126686
rect 113288 126420 113500 126622
rect 113832 126556 114180 126692
rect 114512 126686 114724 126692
rect 114512 126622 114518 126686
rect 114582 126622 114724 126686
rect 114512 126556 114724 126622
rect 115192 126686 116628 126692
rect 115192 126622 115742 126686
rect 115806 126622 116558 126686
rect 116622 126622 116628 126686
rect 115192 126616 116628 126622
rect 115192 126556 115404 126616
rect 113832 126480 115404 126556
rect 113832 126420 114180 126480
rect 113288 126344 114180 126420
rect 114512 126344 114724 126480
rect 115192 126344 115404 126480
rect 115736 126344 115948 126616
rect 116416 126420 116628 126616
rect 116960 126420 117308 126692
rect 116416 126344 117308 126420
rect 117640 126686 117852 126692
rect 117640 126622 117646 126686
rect 117710 126622 117782 126686
rect 117846 126622 117852 126686
rect 117640 126344 117852 126622
rect 118320 126686 118532 126692
rect 118320 126622 118326 126686
rect 118390 126622 118532 126686
rect 118320 126556 118532 126622
rect 118864 126686 119076 126692
rect 118864 126622 119006 126686
rect 119070 126622 119076 126686
rect 118864 126556 119076 126622
rect 118320 126480 119076 126556
rect 118320 126344 118532 126480
rect 118864 126344 119076 126480
rect 119544 126686 120436 126692
rect 119544 126622 119550 126686
rect 119614 126622 120436 126686
rect 119544 126616 120436 126622
rect 119544 126344 119756 126616
rect 120088 126556 120436 126616
rect 120768 126686 120980 126692
rect 120768 126622 120774 126686
rect 120838 126622 120980 126686
rect 120768 126556 120980 126622
rect 120088 126480 120980 126556
rect 120088 126344 120436 126480
rect 120768 126420 120980 126480
rect 121448 126686 121660 126692
rect 121448 126622 121454 126686
rect 121518 126622 121660 126686
rect 121448 126420 121660 126622
rect 120768 126344 121660 126420
rect 121992 126686 122204 126692
rect 121992 126622 121998 126686
rect 122062 126622 122204 126686
rect 121992 126420 122204 126622
rect 122672 126556 122884 126692
rect 122982 126686 123428 126692
rect 122944 126622 122950 126686
rect 123014 126622 123428 126686
rect 122982 126616 123428 126622
rect 123216 126556 123428 126616
rect 122672 126480 123428 126556
rect 122672 126420 122884 126480
rect 121992 126344 122884 126420
rect 123216 126344 123428 126480
rect 123896 126686 124788 126692
rect 123896 126622 123902 126686
rect 123966 126622 124446 126686
rect 124510 126622 124788 126686
rect 123896 126616 124788 126622
rect 123896 126344 124108 126616
rect 124440 126556 124788 126616
rect 125120 126686 125332 126692
rect 125120 126622 125262 126686
rect 125326 126622 125332 126686
rect 125120 126556 125332 126622
rect 124440 126480 125332 126556
rect 124440 126344 124788 126480
rect 125120 126344 125332 126480
rect 125800 126686 126556 126692
rect 125800 126622 125806 126686
rect 125870 126622 126486 126686
rect 126550 126622 126556 126686
rect 125800 126616 126556 126622
rect 125800 126344 126012 126616
rect 126344 126344 126556 126616
rect 127024 126686 127236 126692
rect 127024 126622 127030 126686
rect 127094 126622 127236 126686
rect 127024 126556 127236 126622
rect 127568 126556 127916 126692
rect 127024 126480 127916 126556
rect 127024 126344 127236 126480
rect 127568 126420 127916 126480
rect 128248 126686 129140 126692
rect 128248 126622 128254 126686
rect 128318 126622 128934 126686
rect 128998 126622 129140 126686
rect 128248 126616 129140 126622
rect 128248 126420 128460 126616
rect 127568 126344 128460 126420
rect 128928 126344 129140 126616
rect 129472 126686 129684 126692
rect 129472 126622 129478 126686
rect 129542 126622 129684 126686
rect 129472 126420 129684 126622
rect 130152 126686 130364 126692
rect 130152 126622 130294 126686
rect 130358 126622 130364 126686
rect 130152 126420 130364 126622
rect 129472 126344 130364 126420
rect 130696 126686 131044 126692
rect 130696 126622 130838 126686
rect 130902 126622 131044 126686
rect 130696 126420 131044 126622
rect 131376 126556 131588 126692
rect 132056 126686 132268 126692
rect 132056 126622 132062 126686
rect 132126 126622 132268 126686
rect 132056 126556 132268 126622
rect 131376 126480 132268 126556
rect 131376 126420 131588 126480
rect 130696 126344 131588 126420
rect 132056 126420 132268 126480
rect 132600 126420 132812 126692
rect 132056 126344 132812 126420
rect 133280 126686 133492 126692
rect 133280 126622 133286 126686
rect 133350 126622 133492 126686
rect 133280 126556 133492 126622
rect 133824 126686 134036 126692
rect 133824 126622 133966 126686
rect 134030 126622 134036 126686
rect 133824 126556 134036 126622
rect 133280 126480 134036 126556
rect 133280 126344 133492 126480
rect 133824 126344 134036 126480
rect 134504 126686 134716 126692
rect 134504 126622 134510 126686
rect 134574 126622 134716 126686
rect 134504 126420 134716 126622
rect 135048 126686 135396 126692
rect 135494 126686 135940 126692
rect 135048 126622 135190 126686
rect 135254 126622 135396 126686
rect 135456 126622 135462 126686
rect 135526 126622 135940 126686
rect 135048 126420 135396 126622
rect 135494 126616 135940 126622
rect 134504 126344 135396 126420
rect 135728 126556 135940 126616
rect 136408 126556 136620 126692
rect 135728 126480 136620 126556
rect 135728 126344 135940 126480
rect 136408 126420 136620 126480
rect 136952 126686 137844 126692
rect 136952 126622 137094 126686
rect 137158 126622 137844 126686
rect 136952 126616 137844 126622
rect 136952 126420 137164 126616
rect 136408 126344 137164 126420
rect 137632 126556 137844 126616
rect 138176 126686 138524 126692
rect 138176 126622 138182 126686
rect 138246 126622 138524 126686
rect 138176 126556 138524 126622
rect 138856 126556 139068 126692
rect 137632 126480 139068 126556
rect 137632 126344 137844 126480
rect 138176 126344 138524 126480
rect 138856 126420 139068 126480
rect 139536 126686 139748 126692
rect 139536 126622 139542 126686
rect 139606 126622 139748 126686
rect 139536 126420 139748 126622
rect 140080 126556 140292 126692
rect 140390 126686 140972 126692
rect 140352 126622 140358 126686
rect 140422 126622 140972 126686
rect 140390 126616 140972 126622
rect 140760 126556 140972 126616
rect 140080 126480 140972 126556
rect 140080 126420 140292 126480
rect 138856 126344 140292 126420
rect 140760 126420 140972 126480
rect 141304 126686 141652 126692
rect 141304 126622 141446 126686
rect 141510 126622 141652 126686
rect 141304 126420 141652 126622
rect 140760 126344 141652 126420
rect 141984 126686 142196 126692
rect 141984 126622 141990 126686
rect 142054 126622 142196 126686
rect 141984 126556 142196 126622
rect 142664 126686 142876 126692
rect 142664 126622 142670 126686
rect 142734 126622 142876 126686
rect 142664 126556 142876 126622
rect 143208 126616 144100 126692
rect 143208 126556 143420 126616
rect 141984 126480 143420 126556
rect 141984 126344 142196 126480
rect 142664 126344 142876 126480
rect 143208 126344 143420 126480
rect 143888 126420 144100 126616
rect 144432 126686 144644 126692
rect 144432 126622 144438 126686
rect 144502 126622 144644 126686
rect 144432 126556 144644 126622
rect 145112 126686 145324 126692
rect 145112 126622 145254 126686
rect 145318 126622 145324 126686
rect 145112 126556 145324 126622
rect 144432 126480 145324 126556
rect 144432 126420 144644 126480
rect 143888 126344 144644 126420
rect 145112 126420 145324 126480
rect 145656 126420 146004 126692
rect 146336 126686 146548 126692
rect 146336 126622 146478 126686
rect 146542 126622 146548 126686
rect 146336 126420 146548 126622
rect 145112 126344 146548 126420
rect 147016 126686 147228 126692
rect 147016 126622 147022 126686
rect 147086 126622 147228 126686
rect 147016 126556 147228 126622
rect 147560 126686 147772 126692
rect 147560 126622 147702 126686
rect 147766 126622 147772 126686
rect 147560 126556 147772 126622
rect 147016 126480 147772 126556
rect 147016 126344 147228 126480
rect 147560 126344 147772 126480
rect 148240 126686 148452 126692
rect 148240 126622 148246 126686
rect 148310 126622 148452 126686
rect 148240 126420 148452 126622
rect 148784 126686 149676 126692
rect 148784 126622 149470 126686
rect 149534 126622 149676 126686
rect 148784 126616 149676 126622
rect 148784 126420 149132 126616
rect 148240 126344 149132 126420
rect 149464 126420 149676 126616
rect 150144 126686 150356 126692
rect 150144 126622 150150 126686
rect 150214 126622 150356 126686
rect 150144 126420 150356 126622
rect 150688 126556 150900 126692
rect 151368 126686 151580 126692
rect 151368 126622 151510 126686
rect 151574 126622 151580 126686
rect 151368 126556 151580 126622
rect 150688 126480 151580 126556
rect 150688 126420 150900 126480
rect 149464 126344 150900 126420
rect 151368 126344 151580 126480
rect 151912 126686 152260 126692
rect 151912 126622 151918 126686
rect 151982 126622 152260 126686
rect 151912 126420 152260 126622
rect 152592 126420 152804 126692
rect 153272 126686 154028 126692
rect 153272 126622 153278 126686
rect 153342 126622 153958 126686
rect 154022 126622 154028 126686
rect 153272 126616 154028 126622
rect 153272 126420 153484 126616
rect 151912 126344 153484 126420
rect 153816 126344 154028 126616
rect 154496 126686 154708 126692
rect 154496 126622 154502 126686
rect 154566 126622 154708 126686
rect 154496 126420 154708 126622
rect 155040 126686 155252 126692
rect 155040 126622 155182 126686
rect 155246 126622 155252 126686
rect 155040 126420 155252 126622
rect 154496 126344 155252 126420
rect 155720 126686 155932 126692
rect 155720 126622 155726 126686
rect 155790 126622 155932 126686
rect 155720 126556 155932 126622
rect 156264 126556 156612 126692
rect 156710 126686 157156 126692
rect 156672 126622 156678 126686
rect 156742 126622 157156 126686
rect 156710 126616 157156 126622
rect 155720 126480 156612 126556
rect 155720 126344 155932 126480
rect 156264 126420 156612 126480
rect 156944 126420 157156 126616
rect 157624 126616 158380 126692
rect 157624 126420 157836 126616
rect 158168 126556 158380 126616
rect 157934 126550 158380 126556
rect 157896 126486 157902 126550
rect 157966 126486 158380 126550
rect 157934 126480 158380 126486
rect 156264 126344 157836 126420
rect 158168 126420 158380 126480
rect 158848 126686 159060 126692
rect 158848 126622 158990 126686
rect 159054 126622 159060 126686
rect 158848 126420 159060 126622
rect 159392 126556 159740 126692
rect 160072 126686 160284 126692
rect 160072 126622 160214 126686
rect 160278 126622 160284 126686
rect 160072 126556 160284 126622
rect 159392 126480 160284 126556
rect 159392 126420 159740 126480
rect 158168 126344 159740 126420
rect 160072 126344 160284 126480
rect 160752 126686 160964 126692
rect 160752 126622 160758 126686
rect 160822 126622 160964 126686
rect 160752 126420 160964 126622
rect 161296 126420 161508 126692
rect 161976 126686 162868 126692
rect 161976 126622 161982 126686
rect 162046 126622 162868 126686
rect 161976 126616 162868 126622
rect 161976 126420 162188 126616
rect 160752 126344 162188 126420
rect 162520 126420 162868 126616
rect 163200 126686 163412 126692
rect 163200 126622 163206 126686
rect 163270 126622 163412 126686
rect 163200 126420 163412 126622
rect 163880 126686 164092 126692
rect 163880 126622 163886 126686
rect 163950 126622 164092 126686
rect 163880 126420 164092 126622
rect 162520 126344 164092 126420
rect 164424 126686 164636 126692
rect 164424 126622 164430 126686
rect 164494 126622 164636 126686
rect 164424 126556 164636 126622
rect 165104 126556 165316 126692
rect 165414 126686 165860 126692
rect 165376 126622 165382 126686
rect 165446 126622 165860 126686
rect 165414 126616 165860 126622
rect 164424 126480 165316 126556
rect 164424 126344 164636 126480
rect 165104 126420 165316 126480
rect 165648 126420 165860 126616
rect 165104 126344 165860 126420
rect 166328 126686 167220 126692
rect 166328 126622 166334 126686
rect 166398 126622 166470 126686
rect 166534 126622 167220 126686
rect 166328 126616 167220 126622
rect 166328 126344 166540 126616
rect 166872 126420 167220 126616
rect 167552 126420 167764 126692
rect 168232 126686 168444 126692
rect 168232 126622 168238 126686
rect 168302 126622 168444 126686
rect 168232 126556 168444 126622
rect 168776 126686 168988 126692
rect 168776 126622 168918 126686
rect 168982 126622 168988 126686
rect 168776 126556 168988 126622
rect 168232 126480 168988 126556
rect 168232 126420 168444 126480
rect 166872 126344 168444 126420
rect 168776 126344 168988 126480
rect 169456 126686 169668 126692
rect 169456 126622 169462 126686
rect 169526 126622 169668 126686
rect 169456 126420 169668 126622
rect 170000 126556 170348 126692
rect 170680 126686 171572 126692
rect 170680 126622 170686 126686
rect 170750 126622 171366 126686
rect 171430 126622 171572 126686
rect 170680 126616 171572 126622
rect 170680 126556 170892 126616
rect 170000 126480 170892 126556
rect 170000 126420 170348 126480
rect 169456 126344 170348 126420
rect 170680 126344 170892 126480
rect 171360 126344 171572 126616
rect 171904 126686 172116 126692
rect 171904 126622 171910 126686
rect 171974 126622 172116 126686
rect 171904 126420 172116 126622
rect 172584 126420 172796 126692
rect 173128 126686 173476 126692
rect 173128 126622 173134 126686
rect 173198 126622 173476 126686
rect 173128 126420 173476 126622
rect 173808 126420 174020 126692
rect 174488 126686 174700 126692
rect 174488 126622 174494 126686
rect 174558 126622 174700 126686
rect 174488 126556 174700 126622
rect 175032 126686 175244 126692
rect 175032 126622 175174 126686
rect 175238 126622 175244 126686
rect 175032 126556 175244 126622
rect 174488 126480 175244 126556
rect 174488 126420 174700 126480
rect 171904 126344 174700 126420
rect 175032 126344 175244 126480
rect 175712 126686 175924 126692
rect 175712 126622 175718 126686
rect 175782 126622 175924 126686
rect 175712 126420 175924 126622
rect 176256 126420 176468 126692
rect 176936 126686 177148 126692
rect 176936 126622 176942 126686
rect 177006 126622 177148 126686
rect 176936 126556 177148 126622
rect 177480 126556 177828 126692
rect 176936 126480 177828 126556
rect 176936 126420 177148 126480
rect 175712 126344 177148 126420
rect 177480 126420 177828 126480
rect 178160 126686 178372 126692
rect 178160 126622 178166 126686
rect 178230 126622 178372 126686
rect 178160 126420 178372 126622
rect 178840 126686 179052 126692
rect 178840 126622 178982 126686
rect 179046 126622 179052 126686
rect 178840 126556 179052 126622
rect 179384 126686 180276 126692
rect 179384 126622 180206 126686
rect 180270 126622 180276 126686
rect 179384 126616 180276 126622
rect 179384 126556 179596 126616
rect 178840 126480 179596 126556
rect 178840 126420 179052 126480
rect 177480 126344 179052 126420
rect 179384 126344 179596 126480
rect 180064 126344 180276 126616
rect 180608 126686 181500 126692
rect 180608 126622 180614 126686
rect 180678 126622 181430 126686
rect 181494 126622 181500 126686
rect 180608 126616 181500 126622
rect 180608 126344 180956 126616
rect 181288 126344 181500 126616
rect 181968 126686 182180 126692
rect 181968 126622 181974 126686
rect 182038 126622 182180 126686
rect 181968 126420 182180 126622
rect 182512 126420 182724 126692
rect 183192 126686 183404 126692
rect 183192 126622 183198 126686
rect 183262 126622 183404 126686
rect 183192 126556 183404 126622
rect 183736 126686 184356 126692
rect 183736 126622 184014 126686
rect 184078 126622 184286 126686
rect 184350 126622 184356 126686
rect 183736 126616 184356 126622
rect 184416 126686 185036 126692
rect 184416 126622 184966 126686
rect 185030 126622 185036 126686
rect 184416 126616 185036 126622
rect 185096 126686 185308 126692
rect 185406 126686 185852 126692
rect 185096 126622 185238 126686
rect 185302 126622 185308 126686
rect 185368 126622 185374 126686
rect 185438 126622 185852 126686
rect 183736 126556 184084 126616
rect 183192 126480 184084 126556
rect 183192 126420 183404 126480
rect 181968 126344 183404 126420
rect 183736 126420 184084 126480
rect 184416 126420 184628 126616
rect 183736 126344 184628 126420
rect 185096 126344 185308 126622
rect 185406 126616 185852 126622
rect 185640 126420 185852 126616
rect 186320 126420 186532 126692
rect 186864 126686 187076 126692
rect 186864 126622 187006 126686
rect 187070 126622 187076 126686
rect 186864 126420 187076 126622
rect 187544 126556 187756 126692
rect 188088 126686 188980 126692
rect 188088 126622 188230 126686
rect 188294 126622 188910 126686
rect 188974 126622 188980 126686
rect 188088 126616 188980 126622
rect 188088 126556 188436 126616
rect 187544 126480 188436 126556
rect 187544 126420 187756 126480
rect 185640 126344 187756 126420
rect 188088 126344 188436 126480
rect 188768 126344 188980 126616
rect 189448 126686 189660 126692
rect 189448 126622 189454 126686
rect 189518 126622 189660 126686
rect 189448 126556 189660 126622
rect 189448 126550 191564 126556
rect 189448 126486 191494 126550
rect 191558 126486 191564 126550
rect 189448 126480 191564 126486
rect 216784 126532 216996 126556
rect 189448 126344 189660 126480
rect 216784 126476 216908 126532
rect 216964 126476 216996 126532
rect 216784 126420 216996 126476
rect 190400 126414 190748 126420
rect 190400 126350 190406 126414
rect 190470 126350 190748 126414
rect 28016 126284 28228 126344
rect 28016 126278 28364 126284
rect 28016 126214 28294 126278
rect 28358 126214 28364 126278
rect 28016 126208 28364 126214
rect 190400 126278 190748 126350
rect 216784 126414 217540 126420
rect 216784 126350 217470 126414
rect 217534 126350 217540 126414
rect 216784 126344 217540 126350
rect 190400 126214 190406 126278
rect 190470 126214 190748 126278
rect 190400 126208 190748 126214
rect 191488 126278 194420 126284
rect 191488 126214 191494 126278
rect 191558 126214 194420 126278
rect 191488 126208 194420 126214
rect 191488 126072 191700 126208
rect 194208 126148 194420 126208
rect 195024 126278 196596 126284
rect 195024 126214 196526 126278
rect 196590 126214 196596 126278
rect 195024 126208 196596 126214
rect 194208 126142 194964 126148
rect 194208 126078 194894 126142
rect 194958 126078 194964 126142
rect 194208 126072 194964 126078
rect 195024 126142 195236 126208
rect 195024 126078 195166 126142
rect 195230 126078 195236 126142
rect 195024 126072 195236 126078
rect 28288 126006 28636 126012
rect 28288 125942 28294 126006
rect 28358 125942 28636 126006
rect 28288 125870 28636 125942
rect 28288 125806 28294 125870
rect 28358 125806 28636 125870
rect 21760 125598 21972 125740
rect 21760 125534 21902 125598
rect 21966 125534 21972 125598
rect 21760 125528 21972 125534
rect 22168 125598 22380 125740
rect 22576 125604 22788 125740
rect 22478 125598 22788 125604
rect 22168 125534 22310 125598
rect 22374 125534 22380 125598
rect 22440 125534 22446 125598
rect 22510 125534 22788 125598
rect 22168 125528 22380 125534
rect 22478 125528 22788 125534
rect 22984 125392 23196 125740
rect 23392 125392 23604 125740
rect 28288 125734 28636 125806
rect 28288 125670 28566 125734
rect 28630 125670 28636 125734
rect 28288 125664 28636 125670
rect 190128 126006 190476 126012
rect 190128 125942 190406 126006
rect 190470 125942 190476 126006
rect 190128 125936 190476 125942
rect 190128 125734 190340 125936
rect 194926 125734 195236 125740
rect 190128 125670 190134 125734
rect 190198 125670 190340 125734
rect 194888 125670 194894 125734
rect 194958 125670 195166 125734
rect 195230 125670 195236 125734
rect 190128 125664 190340 125670
rect 194926 125664 195236 125670
rect 28288 125462 28636 125468
rect 28288 125398 28294 125462
rect 28358 125398 28566 125462
rect 28630 125398 28636 125462
rect 22984 125332 23060 125392
rect 23392 125332 23468 125392
rect 21760 125326 21972 125332
rect 21760 125262 21902 125326
rect 21966 125262 21972 125326
rect 21760 125190 21972 125262
rect 21760 125126 21766 125190
rect 21830 125126 21972 125190
rect 21760 125120 21972 125126
rect 22168 125326 22516 125332
rect 22168 125262 22310 125326
rect 22374 125262 22446 125326
rect 22510 125262 22516 125326
rect 22168 125256 22516 125262
rect 22168 125060 22380 125256
rect 22576 125060 22788 125332
rect 22168 124984 22788 125060
rect 22984 124984 23196 125332
rect 23392 124984 23604 125332
rect 22168 124924 22244 124984
rect 22576 124924 22652 124984
rect 22984 124924 23060 124984
rect 23528 124924 23604 124984
rect 1224 124918 1844 124924
rect 1224 124854 1230 124918
rect 1294 124854 1844 124918
rect 1224 124852 1844 124854
rect 1224 124848 1702 124852
rect 1632 124796 1702 124848
rect 1758 124796 1844 124852
rect 1632 124712 1844 124796
rect 21760 124918 21972 124924
rect 21760 124854 21766 124918
rect 21830 124854 21972 124918
rect 21760 124782 21972 124854
rect 21760 124718 21766 124782
rect 21830 124718 21972 124782
rect 21760 124712 21972 124718
rect 22168 124712 22380 124924
rect 22576 124782 22788 124924
rect 22576 124718 22718 124782
rect 22782 124718 22788 124782
rect 22576 124712 22788 124718
rect 22984 124782 23196 124924
rect 22984 124718 22990 124782
rect 23054 124718 23196 124782
rect 22984 124712 23196 124718
rect 23392 124782 23604 124924
rect 23392 124718 23398 124782
rect 23462 124718 23604 124782
rect 23392 124712 23604 124718
rect 28288 125326 28636 125398
rect 28288 125262 28430 125326
rect 28494 125262 28636 125326
rect 28288 125054 28636 125262
rect 28288 124990 28430 125054
rect 28494 124990 28636 125054
rect 28288 124848 28636 124990
rect 190128 125326 190340 125468
rect 190128 125262 190134 125326
rect 190198 125262 190270 125326
rect 190334 125262 190340 125326
rect 190128 125054 190340 125262
rect 190128 124990 190270 125054
rect 190334 124990 190340 125054
rect 190128 124848 190340 124990
rect 28288 124788 28364 124848
rect 190264 124788 190340 124848
rect 21760 124510 21972 124516
rect 21760 124446 21766 124510
rect 21830 124446 21972 124510
rect 21760 124374 21972 124446
rect 21760 124310 21902 124374
rect 21966 124310 21972 124374
rect 21760 124304 21972 124310
rect 22168 124380 22380 124516
rect 22576 124510 22788 124516
rect 22576 124446 22718 124510
rect 22782 124446 22788 124510
rect 22168 124374 22516 124380
rect 22168 124310 22446 124374
rect 22510 124310 22516 124374
rect 22168 124304 22516 124310
rect 22576 124304 22788 124446
rect 22984 124510 23196 124516
rect 22984 124446 22990 124510
rect 23054 124446 23196 124510
rect 22984 124374 23196 124446
rect 22984 124310 23126 124374
rect 23190 124310 23196 124374
rect 22984 124304 23196 124310
rect 23392 124510 23604 124516
rect 23392 124446 23398 124510
rect 23462 124446 23604 124510
rect 23392 124374 23604 124446
rect 23392 124310 23398 124374
rect 23462 124310 23604 124374
rect 23392 124304 23604 124310
rect 28288 124304 28636 124788
rect 190128 124304 190340 124788
rect 195024 125392 195236 125664
rect 195432 125392 195644 125740
rect 195840 125604 196052 125740
rect 196248 125604 196460 125740
rect 195840 125528 196460 125604
rect 196656 125734 196868 125740
rect 196656 125670 196662 125734
rect 196726 125670 196868 125734
rect 196656 125598 196868 125670
rect 196656 125534 196798 125598
rect 196862 125534 196868 125598
rect 196656 125528 196868 125534
rect 195976 125468 196052 125528
rect 215016 125468 215228 125604
rect 215696 125468 215908 125604
rect 195976 125392 196324 125468
rect 215016 125462 216860 125468
rect 215016 125398 216790 125462
rect 216854 125398 216860 125462
rect 215016 125392 216860 125398
rect 195024 125332 195100 125392
rect 195432 125332 195508 125392
rect 196248 125332 196324 125392
rect 195024 124984 195236 125332
rect 195432 124984 195644 125332
rect 195840 125196 196052 125332
rect 196248 125196 196460 125332
rect 195840 125120 196460 125196
rect 196656 125326 196868 125332
rect 196656 125262 196798 125326
rect 196862 125262 196868 125326
rect 196656 125190 196868 125262
rect 196656 125126 196662 125190
rect 196726 125126 196868 125190
rect 196656 125120 196868 125126
rect 195840 124984 196052 125120
rect 196248 124984 196460 125120
rect 195024 124924 195100 124984
rect 195432 124924 195508 124984
rect 196248 124924 196324 124984
rect 195024 124782 195236 124924
rect 195024 124718 195166 124782
rect 195230 124718 195236 124782
rect 195024 124712 195236 124718
rect 195432 124782 195644 124924
rect 195432 124718 195438 124782
rect 195502 124718 195644 124782
rect 195432 124712 195644 124718
rect 195840 124782 196052 124924
rect 196248 124788 196460 124924
rect 196150 124782 196460 124788
rect 195840 124718 195982 124782
rect 196046 124718 196052 124782
rect 196112 124718 196118 124782
rect 196182 124718 196460 124782
rect 195840 124712 196052 124718
rect 196150 124712 196460 124718
rect 196656 124918 196868 124924
rect 196656 124854 196662 124918
rect 196726 124854 196868 124918
rect 196656 124782 196868 124854
rect 196656 124718 196662 124782
rect 196726 124718 196868 124782
rect 196656 124712 196868 124718
rect 216784 124918 216996 124924
rect 216784 124854 216790 124918
rect 216854 124854 216996 124918
rect 216784 124852 216996 124854
rect 216784 124796 216908 124852
rect 216964 124796 216996 124852
rect 216784 124788 216996 124796
rect 216784 124782 217540 124788
rect 216784 124718 217470 124782
rect 217534 124718 217540 124782
rect 216784 124712 217540 124718
rect 195976 124576 196324 124652
rect 195976 124516 196052 124576
rect 196248 124516 196324 124576
rect 195024 124510 195236 124516
rect 195024 124446 195166 124510
rect 195230 124446 195236 124510
rect 195024 124374 195236 124446
rect 195024 124310 195030 124374
rect 195094 124310 195236 124374
rect 195024 124304 195236 124310
rect 195432 124510 195644 124516
rect 195432 124446 195438 124510
rect 195502 124446 195644 124510
rect 195432 124374 195644 124446
rect 195432 124310 195574 124374
rect 195638 124310 195644 124374
rect 195432 124304 195644 124310
rect 195840 124510 196188 124516
rect 195840 124446 195982 124510
rect 196046 124446 196118 124510
rect 196182 124446 196188 124510
rect 195840 124440 196188 124446
rect 195840 124380 196052 124440
rect 195840 124374 196188 124380
rect 195840 124310 195982 124374
rect 196046 124310 196118 124374
rect 196182 124310 196188 124374
rect 195840 124304 196188 124310
rect 196248 124304 196460 124516
rect 196656 124510 196868 124516
rect 196656 124446 196662 124510
rect 196726 124446 196868 124510
rect 196656 124374 196868 124446
rect 196656 124310 196798 124374
rect 196862 124310 196868 124374
rect 196656 124304 196868 124310
rect 22576 124244 22652 124304
rect 28560 124244 28636 124304
rect 190264 124244 190340 124304
rect 22304 124168 22652 124244
rect 22304 124108 22380 124168
rect 21760 124102 21972 124108
rect 21760 124038 21902 124102
rect 21966 124038 21972 124102
rect 21760 123966 21972 124038
rect 21760 123902 21766 123966
rect 21830 123902 21972 123966
rect 21760 123896 21972 123902
rect 22168 123972 22380 124108
rect 22478 124102 22788 124108
rect 22440 124038 22446 124102
rect 22510 124038 22788 124102
rect 22478 124032 22788 124038
rect 22576 123972 22788 124032
rect 22168 123966 22788 123972
rect 22168 123902 22174 123966
rect 22238 123902 22582 123966
rect 22646 123902 22788 123966
rect 22168 123896 22788 123902
rect 22984 124102 23196 124108
rect 22984 124038 23126 124102
rect 23190 124038 23196 124102
rect 22984 123966 23196 124038
rect 22984 123902 22990 123966
rect 23054 123902 23196 123966
rect 22984 123896 23196 123902
rect 23392 124102 23604 124108
rect 23392 124038 23398 124102
rect 23462 124038 23604 124102
rect 23392 123966 23604 124038
rect 28288 124032 28636 124244
rect 28560 123972 28636 124032
rect 23392 123902 23534 123966
rect 23598 123902 23604 123966
rect 23392 123896 23604 123902
rect 28288 123760 28636 123972
rect 190128 124032 190340 124244
rect 195024 124102 195236 124108
rect 195024 124038 195030 124102
rect 195094 124038 195236 124102
rect 190128 123972 190204 124032
rect 190128 123760 190340 123972
rect 195024 123966 195236 124038
rect 195024 123902 195166 123966
rect 195230 123902 195236 123966
rect 195024 123896 195236 123902
rect 195432 124102 195644 124108
rect 195432 124038 195574 124102
rect 195638 124038 195644 124102
rect 195432 123966 195644 124038
rect 195432 123902 195438 123966
rect 195502 123902 195644 123966
rect 195432 123896 195644 123902
rect 195840 124102 196052 124108
rect 196150 124102 196460 124108
rect 195840 124038 195982 124102
rect 196046 124038 196052 124102
rect 196112 124038 196118 124102
rect 196182 124038 196460 124102
rect 195840 123896 196052 124038
rect 196150 124032 196460 124038
rect 196248 123966 196460 124032
rect 196248 123902 196254 123966
rect 196318 123902 196460 123966
rect 196248 123896 196460 123902
rect 196656 124102 196868 124108
rect 196656 124038 196798 124102
rect 196862 124038 196868 124102
rect 196656 123966 196868 124038
rect 196656 123902 196662 123966
rect 196726 123902 196868 123966
rect 196656 123896 196868 123902
rect 215016 123972 215228 124108
rect 215696 123972 215908 124108
rect 215016 123966 218220 123972
rect 215016 123902 218150 123966
rect 218214 123902 218220 123966
rect 215016 123896 218220 123902
rect 28424 123700 28500 123760
rect 190128 123700 190204 123760
rect 21760 123694 21972 123700
rect 21760 123630 21766 123694
rect 21830 123630 21972 123694
rect 21760 123558 21972 123630
rect 21760 123494 21766 123558
rect 21830 123494 21972 123558
rect 21760 123488 21972 123494
rect 22168 123694 22380 123700
rect 22168 123630 22174 123694
rect 22238 123630 22380 123694
rect 22168 123488 22380 123630
rect 22576 123694 22788 123700
rect 22576 123630 22582 123694
rect 22646 123630 22788 123694
rect 22576 123564 22788 123630
rect 22478 123558 22788 123564
rect 22440 123494 22446 123558
rect 22510 123494 22582 123558
rect 22646 123494 22788 123558
rect 22478 123488 22788 123494
rect 22984 123694 23196 123700
rect 22984 123630 22990 123694
rect 23054 123630 23196 123694
rect 22984 123558 23196 123630
rect 22984 123494 23126 123558
rect 23190 123494 23196 123558
rect 22984 123488 23196 123494
rect 23392 123694 23604 123700
rect 23392 123630 23534 123694
rect 23598 123630 23604 123694
rect 23392 123558 23604 123630
rect 23392 123494 23534 123558
rect 23598 123494 23604 123558
rect 23392 123488 23604 123494
rect 28288 123488 28636 123700
rect 190128 123488 190340 123700
rect 195024 123694 195236 123700
rect 195024 123630 195166 123694
rect 195230 123630 195236 123694
rect 195024 123558 195236 123630
rect 195024 123494 195166 123558
rect 195230 123494 195236 123558
rect 195024 123488 195236 123494
rect 195432 123694 195644 123700
rect 195432 123630 195438 123694
rect 195502 123630 195644 123694
rect 195432 123558 195644 123630
rect 195432 123494 195574 123558
rect 195638 123494 195644 123558
rect 195432 123488 195644 123494
rect 195840 123558 196052 123700
rect 196248 123694 196460 123700
rect 196248 123630 196254 123694
rect 196318 123630 196460 123694
rect 196248 123564 196460 123630
rect 196150 123558 196460 123564
rect 195840 123494 195982 123558
rect 196046 123494 196052 123558
rect 196112 123494 196118 123558
rect 196182 123494 196460 123558
rect 195840 123488 196052 123494
rect 196150 123488 196460 123494
rect 196656 123694 196868 123700
rect 196656 123630 196662 123694
rect 196726 123630 196868 123694
rect 196656 123558 196868 123630
rect 196656 123494 196798 123558
rect 196862 123494 196868 123558
rect 196656 123488 196868 123494
rect 28424 123428 28500 123488
rect 190264 123428 190340 123488
rect 1224 123286 1844 123292
rect 1224 123222 1230 123286
rect 1294 123222 1844 123286
rect 1224 123216 1844 123222
rect 1632 123172 1844 123216
rect 1632 123116 1702 123172
rect 1758 123116 1844 123172
rect 1632 123080 1844 123116
rect 21760 123286 21972 123292
rect 21760 123222 21766 123286
rect 21830 123222 21972 123286
rect 21760 123080 21972 123222
rect 22168 123286 22516 123292
rect 22168 123222 22446 123286
rect 22510 123222 22516 123286
rect 22168 123216 22516 123222
rect 22576 123286 22788 123292
rect 22576 123222 22582 123286
rect 22646 123222 22788 123286
rect 22168 123156 22380 123216
rect 22168 123150 22516 123156
rect 22168 123086 22310 123150
rect 22374 123086 22446 123150
rect 22510 123086 22516 123150
rect 22168 123080 22516 123086
rect 22576 123080 22788 123222
rect 22984 123286 23196 123292
rect 22984 123222 23126 123286
rect 23190 123222 23196 123286
rect 22984 123150 23196 123222
rect 22984 123086 22990 123150
rect 23054 123086 23196 123150
rect 22984 123080 23196 123086
rect 23392 123286 23604 123292
rect 23392 123222 23534 123286
rect 23598 123222 23604 123286
rect 23392 123150 23604 123222
rect 23392 123086 23398 123150
rect 23462 123086 23604 123150
rect 23392 123080 23604 123086
rect 28288 123216 28636 123428
rect 190128 123216 190340 123428
rect 28288 123156 28364 123216
rect 190264 123156 190340 123216
rect 21760 123020 21836 123080
rect 21760 122742 21972 123020
rect 28288 122944 28636 123156
rect 190128 122944 190340 123156
rect 195024 123286 195236 123292
rect 195024 123222 195166 123286
rect 195230 123222 195236 123286
rect 195024 123150 195236 123222
rect 195024 123086 195166 123150
rect 195230 123086 195236 123150
rect 195024 123080 195236 123086
rect 195432 123286 195644 123292
rect 195432 123222 195574 123286
rect 195638 123222 195644 123286
rect 195432 123150 195644 123222
rect 195432 123086 195438 123150
rect 195502 123086 195644 123150
rect 195432 123080 195644 123086
rect 195840 123286 196188 123292
rect 195840 123222 195982 123286
rect 196046 123222 196118 123286
rect 196182 123222 196188 123286
rect 195840 123216 196188 123222
rect 195840 123156 196052 123216
rect 196248 123156 196460 123292
rect 195840 123150 196460 123156
rect 195840 123086 196254 123150
rect 196318 123086 196460 123150
rect 195840 123080 196460 123086
rect 196656 123286 196868 123292
rect 196656 123222 196798 123286
rect 196862 123222 196868 123286
rect 196656 123080 196868 123222
rect 216784 123172 216996 123292
rect 216784 123150 216908 123172
rect 216784 123086 216790 123150
rect 216854 123116 216908 123150
rect 216964 123156 216996 123172
rect 216964 123150 217540 123156
rect 216964 123116 217470 123150
rect 216854 123086 217470 123116
rect 217534 123086 217540 123150
rect 216784 123080 217540 123086
rect 196656 123020 196732 123080
rect 28288 122884 28364 122944
rect 190128 122884 190204 122944
rect 21760 122678 21766 122742
rect 21830 122678 21972 122742
rect 21760 122672 21972 122678
rect 22168 122878 22380 122884
rect 22478 122878 22788 122884
rect 22168 122814 22310 122878
rect 22374 122814 22380 122878
rect 22440 122814 22446 122878
rect 22510 122814 22788 122878
rect 22168 122742 22380 122814
rect 22478 122808 22788 122814
rect 22168 122678 22310 122742
rect 22374 122678 22380 122742
rect 22168 122672 22380 122678
rect 22576 122742 22788 122808
rect 22576 122678 22582 122742
rect 22646 122678 22788 122742
rect 22576 122672 22788 122678
rect 22984 122878 23196 122884
rect 22984 122814 22990 122878
rect 23054 122814 23196 122878
rect 22984 122742 23196 122814
rect 22984 122678 22990 122742
rect 23054 122678 23196 122742
rect 22984 122672 23196 122678
rect 23392 122878 23604 122884
rect 23392 122814 23398 122878
rect 23462 122814 23604 122878
rect 23392 122742 23604 122814
rect 23392 122678 23534 122742
rect 23598 122678 23604 122742
rect 23392 122672 23604 122678
rect 28288 122672 28636 122884
rect 28560 122612 28636 122672
rect 21760 122470 21972 122476
rect 21760 122406 21766 122470
rect 21830 122406 21972 122470
rect 21760 122264 21972 122406
rect 22168 122470 22380 122476
rect 22168 122406 22310 122470
rect 22374 122406 22380 122470
rect 22168 122264 22380 122406
rect 22576 122470 22788 122476
rect 22576 122406 22582 122470
rect 22646 122406 22788 122470
rect 22576 122334 22788 122406
rect 22576 122270 22718 122334
rect 22782 122270 22788 122334
rect 22576 122264 22788 122270
rect 22984 122470 23196 122476
rect 22984 122406 22990 122470
rect 23054 122406 23196 122470
rect 22984 122334 23196 122406
rect 22984 122270 23126 122334
rect 23190 122270 23196 122334
rect 22984 122264 23196 122270
rect 23392 122470 23604 122476
rect 23392 122406 23534 122470
rect 23598 122406 23604 122470
rect 23392 122334 23604 122406
rect 23392 122270 23398 122334
rect 23462 122270 23604 122334
rect 23392 122264 23604 122270
rect 28288 122400 28636 122612
rect 190128 122672 190340 122884
rect 195024 122878 195236 122884
rect 195024 122814 195166 122878
rect 195230 122814 195236 122878
rect 195024 122742 195236 122814
rect 195024 122678 195166 122742
rect 195230 122678 195236 122742
rect 195024 122672 195236 122678
rect 195432 122878 195644 122884
rect 195432 122814 195438 122878
rect 195502 122814 195644 122878
rect 195432 122742 195644 122814
rect 195432 122678 195574 122742
rect 195638 122678 195644 122742
rect 195432 122672 195644 122678
rect 195840 122878 196460 122884
rect 195840 122814 196254 122878
rect 196318 122814 196460 122878
rect 195840 122808 196460 122814
rect 195840 122742 196052 122808
rect 195840 122678 195846 122742
rect 195910 122678 196052 122742
rect 195840 122672 196052 122678
rect 196248 122672 196460 122808
rect 196656 122742 196868 123020
rect 196656 122678 196662 122742
rect 196726 122678 196868 122742
rect 196656 122672 196868 122678
rect 215016 122742 216860 122748
rect 215016 122678 216790 122742
rect 216854 122678 216860 122742
rect 215016 122672 216860 122678
rect 190128 122612 190204 122672
rect 190128 122400 190340 122612
rect 215016 122536 215228 122672
rect 215696 122536 215908 122672
rect 28288 122340 28364 122400
rect 190264 122340 190340 122400
rect 21896 122204 21972 122264
rect 21760 122062 21972 122204
rect 28288 122128 28636 122340
rect 190128 122128 190340 122340
rect 195024 122470 195236 122476
rect 195024 122406 195166 122470
rect 195230 122406 195236 122470
rect 195024 122334 195236 122406
rect 195024 122270 195030 122334
rect 195094 122270 195236 122334
rect 195024 122264 195236 122270
rect 195432 122470 195644 122476
rect 195432 122406 195574 122470
rect 195638 122406 195644 122470
rect 195432 122334 195644 122406
rect 195432 122270 195438 122334
rect 195502 122270 195644 122334
rect 195432 122264 195644 122270
rect 195840 122470 196460 122476
rect 195840 122406 195846 122470
rect 195910 122406 196460 122470
rect 195840 122400 196460 122406
rect 195840 122264 196052 122400
rect 196248 122340 196460 122400
rect 196150 122334 196460 122340
rect 196112 122270 196118 122334
rect 196182 122270 196460 122334
rect 196150 122264 196460 122270
rect 196656 122470 196868 122476
rect 196656 122406 196662 122470
rect 196726 122406 196868 122470
rect 196656 122264 196868 122406
rect 195976 122204 196052 122264
rect 196792 122204 196868 122264
rect 195976 122128 196324 122204
rect 28424 122068 28500 122128
rect 190264 122068 190340 122128
rect 196248 122068 196324 122128
rect 21760 121998 21766 122062
rect 21830 121998 21972 122062
rect 21760 121992 21972 121998
rect 22168 122062 22516 122068
rect 22168 121998 22446 122062
rect 22510 121998 22516 122062
rect 22168 121992 22516 121998
rect 22576 122062 22788 122068
rect 22576 121998 22718 122062
rect 22782 121998 22788 122062
rect 22168 121932 22380 121992
rect 22576 121932 22788 121998
rect 22168 121856 22788 121932
rect 22984 122062 23196 122068
rect 22984 121998 23126 122062
rect 23190 121998 23196 122062
rect 22984 121856 23196 121998
rect 22304 121796 22380 121856
rect 23120 121796 23196 121856
rect 21760 121790 21972 121796
rect 21760 121726 21766 121790
rect 21830 121726 21972 121790
rect 21760 121654 21972 121726
rect 21760 121590 21766 121654
rect 21830 121590 21972 121654
rect 21760 121584 21972 121590
rect 22168 121654 22380 121796
rect 22478 121790 22788 121796
rect 22440 121726 22446 121790
rect 22510 121726 22788 121790
rect 22478 121720 22788 121726
rect 22168 121590 22174 121654
rect 22238 121590 22380 121654
rect 22168 121584 22380 121590
rect 22576 121584 22788 121720
rect 1632 121492 1844 121524
rect 1632 121436 1702 121492
rect 1758 121436 1844 121492
rect 1632 121388 1844 121436
rect 22984 121448 23196 121796
rect 23392 122062 23604 122068
rect 23392 121998 23398 122062
rect 23462 121998 23604 122062
rect 23392 121856 23604 121998
rect 23392 121796 23468 121856
rect 23392 121448 23604 121796
rect 28288 121790 28636 122068
rect 28288 121726 28294 121790
rect 28358 121726 28636 121790
rect 28288 121720 28636 121726
rect 190128 121790 190340 122068
rect 195024 122062 195236 122068
rect 195024 121998 195030 122062
rect 195094 121998 195236 122062
rect 195024 121856 195236 121998
rect 195160 121796 195236 121856
rect 190128 121726 190134 121790
rect 190198 121726 190340 121790
rect 190128 121720 190340 121726
rect 22984 121388 23060 121448
rect 23528 121388 23604 121448
rect 1224 121382 1844 121388
rect 1224 121318 1230 121382
rect 1294 121318 1844 121382
rect 1224 121312 1844 121318
rect 21760 121382 21972 121388
rect 21760 121318 21766 121382
rect 21830 121318 21972 121382
rect 21760 121246 21972 121318
rect 21760 121182 21902 121246
rect 21966 121182 21972 121246
rect 21760 121176 21972 121182
rect 22168 121382 22788 121388
rect 22168 121318 22174 121382
rect 22238 121318 22788 121382
rect 22168 121312 22788 121318
rect 22168 121040 22380 121312
rect 22688 121116 22788 121312
rect 22440 121040 22788 121116
rect 22984 121040 23196 121388
rect 22440 120980 22516 121040
rect 22712 120980 22788 121040
rect 23120 120980 23196 121040
rect 21760 120974 21972 120980
rect 21760 120910 21902 120974
rect 21966 120910 21972 120974
rect 21760 120838 21972 120910
rect 21760 120774 21766 120838
rect 21830 120774 21972 120838
rect 21760 120768 21972 120774
rect 22168 120904 22516 120980
rect 22168 120844 22380 120904
rect 22168 120838 22516 120844
rect 22168 120774 22446 120838
rect 22510 120774 22516 120838
rect 22168 120768 22516 120774
rect 22576 120768 22788 120980
rect 22984 120838 23196 120980
rect 22984 120774 23126 120838
rect 23190 120774 23196 120838
rect 22984 120768 23196 120774
rect 23392 121040 23604 121388
rect 28288 121518 28636 121524
rect 28288 121454 28294 121518
rect 28358 121454 28636 121518
rect 28288 121382 28636 121454
rect 28288 121318 28294 121382
rect 28358 121318 28636 121382
rect 28288 121110 28636 121318
rect 28288 121046 28294 121110
rect 28358 121046 28636 121110
rect 23392 120980 23468 121040
rect 23392 120838 23604 120980
rect 28288 120974 28636 121046
rect 28288 120910 28430 120974
rect 28494 120910 28636 120974
rect 28288 120904 28636 120910
rect 190128 121518 190340 121524
rect 190128 121454 190134 121518
rect 190198 121454 190340 121518
rect 190128 121382 190340 121454
rect 190128 121318 190270 121382
rect 190334 121318 190340 121382
rect 190128 121110 190340 121318
rect 190128 121046 190270 121110
rect 190334 121046 190340 121110
rect 190128 120974 190340 121046
rect 190128 120910 190270 120974
rect 190334 120910 190340 120974
rect 190128 120904 190340 120910
rect 195024 121448 195236 121796
rect 195432 122062 195644 122068
rect 195432 121998 195438 122062
rect 195502 121998 195644 122062
rect 195432 121856 195644 121998
rect 195840 122062 196188 122068
rect 195840 121998 196118 122062
rect 196182 121998 196188 122062
rect 195840 121992 196188 121998
rect 195840 121856 196052 121992
rect 195432 121796 195508 121856
rect 195976 121796 196052 121856
rect 195432 121448 195644 121796
rect 195840 121660 196052 121796
rect 196248 121856 196460 122068
rect 196656 122062 196868 122204
rect 196656 121998 196798 122062
rect 196862 121998 196868 122062
rect 196656 121992 196868 121998
rect 196248 121796 196324 121856
rect 195840 121654 196188 121660
rect 195840 121590 196118 121654
rect 196182 121590 196188 121654
rect 195840 121584 196188 121590
rect 196248 121584 196460 121796
rect 196656 121790 196868 121796
rect 196656 121726 196798 121790
rect 196862 121726 196868 121790
rect 196656 121654 196868 121726
rect 196656 121590 196662 121654
rect 196726 121590 196868 121654
rect 196656 121584 196868 121590
rect 216784 121518 217540 121524
rect 216784 121492 217470 121518
rect 195024 121388 195100 121448
rect 195432 121388 195508 121448
rect 216784 121436 216908 121492
rect 216964 121454 217470 121492
rect 217534 121454 217540 121518
rect 216964 121448 217540 121454
rect 216964 121436 216996 121448
rect 195024 121040 195236 121388
rect 195432 121040 195644 121388
rect 195024 120980 195100 121040
rect 195568 120980 195644 121040
rect 23392 120774 23398 120838
rect 23462 120774 23604 120838
rect 23392 120768 23604 120774
rect 21760 120566 21972 120572
rect 21760 120502 21766 120566
rect 21830 120502 21972 120566
rect 21760 120430 21972 120502
rect 21760 120366 21766 120430
rect 21830 120366 21972 120430
rect 21760 120360 21972 120366
rect 22168 120430 22380 120572
rect 22478 120566 22788 120572
rect 22440 120502 22446 120566
rect 22510 120502 22788 120566
rect 22478 120496 22788 120502
rect 22168 120366 22174 120430
rect 22238 120366 22380 120430
rect 22168 120360 22380 120366
rect 22576 120430 22788 120496
rect 22576 120366 22718 120430
rect 22782 120366 22788 120430
rect 22576 120360 22788 120366
rect 22984 120566 23196 120572
rect 22984 120502 23126 120566
rect 23190 120502 23196 120566
rect 22984 120430 23196 120502
rect 22984 120366 23126 120430
rect 23190 120366 23196 120430
rect 22984 120360 23196 120366
rect 23392 120566 23604 120572
rect 23392 120502 23398 120566
rect 23462 120502 23604 120566
rect 23392 120430 23604 120502
rect 23392 120366 23398 120430
rect 23462 120366 23604 120430
rect 23392 120360 23604 120366
rect 28288 120566 28636 120844
rect 28288 120502 28294 120566
rect 28358 120502 28430 120566
rect 28494 120502 28636 120566
rect 28288 120360 28636 120502
rect 28560 120300 28636 120360
rect 28288 120294 28636 120300
rect 28288 120230 28294 120294
rect 28358 120230 28636 120294
rect 21760 120158 21972 120164
rect 21760 120094 21766 120158
rect 21830 120094 21972 120158
rect 21760 120022 21972 120094
rect 21760 119958 21902 120022
rect 21966 119958 21972 120022
rect 21760 119952 21972 119958
rect 22168 120158 22380 120164
rect 22168 120094 22174 120158
rect 22238 120094 22380 120158
rect 22168 120028 22380 120094
rect 22576 120158 22788 120164
rect 22576 120094 22718 120158
rect 22782 120094 22788 120158
rect 22576 120028 22788 120094
rect 22168 120022 22788 120028
rect 22168 119958 22310 120022
rect 22374 119958 22788 120022
rect 22168 119952 22788 119958
rect 22984 120158 23196 120164
rect 22984 120094 23126 120158
rect 23190 120094 23196 120158
rect 22984 120022 23196 120094
rect 22984 119958 23126 120022
rect 23190 119958 23196 120022
rect 22984 119952 23196 119958
rect 23392 120158 23604 120164
rect 23392 120094 23398 120158
rect 23462 120094 23604 120158
rect 23392 120022 23604 120094
rect 28288 120088 28636 120230
rect 190128 120566 190340 120844
rect 195024 120838 195236 120980
rect 195024 120774 195166 120838
rect 195230 120774 195236 120838
rect 195024 120768 195236 120774
rect 195432 120838 195644 120980
rect 195432 120774 195438 120838
rect 195502 120774 195644 120838
rect 195432 120768 195644 120774
rect 195840 121252 196052 121388
rect 196150 121382 196460 121388
rect 196112 121318 196118 121382
rect 196182 121318 196460 121382
rect 196150 121312 196460 121318
rect 196248 121252 196460 121312
rect 195840 121176 196460 121252
rect 196656 121382 196868 121388
rect 196656 121318 196662 121382
rect 196726 121318 196868 121382
rect 196656 121246 196868 121318
rect 196656 121182 196798 121246
rect 196862 121182 196868 121246
rect 196656 121176 196868 121182
rect 215016 121312 215908 121388
rect 216784 121312 216996 121436
rect 195840 121116 196052 121176
rect 195840 121040 196188 121116
rect 196248 121040 196460 121176
rect 215016 121040 215228 121312
rect 215696 121116 215908 121312
rect 215696 121110 218220 121116
rect 215696 121046 218150 121110
rect 218214 121046 218220 121110
rect 215696 121040 218220 121046
rect 195840 120980 195916 121040
rect 196112 120980 196188 121040
rect 195840 120838 196052 120980
rect 196112 120904 196460 120980
rect 195840 120774 195846 120838
rect 195910 120774 196052 120838
rect 195840 120768 196052 120774
rect 196248 120768 196460 120904
rect 196656 120974 196868 120980
rect 196656 120910 196798 120974
rect 196862 120910 196868 120974
rect 196656 120838 196868 120910
rect 196656 120774 196662 120838
rect 196726 120774 196868 120838
rect 196656 120768 196868 120774
rect 190128 120502 190134 120566
rect 190198 120502 190270 120566
rect 190334 120502 190340 120566
rect 190128 120360 190340 120502
rect 195024 120566 195236 120572
rect 195024 120502 195166 120566
rect 195230 120502 195236 120566
rect 195024 120430 195236 120502
rect 195024 120366 195166 120430
rect 195230 120366 195236 120430
rect 195024 120360 195236 120366
rect 195432 120566 195644 120572
rect 195432 120502 195438 120566
rect 195502 120502 195644 120566
rect 195432 120430 195644 120502
rect 195432 120366 195574 120430
rect 195638 120366 195644 120430
rect 195432 120360 195644 120366
rect 195840 120566 196052 120572
rect 195840 120502 195846 120566
rect 195910 120502 196052 120566
rect 195840 120430 196052 120502
rect 195840 120366 195982 120430
rect 196046 120366 196052 120430
rect 195840 120360 196052 120366
rect 196248 120360 196460 120572
rect 196656 120566 196868 120572
rect 196656 120502 196662 120566
rect 196726 120502 196868 120566
rect 196656 120430 196868 120502
rect 196656 120366 196798 120430
rect 196862 120366 196868 120430
rect 196656 120360 196868 120366
rect 190128 120300 190204 120360
rect 196248 120300 196324 120360
rect 190128 120294 190340 120300
rect 190128 120230 190134 120294
rect 190198 120230 190340 120294
rect 190128 120088 190340 120230
rect 195976 120224 196324 120300
rect 195976 120164 196052 120224
rect 28424 120028 28500 120088
rect 190264 120028 190340 120088
rect 23392 119958 23398 120022
rect 23462 119958 23604 120022
rect 23392 119952 23604 119958
rect 22304 119892 22380 119952
rect 1632 119812 1844 119892
rect 22304 119816 22652 119892
rect 28288 119816 28636 120028
rect 190128 119816 190340 120028
rect 195024 120158 195236 120164
rect 195024 120094 195166 120158
rect 195230 120094 195236 120158
rect 195024 120022 195236 120094
rect 195024 119958 195030 120022
rect 195094 119958 195236 120022
rect 195024 119952 195236 119958
rect 195432 120158 195644 120164
rect 195432 120094 195574 120158
rect 195638 120094 195644 120158
rect 195432 120022 195644 120094
rect 195432 119958 195574 120022
rect 195638 119958 195644 120022
rect 195432 119952 195644 119958
rect 195840 120158 196460 120164
rect 195840 120094 195982 120158
rect 196046 120094 196460 120158
rect 195840 120088 196460 120094
rect 195840 120022 196052 120088
rect 195840 119958 195982 120022
rect 196046 119958 196052 120022
rect 195840 119952 196052 119958
rect 196248 119952 196460 120088
rect 196656 120158 196868 120164
rect 196656 120094 196798 120158
rect 196862 120094 196868 120158
rect 196656 120022 196868 120094
rect 196656 119958 196798 120022
rect 196862 119958 196868 120022
rect 196656 119952 196868 119958
rect 1632 119756 1702 119812
rect 1758 119756 1844 119812
rect 22576 119756 22652 119816
rect 28560 119756 28636 119816
rect 190264 119756 190340 119816
rect 215016 119756 215228 119892
rect 215696 119886 217540 119892
rect 215696 119822 217470 119886
rect 217534 119822 217540 119886
rect 215696 119816 217540 119822
rect 215696 119756 215908 119816
rect 1224 119750 1844 119756
rect 1224 119686 1230 119750
rect 1294 119686 1844 119750
rect 1224 119680 1844 119686
rect 21760 119750 21972 119756
rect 21760 119686 21902 119750
rect 21966 119686 21972 119750
rect 21760 119614 21972 119686
rect 21760 119550 21766 119614
rect 21830 119550 21972 119614
rect 21760 119544 21972 119550
rect 22168 119750 22380 119756
rect 22168 119686 22310 119750
rect 22374 119686 22380 119750
rect 22168 119620 22380 119686
rect 22168 119614 22516 119620
rect 22168 119550 22446 119614
rect 22510 119550 22516 119614
rect 22168 119544 22516 119550
rect 22576 119544 22788 119756
rect 22984 119750 23196 119756
rect 22984 119686 23126 119750
rect 23190 119686 23196 119750
rect 22984 119614 23196 119686
rect 22984 119550 23126 119614
rect 23190 119550 23196 119614
rect 22984 119544 23196 119550
rect 23392 119750 23604 119756
rect 23392 119686 23398 119750
rect 23462 119686 23604 119750
rect 23392 119614 23604 119686
rect 23392 119550 23534 119614
rect 23598 119550 23604 119614
rect 23392 119544 23604 119550
rect 28288 119544 28636 119756
rect 190128 119544 190340 119756
rect 195024 119750 195236 119756
rect 195024 119686 195030 119750
rect 195094 119686 195236 119750
rect 195024 119614 195236 119686
rect 195024 119550 195166 119614
rect 195230 119550 195236 119614
rect 195024 119544 195236 119550
rect 195432 119750 195644 119756
rect 195432 119686 195574 119750
rect 195638 119686 195644 119750
rect 195432 119614 195644 119686
rect 195432 119550 195438 119614
rect 195502 119550 195644 119614
rect 195432 119544 195644 119550
rect 195840 119750 196052 119756
rect 195840 119686 195982 119750
rect 196046 119686 196052 119750
rect 195840 119614 196052 119686
rect 195840 119550 195846 119614
rect 195910 119550 196052 119614
rect 195840 119544 196052 119550
rect 196248 119614 196460 119756
rect 196248 119550 196254 119614
rect 196318 119550 196460 119614
rect 196248 119544 196460 119550
rect 196656 119750 196868 119756
rect 196656 119686 196798 119750
rect 196862 119686 196868 119750
rect 196656 119614 196868 119686
rect 215016 119680 215908 119756
rect 216784 119812 216996 119816
rect 216784 119756 216908 119812
rect 216964 119756 216996 119812
rect 216784 119680 216996 119756
rect 196656 119550 196662 119614
rect 196726 119550 196868 119614
rect 196656 119544 196868 119550
rect 28288 119484 28364 119544
rect 190128 119484 190204 119544
rect 21760 119342 21972 119348
rect 21760 119278 21766 119342
rect 21830 119278 21972 119342
rect 21760 119136 21972 119278
rect 22168 119206 22380 119348
rect 22478 119342 22788 119348
rect 22440 119278 22446 119342
rect 22510 119278 22788 119342
rect 22478 119272 22788 119278
rect 22168 119142 22310 119206
rect 22374 119142 22380 119206
rect 22168 119136 22380 119142
rect 22576 119136 22788 119272
rect 22984 119342 23196 119348
rect 22984 119278 23126 119342
rect 23190 119278 23196 119342
rect 22984 119206 23196 119278
rect 22984 119142 23126 119206
rect 23190 119142 23196 119206
rect 22984 119136 23196 119142
rect 23392 119342 23604 119348
rect 23392 119278 23534 119342
rect 23598 119278 23604 119342
rect 23392 119206 23604 119278
rect 28288 119272 28636 119484
rect 190128 119272 190340 119484
rect 195024 119342 195236 119348
rect 195024 119278 195166 119342
rect 195230 119278 195236 119342
rect 28424 119212 28500 119272
rect 190128 119212 190204 119272
rect 23392 119142 23534 119206
rect 23598 119142 23604 119206
rect 23392 119136 23604 119142
rect 21760 119076 21836 119136
rect 22576 119076 22652 119136
rect 21760 118798 21972 119076
rect 22304 119000 22652 119076
rect 28288 119000 28636 119212
rect 190128 119000 190340 119212
rect 195024 119206 195236 119278
rect 195024 119142 195030 119206
rect 195094 119142 195236 119206
rect 195024 119136 195236 119142
rect 195432 119342 195644 119348
rect 195432 119278 195438 119342
rect 195502 119278 195644 119342
rect 195432 119206 195644 119278
rect 195432 119142 195438 119206
rect 195502 119142 195644 119206
rect 195432 119136 195644 119142
rect 195840 119342 196052 119348
rect 195840 119278 195846 119342
rect 195910 119278 196052 119342
rect 195840 119206 196052 119278
rect 196248 119342 196460 119348
rect 196248 119278 196254 119342
rect 196318 119278 196460 119342
rect 196248 119212 196460 119278
rect 196150 119206 196460 119212
rect 195840 119142 195846 119206
rect 195910 119142 196052 119206
rect 196112 119142 196118 119206
rect 196182 119142 196460 119206
rect 195840 119136 196052 119142
rect 196150 119136 196460 119142
rect 196656 119342 196868 119348
rect 196656 119278 196662 119342
rect 196726 119278 196868 119342
rect 196656 119136 196868 119278
rect 196792 119076 196868 119136
rect 22304 118940 22380 119000
rect 28288 118940 28364 119000
rect 190264 118940 190340 119000
rect 21760 118734 21902 118798
rect 21966 118734 21972 118798
rect 21760 118728 21972 118734
rect 22168 118934 22788 118940
rect 22168 118870 22310 118934
rect 22374 118870 22788 118934
rect 22168 118864 22788 118870
rect 22168 118728 22380 118864
rect 22576 118798 22788 118864
rect 22576 118734 22718 118798
rect 22782 118734 22788 118798
rect 22576 118728 22788 118734
rect 22984 118934 23196 118940
rect 22984 118870 23126 118934
rect 23190 118870 23196 118934
rect 22984 118798 23196 118870
rect 22984 118734 22990 118798
rect 23054 118734 23196 118798
rect 22984 118728 23196 118734
rect 23392 118934 23604 118940
rect 23392 118870 23534 118934
rect 23598 118870 23604 118934
rect 23392 118798 23604 118870
rect 23392 118734 23398 118798
rect 23462 118734 23604 118798
rect 23392 118728 23604 118734
rect 28288 118728 28636 118940
rect 190128 118728 190340 118940
rect 195024 118934 195236 118940
rect 195024 118870 195030 118934
rect 195094 118870 195236 118934
rect 195024 118798 195236 118870
rect 195024 118734 195030 118798
rect 195094 118734 195236 118798
rect 195024 118728 195236 118734
rect 195432 118934 195644 118940
rect 195432 118870 195438 118934
rect 195502 118870 195644 118934
rect 195432 118798 195644 118870
rect 195432 118734 195438 118798
rect 195502 118734 195644 118798
rect 195432 118728 195644 118734
rect 195840 118934 196188 118940
rect 195840 118870 195846 118934
rect 195910 118870 196118 118934
rect 196182 118870 196188 118934
rect 195840 118864 196188 118870
rect 195840 118804 196052 118864
rect 196248 118804 196460 118940
rect 195840 118798 196460 118804
rect 195840 118734 195846 118798
rect 195910 118734 196460 118798
rect 195840 118728 196460 118734
rect 196656 118798 196868 119076
rect 196656 118734 196798 118798
rect 196862 118734 196868 118798
rect 196656 118728 196868 118734
rect 28560 118668 28636 118728
rect 190264 118668 190340 118728
rect 21760 118526 21972 118532
rect 21760 118462 21902 118526
rect 21966 118462 21972 118526
rect 21760 118320 21972 118462
rect 22168 118390 22380 118532
rect 22168 118326 22174 118390
rect 22238 118326 22380 118390
rect 22168 118320 22380 118326
rect 22576 118526 22788 118532
rect 22576 118462 22718 118526
rect 22782 118462 22788 118526
rect 22576 118390 22788 118462
rect 22576 118326 22582 118390
rect 22646 118326 22788 118390
rect 22576 118320 22788 118326
rect 22984 118526 23196 118532
rect 22984 118462 22990 118526
rect 23054 118462 23196 118526
rect 22984 118390 23196 118462
rect 22984 118326 23126 118390
rect 23190 118326 23196 118390
rect 22984 118320 23196 118326
rect 23392 118526 23604 118532
rect 23392 118462 23398 118526
rect 23462 118462 23604 118526
rect 23392 118390 23604 118462
rect 23392 118326 23534 118390
rect 23598 118326 23604 118390
rect 23392 118320 23604 118326
rect 28288 118456 28636 118668
rect 190128 118456 190340 118668
rect 195024 118526 195236 118532
rect 195024 118462 195030 118526
rect 195094 118462 195236 118526
rect 28288 118396 28364 118456
rect 190128 118396 190204 118456
rect 21760 118260 21836 118320
rect 1632 118132 1844 118260
rect 1632 118124 1702 118132
rect 1224 118118 1702 118124
rect 1224 118054 1230 118118
rect 1294 118076 1702 118118
rect 1758 118076 1844 118132
rect 1294 118054 1844 118076
rect 1224 118048 1844 118054
rect 21760 118118 21972 118260
rect 28288 118184 28636 118396
rect 190128 118184 190340 118396
rect 195024 118390 195236 118462
rect 195024 118326 195166 118390
rect 195230 118326 195236 118390
rect 195024 118320 195236 118326
rect 195432 118526 195644 118532
rect 195432 118462 195438 118526
rect 195502 118462 195644 118526
rect 195432 118390 195644 118462
rect 195432 118326 195438 118390
rect 195502 118326 195644 118390
rect 195432 118320 195644 118326
rect 195840 118526 196052 118532
rect 195840 118462 195846 118526
rect 195910 118462 196052 118526
rect 195840 118390 196052 118462
rect 196248 118396 196460 118532
rect 196150 118390 196460 118396
rect 195840 118326 195846 118390
rect 195910 118326 196052 118390
rect 196112 118326 196118 118390
rect 196182 118326 196460 118390
rect 195840 118320 196052 118326
rect 196150 118320 196460 118326
rect 196656 118526 196868 118532
rect 196656 118462 196798 118526
rect 196862 118462 196868 118526
rect 196656 118320 196868 118462
rect 215016 118396 215228 118532
rect 215696 118526 218220 118532
rect 215696 118462 218150 118526
rect 218214 118462 218220 118526
rect 215696 118456 218220 118462
rect 215696 118396 215908 118456
rect 215016 118320 215908 118396
rect 196656 118260 196732 118320
rect 28288 118124 28364 118184
rect 190128 118124 190204 118184
rect 21760 118054 21766 118118
rect 21830 118054 21972 118118
rect 21760 118048 21972 118054
rect 22168 118118 22380 118124
rect 22168 118054 22174 118118
rect 22238 118054 22380 118118
rect 22168 117912 22380 118054
rect 22576 118118 22788 118124
rect 22576 118054 22582 118118
rect 22646 118054 22788 118118
rect 22576 117988 22788 118054
rect 22478 117982 22788 117988
rect 22440 117918 22446 117982
rect 22510 117918 22788 117982
rect 22478 117912 22788 117918
rect 22984 118118 23196 118124
rect 22984 118054 23126 118118
rect 23190 118054 23196 118118
rect 22984 117982 23196 118054
rect 22984 117918 23126 117982
rect 23190 117918 23196 117982
rect 22984 117912 23196 117918
rect 23392 118118 23604 118124
rect 23392 118054 23534 118118
rect 23598 118054 23604 118118
rect 23392 117982 23604 118054
rect 23392 117918 23398 117982
rect 23462 117918 23604 117982
rect 23392 117912 23604 117918
rect 22304 117852 22380 117912
rect 21760 117846 21972 117852
rect 21760 117782 21766 117846
rect 21830 117782 21972 117846
rect 21760 117504 21972 117782
rect 22168 117776 22788 117852
rect 22168 117716 22380 117776
rect 22168 117710 22516 117716
rect 22168 117646 22446 117710
rect 22510 117646 22516 117710
rect 22168 117640 22516 117646
rect 22168 117504 22380 117640
rect 22576 117574 22788 117776
rect 22576 117510 22582 117574
rect 22646 117510 22788 117574
rect 22576 117504 22788 117510
rect 22984 117710 23196 117716
rect 22984 117646 23126 117710
rect 23190 117646 23196 117710
rect 22984 117504 23196 117646
rect 23392 117710 23604 117716
rect 23392 117646 23398 117710
rect 23462 117646 23604 117710
rect 23392 117504 23604 117646
rect 28288 117710 28636 118124
rect 28288 117646 28294 117710
rect 28358 117646 28636 117710
rect 28288 117640 28636 117646
rect 190128 117640 190340 118124
rect 195024 118118 195236 118124
rect 195024 118054 195166 118118
rect 195230 118054 195236 118118
rect 195024 117982 195236 118054
rect 195024 117918 195030 117982
rect 195094 117918 195236 117982
rect 195024 117912 195236 117918
rect 195432 118118 195644 118124
rect 195432 118054 195438 118118
rect 195502 118054 195644 118118
rect 195432 117982 195644 118054
rect 195432 117918 195438 117982
rect 195502 117918 195644 117982
rect 195432 117912 195644 117918
rect 195840 118118 196188 118124
rect 195840 118054 195846 118118
rect 195910 118054 196118 118118
rect 196182 118054 196188 118118
rect 195840 118048 196188 118054
rect 195840 117912 196052 118048
rect 196248 117988 196460 118124
rect 196656 118118 196868 118260
rect 196656 118054 196662 118118
rect 196726 118054 196868 118118
rect 196656 118048 196868 118054
rect 216784 118254 217540 118260
rect 216784 118190 217470 118254
rect 217534 118190 217540 118254
rect 216784 118184 217540 118190
rect 216784 118132 216996 118184
rect 216784 118076 216908 118132
rect 216964 118076 216996 118132
rect 216784 118048 216996 118076
rect 195976 117852 196052 117912
rect 196112 117912 196460 117988
rect 196112 117852 196188 117912
rect 195840 117776 196188 117852
rect 195024 117710 195236 117716
rect 195024 117646 195030 117710
rect 195094 117646 195236 117710
rect 28424 117580 28500 117640
rect 190128 117580 190204 117640
rect 21760 117444 21836 117504
rect 22984 117444 23060 117504
rect 23392 117444 23468 117504
rect 21760 117302 21972 117444
rect 21760 117238 21766 117302
rect 21830 117238 21972 117302
rect 21760 117232 21972 117238
rect 22168 117096 22380 117308
rect 22576 117302 22788 117308
rect 22576 117238 22582 117302
rect 22646 117238 22788 117302
rect 22576 117096 22788 117238
rect 22984 117096 23196 117444
rect 23392 117096 23604 117444
rect 22168 117036 22244 117096
rect 22576 117036 22652 117096
rect 22984 117036 23060 117096
rect 23528 117036 23604 117096
rect 21760 117030 21972 117036
rect 21760 116966 21766 117030
rect 21830 116966 21972 117030
rect 21760 116894 21972 116966
rect 21760 116830 21902 116894
rect 21966 116830 21972 116894
rect 21760 116824 21972 116830
rect 22168 116894 22380 117036
rect 22576 116900 22788 117036
rect 22478 116894 22788 116900
rect 22168 116830 22310 116894
rect 22374 116830 22380 116894
rect 22440 116830 22446 116894
rect 22510 116830 22788 116894
rect 22168 116824 22380 116830
rect 22478 116824 22788 116830
rect 22984 116688 23196 117036
rect 23392 116688 23604 117036
rect 28288 117438 28636 117580
rect 28288 117374 28294 117438
rect 28358 117374 28430 117438
rect 28494 117374 28636 117438
rect 28288 117166 28636 117374
rect 28288 117102 28430 117166
rect 28494 117102 28636 117166
rect 28288 117030 28636 117102
rect 28288 116966 28566 117030
rect 28630 116966 28636 117030
rect 28288 116960 28636 116966
rect 190128 117438 190340 117580
rect 195024 117504 195236 117646
rect 195160 117444 195236 117504
rect 190128 117374 190134 117438
rect 190198 117374 190340 117438
rect 190128 117166 190340 117374
rect 190128 117102 190134 117166
rect 190198 117102 190340 117166
rect 190128 117030 190340 117102
rect 190128 116966 190270 117030
rect 190334 116966 190340 117030
rect 190128 116960 190340 116966
rect 195024 117096 195236 117444
rect 195432 117710 195644 117716
rect 195432 117646 195438 117710
rect 195502 117646 195644 117710
rect 195432 117504 195644 117646
rect 195840 117580 196052 117776
rect 196248 117580 196460 117852
rect 195840 117574 196460 117580
rect 195840 117510 195846 117574
rect 195910 117510 196460 117574
rect 195840 117504 196460 117510
rect 196656 117846 196868 117852
rect 196656 117782 196662 117846
rect 196726 117782 196868 117846
rect 196656 117504 196868 117782
rect 216492 117674 216558 117675
rect 216450 117610 216493 117674
rect 216557 117610 216600 117674
rect 216492 117609 216558 117610
rect 195432 117444 195508 117504
rect 196656 117444 196732 117504
rect 195432 117096 195644 117444
rect 195024 117036 195100 117096
rect 195568 117036 195644 117096
rect 22984 116628 23060 116688
rect 23528 116628 23604 116688
rect 21760 116622 21972 116628
rect 21760 116558 21902 116622
rect 21966 116558 21972 116622
rect 1224 116486 1844 116492
rect 1224 116422 1230 116486
rect 1294 116452 1844 116486
rect 1294 116422 1702 116452
rect 1224 116416 1702 116422
rect 1632 116396 1702 116416
rect 1758 116396 1844 116452
rect 21760 116486 21972 116558
rect 21760 116422 21902 116486
rect 21966 116422 21972 116486
rect 21760 116416 21972 116422
rect 22168 116622 22516 116628
rect 22168 116558 22310 116622
rect 22374 116558 22446 116622
rect 22510 116558 22516 116622
rect 22168 116552 22516 116558
rect 1632 116280 1844 116396
rect 22168 116356 22380 116552
rect 22576 116356 22788 116628
rect 22984 116486 23196 116628
rect 22984 116422 23126 116486
rect 23190 116422 23196 116486
rect 22984 116416 23196 116422
rect 23392 116486 23604 116628
rect 23392 116422 23534 116486
rect 23598 116422 23604 116486
rect 23392 116416 23604 116422
rect 28288 116758 28636 116764
rect 28288 116694 28566 116758
rect 28630 116694 28636 116758
rect 28288 116622 28636 116694
rect 28288 116558 28430 116622
rect 28494 116558 28636 116622
rect 28288 116416 28636 116558
rect 190128 116758 190340 116764
rect 190128 116694 190270 116758
rect 190334 116694 190340 116758
rect 190128 116622 190340 116694
rect 190128 116558 190270 116622
rect 190334 116558 190340 116622
rect 190128 116416 190340 116558
rect 195024 116688 195236 117036
rect 195432 116688 195644 117036
rect 195840 117302 196052 117308
rect 195840 117238 195846 117302
rect 195910 117238 196052 117302
rect 195840 117096 196052 117238
rect 196248 117096 196460 117308
rect 196656 117302 196868 117444
rect 196656 117238 196662 117302
rect 196726 117238 196868 117302
rect 196656 117232 196868 117238
rect 195840 117036 195916 117096
rect 196248 117036 196324 117096
rect 195840 116894 196052 117036
rect 196248 116900 196460 117036
rect 196150 116894 196460 116900
rect 195840 116830 195846 116894
rect 195910 116830 196052 116894
rect 196112 116830 196118 116894
rect 196182 116830 196460 116894
rect 195840 116824 196052 116830
rect 196150 116824 196460 116830
rect 196656 117030 196868 117036
rect 196656 116966 196662 117030
rect 196726 116966 196868 117030
rect 196656 116894 196868 116966
rect 196656 116830 196798 116894
rect 196862 116830 196868 116894
rect 196656 116824 196868 116830
rect 215016 116960 215908 117036
rect 215016 116824 215228 116960
rect 215696 116900 215908 116960
rect 215696 116894 216860 116900
rect 215696 116830 216790 116894
rect 216854 116830 216860 116894
rect 215696 116824 216860 116830
rect 195024 116628 195100 116688
rect 195568 116628 195644 116688
rect 195024 116486 195236 116628
rect 195024 116422 195166 116486
rect 195230 116422 195236 116486
rect 195024 116416 195236 116422
rect 195432 116486 195644 116628
rect 195432 116422 195438 116486
rect 195502 116422 195644 116486
rect 195432 116416 195644 116422
rect 195840 116622 196188 116628
rect 195840 116558 195846 116622
rect 195910 116558 196118 116622
rect 196182 116558 196188 116622
rect 195840 116552 196188 116558
rect 195840 116492 196052 116552
rect 196248 116492 196460 116628
rect 195840 116416 196460 116492
rect 196656 116622 196868 116628
rect 196656 116558 196798 116622
rect 196862 116558 196868 116622
rect 196656 116486 196868 116558
rect 196656 116422 196798 116486
rect 196862 116422 196868 116486
rect 196656 116416 196868 116422
rect 216784 116486 216996 116492
rect 216784 116422 216790 116486
rect 216854 116452 216996 116486
rect 216854 116422 216908 116452
rect 22168 116280 22788 116356
rect 22712 116220 22788 116280
rect 28288 116356 28364 116416
rect 190264 116356 190340 116416
rect 28288 116350 28636 116356
rect 28288 116286 28430 116350
rect 28494 116286 28636 116350
rect 21760 116214 21972 116220
rect 21760 116150 21902 116214
rect 21966 116150 21972 116214
rect 21760 116078 21972 116150
rect 21760 116014 21902 116078
rect 21966 116014 21972 116078
rect 21760 116008 21972 116014
rect 22168 116078 22380 116220
rect 22168 116014 22174 116078
rect 22238 116014 22380 116078
rect 22168 116008 22380 116014
rect 22576 116078 22788 116220
rect 22576 116014 22582 116078
rect 22646 116014 22788 116078
rect 22576 116008 22788 116014
rect 22984 116214 23196 116220
rect 22984 116150 23126 116214
rect 23190 116150 23196 116214
rect 22984 116078 23196 116150
rect 22984 116014 22990 116078
rect 23054 116014 23196 116078
rect 22984 116008 23196 116014
rect 23392 116214 23604 116220
rect 23392 116150 23534 116214
rect 23598 116150 23604 116214
rect 23392 116078 23604 116150
rect 23392 116014 23398 116078
rect 23462 116014 23604 116078
rect 23392 116008 23604 116014
rect 28288 116144 28636 116286
rect 190128 116350 190340 116356
rect 190128 116286 190270 116350
rect 190334 116286 190340 116350
rect 190128 116144 190340 116286
rect 195840 116280 196052 116416
rect 196248 116280 196460 116416
rect 216784 116396 216908 116422
rect 216964 116396 216996 116452
rect 216784 116356 216996 116396
rect 216784 116350 217540 116356
rect 216784 116286 217470 116350
rect 217534 116286 217540 116350
rect 216784 116280 217540 116286
rect 196248 116220 196324 116280
rect 195024 116214 195236 116220
rect 195024 116150 195166 116214
rect 195230 116150 195236 116214
rect 28288 116084 28364 116144
rect 190128 116084 190204 116144
rect 28288 115872 28636 116084
rect 28560 115812 28636 115872
rect 21760 115806 21972 115812
rect 21760 115742 21902 115806
rect 21966 115742 21972 115806
rect 21760 115670 21972 115742
rect 21760 115606 21902 115670
rect 21966 115606 21972 115670
rect 21760 115600 21972 115606
rect 22168 115806 22788 115812
rect 22168 115742 22174 115806
rect 22238 115742 22582 115806
rect 22646 115742 22788 115806
rect 22168 115736 22788 115742
rect 22168 115676 22380 115736
rect 22168 115670 22516 115676
rect 22168 115606 22310 115670
rect 22374 115606 22446 115670
rect 22510 115606 22516 115670
rect 22168 115600 22516 115606
rect 22576 115600 22788 115736
rect 22984 115806 23196 115812
rect 22984 115742 22990 115806
rect 23054 115742 23196 115806
rect 22984 115670 23196 115742
rect 22984 115606 22990 115670
rect 23054 115606 23196 115670
rect 22984 115600 23196 115606
rect 23392 115806 23604 115812
rect 23392 115742 23398 115806
rect 23462 115742 23604 115806
rect 23392 115670 23604 115742
rect 23392 115606 23398 115670
rect 23462 115606 23604 115670
rect 23392 115600 23604 115606
rect 28288 115600 28636 115812
rect 190128 115872 190340 116084
rect 195024 116078 195236 116150
rect 195024 116014 195166 116078
rect 195230 116014 195236 116078
rect 195024 116008 195236 116014
rect 195432 116214 195644 116220
rect 195432 116150 195438 116214
rect 195502 116150 195644 116214
rect 195432 116078 195644 116150
rect 195432 116014 195438 116078
rect 195502 116014 195644 116078
rect 195432 116008 195644 116014
rect 195840 116078 196052 116220
rect 196248 116084 196460 116220
rect 196150 116078 196460 116084
rect 195840 116014 195982 116078
rect 196046 116014 196052 116078
rect 196112 116014 196118 116078
rect 196182 116014 196460 116078
rect 195840 116008 196052 116014
rect 196150 116008 196460 116014
rect 196656 116214 196868 116220
rect 196656 116150 196798 116214
rect 196862 116150 196868 116214
rect 196656 116078 196868 116150
rect 196656 116014 196798 116078
rect 196862 116014 196868 116078
rect 196656 116008 196868 116014
rect 190128 115812 190204 115872
rect 190128 115600 190340 115812
rect 195024 115806 195236 115812
rect 195024 115742 195166 115806
rect 195230 115742 195236 115806
rect 195024 115670 195236 115742
rect 195024 115606 195030 115670
rect 195094 115606 195236 115670
rect 195024 115600 195236 115606
rect 195432 115806 195644 115812
rect 195432 115742 195438 115806
rect 195502 115742 195644 115806
rect 195432 115670 195644 115742
rect 195432 115606 195438 115670
rect 195502 115606 195644 115670
rect 195432 115600 195644 115606
rect 195840 115806 196188 115812
rect 195840 115742 195982 115806
rect 196046 115742 196118 115806
rect 196182 115742 196188 115806
rect 195840 115736 196188 115742
rect 195840 115676 196052 115736
rect 196248 115676 196460 115812
rect 195840 115670 196460 115676
rect 195840 115606 196390 115670
rect 196454 115606 196460 115670
rect 195840 115600 196460 115606
rect 196656 115806 196868 115812
rect 196656 115742 196798 115806
rect 196862 115742 196868 115806
rect 196656 115670 196868 115742
rect 196656 115606 196798 115670
rect 196862 115606 196868 115670
rect 196656 115600 196868 115606
rect 28560 115540 28636 115600
rect 190264 115540 190340 115600
rect 21760 115398 21972 115404
rect 21760 115334 21902 115398
rect 21966 115334 21972 115398
rect 21760 115262 21972 115334
rect 21760 115198 21766 115262
rect 21830 115198 21972 115262
rect 21760 115192 21972 115198
rect 22168 115398 22380 115404
rect 22478 115398 22788 115404
rect 22168 115334 22310 115398
rect 22374 115334 22380 115398
rect 22440 115334 22446 115398
rect 22510 115334 22788 115398
rect 22168 115268 22380 115334
rect 22478 115328 22788 115334
rect 22168 115262 22516 115268
rect 22168 115198 22174 115262
rect 22238 115198 22446 115262
rect 22510 115198 22516 115262
rect 22168 115192 22516 115198
rect 22576 115192 22788 115328
rect 22984 115398 23196 115404
rect 22984 115334 22990 115398
rect 23054 115334 23196 115398
rect 22984 115262 23196 115334
rect 22984 115198 23126 115262
rect 23190 115198 23196 115262
rect 22984 115192 23196 115198
rect 23392 115398 23604 115404
rect 23392 115334 23398 115398
rect 23462 115334 23604 115398
rect 23392 115262 23604 115334
rect 28288 115328 28636 115540
rect 28560 115268 28636 115328
rect 23392 115198 23534 115262
rect 23598 115198 23604 115262
rect 23392 115192 23604 115198
rect 28288 115056 28636 115268
rect 190128 115328 190340 115540
rect 195024 115398 195236 115404
rect 195024 115334 195030 115398
rect 195094 115334 195236 115398
rect 190128 115268 190204 115328
rect 190128 115056 190340 115268
rect 195024 115262 195236 115334
rect 195024 115198 195166 115262
rect 195230 115198 195236 115262
rect 195024 115192 195236 115198
rect 195432 115398 195644 115404
rect 195432 115334 195438 115398
rect 195502 115334 195644 115398
rect 195432 115262 195644 115334
rect 195432 115198 195438 115262
rect 195502 115198 195644 115262
rect 195432 115192 195644 115198
rect 195840 115262 196052 115404
rect 195840 115198 195846 115262
rect 195910 115198 196052 115262
rect 195840 115192 196052 115198
rect 196248 115398 196460 115404
rect 196248 115334 196390 115398
rect 196454 115334 196460 115398
rect 196248 115262 196460 115334
rect 196248 115198 196254 115262
rect 196318 115198 196460 115262
rect 196248 115192 196460 115198
rect 196656 115398 196868 115404
rect 196656 115334 196798 115398
rect 196862 115334 196868 115398
rect 196656 115262 196868 115334
rect 196656 115198 196662 115262
rect 196726 115198 196868 115262
rect 196656 115192 196868 115198
rect 28424 114996 28500 115056
rect 190128 114996 190204 115056
rect 21760 114990 21972 114996
rect 21760 114926 21766 114990
rect 21830 114926 21972 114990
rect 1632 114772 1844 114860
rect 21760 114854 21972 114926
rect 21760 114790 21766 114854
rect 21830 114790 21972 114854
rect 21760 114784 21972 114790
rect 22168 114990 22380 114996
rect 22478 114990 22788 114996
rect 22168 114926 22174 114990
rect 22238 114926 22380 114990
rect 22440 114926 22446 114990
rect 22510 114926 22788 114990
rect 22168 114784 22380 114926
rect 22478 114920 22788 114926
rect 22576 114860 22788 114920
rect 22478 114854 22788 114860
rect 22440 114790 22446 114854
rect 22510 114790 22788 114854
rect 22478 114784 22788 114790
rect 22984 114990 23196 114996
rect 22984 114926 23126 114990
rect 23190 114926 23196 114990
rect 22984 114854 23196 114926
rect 22984 114790 23126 114854
rect 23190 114790 23196 114854
rect 22984 114784 23196 114790
rect 23392 114990 23604 114996
rect 23392 114926 23534 114990
rect 23598 114926 23604 114990
rect 23392 114854 23604 114926
rect 23392 114790 23398 114854
rect 23462 114790 23604 114854
rect 23392 114784 23604 114790
rect 28288 114784 28636 114996
rect 190128 114784 190340 114996
rect 195024 114990 195236 114996
rect 195024 114926 195166 114990
rect 195230 114926 195236 114990
rect 195024 114854 195236 114926
rect 195024 114790 195030 114854
rect 195094 114790 195236 114854
rect 195024 114784 195236 114790
rect 195432 114990 195644 114996
rect 195432 114926 195438 114990
rect 195502 114926 195644 114990
rect 195432 114854 195644 114926
rect 195432 114790 195574 114854
rect 195638 114790 195644 114854
rect 195432 114784 195644 114790
rect 195840 114990 196052 114996
rect 195840 114926 195846 114990
rect 195910 114926 196052 114990
rect 195840 114854 196052 114926
rect 195840 114790 195982 114854
rect 196046 114790 196052 114854
rect 195840 114784 196052 114790
rect 196248 114990 196460 114996
rect 196248 114926 196254 114990
rect 196318 114926 196460 114990
rect 196248 114784 196460 114926
rect 196656 114990 196868 114996
rect 196656 114926 196662 114990
rect 196726 114926 196868 114990
rect 196656 114854 196868 114926
rect 196656 114790 196798 114854
rect 196862 114790 196868 114854
rect 196656 114784 196868 114790
rect 216784 114854 217540 114860
rect 216784 114790 217470 114854
rect 217534 114790 217540 114854
rect 216784 114784 217540 114790
rect 1632 114724 1702 114772
rect 1224 114718 1702 114724
rect 1224 114654 1230 114718
rect 1294 114716 1702 114718
rect 1758 114716 1844 114772
rect 28424 114724 28500 114784
rect 190128 114724 190204 114784
rect 196248 114724 196324 114784
rect 1294 114654 1844 114716
rect 1224 114648 1844 114654
rect 21760 114582 21972 114588
rect 21760 114518 21766 114582
rect 21830 114518 21972 114582
rect 21760 114376 21972 114518
rect 22168 114582 22516 114588
rect 22168 114518 22446 114582
rect 22510 114518 22516 114582
rect 22168 114512 22516 114518
rect 22168 114452 22380 114512
rect 22576 114452 22788 114588
rect 22168 114446 22788 114452
rect 22168 114382 22174 114446
rect 22238 114382 22788 114446
rect 22168 114376 22788 114382
rect 22984 114582 23196 114588
rect 22984 114518 23126 114582
rect 23190 114518 23196 114582
rect 22984 114446 23196 114518
rect 22984 114382 22990 114446
rect 23054 114382 23196 114446
rect 22984 114376 23196 114382
rect 23392 114582 23604 114588
rect 23392 114518 23398 114582
rect 23462 114518 23604 114582
rect 23392 114446 23604 114518
rect 23392 114382 23534 114446
rect 23598 114382 23604 114446
rect 23392 114376 23604 114382
rect 28288 114512 28636 114724
rect 190128 114512 190340 114724
rect 195976 114648 196324 114724
rect 216784 114772 216996 114784
rect 216784 114716 216908 114772
rect 216964 114716 216996 114772
rect 216784 114648 216996 114716
rect 195976 114588 196052 114648
rect 28288 114452 28364 114512
rect 190264 114452 190340 114512
rect 21760 114316 21836 114376
rect 21760 113968 21972 114316
rect 28288 114310 28636 114452
rect 28288 114246 28566 114310
rect 28630 114246 28636 114310
rect 28288 114240 28636 114246
rect 190128 114310 190340 114452
rect 195024 114582 195236 114588
rect 195024 114518 195030 114582
rect 195094 114518 195236 114582
rect 195024 114446 195236 114518
rect 195024 114382 195030 114446
rect 195094 114382 195236 114446
rect 195024 114376 195236 114382
rect 195432 114582 195644 114588
rect 195432 114518 195574 114582
rect 195638 114518 195644 114582
rect 195432 114446 195644 114518
rect 195432 114382 195438 114446
rect 195502 114382 195644 114446
rect 195432 114376 195644 114382
rect 195840 114582 196460 114588
rect 195840 114518 195982 114582
rect 196046 114518 196460 114582
rect 195840 114512 196460 114518
rect 195840 114376 196052 114512
rect 196248 114446 196460 114512
rect 196248 114382 196390 114446
rect 196454 114382 196460 114446
rect 196248 114376 196460 114382
rect 196656 114582 196868 114588
rect 196656 114518 196798 114582
rect 196862 114518 196868 114582
rect 196656 114376 196868 114518
rect 196792 114316 196868 114376
rect 190128 114246 190270 114310
rect 190334 114246 190340 114310
rect 190128 114240 190340 114246
rect 28288 114180 28364 114240
rect 190264 114180 190340 114240
rect 22168 114174 22380 114180
rect 22168 114110 22174 114174
rect 22238 114110 22380 114174
rect 22168 113968 22380 114110
rect 22576 114044 22788 114180
rect 22440 113968 22788 114044
rect 22984 114174 23196 114180
rect 22984 114110 22990 114174
rect 23054 114110 23196 114174
rect 22984 114038 23196 114110
rect 22984 113974 23126 114038
rect 23190 113974 23196 114038
rect 22984 113968 23196 113974
rect 23392 114174 23604 114180
rect 23392 114110 23534 114174
rect 23598 114110 23604 114174
rect 23392 114038 23604 114110
rect 23392 113974 23534 114038
rect 23598 113974 23604 114038
rect 23392 113968 23604 113974
rect 28288 114038 28636 114180
rect 28288 113974 28566 114038
rect 28630 113974 28636 114038
rect 21760 113908 21836 113968
rect 22168 113908 22244 113968
rect 22440 113908 22516 113968
rect 22712 113908 22788 113968
rect 21760 113560 21972 113908
rect 22168 113832 22516 113908
rect 22168 113630 22380 113832
rect 22168 113566 22174 113630
rect 22238 113566 22380 113630
rect 22168 113560 22380 113566
rect 22576 113560 22788 113908
rect 22984 113766 23196 113772
rect 22984 113702 23126 113766
rect 23190 113702 23196 113766
rect 22984 113560 23196 113702
rect 23392 113766 23604 113772
rect 23392 113702 23534 113766
rect 23598 113702 23604 113766
rect 23392 113560 23604 113702
rect 28288 113766 28636 113974
rect 28288 113702 28294 113766
rect 28358 113702 28636 113766
rect 28288 113696 28636 113702
rect 190128 114038 190340 114180
rect 190128 113974 190270 114038
rect 190334 113974 190340 114038
rect 190128 113696 190340 113974
rect 195024 114174 195236 114180
rect 195024 114110 195030 114174
rect 195094 114110 195236 114174
rect 195024 114038 195236 114110
rect 195024 113974 195166 114038
rect 195230 113974 195236 114038
rect 195024 113968 195236 113974
rect 195432 114174 195644 114180
rect 195432 114110 195438 114174
rect 195502 114110 195644 114174
rect 195432 114038 195644 114110
rect 195432 113974 195574 114038
rect 195638 113974 195644 114038
rect 195432 113968 195644 113974
rect 195840 113968 196052 114180
rect 196248 114174 196460 114180
rect 196248 114110 196390 114174
rect 196454 114110 196460 114174
rect 196248 113968 196460 114110
rect 196656 113968 196868 114316
rect 195840 113908 195916 113968
rect 196384 113908 196460 113968
rect 196792 113908 196868 113968
rect 28560 113636 28636 113696
rect 190264 113636 190340 113696
rect 21896 113500 21972 113560
rect 21760 113358 21972 113500
rect 22984 113500 23060 113560
rect 23392 113500 23468 113560
rect 21760 113294 21766 113358
rect 21830 113294 21972 113358
rect 21760 113288 21972 113294
rect 22168 113358 22380 113364
rect 22168 113294 22174 113358
rect 22238 113294 22380 113358
rect 22168 113228 22380 113294
rect 22576 113228 22788 113364
rect 1632 113092 1844 113228
rect 22168 113152 22788 113228
rect 22984 113152 23196 113500
rect 23392 113152 23604 113500
rect 28288 113494 28636 113636
rect 28288 113430 28294 113494
rect 28358 113430 28636 113494
rect 22168 113092 22244 113152
rect 22576 113092 22652 113152
rect 22984 113092 23060 113152
rect 23392 113092 23468 113152
rect 1224 113086 1702 113092
rect 1224 113022 1230 113086
rect 1294 113036 1702 113086
rect 1758 113036 1844 113092
rect 1294 113022 1844 113036
rect 1224 113016 1844 113022
rect 1632 112880 1844 113016
rect 21760 113086 21972 113092
rect 21760 113022 21766 113086
rect 21830 113022 21972 113086
rect 21760 112950 21972 113022
rect 21760 112886 21766 112950
rect 21830 112886 21972 112950
rect 21760 112880 21972 112886
rect 22168 112880 22380 113092
rect 22576 112950 22788 113092
rect 22576 112886 22582 112950
rect 22646 112886 22788 112950
rect 22576 112880 22788 112886
rect 22984 112744 23196 113092
rect 23392 112744 23604 113092
rect 28288 113086 28636 113430
rect 28288 113022 28430 113086
rect 28494 113022 28636 113086
rect 28288 113016 28636 113022
rect 190128 113494 190340 113636
rect 190128 113430 190134 113494
rect 190198 113430 190340 113494
rect 190128 113222 190340 113430
rect 190128 113158 190134 113222
rect 190198 113158 190270 113222
rect 190334 113158 190340 113222
rect 190128 113086 190340 113158
rect 195024 113766 195236 113772
rect 195024 113702 195166 113766
rect 195230 113702 195236 113766
rect 195024 113560 195236 113702
rect 195432 113766 195644 113772
rect 195432 113702 195574 113766
rect 195638 113702 195644 113766
rect 195432 113560 195644 113702
rect 195840 113630 196052 113908
rect 196248 113636 196460 113908
rect 196150 113630 196460 113636
rect 195840 113566 195982 113630
rect 196046 113566 196052 113630
rect 196112 113566 196118 113630
rect 196182 113566 196460 113630
rect 195840 113560 196052 113566
rect 196150 113560 196460 113566
rect 196656 113560 196868 113908
rect 195024 113500 195100 113560
rect 195432 113500 195508 113560
rect 196656 113500 196732 113560
rect 195024 113152 195236 113500
rect 195160 113092 195236 113152
rect 190128 113022 190134 113086
rect 190198 113022 190340 113086
rect 190128 113016 190340 113022
rect 22984 112684 23060 112744
rect 23528 112684 23604 112744
rect 21760 112678 21972 112684
rect 21760 112614 21766 112678
rect 21830 112614 21972 112678
rect 21760 112542 21972 112614
rect 21760 112478 21902 112542
rect 21966 112478 21972 112542
rect 21760 112472 21972 112478
rect 22168 112336 22380 112684
rect 22304 112276 22380 112336
rect 22576 112678 22788 112684
rect 22576 112614 22582 112678
rect 22646 112614 22788 112678
rect 22576 112336 22788 112614
rect 22984 112542 23196 112684
rect 22984 112478 23126 112542
rect 23190 112478 23196 112542
rect 22984 112472 23196 112478
rect 23392 112542 23604 112684
rect 23392 112478 23398 112542
rect 23462 112478 23604 112542
rect 23392 112472 23604 112478
rect 28288 112814 28636 112820
rect 28288 112750 28430 112814
rect 28494 112750 28636 112814
rect 28288 112472 28636 112750
rect 190128 112814 190340 112820
rect 190128 112750 190270 112814
rect 190334 112750 190340 112814
rect 190128 112678 190340 112750
rect 190128 112614 190134 112678
rect 190198 112614 190340 112678
rect 190128 112472 190340 112614
rect 195024 112744 195236 113092
rect 195432 113152 195644 113500
rect 195840 113358 196188 113364
rect 195840 113294 195982 113358
rect 196046 113294 196118 113358
rect 196182 113294 196188 113358
rect 195840 113288 196188 113294
rect 195840 113228 196052 113288
rect 196248 113228 196460 113364
rect 196656 113358 196868 113500
rect 196656 113294 196662 113358
rect 196726 113294 196868 113358
rect 196656 113288 196868 113294
rect 195840 113152 196460 113228
rect 195432 113092 195508 113152
rect 195976 113092 196052 113152
rect 196384 113092 196460 113152
rect 216784 113092 216996 113228
rect 195432 112744 195644 113092
rect 195840 112950 196052 113092
rect 195840 112886 195982 112950
rect 196046 112886 196052 112950
rect 195840 112880 196052 112886
rect 196248 112880 196460 113092
rect 196656 113086 196868 113092
rect 196656 113022 196662 113086
rect 196726 113022 196868 113086
rect 196656 112950 196868 113022
rect 196656 112886 196662 112950
rect 196726 112886 196868 112950
rect 196656 112880 196868 112886
rect 216784 113036 216908 113092
rect 216964 113036 216996 113092
rect 216784 112956 216996 113036
rect 216784 112950 217540 112956
rect 216784 112886 217470 112950
rect 217534 112886 217540 112950
rect 216784 112880 217540 112886
rect 195024 112684 195100 112744
rect 195432 112684 195508 112744
rect 195024 112542 195236 112684
rect 195024 112478 195030 112542
rect 195094 112478 195236 112542
rect 195024 112472 195236 112478
rect 195432 112542 195644 112684
rect 195432 112478 195574 112542
rect 195638 112478 195644 112542
rect 195432 112472 195644 112478
rect 195840 112678 196052 112684
rect 195840 112614 195982 112678
rect 196046 112614 196052 112678
rect 28288 112412 28364 112472
rect 190264 112412 190340 112472
rect 22576 112276 22652 112336
rect 21760 112270 21972 112276
rect 21760 112206 21902 112270
rect 21966 112206 21972 112270
rect 21760 112134 21972 112206
rect 21760 112070 21902 112134
rect 21966 112070 21972 112134
rect 21760 112064 21972 112070
rect 22168 112200 22788 112276
rect 22168 112140 22380 112200
rect 22168 112134 22516 112140
rect 22168 112070 22310 112134
rect 22374 112070 22446 112134
rect 22510 112070 22516 112134
rect 22168 112064 22516 112070
rect 22576 112064 22788 112200
rect 22984 112270 23196 112276
rect 22984 112206 23126 112270
rect 23190 112206 23196 112270
rect 22984 112134 23196 112206
rect 22984 112070 22990 112134
rect 23054 112070 23196 112134
rect 22984 112064 23196 112070
rect 23392 112270 23604 112276
rect 23392 112206 23398 112270
rect 23462 112206 23604 112270
rect 23392 112134 23604 112206
rect 28288 112200 28636 112412
rect 190128 112200 190340 112412
rect 195840 112412 196052 112614
rect 195840 112336 196188 112412
rect 196112 112276 196188 112336
rect 196248 112336 196460 112684
rect 196656 112678 196868 112684
rect 196656 112614 196662 112678
rect 196726 112614 196868 112678
rect 196656 112542 196868 112614
rect 196656 112478 196798 112542
rect 196862 112478 196868 112542
rect 196656 112472 196868 112478
rect 196248 112276 196324 112336
rect 28424 112140 28500 112200
rect 190264 112140 190340 112200
rect 23392 112070 23398 112134
rect 23462 112070 23604 112134
rect 23392 112064 23604 112070
rect 21760 111862 21972 111868
rect 21760 111798 21902 111862
rect 21966 111798 21972 111862
rect 21760 111726 21972 111798
rect 21760 111662 21902 111726
rect 21966 111662 21972 111726
rect 21760 111656 21972 111662
rect 22168 111862 22380 111868
rect 22478 111862 22788 111868
rect 22168 111798 22310 111862
rect 22374 111798 22380 111862
rect 22440 111798 22446 111862
rect 22510 111798 22788 111862
rect 22168 111726 22380 111798
rect 22478 111792 22788 111798
rect 22168 111662 22174 111726
rect 22238 111662 22380 111726
rect 22168 111656 22380 111662
rect 22576 111726 22788 111792
rect 22576 111662 22582 111726
rect 22646 111662 22788 111726
rect 22576 111656 22788 111662
rect 22984 111862 23196 111868
rect 22984 111798 22990 111862
rect 23054 111798 23196 111862
rect 22984 111726 23196 111798
rect 22984 111662 23126 111726
rect 23190 111662 23196 111726
rect 22984 111656 23196 111662
rect 23392 111862 23604 111868
rect 23392 111798 23398 111862
rect 23462 111798 23604 111862
rect 23392 111726 23604 111798
rect 23392 111662 23534 111726
rect 23598 111662 23604 111726
rect 23392 111656 23604 111662
rect 28288 111862 28636 112140
rect 28288 111798 28294 111862
rect 28358 111798 28636 111862
rect 28288 111656 28636 111798
rect 28560 111596 28636 111656
rect 28288 111590 28636 111596
rect 28288 111526 28294 111590
rect 28358 111526 28636 111590
rect 1632 111412 1844 111460
rect 1632 111356 1702 111412
rect 1758 111356 1844 111412
rect 1632 111324 1844 111356
rect 1224 111318 1844 111324
rect 1224 111254 1230 111318
rect 1294 111254 1844 111318
rect 1224 111248 1844 111254
rect 21760 111454 21972 111460
rect 21760 111390 21902 111454
rect 21966 111390 21972 111454
rect 21760 111318 21972 111390
rect 21760 111254 21902 111318
rect 21966 111254 21972 111318
rect 21760 111248 21972 111254
rect 22168 111454 22380 111460
rect 22168 111390 22174 111454
rect 22238 111390 22380 111454
rect 22168 111324 22380 111390
rect 22576 111454 22788 111460
rect 22576 111390 22582 111454
rect 22646 111390 22788 111454
rect 22168 111318 22516 111324
rect 22168 111254 22446 111318
rect 22510 111254 22516 111318
rect 22168 111248 22516 111254
rect 22576 111248 22788 111390
rect 22984 111454 23196 111460
rect 22984 111390 23126 111454
rect 23190 111390 23196 111454
rect 22984 111318 23196 111390
rect 22984 111254 23126 111318
rect 23190 111254 23196 111318
rect 22984 111248 23196 111254
rect 23392 111454 23604 111460
rect 23392 111390 23534 111454
rect 23598 111390 23604 111454
rect 23392 111318 23604 111390
rect 28288 111384 28636 111526
rect 190128 111656 190340 112140
rect 195024 112270 195236 112276
rect 195024 112206 195030 112270
rect 195094 112206 195236 112270
rect 195024 112134 195236 112206
rect 195024 112070 195030 112134
rect 195094 112070 195236 112134
rect 195024 112064 195236 112070
rect 195432 112270 195644 112276
rect 195432 112206 195574 112270
rect 195638 112206 195644 112270
rect 195432 112134 195644 112206
rect 195432 112070 195438 112134
rect 195502 112070 195644 112134
rect 195432 112064 195644 112070
rect 195840 112140 196052 112276
rect 196112 112200 196460 112276
rect 196248 112140 196460 112200
rect 195840 112064 196460 112140
rect 196656 112270 196868 112276
rect 196656 112206 196798 112270
rect 196862 112206 196868 112270
rect 196656 112134 196868 112206
rect 196656 112070 196662 112134
rect 196726 112070 196868 112134
rect 196656 112064 196868 112070
rect 196248 112004 196324 112064
rect 196112 111928 196324 112004
rect 196112 111868 196188 111928
rect 195024 111862 195236 111868
rect 195024 111798 195030 111862
rect 195094 111798 195236 111862
rect 195024 111726 195236 111798
rect 195024 111662 195030 111726
rect 195094 111662 195236 111726
rect 195024 111656 195236 111662
rect 195432 111862 195644 111868
rect 195432 111798 195438 111862
rect 195502 111798 195644 111862
rect 195432 111726 195644 111798
rect 195432 111662 195574 111726
rect 195638 111662 195644 111726
rect 195432 111656 195644 111662
rect 195840 111792 196188 111868
rect 195840 111726 196052 111792
rect 195840 111662 195982 111726
rect 196046 111662 196052 111726
rect 195840 111656 196052 111662
rect 196248 111656 196460 111868
rect 196656 111862 196868 111868
rect 196656 111798 196662 111862
rect 196726 111798 196868 111862
rect 196656 111726 196868 111798
rect 196656 111662 196662 111726
rect 196726 111662 196868 111726
rect 196656 111656 196868 111662
rect 190128 111596 190204 111656
rect 196248 111596 196324 111656
rect 190128 111384 190340 111596
rect 195976 111520 196324 111596
rect 195976 111460 196052 111520
rect 28424 111324 28500 111384
rect 190264 111324 190340 111384
rect 23392 111254 23398 111318
rect 23462 111254 23604 111318
rect 23392 111248 23604 111254
rect 28288 111112 28636 111324
rect 190128 111112 190340 111324
rect 195024 111454 195236 111460
rect 195024 111390 195030 111454
rect 195094 111390 195236 111454
rect 195024 111318 195236 111390
rect 195024 111254 195030 111318
rect 195094 111254 195236 111318
rect 195024 111248 195236 111254
rect 195432 111454 195644 111460
rect 195432 111390 195574 111454
rect 195638 111390 195644 111454
rect 195432 111318 195644 111390
rect 195432 111254 195438 111318
rect 195502 111254 195644 111318
rect 195432 111248 195644 111254
rect 195840 111454 196460 111460
rect 195840 111390 195982 111454
rect 196046 111390 196460 111454
rect 195840 111384 196460 111390
rect 195840 111248 196052 111384
rect 196248 111318 196460 111384
rect 196248 111254 196390 111318
rect 196454 111254 196460 111318
rect 196248 111248 196460 111254
rect 196656 111454 196868 111460
rect 196656 111390 196662 111454
rect 196726 111390 196868 111454
rect 196656 111318 196868 111390
rect 196656 111254 196798 111318
rect 196862 111254 196868 111318
rect 196656 111248 196868 111254
rect 216784 111454 217540 111460
rect 216784 111412 217470 111454
rect 216784 111356 216908 111412
rect 216964 111390 217470 111412
rect 217534 111390 217540 111454
rect 216964 111384 217540 111390
rect 216964 111356 216996 111384
rect 216784 111248 216996 111356
rect 28560 111052 28636 111112
rect 190264 111052 190340 111112
rect 21760 111046 21972 111052
rect 21760 110982 21902 111046
rect 21966 110982 21972 111046
rect 21760 110910 21972 110982
rect 21760 110846 21766 110910
rect 21830 110846 21972 110910
rect 21760 110840 21972 110846
rect 22168 110910 22380 111052
rect 22478 111046 22788 111052
rect 22440 110982 22446 111046
rect 22510 110982 22788 111046
rect 22478 110976 22788 110982
rect 22168 110846 22174 110910
rect 22238 110846 22380 110910
rect 22168 110840 22380 110846
rect 22576 110910 22788 110976
rect 22576 110846 22582 110910
rect 22646 110846 22788 110910
rect 22576 110840 22788 110846
rect 22984 111046 23196 111052
rect 22984 110982 23126 111046
rect 23190 110982 23196 111046
rect 22984 110910 23196 110982
rect 22984 110846 23126 110910
rect 23190 110846 23196 110910
rect 22984 110840 23196 110846
rect 23392 111046 23604 111052
rect 23392 110982 23398 111046
rect 23462 110982 23604 111046
rect 23392 110910 23604 110982
rect 23392 110846 23534 110910
rect 23598 110846 23604 110910
rect 23392 110840 23604 110846
rect 28288 110840 28636 111052
rect 190128 110840 190340 111052
rect 195024 111046 195236 111052
rect 195024 110982 195030 111046
rect 195094 110982 195236 111046
rect 195024 110910 195236 110982
rect 195024 110846 195166 110910
rect 195230 110846 195236 110910
rect 195024 110840 195236 110846
rect 195432 111046 195644 111052
rect 195432 110982 195438 111046
rect 195502 110982 195644 111046
rect 195432 110910 195644 110982
rect 195432 110846 195574 110910
rect 195638 110846 195644 110910
rect 195432 110840 195644 110846
rect 195840 111046 196460 111052
rect 195840 110982 196390 111046
rect 196454 110982 196460 111046
rect 195840 110976 196460 110982
rect 195840 110840 196052 110976
rect 196248 110910 196460 110976
rect 196248 110846 196254 110910
rect 196318 110846 196460 110910
rect 196248 110840 196460 110846
rect 196656 111046 196868 111052
rect 196656 110982 196798 111046
rect 196862 110982 196868 111046
rect 196656 110910 196868 110982
rect 196656 110846 196662 110910
rect 196726 110846 196868 110910
rect 196656 110840 196868 110846
rect 28288 110780 28364 110840
rect 190128 110780 190204 110840
rect 21760 110638 21972 110644
rect 21760 110574 21766 110638
rect 21830 110574 21972 110638
rect 21760 110432 21972 110574
rect 22168 110638 22380 110644
rect 22168 110574 22174 110638
rect 22238 110574 22380 110638
rect 22168 110502 22380 110574
rect 22576 110638 22788 110644
rect 22576 110574 22582 110638
rect 22646 110574 22788 110638
rect 22576 110508 22788 110574
rect 22478 110502 22788 110508
rect 22168 110438 22174 110502
rect 22238 110438 22380 110502
rect 22440 110438 22446 110502
rect 22510 110438 22788 110502
rect 22168 110432 22380 110438
rect 22478 110432 22788 110438
rect 22984 110638 23196 110644
rect 22984 110574 23126 110638
rect 23190 110574 23196 110638
rect 22984 110502 23196 110574
rect 22984 110438 23126 110502
rect 23190 110438 23196 110502
rect 22984 110432 23196 110438
rect 23392 110638 23604 110644
rect 23392 110574 23534 110638
rect 23598 110574 23604 110638
rect 23392 110502 23604 110574
rect 28288 110568 28636 110780
rect 190128 110568 190340 110780
rect 195024 110638 195236 110644
rect 195024 110574 195166 110638
rect 195230 110574 195236 110638
rect 28424 110508 28500 110568
rect 190128 110508 190204 110568
rect 23392 110438 23534 110502
rect 23598 110438 23604 110502
rect 23392 110432 23604 110438
rect 21760 110372 21836 110432
rect 21760 110024 21972 110372
rect 28288 110296 28636 110508
rect 190128 110366 190340 110508
rect 195024 110502 195236 110574
rect 195024 110438 195166 110502
rect 195230 110438 195236 110502
rect 195024 110432 195236 110438
rect 195432 110638 195644 110644
rect 195432 110574 195574 110638
rect 195638 110574 195644 110638
rect 195432 110502 195644 110574
rect 195432 110438 195438 110502
rect 195502 110438 195644 110502
rect 195432 110432 195644 110438
rect 195840 110502 196052 110644
rect 195840 110438 195846 110502
rect 195910 110438 196052 110502
rect 195840 110432 196052 110438
rect 196248 110638 196460 110644
rect 196248 110574 196254 110638
rect 196318 110574 196460 110638
rect 196248 110432 196460 110574
rect 196656 110638 196868 110644
rect 196656 110574 196662 110638
rect 196726 110574 196868 110638
rect 196656 110432 196868 110574
rect 196248 110372 196324 110432
rect 190128 110302 190270 110366
rect 190334 110302 190340 110366
rect 190128 110296 190340 110302
rect 28288 110236 28364 110296
rect 190264 110236 190340 110296
rect 195976 110296 196324 110372
rect 196656 110372 196732 110432
rect 195976 110236 196052 110296
rect 22168 110230 22516 110236
rect 22168 110166 22174 110230
rect 22238 110166 22446 110230
rect 22510 110166 22516 110230
rect 22168 110160 22516 110166
rect 22168 110024 22380 110160
rect 22576 110100 22788 110236
rect 22478 110094 22788 110100
rect 22440 110030 22446 110094
rect 22510 110030 22788 110094
rect 22478 110024 22788 110030
rect 22984 110230 23196 110236
rect 22984 110166 23126 110230
rect 23190 110166 23196 110230
rect 22984 110094 23196 110166
rect 22984 110030 22990 110094
rect 23054 110030 23196 110094
rect 22984 110024 23196 110030
rect 23392 110230 23604 110236
rect 23392 110166 23534 110230
rect 23598 110166 23604 110230
rect 23392 110094 23604 110166
rect 23392 110030 23398 110094
rect 23462 110030 23604 110094
rect 23392 110024 23604 110030
rect 21760 109964 21836 110024
rect 22168 109964 22244 110024
rect 1632 109732 1844 109828
rect 1632 109692 1702 109732
rect 1224 109686 1702 109692
rect 1224 109622 1230 109686
rect 1294 109676 1702 109686
rect 1758 109676 1844 109732
rect 1294 109622 1844 109676
rect 1224 109616 1844 109622
rect 21760 109616 21972 109964
rect 22168 109888 22788 109964
rect 22168 109828 22380 109888
rect 22168 109822 22516 109828
rect 22168 109758 22446 109822
rect 22510 109758 22516 109822
rect 22168 109752 22516 109758
rect 22168 109616 22380 109752
rect 22576 109686 22788 109888
rect 22576 109622 22582 109686
rect 22646 109622 22788 109686
rect 22576 109616 22788 109622
rect 22984 109822 23196 109828
rect 22984 109758 22990 109822
rect 23054 109758 23196 109822
rect 22984 109686 23196 109758
rect 22984 109622 22990 109686
rect 23054 109622 23196 109686
rect 22984 109616 23196 109622
rect 23392 109822 23604 109828
rect 23392 109758 23398 109822
rect 23462 109758 23604 109822
rect 23392 109686 23604 109758
rect 23392 109622 23534 109686
rect 23598 109622 23604 109686
rect 23392 109616 23604 109622
rect 28288 109752 28636 110236
rect 190128 110094 190340 110236
rect 190128 110030 190134 110094
rect 190198 110030 190270 110094
rect 190334 110030 190340 110094
rect 190128 109752 190340 110030
rect 195024 110230 195236 110236
rect 195024 110166 195166 110230
rect 195230 110166 195236 110230
rect 195024 110094 195236 110166
rect 195024 110030 195030 110094
rect 195094 110030 195236 110094
rect 195024 110024 195236 110030
rect 195432 110230 195644 110236
rect 195432 110166 195438 110230
rect 195502 110166 195644 110230
rect 195432 110094 195644 110166
rect 195432 110030 195574 110094
rect 195638 110030 195644 110094
rect 195432 110024 195644 110030
rect 195840 110230 196460 110236
rect 195840 110166 195846 110230
rect 195910 110166 196460 110230
rect 195840 110160 196460 110166
rect 195840 110100 196052 110160
rect 195840 110024 196188 110100
rect 196248 110024 196460 110160
rect 196656 110024 196868 110372
rect 195840 109964 195916 110024
rect 196112 109964 196188 110024
rect 196792 109964 196868 110024
rect 195024 109822 195236 109828
rect 195024 109758 195030 109822
rect 195094 109758 195236 109822
rect 28288 109692 28364 109752
rect 21760 109556 21836 109616
rect 21760 109414 21972 109556
rect 28288 109480 28636 109692
rect 190128 109686 190340 109692
rect 190128 109622 190134 109686
rect 190198 109622 190340 109686
rect 190128 109550 190340 109622
rect 195024 109686 195236 109758
rect 195024 109622 195166 109686
rect 195230 109622 195236 109686
rect 195024 109616 195236 109622
rect 195432 109822 195644 109828
rect 195432 109758 195574 109822
rect 195638 109758 195644 109822
rect 195432 109686 195644 109758
rect 195432 109622 195574 109686
rect 195638 109622 195644 109686
rect 195432 109616 195644 109622
rect 195840 109692 196052 109964
rect 196112 109888 196460 109964
rect 195840 109686 196188 109692
rect 195840 109622 196118 109686
rect 196182 109622 196188 109686
rect 195840 109616 196188 109622
rect 196248 109616 196460 109888
rect 196656 109616 196868 109964
rect 216784 109822 217540 109828
rect 216784 109758 217470 109822
rect 217534 109758 217540 109822
rect 216784 109752 217540 109758
rect 216784 109732 216996 109752
rect 216784 109676 216908 109732
rect 216964 109676 216996 109732
rect 216784 109616 216996 109676
rect 190128 109486 190270 109550
rect 190334 109486 190340 109550
rect 190128 109480 190340 109486
rect 196656 109556 196732 109616
rect 28288 109420 28364 109480
rect 190128 109420 190204 109480
rect 21760 109350 21766 109414
rect 21830 109350 21972 109414
rect 21760 109344 21972 109350
rect 22168 109208 22380 109420
rect 22576 109414 22788 109420
rect 22576 109350 22582 109414
rect 22646 109350 22788 109414
rect 22576 109284 22788 109350
rect 22304 109148 22380 109208
rect 22440 109208 22788 109284
rect 22984 109414 23196 109420
rect 22984 109350 22990 109414
rect 23054 109350 23196 109414
rect 22984 109208 23196 109350
rect 23392 109414 23604 109420
rect 23392 109350 23534 109414
rect 23598 109350 23604 109414
rect 23392 109208 23604 109350
rect 22440 109148 22516 109208
rect 22984 109148 23060 109208
rect 23528 109148 23604 109208
rect 21760 109142 21972 109148
rect 21760 109078 21766 109142
rect 21830 109078 21972 109142
rect 21760 109006 21972 109078
rect 21760 108942 21766 109006
rect 21830 108942 21972 109006
rect 21760 108936 21972 108942
rect 22168 109072 22516 109148
rect 22168 109012 22380 109072
rect 22168 109006 22516 109012
rect 22168 108942 22446 109006
rect 22510 108942 22516 109006
rect 22168 108936 22516 108942
rect 22576 108936 22788 109148
rect 22304 108876 22380 108936
rect 22576 108876 22652 108936
rect 22304 108800 22652 108876
rect 22984 108800 23196 109148
rect 23120 108740 23196 108800
rect 21760 108734 21972 108740
rect 21760 108670 21766 108734
rect 21830 108670 21972 108734
rect 21760 108598 21972 108670
rect 21760 108534 21766 108598
rect 21830 108534 21972 108598
rect 21760 108528 21972 108534
rect 22168 108392 22380 108740
rect 22478 108734 22788 108740
rect 22440 108670 22446 108734
rect 22510 108670 22788 108734
rect 22478 108664 22788 108670
rect 22576 108392 22788 108664
rect 22984 108392 23196 108740
rect 23392 108800 23604 109148
rect 28288 109142 28636 109420
rect 28288 109078 28430 109142
rect 28494 109078 28636 109142
rect 28288 109072 28636 109078
rect 190128 109278 190340 109420
rect 190128 109214 190270 109278
rect 190334 109214 190340 109278
rect 190128 109142 190340 109214
rect 190128 109078 190270 109142
rect 190334 109078 190340 109142
rect 190128 109072 190340 109078
rect 195024 109414 195236 109420
rect 195024 109350 195166 109414
rect 195230 109350 195236 109414
rect 195024 109208 195236 109350
rect 195432 109414 195644 109420
rect 195432 109350 195574 109414
rect 195638 109350 195644 109414
rect 195432 109208 195644 109350
rect 195840 109284 196052 109420
rect 196150 109414 196460 109420
rect 196112 109350 196118 109414
rect 196182 109350 196460 109414
rect 196150 109344 196460 109350
rect 196656 109414 196868 109556
rect 196656 109350 196798 109414
rect 196862 109350 196868 109414
rect 196656 109344 196868 109350
rect 195840 109208 196188 109284
rect 195024 109148 195100 109208
rect 195432 109148 195508 109208
rect 195976 109148 196052 109208
rect 28288 108870 28636 108876
rect 28288 108806 28430 108870
rect 28494 108806 28636 108870
rect 23392 108740 23468 108800
rect 23392 108392 23604 108740
rect 28288 108734 28636 108806
rect 28288 108670 28294 108734
rect 28358 108670 28636 108734
rect 28288 108664 28636 108670
rect 190128 108870 190340 108876
rect 190128 108806 190270 108870
rect 190334 108806 190340 108870
rect 190128 108734 190340 108806
rect 195024 108800 195236 109148
rect 195160 108740 195236 108800
rect 190128 108670 190134 108734
rect 190198 108670 190340 108734
rect 28404 108468 28502 108664
rect 22168 108332 22244 108392
rect 22576 108332 22652 108392
rect 23120 108332 23196 108392
rect 23528 108332 23604 108392
rect 21760 108326 21972 108332
rect 21760 108262 21766 108326
rect 21830 108262 21972 108326
rect 1224 108190 1844 108196
rect 1224 108126 1230 108190
rect 1294 108126 1844 108190
rect 1224 108120 1844 108126
rect 21760 108190 21972 108262
rect 21760 108126 21902 108190
rect 21966 108126 21972 108190
rect 21760 108120 21972 108126
rect 22168 108256 22788 108332
rect 22168 108120 22380 108256
rect 22576 108190 22788 108256
rect 22576 108126 22718 108190
rect 22782 108126 22788 108190
rect 22576 108120 22788 108126
rect 22984 108190 23196 108332
rect 22984 108126 23126 108190
rect 23190 108126 23196 108190
rect 22984 108120 23196 108126
rect 23392 108190 23604 108332
rect 23392 108126 23398 108190
rect 23462 108126 23604 108190
rect 23392 108120 23604 108126
rect 28288 108462 28636 108468
rect 28288 108398 28294 108462
rect 28358 108398 28636 108462
rect 28288 108256 28636 108398
rect 190128 108462 190340 108670
rect 190128 108398 190134 108462
rect 190198 108398 190340 108462
rect 190128 108326 190340 108398
rect 195024 108392 195236 108740
rect 195432 108800 195644 109148
rect 195840 108936 196052 109148
rect 196112 109148 196188 109208
rect 196248 109208 196460 109344
rect 196248 109148 196324 109208
rect 196112 109072 196460 109148
rect 196248 109012 196460 109072
rect 196150 109006 196460 109012
rect 196112 108942 196118 109006
rect 196182 108942 196460 109006
rect 196150 108936 196460 108942
rect 196656 109142 196868 109148
rect 196656 109078 196798 109142
rect 196862 109078 196868 109142
rect 196656 109006 196868 109078
rect 196656 108942 196798 109006
rect 196862 108942 196868 109006
rect 196656 108936 196868 108942
rect 195432 108740 195508 108800
rect 195432 108392 195644 108740
rect 195840 108734 196188 108740
rect 195840 108670 196118 108734
rect 196182 108670 196188 108734
rect 195840 108664 196188 108670
rect 195840 108468 196052 108664
rect 196248 108468 196460 108740
rect 196656 108734 196868 108740
rect 196656 108670 196798 108734
rect 196862 108670 196868 108734
rect 196656 108598 196868 108670
rect 196656 108534 196662 108598
rect 196726 108534 196868 108598
rect 196656 108528 196868 108534
rect 195840 108462 196460 108468
rect 195840 108398 196254 108462
rect 196318 108398 196460 108462
rect 195840 108392 196460 108398
rect 195160 108332 195236 108392
rect 195568 108332 195644 108392
rect 196248 108332 196324 108392
rect 190128 108262 190134 108326
rect 190198 108262 190340 108326
rect 190128 108256 190340 108262
rect 28288 108196 28364 108256
rect 1632 108052 1844 108120
rect 1632 107996 1702 108052
rect 1758 107996 1844 108052
rect 1632 107848 1844 107996
rect 21760 107918 21972 107924
rect 21760 107854 21902 107918
rect 21966 107854 21972 107918
rect 21760 107782 21972 107854
rect 21760 107718 21902 107782
rect 21966 107718 21972 107782
rect 21760 107712 21972 107718
rect 22168 107918 22788 107924
rect 22168 107854 22718 107918
rect 22782 107854 22788 107918
rect 22168 107848 22788 107854
rect 22168 107788 22380 107848
rect 22168 107782 22516 107788
rect 22168 107718 22446 107782
rect 22510 107718 22516 107782
rect 22168 107712 22516 107718
rect 22576 107712 22788 107848
rect 22984 107918 23196 107924
rect 22984 107854 23126 107918
rect 23190 107854 23196 107918
rect 22984 107782 23196 107854
rect 22984 107718 22990 107782
rect 23054 107718 23196 107782
rect 22984 107712 23196 107718
rect 23392 107918 23604 107924
rect 23392 107854 23398 107918
rect 23462 107854 23604 107918
rect 23392 107782 23604 107854
rect 23392 107718 23398 107782
rect 23462 107718 23604 107782
rect 23392 107712 23604 107718
rect 28288 107918 28636 108196
rect 28288 107854 28430 107918
rect 28494 107854 28636 107918
rect 28288 107712 28636 107854
rect 190128 107918 190340 108196
rect 195024 108190 195236 108332
rect 195024 108126 195030 108190
rect 195094 108126 195236 108190
rect 195024 108120 195236 108126
rect 195432 108190 195644 108332
rect 195432 108126 195438 108190
rect 195502 108126 195644 108190
rect 195432 108120 195644 108126
rect 195840 108326 196188 108332
rect 195840 108262 196118 108326
rect 196182 108262 196188 108326
rect 195840 108256 196188 108262
rect 195840 108120 196052 108256
rect 196248 108196 196460 108332
rect 196150 108190 196460 108196
rect 196112 108126 196118 108190
rect 196182 108126 196460 108190
rect 196150 108120 196460 108126
rect 196656 108326 196868 108332
rect 196656 108262 196662 108326
rect 196726 108262 196868 108326
rect 196656 108190 196868 108262
rect 196656 108126 196798 108190
rect 196862 108126 196868 108190
rect 196656 108120 196868 108126
rect 216784 108190 217540 108196
rect 216784 108126 217470 108190
rect 217534 108126 217540 108190
rect 216784 108120 217540 108126
rect 195976 108060 196052 108120
rect 195976 107984 196324 108060
rect 196248 107924 196324 107984
rect 216784 108052 216996 108120
rect 216784 107996 216908 108052
rect 216964 107996 216996 108052
rect 190128 107854 190134 107918
rect 190198 107854 190270 107918
rect 190334 107854 190340 107918
rect 190128 107712 190340 107854
rect 195024 107918 195236 107924
rect 195024 107854 195030 107918
rect 195094 107854 195236 107918
rect 195024 107782 195236 107854
rect 195024 107718 195166 107782
rect 195230 107718 195236 107782
rect 195024 107712 195236 107718
rect 195432 107918 195644 107924
rect 195432 107854 195438 107918
rect 195502 107854 195644 107918
rect 195432 107782 195644 107854
rect 195432 107718 195574 107782
rect 195638 107718 195644 107782
rect 195432 107712 195644 107718
rect 195840 107918 196188 107924
rect 195840 107854 196118 107918
rect 196182 107854 196188 107918
rect 195840 107848 196188 107854
rect 195840 107712 196052 107848
rect 196248 107782 196460 107924
rect 196248 107718 196390 107782
rect 196454 107718 196460 107782
rect 196248 107712 196460 107718
rect 196656 107918 196868 107924
rect 196656 107854 196798 107918
rect 196862 107854 196868 107918
rect 196656 107782 196868 107854
rect 216784 107848 216996 107996
rect 196656 107718 196798 107782
rect 196862 107718 196868 107782
rect 196656 107712 196868 107718
rect 28424 107652 28500 107712
rect 190128 107652 190204 107712
rect 28288 107646 28636 107652
rect 28288 107582 28430 107646
rect 28494 107582 28636 107646
rect 21760 107510 21972 107516
rect 21760 107446 21902 107510
rect 21966 107446 21972 107510
rect 21760 107374 21972 107446
rect 21760 107310 21902 107374
rect 21966 107310 21972 107374
rect 21760 107304 21972 107310
rect 22168 107374 22380 107516
rect 22478 107510 22788 107516
rect 22440 107446 22446 107510
rect 22510 107446 22788 107510
rect 22478 107440 22788 107446
rect 22168 107310 22174 107374
rect 22238 107310 22380 107374
rect 22168 107304 22380 107310
rect 22576 107374 22788 107440
rect 22576 107310 22582 107374
rect 22646 107310 22788 107374
rect 22576 107304 22788 107310
rect 22984 107510 23196 107516
rect 22984 107446 22990 107510
rect 23054 107446 23196 107510
rect 22984 107374 23196 107446
rect 22984 107310 22990 107374
rect 23054 107310 23196 107374
rect 22984 107304 23196 107310
rect 23392 107510 23604 107516
rect 23392 107446 23398 107510
rect 23462 107446 23604 107510
rect 23392 107374 23604 107446
rect 23392 107310 23398 107374
rect 23462 107310 23604 107374
rect 23392 107304 23604 107310
rect 28288 107440 28636 107582
rect 190128 107646 190340 107652
rect 190128 107582 190270 107646
rect 190334 107582 190340 107646
rect 190128 107440 190340 107582
rect 195024 107510 195236 107516
rect 195024 107446 195166 107510
rect 195230 107446 195236 107510
rect 28288 107380 28364 107440
rect 190128 107380 190204 107440
rect 28288 107168 28636 107380
rect 190128 107168 190340 107380
rect 195024 107374 195236 107446
rect 195024 107310 195030 107374
rect 195094 107310 195236 107374
rect 195024 107304 195236 107310
rect 195432 107510 195644 107516
rect 195432 107446 195574 107510
rect 195638 107446 195644 107510
rect 195432 107374 195644 107446
rect 195432 107310 195438 107374
rect 195502 107310 195644 107374
rect 195432 107304 195644 107310
rect 195840 107374 196052 107516
rect 195840 107310 195982 107374
rect 196046 107310 196052 107374
rect 195840 107304 196052 107310
rect 196248 107510 196460 107516
rect 196248 107446 196390 107510
rect 196454 107446 196460 107510
rect 196248 107374 196460 107446
rect 196248 107310 196254 107374
rect 196318 107310 196460 107374
rect 196248 107304 196460 107310
rect 196656 107510 196868 107516
rect 196656 107446 196798 107510
rect 196862 107446 196868 107510
rect 196656 107374 196868 107446
rect 196656 107310 196798 107374
rect 196862 107310 196868 107374
rect 196656 107304 196868 107310
rect 28560 107108 28636 107168
rect 190264 107108 190340 107168
rect 21760 107102 21972 107108
rect 21760 107038 21902 107102
rect 21966 107038 21972 107102
rect 21760 106966 21972 107038
rect 21760 106902 21902 106966
rect 21966 106902 21972 106966
rect 21760 106896 21972 106902
rect 22168 107102 22380 107108
rect 22168 107038 22174 107102
rect 22238 107038 22380 107102
rect 22168 106972 22380 107038
rect 22576 107102 22788 107108
rect 22576 107038 22582 107102
rect 22646 107038 22788 107102
rect 22576 106972 22788 107038
rect 22168 106966 22788 106972
rect 22168 106902 22310 106966
rect 22374 106902 22788 106966
rect 22168 106896 22788 106902
rect 22984 107102 23196 107108
rect 22984 107038 22990 107102
rect 23054 107038 23196 107102
rect 22984 106966 23196 107038
rect 22984 106902 23126 106966
rect 23190 106902 23196 106966
rect 22984 106896 23196 106902
rect 23392 107102 23604 107108
rect 23392 107038 23398 107102
rect 23462 107038 23604 107102
rect 23392 106966 23604 107038
rect 23392 106902 23398 106966
rect 23462 106902 23604 106966
rect 23392 106896 23604 106902
rect 28288 106896 28636 107108
rect 190128 106896 190340 107108
rect 195024 107102 195236 107108
rect 195024 107038 195030 107102
rect 195094 107038 195236 107102
rect 195024 106966 195236 107038
rect 195024 106902 195030 106966
rect 195094 106902 195236 106966
rect 195024 106896 195236 106902
rect 195432 107102 195644 107108
rect 195432 107038 195438 107102
rect 195502 107038 195644 107102
rect 195432 106966 195644 107038
rect 195432 106902 195438 106966
rect 195502 106902 195644 106966
rect 195432 106896 195644 106902
rect 195840 107102 196460 107108
rect 195840 107038 195982 107102
rect 196046 107038 196254 107102
rect 196318 107038 196460 107102
rect 195840 107032 196460 107038
rect 195840 106972 196052 107032
rect 195840 106966 196188 106972
rect 195840 106902 196118 106966
rect 196182 106902 196188 106966
rect 195840 106896 196188 106902
rect 196248 106896 196460 107032
rect 196656 107102 196868 107108
rect 196656 107038 196798 107102
rect 196862 107038 196868 107102
rect 196656 106966 196868 107038
rect 196656 106902 196798 106966
rect 196862 106902 196868 106966
rect 196656 106896 196868 106902
rect 22304 106836 22380 106896
rect 28560 106836 28636 106896
rect 190264 106836 190340 106896
rect 22304 106760 22652 106836
rect 22576 106700 22652 106760
rect 21760 106694 21972 106700
rect 21760 106630 21902 106694
rect 21966 106630 21972 106694
rect 21760 106488 21972 106630
rect 22168 106694 22380 106700
rect 22168 106630 22310 106694
rect 22374 106630 22380 106694
rect 22168 106558 22380 106630
rect 22168 106494 22174 106558
rect 22238 106494 22380 106558
rect 22168 106488 22380 106494
rect 22576 106488 22788 106700
rect 22984 106694 23196 106700
rect 22984 106630 23126 106694
rect 23190 106630 23196 106694
rect 22984 106558 23196 106630
rect 22984 106494 23126 106558
rect 23190 106494 23196 106558
rect 22984 106488 23196 106494
rect 23392 106694 23604 106700
rect 23392 106630 23398 106694
rect 23462 106630 23604 106694
rect 23392 106558 23604 106630
rect 28288 106624 28636 106836
rect 190128 106624 190340 106836
rect 28560 106564 28636 106624
rect 190264 106564 190340 106624
rect 23392 106494 23534 106558
rect 23598 106494 23604 106558
rect 23392 106488 23604 106494
rect 21760 106428 21836 106488
rect 1224 106422 1844 106428
rect 1224 106358 1230 106422
rect 1294 106372 1844 106422
rect 1294 106358 1702 106372
rect 1224 106352 1702 106358
rect 1632 106316 1702 106352
rect 1758 106316 1844 106372
rect 1632 106216 1844 106316
rect 21760 106080 21972 106428
rect 28288 106352 28636 106564
rect 190128 106352 190340 106564
rect 195024 106694 195236 106700
rect 195024 106630 195030 106694
rect 195094 106630 195236 106694
rect 195024 106558 195236 106630
rect 195024 106494 195166 106558
rect 195230 106494 195236 106558
rect 195024 106488 195236 106494
rect 195432 106694 195644 106700
rect 195432 106630 195438 106694
rect 195502 106630 195644 106694
rect 195432 106558 195644 106630
rect 195432 106494 195574 106558
rect 195638 106494 195644 106558
rect 195432 106488 195644 106494
rect 195840 106558 196052 106700
rect 196150 106694 196460 106700
rect 196112 106630 196118 106694
rect 196182 106630 196460 106694
rect 196150 106624 196460 106630
rect 195840 106494 195846 106558
rect 195910 106494 196052 106558
rect 195840 106488 196052 106494
rect 196248 106558 196460 106624
rect 196248 106494 196254 106558
rect 196318 106494 196460 106558
rect 196248 106488 196460 106494
rect 196656 106694 196868 106700
rect 196656 106630 196798 106694
rect 196862 106630 196868 106694
rect 196656 106488 196868 106630
rect 196656 106428 196732 106488
rect 28424 106292 28500 106352
rect 190128 106292 190204 106352
rect 22168 106286 22380 106292
rect 22168 106222 22174 106286
rect 22238 106222 22380 106286
rect 22168 106080 22380 106222
rect 22576 106156 22788 106292
rect 21760 106020 21836 106080
rect 22304 106020 22380 106080
rect 22440 106080 22788 106156
rect 22984 106286 23196 106292
rect 22984 106222 23126 106286
rect 23190 106222 23196 106286
rect 22984 106150 23196 106222
rect 22984 106086 23126 106150
rect 23190 106086 23196 106150
rect 22984 106080 23196 106086
rect 23392 106286 23604 106292
rect 23392 106222 23534 106286
rect 23598 106222 23604 106286
rect 23392 106150 23604 106222
rect 23392 106086 23534 106150
rect 23598 106086 23604 106150
rect 23392 106080 23604 106086
rect 28288 106080 28636 106292
rect 190128 106080 190340 106292
rect 195024 106286 195236 106292
rect 195024 106222 195166 106286
rect 195230 106222 195236 106286
rect 195024 106150 195236 106222
rect 195024 106086 195166 106150
rect 195230 106086 195236 106150
rect 195024 106080 195236 106086
rect 195432 106286 195644 106292
rect 195432 106222 195574 106286
rect 195638 106222 195644 106286
rect 195432 106150 195644 106222
rect 195432 106086 195574 106150
rect 195638 106086 195644 106150
rect 195432 106080 195644 106086
rect 195840 106286 196052 106292
rect 195840 106222 195846 106286
rect 195910 106222 196052 106286
rect 195840 106080 196052 106222
rect 196248 106286 196460 106292
rect 196248 106222 196254 106286
rect 196318 106222 196460 106286
rect 196248 106156 196460 106222
rect 196112 106080 196460 106156
rect 196656 106080 196868 106428
rect 216784 106372 216996 106428
rect 216784 106316 216908 106372
rect 216964 106316 216996 106372
rect 216784 106292 216996 106316
rect 216784 106286 217540 106292
rect 216784 106222 217470 106286
rect 217534 106222 217540 106286
rect 216784 106216 217540 106222
rect 22440 106020 22516 106080
rect 28424 106020 28500 106080
rect 190128 106020 190204 106080
rect 195840 106020 195916 106080
rect 196112 106020 196188 106080
rect 196792 106020 196868 106080
rect 21760 105672 21972 106020
rect 22168 105944 22516 106020
rect 22576 105944 22788 106020
rect 22168 105748 22380 105944
rect 22688 105748 22788 105944
rect 22168 105742 22788 105748
rect 22168 105678 22174 105742
rect 22238 105678 22582 105742
rect 22646 105678 22788 105742
rect 22168 105672 22788 105678
rect 22984 105878 23196 105884
rect 22984 105814 23126 105878
rect 23190 105814 23196 105878
rect 22984 105742 23196 105814
rect 22984 105678 23126 105742
rect 23190 105678 23196 105742
rect 22984 105672 23196 105678
rect 23392 105878 23604 105884
rect 23392 105814 23534 105878
rect 23598 105814 23604 105878
rect 23392 105742 23604 105814
rect 23392 105678 23534 105742
rect 23598 105678 23604 105742
rect 23392 105672 23604 105678
rect 28288 105808 28636 106020
rect 190128 105808 190340 106020
rect 195840 105944 196188 106020
rect 28288 105748 28364 105808
rect 190264 105748 190340 105808
rect 21896 105612 21972 105672
rect 21760 105470 21972 105612
rect 28288 105606 28636 105748
rect 28288 105542 28566 105606
rect 28630 105542 28636 105606
rect 28288 105536 28636 105542
rect 190128 105606 190340 105748
rect 195024 105878 195236 105884
rect 195024 105814 195166 105878
rect 195230 105814 195236 105878
rect 195024 105742 195236 105814
rect 195024 105678 195166 105742
rect 195230 105678 195236 105742
rect 195024 105672 195236 105678
rect 195432 105878 195644 105884
rect 195432 105814 195574 105878
rect 195638 105814 195644 105878
rect 195432 105742 195644 105814
rect 195432 105678 195438 105742
rect 195502 105678 195644 105742
rect 195432 105672 195644 105678
rect 195840 105748 196052 105944
rect 196248 105748 196460 106020
rect 195840 105742 196460 105748
rect 195840 105678 196254 105742
rect 196318 105678 196460 105742
rect 195840 105672 196460 105678
rect 196656 105672 196868 106020
rect 196792 105612 196868 105672
rect 190128 105542 190270 105606
rect 190334 105542 190340 105606
rect 190128 105536 190340 105542
rect 28288 105476 28364 105536
rect 190264 105476 190340 105536
rect 21760 105406 21766 105470
rect 21830 105406 21972 105470
rect 21760 105400 21972 105406
rect 22168 105470 22380 105476
rect 22168 105406 22174 105470
rect 22238 105406 22380 105470
rect 22168 105264 22380 105406
rect 22576 105470 22788 105476
rect 22576 105406 22582 105470
rect 22646 105406 22788 105470
rect 22576 105264 22788 105406
rect 22984 105470 23196 105476
rect 22984 105406 23126 105470
rect 23190 105406 23196 105470
rect 22984 105264 23196 105406
rect 23392 105470 23604 105476
rect 23392 105406 23534 105470
rect 23598 105406 23604 105470
rect 23392 105264 23604 105406
rect 22168 105204 22244 105264
rect 22576 105204 22652 105264
rect 22984 105204 23060 105264
rect 23528 105204 23604 105264
rect 21760 105198 21972 105204
rect 21760 105134 21766 105198
rect 21830 105134 21972 105198
rect 21760 105062 21972 105134
rect 21760 104998 21766 105062
rect 21830 104998 21972 105062
rect 21760 104992 21972 104998
rect 22168 104992 22380 105204
rect 22576 105068 22788 105204
rect 22478 105062 22788 105068
rect 22440 104998 22446 105062
rect 22510 104998 22582 105062
rect 22646 104998 22788 105062
rect 22478 104992 22788 104998
rect 22984 104856 23196 105204
rect 23120 104796 23196 104856
rect 1224 104790 1844 104796
rect 1224 104726 1230 104790
rect 1294 104726 1844 104790
rect 1224 104720 1844 104726
rect 1632 104692 1844 104720
rect 1632 104636 1702 104692
rect 1758 104636 1844 104692
rect 1632 104584 1844 104636
rect 21760 104790 21972 104796
rect 21760 104726 21766 104790
rect 21830 104726 21972 104790
rect 21760 104654 21972 104726
rect 21760 104590 21766 104654
rect 21830 104590 21972 104654
rect 21760 104584 21972 104590
rect 22168 104790 22516 104796
rect 22168 104726 22446 104790
rect 22510 104726 22516 104790
rect 22168 104720 22516 104726
rect 22576 104790 22788 104796
rect 22576 104726 22582 104790
rect 22646 104726 22788 104790
rect 22168 104448 22380 104720
rect 22576 104448 22788 104726
rect 22984 104448 23196 104796
rect 23392 104856 23604 105204
rect 28288 105334 28636 105476
rect 28288 105270 28566 105334
rect 28630 105270 28636 105334
rect 28288 105198 28636 105270
rect 28288 105134 28430 105198
rect 28494 105134 28636 105198
rect 28288 105128 28636 105134
rect 190128 105334 190340 105476
rect 190128 105270 190270 105334
rect 190334 105270 190340 105334
rect 190128 105198 190340 105270
rect 195024 105470 195236 105476
rect 195024 105406 195166 105470
rect 195230 105406 195236 105470
rect 195024 105264 195236 105406
rect 195432 105470 195644 105476
rect 195432 105406 195438 105470
rect 195502 105406 195644 105470
rect 195432 105264 195644 105406
rect 195160 105204 195236 105264
rect 195568 105204 195644 105264
rect 190128 105134 190270 105198
rect 190334 105134 190340 105198
rect 190128 105128 190340 105134
rect 28288 104926 28636 104932
rect 28288 104862 28430 104926
rect 28494 104862 28636 104926
rect 23392 104796 23468 104856
rect 23392 104448 23604 104796
rect 22168 104388 22244 104448
rect 22576 104388 22652 104448
rect 23120 104388 23196 104448
rect 23528 104388 23604 104448
rect 21760 104382 21972 104388
rect 21760 104318 21766 104382
rect 21830 104318 21972 104382
rect 21760 104246 21972 104318
rect 21760 104182 21766 104246
rect 21830 104182 21972 104246
rect 21760 104176 21972 104182
rect 22168 104176 22380 104388
rect 22576 104246 22788 104388
rect 22576 104182 22582 104246
rect 22646 104182 22788 104246
rect 22576 104176 22788 104182
rect 22984 104246 23196 104388
rect 22984 104182 22990 104246
rect 23054 104182 23196 104246
rect 22984 104176 23196 104182
rect 23392 104246 23604 104388
rect 28288 104312 28636 104862
rect 190128 104926 190340 104932
rect 190128 104862 190270 104926
rect 190334 104862 190340 104926
rect 190128 104518 190340 104862
rect 190128 104454 190270 104518
rect 190334 104454 190340 104518
rect 190128 104312 190340 104454
rect 195024 104856 195236 105204
rect 195432 104856 195644 105204
rect 195840 105264 196052 105476
rect 196248 105470 196460 105476
rect 196248 105406 196254 105470
rect 196318 105406 196460 105470
rect 196248 105264 196460 105406
rect 196656 105470 196868 105612
rect 196656 105406 196662 105470
rect 196726 105406 196868 105470
rect 196656 105400 196868 105406
rect 195840 105204 195916 105264
rect 196248 105204 196324 105264
rect 195840 105062 196052 105204
rect 196248 105068 196460 105204
rect 196150 105062 196460 105068
rect 195840 104998 195846 105062
rect 195910 104998 196052 105062
rect 196112 104998 196118 105062
rect 196182 104998 196460 105062
rect 195840 104992 196052 104998
rect 196150 104992 196460 104998
rect 196656 105198 196868 105204
rect 196656 105134 196662 105198
rect 196726 105134 196868 105198
rect 196656 105062 196868 105134
rect 196656 104998 196798 105062
rect 196862 104998 196868 105062
rect 196656 104992 196868 104998
rect 195024 104796 195100 104856
rect 195432 104796 195508 104856
rect 195024 104448 195236 104796
rect 195432 104448 195644 104796
rect 195160 104388 195236 104448
rect 195568 104388 195644 104448
rect 28424 104252 28500 104312
rect 190264 104252 190340 104312
rect 23392 104182 23534 104246
rect 23598 104182 23604 104246
rect 23392 104176 23604 104182
rect 21760 103974 21972 103980
rect 21760 103910 21766 103974
rect 21830 103910 21972 103974
rect 21760 103838 21972 103910
rect 21760 103774 21902 103838
rect 21966 103774 21972 103838
rect 21760 103768 21972 103774
rect 22168 103844 22380 103980
rect 22576 103974 22788 103980
rect 22576 103910 22582 103974
rect 22646 103910 22788 103974
rect 22576 103844 22788 103910
rect 22168 103768 22788 103844
rect 22984 103974 23196 103980
rect 22984 103910 22990 103974
rect 23054 103910 23196 103974
rect 22984 103838 23196 103910
rect 22984 103774 22990 103838
rect 23054 103774 23196 103838
rect 22984 103768 23196 103774
rect 23392 103974 23604 103980
rect 23392 103910 23534 103974
rect 23598 103910 23604 103974
rect 23392 103838 23604 103910
rect 23392 103774 23398 103838
rect 23462 103774 23604 103838
rect 23392 103768 23604 103774
rect 28288 103768 28636 104252
rect 190128 104246 190340 104252
rect 190128 104182 190270 104246
rect 190334 104182 190340 104246
rect 190128 103768 190340 104182
rect 195024 104246 195236 104388
rect 195024 104182 195166 104246
rect 195230 104182 195236 104246
rect 195024 104176 195236 104182
rect 195432 104246 195644 104388
rect 195432 104182 195574 104246
rect 195638 104182 195644 104246
rect 195432 104176 195644 104182
rect 195840 104790 196188 104796
rect 195840 104726 195846 104790
rect 195910 104726 196118 104790
rect 196182 104726 196188 104790
rect 195840 104720 196188 104726
rect 195840 104524 196052 104720
rect 196248 104524 196460 104796
rect 196656 104790 196868 104796
rect 196656 104726 196798 104790
rect 196862 104726 196868 104790
rect 196656 104654 196868 104726
rect 196656 104590 196662 104654
rect 196726 104590 196868 104654
rect 196656 104584 196868 104590
rect 216784 104692 216996 104796
rect 216784 104636 216908 104692
rect 216964 104660 216996 104692
rect 216964 104654 217540 104660
rect 216964 104636 217470 104654
rect 216784 104590 217470 104636
rect 217534 104590 217540 104654
rect 216784 104584 217540 104590
rect 195840 104448 196460 104524
rect 195840 104388 195916 104448
rect 196248 104388 196324 104448
rect 195840 104246 196052 104388
rect 195840 104182 195846 104246
rect 195910 104182 196052 104246
rect 195840 104176 196052 104182
rect 196248 104176 196460 104388
rect 196656 104382 196868 104388
rect 196656 104318 196662 104382
rect 196726 104318 196868 104382
rect 196656 104246 196868 104318
rect 196656 104182 196662 104246
rect 196726 104182 196868 104246
rect 196656 104176 196868 104182
rect 195024 103974 195236 103980
rect 195024 103910 195166 103974
rect 195230 103910 195236 103974
rect 195024 103838 195236 103910
rect 195024 103774 195030 103838
rect 195094 103774 195236 103838
rect 195024 103768 195236 103774
rect 195432 103974 195644 103980
rect 195432 103910 195574 103974
rect 195638 103910 195644 103974
rect 195432 103838 195644 103910
rect 195432 103774 195438 103838
rect 195502 103774 195644 103838
rect 195432 103768 195644 103774
rect 195840 103974 196052 103980
rect 195840 103910 195846 103974
rect 195910 103910 196052 103974
rect 195840 103844 196052 103910
rect 196248 103844 196460 103980
rect 195840 103768 196460 103844
rect 196656 103974 196868 103980
rect 196656 103910 196662 103974
rect 196726 103910 196868 103974
rect 196656 103838 196868 103910
rect 196656 103774 196798 103838
rect 196862 103774 196868 103838
rect 196656 103768 196868 103774
rect 22304 103708 22380 103768
rect 28288 103708 28364 103768
rect 190264 103708 190340 103768
rect 22304 103632 22652 103708
rect 22576 103572 22652 103632
rect 21760 103566 21972 103572
rect 21760 103502 21902 103566
rect 21966 103502 21972 103566
rect 21760 103430 21972 103502
rect 21760 103366 21766 103430
rect 21830 103366 21972 103430
rect 21760 103360 21972 103366
rect 22168 103496 22788 103572
rect 22168 103436 22380 103496
rect 22168 103430 22516 103436
rect 22168 103366 22446 103430
rect 22510 103366 22516 103430
rect 22168 103360 22516 103366
rect 22576 103360 22788 103496
rect 22984 103566 23196 103572
rect 22984 103502 22990 103566
rect 23054 103502 23196 103566
rect 22984 103430 23196 103502
rect 22984 103366 23126 103430
rect 23190 103366 23196 103430
rect 22984 103360 23196 103366
rect 23392 103566 23604 103572
rect 23392 103502 23398 103566
rect 23462 103502 23604 103566
rect 23392 103430 23604 103502
rect 28288 103496 28636 103708
rect 190128 103496 190340 103708
rect 195976 103708 196052 103768
rect 195976 103632 196324 103708
rect 196248 103572 196324 103632
rect 28424 103436 28500 103496
rect 190264 103436 190340 103496
rect 23392 103366 23398 103430
rect 23462 103366 23604 103430
rect 23392 103360 23604 103366
rect 28288 103224 28636 103436
rect 190128 103224 190340 103436
rect 195024 103566 195236 103572
rect 195024 103502 195030 103566
rect 195094 103502 195236 103566
rect 195024 103430 195236 103502
rect 195024 103366 195166 103430
rect 195230 103366 195236 103430
rect 195024 103360 195236 103366
rect 195432 103566 195644 103572
rect 195432 103502 195438 103566
rect 195502 103502 195644 103566
rect 195432 103430 195644 103502
rect 195432 103366 195574 103430
rect 195638 103366 195644 103430
rect 195432 103360 195644 103366
rect 195840 103496 196460 103572
rect 195840 103430 196052 103496
rect 195840 103366 195846 103430
rect 195910 103366 196052 103430
rect 195840 103360 196052 103366
rect 196248 103360 196460 103496
rect 196656 103566 196868 103572
rect 196656 103502 196798 103566
rect 196862 103502 196868 103566
rect 196656 103430 196868 103502
rect 196656 103366 196798 103430
rect 196862 103366 196868 103430
rect 196656 103360 196868 103366
rect 28288 103164 28364 103224
rect 190128 103164 190204 103224
rect 1224 103158 1844 103164
rect 1224 103094 1230 103158
rect 1294 103094 1844 103158
rect 1224 103088 1844 103094
rect 1632 103012 1844 103088
rect 1632 102956 1702 103012
rect 1758 102956 1844 103012
rect 1632 102816 1844 102956
rect 21760 103158 21972 103164
rect 21760 103094 21766 103158
rect 21830 103094 21972 103158
rect 21760 103022 21972 103094
rect 21760 102958 21902 103022
rect 21966 102958 21972 103022
rect 21760 102952 21972 102958
rect 22168 103022 22380 103164
rect 22478 103158 22788 103164
rect 22440 103094 22446 103158
rect 22510 103094 22788 103158
rect 22478 103088 22788 103094
rect 22168 102958 22310 103022
rect 22374 102958 22380 103022
rect 22168 102952 22380 102958
rect 22576 103022 22788 103088
rect 22576 102958 22718 103022
rect 22782 102958 22788 103022
rect 22576 102952 22788 102958
rect 22984 103158 23196 103164
rect 22984 103094 23126 103158
rect 23190 103094 23196 103158
rect 22984 103022 23196 103094
rect 22984 102958 22990 103022
rect 23054 102958 23196 103022
rect 22984 102952 23196 102958
rect 23392 103158 23604 103164
rect 23392 103094 23398 103158
rect 23462 103094 23604 103158
rect 23392 103022 23604 103094
rect 23392 102958 23398 103022
rect 23462 102958 23604 103022
rect 23392 102952 23604 102958
rect 28288 102952 28636 103164
rect 28560 102892 28636 102952
rect 21760 102750 21972 102756
rect 21760 102686 21902 102750
rect 21966 102686 21972 102750
rect 21760 102544 21972 102686
rect 22168 102750 22380 102756
rect 22168 102686 22310 102750
rect 22374 102686 22380 102750
rect 22168 102620 22380 102686
rect 22576 102750 22788 102756
rect 22576 102686 22718 102750
rect 22782 102686 22788 102750
rect 22168 102614 22516 102620
rect 22168 102550 22446 102614
rect 22510 102550 22516 102614
rect 22168 102544 22516 102550
rect 22576 102544 22788 102686
rect 22984 102750 23196 102756
rect 22984 102686 22990 102750
rect 23054 102686 23196 102750
rect 22984 102614 23196 102686
rect 22984 102550 22990 102614
rect 23054 102550 23196 102614
rect 22984 102544 23196 102550
rect 23392 102750 23604 102756
rect 23392 102686 23398 102750
rect 23462 102686 23604 102750
rect 23392 102614 23604 102686
rect 28288 102680 28636 102892
rect 190128 102952 190340 103164
rect 195024 103158 195236 103164
rect 195024 103094 195166 103158
rect 195230 103094 195236 103158
rect 195024 103022 195236 103094
rect 195024 102958 195166 103022
rect 195230 102958 195236 103022
rect 195024 102952 195236 102958
rect 195432 103158 195644 103164
rect 195432 103094 195574 103158
rect 195638 103094 195644 103158
rect 195432 103022 195644 103094
rect 195432 102958 195438 103022
rect 195502 102958 195644 103022
rect 195432 102952 195644 102958
rect 195840 103158 196460 103164
rect 195840 103094 195846 103158
rect 195910 103094 196460 103158
rect 195840 103088 196460 103094
rect 195840 102952 196052 103088
rect 196248 102952 196460 103088
rect 196656 103158 196868 103164
rect 196656 103094 196798 103158
rect 196862 103094 196868 103158
rect 196656 103022 196868 103094
rect 196656 102958 196798 103022
rect 196862 102958 196868 103022
rect 196656 102952 196868 102958
rect 216784 103028 216996 103164
rect 216784 103022 217540 103028
rect 216784 103012 217470 103022
rect 216784 102956 216908 103012
rect 216964 102958 217470 103012
rect 217534 102958 217540 103022
rect 216964 102956 217540 102958
rect 216784 102952 217540 102956
rect 190128 102892 190204 102952
rect 196248 102892 196324 102952
rect 190128 102680 190340 102892
rect 195976 102816 196324 102892
rect 216784 102816 216996 102952
rect 195976 102756 196052 102816
rect 28424 102620 28500 102680
rect 190264 102620 190340 102680
rect 23392 102550 23398 102614
rect 23462 102550 23604 102614
rect 23392 102544 23604 102550
rect 21896 102484 21972 102544
rect 22576 102484 22652 102544
rect 21760 102206 21972 102484
rect 22304 102408 22652 102484
rect 28288 102408 28636 102620
rect 190128 102408 190340 102620
rect 195024 102750 195236 102756
rect 195024 102686 195166 102750
rect 195230 102686 195236 102750
rect 195024 102614 195236 102686
rect 195024 102550 195030 102614
rect 195094 102550 195236 102614
rect 195024 102544 195236 102550
rect 195432 102750 195644 102756
rect 195432 102686 195438 102750
rect 195502 102686 195644 102750
rect 195432 102614 195644 102686
rect 195432 102550 195574 102614
rect 195638 102550 195644 102614
rect 195432 102544 195644 102550
rect 195840 102680 196460 102756
rect 195840 102614 196052 102680
rect 195840 102550 195982 102614
rect 196046 102550 196052 102614
rect 195840 102544 196052 102550
rect 196248 102614 196460 102680
rect 196248 102550 196390 102614
rect 196454 102550 196460 102614
rect 196248 102544 196460 102550
rect 196656 102750 196868 102756
rect 196656 102686 196798 102750
rect 196862 102686 196868 102750
rect 196656 102544 196868 102686
rect 196792 102484 196868 102544
rect 22304 102348 22380 102408
rect 28560 102348 28636 102408
rect 190264 102348 190340 102408
rect 21760 102142 21902 102206
rect 21966 102142 21972 102206
rect 21760 102136 21972 102142
rect 22168 102212 22380 102348
rect 22478 102342 22788 102348
rect 22440 102278 22446 102342
rect 22510 102278 22788 102342
rect 22478 102272 22788 102278
rect 22576 102212 22788 102272
rect 22168 102136 22788 102212
rect 22984 102342 23196 102348
rect 22984 102278 22990 102342
rect 23054 102278 23196 102342
rect 22984 102206 23196 102278
rect 22984 102142 23126 102206
rect 23190 102142 23196 102206
rect 22984 102136 23196 102142
rect 23392 102342 23604 102348
rect 23392 102278 23398 102342
rect 23462 102278 23604 102342
rect 23392 102206 23604 102278
rect 23392 102142 23534 102206
rect 23598 102142 23604 102206
rect 23392 102136 23604 102142
rect 28288 102136 28636 102348
rect 190128 102136 190340 102348
rect 195024 102342 195236 102348
rect 195024 102278 195030 102342
rect 195094 102278 195236 102342
rect 195024 102206 195236 102278
rect 195024 102142 195166 102206
rect 195230 102142 195236 102206
rect 195024 102136 195236 102142
rect 195432 102342 195644 102348
rect 195432 102278 195574 102342
rect 195638 102278 195644 102342
rect 195432 102206 195644 102278
rect 195432 102142 195438 102206
rect 195502 102142 195644 102206
rect 195432 102136 195644 102142
rect 195840 102342 196052 102348
rect 195840 102278 195982 102342
rect 196046 102278 196052 102342
rect 195840 102212 196052 102278
rect 196248 102342 196460 102348
rect 196248 102278 196390 102342
rect 196454 102278 196460 102342
rect 195840 102206 196188 102212
rect 195840 102142 196118 102206
rect 196182 102142 196188 102206
rect 195840 102136 196188 102142
rect 196248 102136 196460 102278
rect 196656 102206 196868 102484
rect 196656 102142 196662 102206
rect 196726 102142 196868 102206
rect 196656 102136 196868 102142
rect 22576 102076 22652 102136
rect 22440 102000 22652 102076
rect 28288 102076 28364 102136
rect 190128 102076 190204 102136
rect 22440 101940 22516 102000
rect 21760 101934 21972 101940
rect 21760 101870 21902 101934
rect 21966 101870 21972 101934
rect 21760 101728 21972 101870
rect 22168 101864 22516 101940
rect 22168 101798 22380 101864
rect 22576 101804 22788 101940
rect 22478 101798 22788 101804
rect 22168 101734 22310 101798
rect 22374 101734 22380 101798
rect 22440 101734 22446 101798
rect 22510 101734 22788 101798
rect 22168 101728 22380 101734
rect 22478 101728 22788 101734
rect 22984 101934 23196 101940
rect 22984 101870 23126 101934
rect 23190 101870 23196 101934
rect 22984 101798 23196 101870
rect 22984 101734 23126 101798
rect 23190 101734 23196 101798
rect 22984 101728 23196 101734
rect 23392 101934 23604 101940
rect 23392 101870 23534 101934
rect 23598 101870 23604 101934
rect 23392 101798 23604 101870
rect 28288 101864 28636 102076
rect 190128 101864 190340 102076
rect 195024 101934 195236 101940
rect 195024 101870 195166 101934
rect 195230 101870 195236 101934
rect 28424 101804 28500 101864
rect 190128 101804 190204 101864
rect 23392 101734 23534 101798
rect 23598 101734 23604 101798
rect 23392 101728 23604 101734
rect 21896 101668 21972 101728
rect 21760 101526 21972 101668
rect 22304 101592 22652 101668
rect 28288 101662 28636 101804
rect 28288 101598 28430 101662
rect 28494 101598 28636 101662
rect 28288 101592 28636 101598
rect 190128 101592 190340 101804
rect 195024 101798 195236 101870
rect 195024 101734 195030 101798
rect 195094 101734 195236 101798
rect 195024 101728 195236 101734
rect 195432 101934 195644 101940
rect 195432 101870 195438 101934
rect 195502 101870 195644 101934
rect 195432 101798 195644 101870
rect 195432 101734 195438 101798
rect 195502 101734 195644 101798
rect 195432 101728 195644 101734
rect 195840 101798 196052 101940
rect 196150 101934 196460 101940
rect 196112 101870 196118 101934
rect 196182 101870 196460 101934
rect 196150 101864 196460 101870
rect 195840 101734 195846 101798
rect 195910 101734 196052 101798
rect 195840 101728 196052 101734
rect 196248 101728 196460 101864
rect 196656 101934 196868 101940
rect 196656 101870 196662 101934
rect 196726 101870 196868 101934
rect 196656 101728 196868 101870
rect 196248 101668 196324 101728
rect 22304 101532 22380 101592
rect 22576 101532 22652 101592
rect 28424 101532 28500 101592
rect 190264 101532 190340 101592
rect 195976 101592 196324 101668
rect 196656 101668 196732 101728
rect 195976 101532 196052 101592
rect 21760 101462 21902 101526
rect 21966 101462 21972 101526
rect 21760 101456 21972 101462
rect 22168 101526 22516 101532
rect 22168 101462 22310 101526
rect 22374 101462 22446 101526
rect 22510 101462 22516 101526
rect 22168 101456 22516 101462
rect 22168 101396 22380 101456
rect 1632 101332 1844 101396
rect 1632 101276 1702 101332
rect 1758 101276 1844 101332
rect 22168 101320 22516 101396
rect 22576 101320 22788 101532
rect 22984 101526 23196 101532
rect 22984 101462 23126 101526
rect 23190 101462 23196 101526
rect 22984 101390 23196 101462
rect 22984 101326 22990 101390
rect 23054 101326 23196 101390
rect 22984 101320 23196 101326
rect 23392 101526 23604 101532
rect 23392 101462 23534 101526
rect 23598 101462 23604 101526
rect 23392 101390 23604 101462
rect 23392 101326 23534 101390
rect 23598 101326 23604 101390
rect 23392 101320 23604 101326
rect 28288 101390 28636 101532
rect 28288 101326 28430 101390
rect 28494 101326 28636 101390
rect 1632 101260 1844 101276
rect 22304 101260 22380 101320
rect 1224 101254 1844 101260
rect 1224 101190 1230 101254
rect 1294 101190 1844 101254
rect 1224 101184 1844 101190
rect 21760 101254 21972 101260
rect 21760 101190 21902 101254
rect 21966 101190 21972 101254
rect 21760 100912 21972 101190
rect 22168 100982 22380 101260
rect 22440 101260 22516 101320
rect 22440 101184 22788 101260
rect 22168 100918 22174 100982
rect 22238 100918 22380 100982
rect 22168 100912 22380 100918
rect 22576 100982 22788 101184
rect 22576 100918 22582 100982
rect 22646 100918 22788 100982
rect 22576 100912 22788 100918
rect 22984 101118 23196 101124
rect 22984 101054 22990 101118
rect 23054 101054 23196 101118
rect 22984 100912 23196 101054
rect 23392 101118 23604 101124
rect 23392 101054 23534 101118
rect 23598 101054 23604 101118
rect 23392 100912 23604 101054
rect 28288 101048 28636 101326
rect 28560 100988 28636 101048
rect 21760 100852 21836 100912
rect 22984 100852 23060 100912
rect 23528 100852 23604 100912
rect 21760 100710 21972 100852
rect 21760 100646 21766 100710
rect 21830 100646 21972 100710
rect 21760 100640 21972 100646
rect 22168 100710 22380 100716
rect 22168 100646 22174 100710
rect 22238 100646 22380 100710
rect 22168 100504 22380 100646
rect 22576 100710 22788 100716
rect 22576 100646 22582 100710
rect 22646 100646 22788 100710
rect 22576 100504 22788 100646
rect 22304 100444 22380 100504
rect 22712 100444 22788 100504
rect 21760 100438 21972 100444
rect 21760 100374 21766 100438
rect 21830 100374 21972 100438
rect 21760 100302 21972 100374
rect 21760 100238 21766 100302
rect 21830 100238 21972 100302
rect 21760 100232 21972 100238
rect 22168 100308 22380 100444
rect 22168 100302 22516 100308
rect 22168 100238 22446 100302
rect 22510 100238 22516 100302
rect 22168 100232 22516 100238
rect 22576 100232 22788 100444
rect 22984 100504 23196 100852
rect 23392 100504 23604 100852
rect 22984 100444 23060 100504
rect 23392 100444 23468 100504
rect 22984 100302 23196 100444
rect 22984 100238 23126 100302
rect 23190 100238 23196 100302
rect 22984 100232 23196 100238
rect 23392 100302 23604 100444
rect 28288 100368 28636 100988
rect 28560 100308 28636 100368
rect 23392 100238 23398 100302
rect 23462 100238 23604 100302
rect 23392 100232 23604 100238
rect 21760 100030 21972 100036
rect 21760 99966 21766 100030
rect 21830 99966 21972 100030
rect 21760 99894 21972 99966
rect 21760 99830 21766 99894
rect 21830 99830 21972 99894
rect 21760 99824 21972 99830
rect 1632 99652 1844 99764
rect 1632 99628 1702 99652
rect 1224 99622 1702 99628
rect 1224 99558 1230 99622
rect 1294 99596 1702 99622
rect 1758 99596 1844 99652
rect 22168 99688 22380 100036
rect 22478 100030 22788 100036
rect 22440 99966 22446 100030
rect 22510 99966 22788 100030
rect 22478 99960 22788 99966
rect 22688 99764 22788 99960
rect 22984 100030 23196 100036
rect 22984 99966 23126 100030
rect 23190 99966 23196 100030
rect 22984 99894 23196 99966
rect 22984 99830 23126 99894
rect 23190 99830 23196 99894
rect 22984 99824 23196 99830
rect 23392 100030 23604 100036
rect 23392 99966 23398 100030
rect 23462 99966 23604 100030
rect 23392 99894 23604 99966
rect 23392 99830 23534 99894
rect 23598 99830 23604 99894
rect 23392 99824 23604 99830
rect 28288 99824 28636 100308
rect 190128 101390 190340 101532
rect 190128 101326 190270 101390
rect 190334 101326 190340 101390
rect 190128 101048 190340 101326
rect 195024 101526 195236 101532
rect 195024 101462 195030 101526
rect 195094 101462 195236 101526
rect 195024 101390 195236 101462
rect 195024 101326 195030 101390
rect 195094 101326 195236 101390
rect 195024 101320 195236 101326
rect 195432 101526 195644 101532
rect 195432 101462 195438 101526
rect 195502 101462 195644 101526
rect 195432 101390 195644 101462
rect 195432 101326 195438 101390
rect 195502 101326 195644 101390
rect 195432 101320 195644 101326
rect 195840 101526 196460 101532
rect 195840 101462 195846 101526
rect 195910 101462 196460 101526
rect 195840 101456 196460 101462
rect 196656 101526 196868 101668
rect 196656 101462 196798 101526
rect 196862 101462 196868 101526
rect 196656 101456 196868 101462
rect 195840 101396 196052 101456
rect 195840 101320 196188 101396
rect 196248 101320 196460 101456
rect 216784 101390 217540 101396
rect 216784 101332 217470 101390
rect 196112 101260 196188 101320
rect 216784 101276 216908 101332
rect 216964 101326 217470 101332
rect 217534 101326 217540 101390
rect 216964 101320 217540 101326
rect 216964 101276 216996 101320
rect 195024 101118 195236 101124
rect 195024 101054 195030 101118
rect 195094 101054 195236 101118
rect 190128 100988 190204 101048
rect 190128 100982 190340 100988
rect 190128 100918 190270 100982
rect 190334 100918 190340 100982
rect 190128 100368 190340 100918
rect 195024 100912 195236 101054
rect 195432 101118 195644 101124
rect 195432 101054 195438 101118
rect 195502 101054 195644 101118
rect 195432 100912 195644 101054
rect 195840 100982 196052 101260
rect 196112 101184 196460 101260
rect 195840 100918 195846 100982
rect 195910 100918 196052 100982
rect 195840 100912 196052 100918
rect 196248 100982 196460 101184
rect 196248 100918 196254 100982
rect 196318 100918 196460 100982
rect 196248 100912 196460 100918
rect 196656 101254 196868 101260
rect 196656 101190 196798 101254
rect 196862 101190 196868 101254
rect 196656 100912 196868 101190
rect 216784 101184 216996 101276
rect 195024 100852 195100 100912
rect 195568 100852 195644 100912
rect 196656 100852 196732 100912
rect 195024 100504 195236 100852
rect 195432 100776 196868 100852
rect 195432 100504 195644 100776
rect 195840 100710 196052 100716
rect 195840 100646 195846 100710
rect 195910 100646 196052 100710
rect 195840 100504 196052 100646
rect 196248 100710 196460 100716
rect 196248 100646 196254 100710
rect 196318 100646 196460 100710
rect 196248 100504 196460 100646
rect 196656 100710 196868 100776
rect 196656 100646 196662 100710
rect 196726 100646 196868 100710
rect 196656 100640 196868 100646
rect 195024 100444 195100 100504
rect 195432 100444 195508 100504
rect 195976 100444 196052 100504
rect 196384 100444 196460 100504
rect 190128 100308 190204 100368
rect 190128 99824 190340 100308
rect 195024 100302 195236 100444
rect 195024 100238 195030 100302
rect 195094 100238 195236 100302
rect 195024 100232 195236 100238
rect 195432 100302 195644 100444
rect 195432 100238 195574 100302
rect 195638 100238 195644 100302
rect 195432 100232 195644 100238
rect 195840 100368 196460 100444
rect 195840 100302 196052 100368
rect 195840 100238 195846 100302
rect 195910 100238 196052 100302
rect 195840 100232 196052 100238
rect 196248 100232 196460 100368
rect 196656 100438 196868 100444
rect 196656 100374 196662 100438
rect 196726 100374 196868 100438
rect 196656 100302 196868 100374
rect 196656 100238 196798 100302
rect 196862 100238 196868 100302
rect 196656 100232 196868 100238
rect 195024 100030 195236 100036
rect 195024 99966 195030 100030
rect 195094 99966 195236 100030
rect 195024 99894 195236 99966
rect 195024 99830 195166 99894
rect 195230 99830 195236 99894
rect 195024 99824 195236 99830
rect 195432 100030 195644 100036
rect 195432 99966 195574 100030
rect 195638 99966 195644 100030
rect 195432 99894 195644 99966
rect 195432 99830 195574 99894
rect 195638 99830 195644 99894
rect 195432 99824 195644 99830
rect 195840 100030 196052 100036
rect 195840 99966 195846 100030
rect 195910 99966 196052 100030
rect 22576 99688 22788 99764
rect 28288 99764 28364 99824
rect 190128 99764 190204 99824
rect 22168 99628 22244 99688
rect 22576 99628 22652 99688
rect 1294 99558 1844 99596
rect 1224 99552 1844 99558
rect 21760 99622 21972 99628
rect 21760 99558 21766 99622
rect 21830 99558 21972 99622
rect 21760 99486 21972 99558
rect 21760 99422 21902 99486
rect 21966 99422 21972 99486
rect 21760 99416 21972 99422
rect 22168 99552 22788 99628
rect 22168 99416 22380 99552
rect 22576 99486 22788 99552
rect 22576 99422 22718 99486
rect 22782 99422 22788 99486
rect 22576 99416 22788 99422
rect 22984 99622 23196 99628
rect 22984 99558 23126 99622
rect 23190 99558 23196 99622
rect 22984 99486 23196 99558
rect 22984 99422 23126 99486
rect 23190 99422 23196 99486
rect 22984 99416 23196 99422
rect 23392 99622 23604 99628
rect 23392 99558 23534 99622
rect 23598 99558 23604 99622
rect 23392 99486 23604 99558
rect 23392 99422 23398 99486
rect 23462 99422 23604 99486
rect 23392 99416 23604 99422
rect 28288 99552 28636 99764
rect 190128 99552 190340 99764
rect 195840 99688 196052 99966
rect 196248 99764 196460 100036
rect 196656 100030 196868 100036
rect 196656 99966 196798 100030
rect 196862 99966 196868 100030
rect 196656 99894 196868 99966
rect 196656 99830 196662 99894
rect 196726 99830 196868 99894
rect 196656 99824 196868 99830
rect 195976 99628 196052 99688
rect 196112 99688 196460 99764
rect 216784 99758 217540 99764
rect 216784 99694 217470 99758
rect 217534 99694 217540 99758
rect 216784 99688 217540 99694
rect 196112 99628 196188 99688
rect 216784 99652 216996 99688
rect 28288 99492 28364 99552
rect 190264 99492 190340 99552
rect 28288 99280 28636 99492
rect 190128 99280 190340 99492
rect 195024 99622 195236 99628
rect 195024 99558 195166 99622
rect 195230 99558 195236 99622
rect 195024 99486 195236 99558
rect 195024 99422 195030 99486
rect 195094 99422 195236 99486
rect 195024 99416 195236 99422
rect 195432 99622 195644 99628
rect 195432 99558 195574 99622
rect 195638 99558 195644 99622
rect 195432 99486 195644 99558
rect 195432 99422 195574 99486
rect 195638 99422 195644 99486
rect 195432 99416 195644 99422
rect 195840 99552 196188 99628
rect 195840 99492 196052 99552
rect 196248 99492 196460 99628
rect 195840 99416 196460 99492
rect 196656 99622 196868 99628
rect 196656 99558 196662 99622
rect 196726 99558 196868 99622
rect 196656 99486 196868 99558
rect 216784 99596 216908 99652
rect 216964 99596 216996 99652
rect 216784 99552 216996 99596
rect 196656 99422 196798 99486
rect 196862 99422 196868 99486
rect 196656 99416 196868 99422
rect 195976 99356 196052 99416
rect 195976 99280 196324 99356
rect 28560 99220 28636 99280
rect 190264 99220 190340 99280
rect 196248 99220 196324 99280
rect 21760 99214 21972 99220
rect 21760 99150 21902 99214
rect 21966 99150 21972 99214
rect 21760 99078 21972 99150
rect 21760 99014 21766 99078
rect 21830 99014 21972 99078
rect 21760 99008 21972 99014
rect 22168 99084 22380 99220
rect 22576 99214 22788 99220
rect 22576 99150 22718 99214
rect 22782 99150 22788 99214
rect 22576 99084 22788 99150
rect 22168 99008 22788 99084
rect 22984 99214 23196 99220
rect 22984 99150 23126 99214
rect 23190 99150 23196 99214
rect 22984 99078 23196 99150
rect 22984 99014 23126 99078
rect 23190 99014 23196 99078
rect 22984 99008 23196 99014
rect 23392 99214 23604 99220
rect 23392 99150 23398 99214
rect 23462 99150 23604 99214
rect 23392 99078 23604 99150
rect 23392 99014 23534 99078
rect 23598 99014 23604 99078
rect 23392 99008 23604 99014
rect 28288 99008 28636 99220
rect 190128 99008 190340 99220
rect 195024 99214 195236 99220
rect 195024 99150 195030 99214
rect 195094 99150 195236 99214
rect 195024 99078 195236 99150
rect 195024 99014 195030 99078
rect 195094 99014 195236 99078
rect 195024 99008 195236 99014
rect 195432 99214 195644 99220
rect 195432 99150 195574 99214
rect 195638 99150 195644 99214
rect 195432 99078 195644 99150
rect 195432 99014 195574 99078
rect 195638 99014 195644 99078
rect 195432 99008 195644 99014
rect 195840 99144 196460 99220
rect 195840 99084 196052 99144
rect 195840 99078 196188 99084
rect 195840 99014 196118 99078
rect 196182 99014 196188 99078
rect 195840 99008 196188 99014
rect 196248 99008 196460 99144
rect 196656 99214 196868 99220
rect 196656 99150 196798 99214
rect 196862 99150 196868 99214
rect 196656 99078 196868 99150
rect 196656 99014 196798 99078
rect 196862 99014 196868 99078
rect 196656 99008 196868 99014
rect 22304 98948 22380 99008
rect 28424 98948 28500 99008
rect 190264 98948 190340 99008
rect 22304 98872 22652 98948
rect 22576 98812 22652 98872
rect 21760 98806 21972 98812
rect 21760 98742 21766 98806
rect 21830 98742 21972 98806
rect 21760 98670 21972 98742
rect 21760 98606 21766 98670
rect 21830 98606 21972 98670
rect 21760 98600 21972 98606
rect 22168 98670 22380 98812
rect 22168 98606 22174 98670
rect 22238 98606 22380 98670
rect 22168 98600 22380 98606
rect 22576 98670 22788 98812
rect 22576 98606 22718 98670
rect 22782 98606 22788 98670
rect 22576 98600 22788 98606
rect 22984 98806 23196 98812
rect 22984 98742 23126 98806
rect 23190 98742 23196 98806
rect 22984 98670 23196 98742
rect 22984 98606 22990 98670
rect 23054 98606 23196 98670
rect 22984 98600 23196 98606
rect 23392 98806 23604 98812
rect 23392 98742 23534 98806
rect 23598 98742 23604 98806
rect 23392 98670 23604 98742
rect 23392 98606 23534 98670
rect 23598 98606 23604 98670
rect 23392 98600 23604 98606
rect 28288 98736 28636 98948
rect 190128 98736 190340 98948
rect 195024 98806 195236 98812
rect 195024 98742 195030 98806
rect 195094 98742 195236 98806
rect 28288 98676 28364 98736
rect 190128 98676 190204 98736
rect 28288 98464 28636 98676
rect 190128 98464 190340 98676
rect 195024 98670 195236 98742
rect 195024 98606 195030 98670
rect 195094 98606 195236 98670
rect 195024 98600 195236 98606
rect 195432 98806 195644 98812
rect 195432 98742 195574 98806
rect 195638 98742 195644 98806
rect 195432 98670 195644 98742
rect 195432 98606 195574 98670
rect 195638 98606 195644 98670
rect 195432 98600 195644 98606
rect 195840 98670 196052 98812
rect 196150 98806 196460 98812
rect 196112 98742 196118 98806
rect 196182 98742 196460 98806
rect 196150 98736 196460 98742
rect 195840 98606 195982 98670
rect 196046 98606 196052 98670
rect 195840 98600 196052 98606
rect 196248 98600 196460 98736
rect 196656 98806 196868 98812
rect 196656 98742 196798 98806
rect 196862 98742 196868 98806
rect 196656 98670 196868 98742
rect 196656 98606 196662 98670
rect 196726 98606 196868 98670
rect 196656 98600 196868 98606
rect 196248 98540 196324 98600
rect 195976 98464 196324 98540
rect 28424 98404 28500 98464
rect 190128 98404 190204 98464
rect 195976 98404 196052 98464
rect 21760 98398 21972 98404
rect 21760 98334 21766 98398
rect 21830 98334 21972 98398
rect 21760 98262 21972 98334
rect 21760 98198 21902 98262
rect 21966 98198 21972 98262
rect 21760 98192 21972 98198
rect 22168 98398 22788 98404
rect 22168 98334 22174 98398
rect 22238 98334 22718 98398
rect 22782 98334 22788 98398
rect 22168 98328 22788 98334
rect 22168 98268 22380 98328
rect 22168 98262 22516 98268
rect 22168 98198 22310 98262
rect 22374 98198 22446 98262
rect 22510 98198 22516 98262
rect 22168 98192 22516 98198
rect 22576 98192 22788 98328
rect 22984 98398 23196 98404
rect 22984 98334 22990 98398
rect 23054 98334 23196 98398
rect 22984 98262 23196 98334
rect 22984 98198 23126 98262
rect 23190 98198 23196 98262
rect 22984 98192 23196 98198
rect 23392 98398 23604 98404
rect 23392 98334 23534 98398
rect 23598 98334 23604 98398
rect 23392 98262 23604 98334
rect 23392 98198 23398 98262
rect 23462 98198 23604 98262
rect 23392 98192 23604 98198
rect 28288 98192 28636 98404
rect 190128 98192 190340 98404
rect 195024 98398 195236 98404
rect 195024 98334 195030 98398
rect 195094 98334 195236 98398
rect 195024 98262 195236 98334
rect 195024 98198 195030 98262
rect 195094 98198 195236 98262
rect 195024 98192 195236 98198
rect 195432 98398 195644 98404
rect 195432 98334 195574 98398
rect 195638 98334 195644 98398
rect 195432 98262 195644 98334
rect 195432 98198 195574 98262
rect 195638 98198 195644 98262
rect 195432 98192 195644 98198
rect 195840 98398 196460 98404
rect 195840 98334 195982 98398
rect 196046 98334 196460 98398
rect 195840 98328 196460 98334
rect 195840 98192 196052 98328
rect 196248 98262 196460 98328
rect 196248 98198 196390 98262
rect 196454 98198 196460 98262
rect 196248 98192 196460 98198
rect 196656 98398 196868 98404
rect 196656 98334 196662 98398
rect 196726 98334 196868 98398
rect 196656 98262 196868 98334
rect 196656 98198 196798 98262
rect 196862 98198 196868 98262
rect 196656 98192 196868 98198
rect 28424 98132 28500 98192
rect 190264 98132 190340 98192
rect 1224 97990 1844 97996
rect 1224 97926 1230 97990
rect 1294 97972 1844 97990
rect 1294 97926 1702 97972
rect 1224 97920 1702 97926
rect 1632 97916 1702 97920
rect 1758 97916 1844 97972
rect 1632 97784 1844 97916
rect 21760 97990 21972 97996
rect 21760 97926 21902 97990
rect 21966 97926 21972 97990
rect 21760 97784 21972 97926
rect 22168 97990 22380 97996
rect 22478 97990 22788 97996
rect 22168 97926 22310 97990
rect 22374 97926 22380 97990
rect 22440 97926 22446 97990
rect 22510 97926 22788 97990
rect 22168 97854 22380 97926
rect 22478 97920 22788 97926
rect 22168 97790 22174 97854
rect 22238 97790 22380 97854
rect 22168 97784 22380 97790
rect 22576 97784 22788 97920
rect 22984 97990 23196 97996
rect 22984 97926 23126 97990
rect 23190 97926 23196 97990
rect 22984 97854 23196 97926
rect 22984 97790 22990 97854
rect 23054 97790 23196 97854
rect 22984 97784 23196 97790
rect 23392 97990 23604 97996
rect 23392 97926 23398 97990
rect 23462 97926 23604 97990
rect 23392 97854 23604 97926
rect 28288 97920 28636 98132
rect 190128 97920 190340 98132
rect 28560 97860 28636 97920
rect 190264 97860 190340 97920
rect 23392 97790 23534 97854
rect 23598 97790 23604 97854
rect 23392 97784 23604 97790
rect 21760 97724 21836 97784
rect 21760 97376 21972 97724
rect 28288 97648 28636 97860
rect 190128 97648 190340 97860
rect 195024 97990 195236 97996
rect 195024 97926 195030 97990
rect 195094 97926 195236 97990
rect 195024 97854 195236 97926
rect 195024 97790 195166 97854
rect 195230 97790 195236 97854
rect 195024 97784 195236 97790
rect 195432 97990 195644 97996
rect 195432 97926 195574 97990
rect 195638 97926 195644 97990
rect 195432 97854 195644 97926
rect 195432 97790 195438 97854
rect 195502 97790 195644 97854
rect 195432 97784 195644 97790
rect 195840 97854 196052 97996
rect 195840 97790 195846 97854
rect 195910 97790 196052 97854
rect 195840 97784 196052 97790
rect 196248 97990 196460 97996
rect 196248 97926 196390 97990
rect 196454 97926 196460 97990
rect 196248 97854 196460 97926
rect 196248 97790 196254 97854
rect 196318 97790 196460 97854
rect 196248 97784 196460 97790
rect 196656 97990 196868 97996
rect 196656 97926 196798 97990
rect 196862 97926 196868 97990
rect 196656 97784 196868 97926
rect 216784 97972 216996 97996
rect 216784 97916 216908 97972
rect 216964 97916 216996 97972
rect 216784 97860 216996 97916
rect 216784 97854 217540 97860
rect 216784 97790 217470 97854
rect 217534 97790 217540 97854
rect 216784 97784 217540 97790
rect 196792 97724 196868 97784
rect 28424 97588 28500 97648
rect 190128 97588 190204 97648
rect 22168 97582 22380 97588
rect 22168 97518 22174 97582
rect 22238 97518 22380 97582
rect 22168 97376 22380 97518
rect 22576 97452 22788 97588
rect 21760 97316 21836 97376
rect 22304 97316 22380 97376
rect 22440 97376 22788 97452
rect 22984 97582 23196 97588
rect 22984 97518 22990 97582
rect 23054 97518 23196 97582
rect 22984 97446 23196 97518
rect 22984 97382 22990 97446
rect 23054 97382 23196 97446
rect 22984 97376 23196 97382
rect 23392 97582 23604 97588
rect 23392 97518 23534 97582
rect 23598 97518 23604 97582
rect 23392 97446 23604 97518
rect 23392 97382 23534 97446
rect 23598 97382 23604 97446
rect 23392 97376 23604 97382
rect 22440 97316 22516 97376
rect 21760 96968 21972 97316
rect 22168 97240 22516 97316
rect 22168 97044 22380 97240
rect 22576 97044 22788 97316
rect 22168 97038 22788 97044
rect 22168 96974 22718 97038
rect 22782 96974 22788 97038
rect 22168 96968 22788 96974
rect 22984 97174 23196 97180
rect 22984 97110 22990 97174
rect 23054 97110 23196 97174
rect 22984 96968 23196 97110
rect 23392 97174 23604 97180
rect 23392 97110 23534 97174
rect 23598 97110 23604 97174
rect 23392 96968 23604 97110
rect 21896 96908 21972 96968
rect 23120 96908 23196 96968
rect 23528 96908 23604 96968
rect 21760 96766 21972 96908
rect 21760 96702 21766 96766
rect 21830 96702 21972 96766
rect 21760 96696 21972 96702
rect 22168 96560 22380 96772
rect 22576 96766 22788 96772
rect 22576 96702 22718 96766
rect 22782 96702 22788 96766
rect 22576 96560 22788 96702
rect 22984 96560 23196 96908
rect 23392 96560 23604 96908
rect 22168 96500 22244 96560
rect 22576 96500 22652 96560
rect 22984 96500 23060 96560
rect 23528 96500 23604 96560
rect 21760 96494 21972 96500
rect 21760 96430 21766 96494
rect 21830 96430 21972 96494
rect 1632 96292 1844 96364
rect 1632 96236 1702 96292
rect 1758 96236 1844 96292
rect 21760 96358 21972 96430
rect 21760 96294 21766 96358
rect 21830 96294 21972 96358
rect 21760 96288 21972 96294
rect 22168 96358 22380 96500
rect 22168 96294 22310 96358
rect 22374 96294 22380 96358
rect 22168 96288 22380 96294
rect 22576 96288 22788 96500
rect 1632 96228 1844 96236
rect 22576 96228 22652 96288
rect 1224 96222 1844 96228
rect 1224 96158 1230 96222
rect 1294 96158 1844 96222
rect 1224 96152 1844 96158
rect 22304 96152 22652 96228
rect 22984 96152 23196 96500
rect 23392 96152 23604 96500
rect 28288 97104 28636 97588
rect 190128 97104 190340 97588
rect 195024 97582 195236 97588
rect 195024 97518 195166 97582
rect 195230 97518 195236 97582
rect 195024 97446 195236 97518
rect 195024 97382 195030 97446
rect 195094 97382 195236 97446
rect 195024 97376 195236 97382
rect 195432 97582 195644 97588
rect 195432 97518 195438 97582
rect 195502 97518 195644 97582
rect 195432 97446 195644 97518
rect 195432 97382 195574 97446
rect 195638 97382 195644 97446
rect 195432 97376 195644 97382
rect 195840 97582 196052 97588
rect 195840 97518 195846 97582
rect 195910 97518 196052 97582
rect 195840 97376 196052 97518
rect 196248 97582 196460 97588
rect 196248 97518 196254 97582
rect 196318 97518 196460 97582
rect 196248 97376 196460 97518
rect 196656 97376 196868 97724
rect 195840 97316 195916 97376
rect 196248 97316 196324 97376
rect 196792 97316 196868 97376
rect 195024 97174 195236 97180
rect 195024 97110 195030 97174
rect 195094 97110 195236 97174
rect 28288 97044 28364 97104
rect 190128 97044 190204 97104
rect 28288 96902 28636 97044
rect 28288 96838 28566 96902
rect 28630 96838 28636 96902
rect 28288 96630 28636 96838
rect 28288 96566 28566 96630
rect 28630 96566 28636 96630
rect 28288 96494 28636 96566
rect 28288 96430 28430 96494
rect 28494 96430 28636 96494
rect 28288 96424 28636 96430
rect 190128 96494 190340 97044
rect 190128 96430 190134 96494
rect 190198 96430 190340 96494
rect 190128 96424 190340 96430
rect 195024 96968 195236 97110
rect 195432 97174 195644 97180
rect 195432 97110 195574 97174
rect 195638 97110 195644 97174
rect 195432 96968 195644 97110
rect 195840 97044 196052 97316
rect 196248 97044 196460 97316
rect 195840 97038 196460 97044
rect 195840 96974 196254 97038
rect 196318 96974 196460 97038
rect 195840 96968 196460 96974
rect 196656 96968 196868 97316
rect 195024 96908 195100 96968
rect 195568 96908 195644 96968
rect 196792 96908 196868 96968
rect 195024 96560 195236 96908
rect 195432 96560 195644 96908
rect 195840 96560 196052 96772
rect 196248 96766 196460 96772
rect 196248 96702 196254 96766
rect 196318 96702 196460 96766
rect 196248 96560 196460 96702
rect 196656 96766 196868 96908
rect 196656 96702 196662 96766
rect 196726 96702 196868 96766
rect 196656 96696 196868 96702
rect 195024 96500 195100 96560
rect 195432 96500 195508 96560
rect 195840 96500 195916 96560
rect 196248 96500 196324 96560
rect 28288 96222 28636 96228
rect 28288 96158 28430 96222
rect 28494 96158 28636 96222
rect 22304 96092 22380 96152
rect 22984 96092 23060 96152
rect 23392 96092 23468 96152
rect 21760 96086 21972 96092
rect 21760 96022 21766 96086
rect 21830 96022 21972 96086
rect 21760 95950 21972 96022
rect 21760 95886 21766 95950
rect 21830 95886 21972 95950
rect 21760 95880 21972 95886
rect 22168 96086 22788 96092
rect 22168 96022 22310 96086
rect 22374 96022 22788 96086
rect 22168 96016 22788 96022
rect 22168 95744 22380 96016
rect 22576 95744 22788 96016
rect 22984 95950 23196 96092
rect 22984 95886 22990 95950
rect 23054 95886 23196 95950
rect 22984 95880 23196 95886
rect 23392 95950 23604 96092
rect 23392 95886 23398 95950
rect 23462 95886 23604 95950
rect 23392 95880 23604 95886
rect 28288 96086 28636 96158
rect 28288 96022 28430 96086
rect 28494 96022 28636 96086
rect 28288 95880 28636 96022
rect 190128 96222 190340 96228
rect 190128 96158 190134 96222
rect 190198 96158 190340 96222
rect 190128 95880 190340 96158
rect 195024 96152 195236 96500
rect 195432 96152 195644 96500
rect 195840 96358 196052 96500
rect 196248 96364 196460 96500
rect 196150 96358 196460 96364
rect 195840 96294 195982 96358
rect 196046 96294 196052 96358
rect 196112 96294 196118 96358
rect 196182 96294 196460 96358
rect 195840 96288 196052 96294
rect 196150 96288 196460 96294
rect 196656 96494 196868 96500
rect 196656 96430 196662 96494
rect 196726 96430 196868 96494
rect 196656 96358 196868 96430
rect 196656 96294 196662 96358
rect 196726 96294 196868 96358
rect 196656 96288 196868 96294
rect 216784 96358 217540 96364
rect 216784 96294 217470 96358
rect 217534 96294 217540 96358
rect 216784 96292 217540 96294
rect 216784 96236 216908 96292
rect 216964 96288 217540 96292
rect 216964 96236 216996 96288
rect 216784 96152 216996 96236
rect 195024 96092 195100 96152
rect 195432 96092 195508 96152
rect 195024 95950 195236 96092
rect 195024 95886 195030 95950
rect 195094 95886 195236 95950
rect 195024 95880 195236 95886
rect 195432 95950 195644 96092
rect 195432 95886 195574 95950
rect 195638 95886 195644 95950
rect 195432 95880 195644 95886
rect 195840 96086 196188 96092
rect 195840 96022 195982 96086
rect 196046 96022 196118 96086
rect 196182 96022 196188 96086
rect 195840 96016 196188 96022
rect 28424 95820 28500 95880
rect 190264 95820 190340 95880
rect 22168 95684 22244 95744
rect 22712 95684 22788 95744
rect 28288 95814 28636 95820
rect 28288 95750 28430 95814
rect 28494 95750 28636 95814
rect 21760 95678 21972 95684
rect 21760 95614 21766 95678
rect 21830 95614 21972 95678
rect 21760 95542 21972 95614
rect 21760 95478 21766 95542
rect 21830 95478 21972 95542
rect 21760 95472 21972 95478
rect 22168 95472 22380 95684
rect 22576 95542 22788 95684
rect 22576 95478 22582 95542
rect 22646 95478 22788 95542
rect 22576 95472 22788 95478
rect 22984 95678 23196 95684
rect 22984 95614 22990 95678
rect 23054 95614 23196 95678
rect 22984 95542 23196 95614
rect 22984 95478 22990 95542
rect 23054 95478 23196 95542
rect 22984 95472 23196 95478
rect 23392 95678 23604 95684
rect 23392 95614 23398 95678
rect 23462 95614 23604 95678
rect 23392 95542 23604 95614
rect 28288 95608 28636 95750
rect 190128 95608 190340 95820
rect 195840 95820 196052 96016
rect 196248 95820 196460 96092
rect 196656 96086 196868 96092
rect 196656 96022 196662 96086
rect 196726 96022 196868 96086
rect 196656 95950 196868 96022
rect 196656 95886 196798 95950
rect 196862 95886 196868 95950
rect 196656 95880 196868 95886
rect 195840 95814 196460 95820
rect 195840 95750 196254 95814
rect 196318 95750 196460 95814
rect 195840 95744 196460 95750
rect 196248 95684 196324 95744
rect 28424 95548 28500 95608
rect 190264 95548 190340 95608
rect 23392 95478 23534 95542
rect 23598 95478 23604 95542
rect 23392 95472 23604 95478
rect 21760 95270 21972 95276
rect 21760 95206 21766 95270
rect 21830 95206 21972 95270
rect 21760 95134 21972 95206
rect 21760 95070 21902 95134
rect 21966 95070 21972 95134
rect 21760 95064 21972 95070
rect 22168 95140 22380 95276
rect 22576 95270 22788 95276
rect 22576 95206 22582 95270
rect 22646 95206 22788 95270
rect 22576 95140 22788 95206
rect 22168 95134 22788 95140
rect 22168 95070 22718 95134
rect 22782 95070 22788 95134
rect 22168 95064 22788 95070
rect 22984 95270 23196 95276
rect 22984 95206 22990 95270
rect 23054 95206 23196 95270
rect 22984 95134 23196 95206
rect 22984 95070 23126 95134
rect 23190 95070 23196 95134
rect 22984 95064 23196 95070
rect 23392 95270 23604 95276
rect 23392 95206 23534 95270
rect 23598 95206 23604 95270
rect 23392 95134 23604 95206
rect 23392 95070 23398 95134
rect 23462 95070 23604 95134
rect 23392 95064 23604 95070
rect 28288 95064 28636 95548
rect 190128 95270 190340 95548
rect 195024 95678 195236 95684
rect 195024 95614 195030 95678
rect 195094 95614 195236 95678
rect 195024 95542 195236 95614
rect 195024 95478 195166 95542
rect 195230 95478 195236 95542
rect 195024 95472 195236 95478
rect 195432 95678 195644 95684
rect 195432 95614 195574 95678
rect 195638 95614 195644 95678
rect 195432 95542 195644 95614
rect 195432 95478 195574 95542
rect 195638 95478 195644 95542
rect 195432 95472 195644 95478
rect 195840 95678 196188 95684
rect 195840 95614 196118 95678
rect 196182 95614 196188 95678
rect 195840 95608 196188 95614
rect 195840 95548 196052 95608
rect 195840 95542 196188 95548
rect 195840 95478 196118 95542
rect 196182 95478 196188 95542
rect 195840 95472 196188 95478
rect 196248 95472 196460 95684
rect 196656 95678 196868 95684
rect 196656 95614 196798 95678
rect 196862 95614 196868 95678
rect 196656 95542 196868 95614
rect 196656 95478 196662 95542
rect 196726 95478 196868 95542
rect 196656 95472 196868 95478
rect 190128 95206 190270 95270
rect 190334 95206 190340 95270
rect 190128 95064 190340 95206
rect 195024 95270 195236 95276
rect 195024 95206 195166 95270
rect 195230 95206 195236 95270
rect 195024 95134 195236 95206
rect 195024 95070 195030 95134
rect 195094 95070 195236 95134
rect 195024 95064 195236 95070
rect 195432 95270 195644 95276
rect 195432 95206 195574 95270
rect 195638 95206 195644 95270
rect 195432 95134 195644 95206
rect 195432 95070 195574 95134
rect 195638 95070 195644 95134
rect 195432 95064 195644 95070
rect 195840 95134 196052 95276
rect 196150 95270 196460 95276
rect 196112 95206 196118 95270
rect 196182 95206 196460 95270
rect 196150 95200 196460 95206
rect 195840 95070 195982 95134
rect 196046 95070 196052 95134
rect 195840 95064 196052 95070
rect 196248 95064 196460 95200
rect 196656 95270 196868 95276
rect 196656 95206 196662 95270
rect 196726 95206 196868 95270
rect 196656 95134 196868 95206
rect 196656 95070 196798 95134
rect 196862 95070 196868 95134
rect 196656 95064 196868 95070
rect 28560 95004 28636 95064
rect 190264 95004 190340 95064
rect 196248 95004 196324 95064
rect 21760 94862 21972 94868
rect 21760 94798 21902 94862
rect 21966 94798 21972 94862
rect 1224 94726 1844 94732
rect 1224 94662 1230 94726
rect 1294 94662 1844 94726
rect 1224 94656 1844 94662
rect 21760 94726 21972 94798
rect 21760 94662 21766 94726
rect 21830 94662 21972 94726
rect 21760 94656 21972 94662
rect 22168 94862 22788 94868
rect 22168 94798 22718 94862
rect 22782 94798 22788 94862
rect 22168 94792 22788 94798
rect 22168 94732 22380 94792
rect 22168 94726 22516 94732
rect 22168 94662 22310 94726
rect 22374 94662 22446 94726
rect 22510 94662 22516 94726
rect 22168 94656 22516 94662
rect 22576 94656 22788 94792
rect 22984 94862 23196 94868
rect 22984 94798 23126 94862
rect 23190 94798 23196 94862
rect 22984 94726 23196 94798
rect 22984 94662 22990 94726
rect 23054 94662 23196 94726
rect 22984 94656 23196 94662
rect 23392 94862 23604 94868
rect 23392 94798 23398 94862
rect 23462 94798 23604 94862
rect 23392 94726 23604 94798
rect 28288 94792 28636 95004
rect 190128 94998 190340 95004
rect 190128 94934 190270 94998
rect 190334 94934 190340 94998
rect 190128 94792 190340 94934
rect 195976 94928 196324 95004
rect 195976 94868 196052 94928
rect 28424 94732 28500 94792
rect 190264 94732 190340 94792
rect 23392 94662 23534 94726
rect 23598 94662 23604 94726
rect 23392 94656 23604 94662
rect 1632 94612 1844 94656
rect 1632 94556 1702 94612
rect 1758 94556 1844 94612
rect 1632 94520 1844 94556
rect 28288 94520 28636 94732
rect 190128 94520 190340 94732
rect 195024 94862 195236 94868
rect 195024 94798 195030 94862
rect 195094 94798 195236 94862
rect 195024 94726 195236 94798
rect 195024 94662 195030 94726
rect 195094 94662 195236 94726
rect 195024 94656 195236 94662
rect 195432 94862 195644 94868
rect 195432 94798 195574 94862
rect 195638 94798 195644 94862
rect 195432 94726 195644 94798
rect 195432 94662 195574 94726
rect 195638 94662 195644 94726
rect 195432 94656 195644 94662
rect 195840 94862 196460 94868
rect 195840 94798 195982 94862
rect 196046 94798 196460 94862
rect 195840 94792 196460 94798
rect 195840 94732 196052 94792
rect 195840 94726 196188 94732
rect 195840 94662 196118 94726
rect 196182 94662 196188 94726
rect 195840 94656 196188 94662
rect 196248 94656 196460 94792
rect 196656 94862 196868 94868
rect 196656 94798 196798 94862
rect 196862 94798 196868 94862
rect 196656 94726 196868 94798
rect 196656 94662 196662 94726
rect 196726 94662 196868 94726
rect 196656 94656 196868 94662
rect 216784 94612 216996 94732
rect 216784 94556 216908 94612
rect 216964 94596 216996 94612
rect 216964 94590 217540 94596
rect 216964 94556 217470 94590
rect 216784 94526 217470 94556
rect 217534 94526 217540 94590
rect 216784 94520 217540 94526
rect 28288 94460 28364 94520
rect 190128 94460 190204 94520
rect 21760 94454 21972 94460
rect 21760 94390 21766 94454
rect 21830 94390 21972 94454
rect 21760 94318 21972 94390
rect 21760 94254 21766 94318
rect 21830 94254 21972 94318
rect 21760 94248 21972 94254
rect 22168 94454 22380 94460
rect 22478 94454 22788 94460
rect 22168 94390 22310 94454
rect 22374 94390 22380 94454
rect 22440 94390 22446 94454
rect 22510 94390 22788 94454
rect 22168 94248 22380 94390
rect 22478 94384 22788 94390
rect 22576 94318 22788 94384
rect 22576 94254 22718 94318
rect 22782 94254 22788 94318
rect 22576 94248 22788 94254
rect 22984 94454 23196 94460
rect 22984 94390 22990 94454
rect 23054 94390 23196 94454
rect 22984 94318 23196 94390
rect 22984 94254 22990 94318
rect 23054 94254 23196 94318
rect 22984 94248 23196 94254
rect 23392 94454 23604 94460
rect 23392 94390 23534 94454
rect 23598 94390 23604 94454
rect 23392 94318 23604 94390
rect 23392 94254 23534 94318
rect 23598 94254 23604 94318
rect 23392 94248 23604 94254
rect 28288 94248 28636 94460
rect 28560 94188 28636 94248
rect 21760 94046 21972 94052
rect 21760 93982 21766 94046
rect 21830 93982 21972 94046
rect 21760 93840 21972 93982
rect 22168 93916 22380 94052
rect 22576 94046 22788 94052
rect 22576 93982 22718 94046
rect 22782 93982 22788 94046
rect 22576 93916 22788 93982
rect 22168 93910 22788 93916
rect 22168 93846 22310 93910
rect 22374 93846 22788 93910
rect 22168 93840 22788 93846
rect 22984 94046 23196 94052
rect 22984 93982 22990 94046
rect 23054 93982 23196 94046
rect 22984 93910 23196 93982
rect 22984 93846 22990 93910
rect 23054 93846 23196 93910
rect 22984 93840 23196 93846
rect 23392 94046 23604 94052
rect 23392 93982 23534 94046
rect 23598 93982 23604 94046
rect 23392 93910 23604 93982
rect 28288 93976 28636 94188
rect 190128 94248 190340 94460
rect 195024 94454 195236 94460
rect 195024 94390 195030 94454
rect 195094 94390 195236 94454
rect 195024 94318 195236 94390
rect 195024 94254 195030 94318
rect 195094 94254 195236 94318
rect 195024 94248 195236 94254
rect 195432 94454 195644 94460
rect 195432 94390 195574 94454
rect 195638 94390 195644 94454
rect 195432 94318 195644 94390
rect 195432 94254 195438 94318
rect 195502 94254 195644 94318
rect 195432 94248 195644 94254
rect 195840 94318 196052 94460
rect 196150 94454 196460 94460
rect 196112 94390 196118 94454
rect 196182 94390 196460 94454
rect 196150 94384 196460 94390
rect 196248 94324 196460 94384
rect 196150 94318 196460 94324
rect 195840 94254 195982 94318
rect 196046 94254 196052 94318
rect 196112 94254 196118 94318
rect 196182 94254 196254 94318
rect 196318 94254 196460 94318
rect 195840 94248 196052 94254
rect 196150 94248 196460 94254
rect 196656 94454 196868 94460
rect 196656 94390 196662 94454
rect 196726 94390 196868 94454
rect 196656 94318 196868 94390
rect 196656 94254 196662 94318
rect 196726 94254 196868 94318
rect 196656 94248 196868 94254
rect 190128 94188 190204 94248
rect 190128 93976 190340 94188
rect 28424 93916 28500 93976
rect 190264 93916 190340 93976
rect 23392 93846 23398 93910
rect 23462 93846 23604 93910
rect 23392 93840 23604 93846
rect 21896 93780 21972 93840
rect 21760 93432 21972 93780
rect 22304 93780 22380 93840
rect 22304 93704 22652 93780
rect 28288 93774 28636 93916
rect 28288 93710 28294 93774
rect 28358 93710 28636 93774
rect 28288 93704 28636 93710
rect 190128 93704 190340 93916
rect 195024 94046 195236 94052
rect 195024 93982 195030 94046
rect 195094 93982 195236 94046
rect 195024 93910 195236 93982
rect 195024 93846 195030 93910
rect 195094 93846 195236 93910
rect 195024 93840 195236 93846
rect 195432 94046 195644 94052
rect 195432 93982 195438 94046
rect 195502 93982 195644 94046
rect 195432 93910 195644 93982
rect 195432 93846 195438 93910
rect 195502 93846 195644 93910
rect 195432 93840 195644 93846
rect 195840 94046 196188 94052
rect 195840 93982 195982 94046
rect 196046 93982 196118 94046
rect 196182 93982 196188 94046
rect 195840 93976 196188 93982
rect 196248 94046 196460 94052
rect 196248 93982 196254 94046
rect 196318 93982 196460 94046
rect 195840 93910 196052 93976
rect 195840 93846 195982 93910
rect 196046 93846 196052 93910
rect 195840 93840 196052 93846
rect 196248 93840 196460 93982
rect 196656 94046 196868 94052
rect 196656 93982 196662 94046
rect 196726 93982 196868 94046
rect 196656 93840 196868 93982
rect 22576 93644 22652 93704
rect 28560 93644 28636 93704
rect 190264 93644 190340 93704
rect 196656 93780 196732 93840
rect 22168 93638 22380 93644
rect 22168 93574 22310 93638
rect 22374 93574 22380 93638
rect 22168 93432 22380 93574
rect 21896 93372 21972 93432
rect 22304 93372 22380 93432
rect 21760 93024 21972 93372
rect 22168 93024 22380 93372
rect 22576 93432 22788 93644
rect 22984 93638 23196 93644
rect 22984 93574 22990 93638
rect 23054 93574 23196 93638
rect 22984 93502 23196 93574
rect 22984 93438 22990 93502
rect 23054 93438 23196 93502
rect 22984 93432 23196 93438
rect 23392 93638 23604 93644
rect 23392 93574 23398 93638
rect 23462 93574 23604 93638
rect 23392 93502 23604 93574
rect 23392 93438 23534 93502
rect 23598 93438 23604 93502
rect 23392 93432 23604 93438
rect 28288 93502 28636 93644
rect 28288 93438 28294 93502
rect 28358 93438 28636 93502
rect 22576 93372 22652 93432
rect 22576 93024 22788 93372
rect 22984 93230 23196 93236
rect 22984 93166 22990 93230
rect 23054 93166 23196 93230
rect 22984 93094 23196 93166
rect 22984 93030 23126 93094
rect 23190 93030 23196 93094
rect 22984 93024 23196 93030
rect 23392 93230 23604 93236
rect 23392 93166 23534 93230
rect 23598 93166 23604 93230
rect 23392 93094 23604 93166
rect 28288 93160 28636 93438
rect 190128 93160 190340 93644
rect 195024 93638 195236 93644
rect 195024 93574 195030 93638
rect 195094 93574 195236 93638
rect 195024 93502 195236 93574
rect 195024 93438 195166 93502
rect 195230 93438 195236 93502
rect 195024 93432 195236 93438
rect 195432 93638 195644 93644
rect 195432 93574 195438 93638
rect 195502 93574 195644 93638
rect 195432 93502 195644 93574
rect 195432 93438 195574 93502
rect 195638 93438 195644 93502
rect 195432 93432 195644 93438
rect 195840 93638 196460 93644
rect 195840 93574 195982 93638
rect 196046 93574 196460 93638
rect 195840 93568 196460 93574
rect 195840 93432 196052 93568
rect 196248 93432 196460 93568
rect 195840 93372 195916 93432
rect 196384 93372 196460 93432
rect 195024 93230 195236 93236
rect 195024 93166 195166 93230
rect 195230 93166 195236 93230
rect 28424 93100 28500 93160
rect 190128 93100 190204 93160
rect 23392 93030 23398 93094
rect 23462 93030 23604 93094
rect 23392 93024 23604 93030
rect 21760 92964 21836 93024
rect 22576 92964 22652 93024
rect 1632 92932 1844 92964
rect 1632 92876 1702 92932
rect 1758 92876 1844 92932
rect 1632 92828 1844 92876
rect 1224 92822 1844 92828
rect 1224 92758 1230 92822
rect 1294 92758 1844 92822
rect 1224 92752 1844 92758
rect 21760 92822 21972 92964
rect 22304 92888 22652 92964
rect 28288 92888 28636 93100
rect 190128 92958 190340 93100
rect 195024 93094 195236 93166
rect 195024 93030 195030 93094
rect 195094 93030 195236 93094
rect 195024 93024 195236 93030
rect 195432 93230 195644 93236
rect 195432 93166 195574 93230
rect 195638 93166 195644 93230
rect 195432 93094 195644 93166
rect 195432 93030 195574 93094
rect 195638 93030 195644 93094
rect 195432 93024 195644 93030
rect 195840 93024 196052 93372
rect 196248 93024 196460 93372
rect 196656 93432 196868 93780
rect 196656 93372 196732 93432
rect 196656 93024 196868 93372
rect 196248 92964 196324 93024
rect 196792 92964 196868 93024
rect 190128 92894 190270 92958
rect 190334 92894 190340 92958
rect 190128 92888 190340 92894
rect 22304 92828 22380 92888
rect 28424 92828 28500 92888
rect 190264 92828 190340 92888
rect 195976 92888 196324 92964
rect 195976 92828 196052 92888
rect 21760 92758 21902 92822
rect 21966 92758 21972 92822
rect 21760 92752 21972 92758
rect 22168 92752 22788 92828
rect 22168 92616 22380 92752
rect 22576 92616 22788 92752
rect 22168 92556 22244 92616
rect 22712 92556 22788 92616
rect 21760 92550 21972 92556
rect 21760 92486 21902 92550
rect 21966 92486 21972 92550
rect 21760 92414 21972 92486
rect 21760 92350 21766 92414
rect 21830 92350 21972 92414
rect 21760 92344 21972 92350
rect 22168 92420 22380 92556
rect 22168 92414 22516 92420
rect 22168 92350 22446 92414
rect 22510 92350 22516 92414
rect 22168 92344 22516 92350
rect 22576 92344 22788 92556
rect 22984 92822 23196 92828
rect 22984 92758 23126 92822
rect 23190 92758 23196 92822
rect 22984 92616 23196 92758
rect 23392 92822 23604 92828
rect 23392 92758 23398 92822
rect 23462 92758 23604 92822
rect 23392 92616 23604 92758
rect 22984 92556 23060 92616
rect 23392 92556 23468 92616
rect 22984 92208 23196 92556
rect 23392 92208 23604 92556
rect 28288 92550 28636 92828
rect 28288 92486 28566 92550
rect 28630 92486 28636 92550
rect 28288 92480 28636 92486
rect 190128 92686 190340 92828
rect 190128 92622 190270 92686
rect 190334 92622 190340 92686
rect 190128 92550 190340 92622
rect 190128 92486 190134 92550
rect 190198 92486 190340 92550
rect 190128 92480 190340 92486
rect 195024 92822 195236 92828
rect 195024 92758 195030 92822
rect 195094 92758 195236 92822
rect 195024 92616 195236 92758
rect 195432 92822 195644 92828
rect 195432 92758 195574 92822
rect 195638 92758 195644 92822
rect 195432 92616 195644 92758
rect 195840 92752 196460 92828
rect 196656 92822 196868 92964
rect 196656 92758 196798 92822
rect 196862 92758 196868 92822
rect 196656 92752 196868 92758
rect 216784 92958 217540 92964
rect 216784 92932 217470 92958
rect 216784 92876 216908 92932
rect 216964 92894 217470 92932
rect 217534 92894 217540 92958
rect 216964 92888 217540 92894
rect 216964 92876 216996 92888
rect 216784 92752 216996 92876
rect 195840 92692 196052 92752
rect 195840 92616 196188 92692
rect 196248 92616 196460 92752
rect 195024 92556 195100 92616
rect 195568 92556 195644 92616
rect 195976 92556 196052 92616
rect 23120 92148 23196 92208
rect 23528 92148 23604 92208
rect 21760 92142 21972 92148
rect 21760 92078 21766 92142
rect 21830 92078 21972 92142
rect 21760 92006 21972 92078
rect 21760 91942 21766 92006
rect 21830 91942 21972 92006
rect 21760 91936 21972 91942
rect 22168 91800 22380 92148
rect 22478 92142 22788 92148
rect 22440 92078 22446 92142
rect 22510 92078 22788 92142
rect 22478 92072 22788 92078
rect 22576 91876 22788 92072
rect 22984 92006 23196 92148
rect 22984 91942 22990 92006
rect 23054 91942 23196 92006
rect 22984 91936 23196 91942
rect 23392 92006 23604 92148
rect 23392 91942 23534 92006
rect 23598 91942 23604 92006
rect 23392 91936 23604 91942
rect 28288 92278 28636 92284
rect 28288 92214 28566 92278
rect 28630 92214 28636 92278
rect 28288 91936 28636 92214
rect 190128 92278 190340 92284
rect 190128 92214 190134 92278
rect 190198 92214 190340 92278
rect 190128 91936 190340 92214
rect 195024 92208 195236 92556
rect 195432 92208 195644 92556
rect 195840 92420 196052 92556
rect 196112 92556 196188 92616
rect 196112 92480 196460 92556
rect 195840 92414 196188 92420
rect 195840 92350 196118 92414
rect 196182 92350 196188 92414
rect 195840 92344 196188 92350
rect 196248 92344 196460 92480
rect 196656 92550 196868 92556
rect 196656 92486 196798 92550
rect 196862 92486 196868 92550
rect 196656 92414 196868 92486
rect 196656 92350 196662 92414
rect 196726 92350 196868 92414
rect 196656 92344 196868 92350
rect 195160 92148 195236 92208
rect 195568 92148 195644 92208
rect 195024 92006 195236 92148
rect 195024 91942 195166 92006
rect 195230 91942 195236 92006
rect 195024 91936 195236 91942
rect 195432 92006 195644 92148
rect 195432 91942 195438 92006
rect 195502 91942 195644 92006
rect 195432 91936 195644 91942
rect 22478 91870 22788 91876
rect 22440 91806 22446 91870
rect 22510 91806 22788 91870
rect 22478 91800 22788 91806
rect 28288 91876 28364 91936
rect 190264 91876 190340 91936
rect 22304 91740 22380 91800
rect 21760 91734 21972 91740
rect 21760 91670 21766 91734
rect 21830 91670 21972 91734
rect 21760 91598 21972 91670
rect 21760 91534 21902 91598
rect 21966 91534 21972 91598
rect 21760 91528 21972 91534
rect 22168 91664 22788 91740
rect 22168 91604 22380 91664
rect 22168 91598 22516 91604
rect 22168 91534 22446 91598
rect 22510 91534 22516 91598
rect 22168 91528 22516 91534
rect 22576 91598 22788 91664
rect 22576 91534 22718 91598
rect 22782 91534 22788 91598
rect 22576 91528 22788 91534
rect 22984 91734 23196 91740
rect 22984 91670 22990 91734
rect 23054 91670 23196 91734
rect 22984 91598 23196 91670
rect 22984 91534 23126 91598
rect 23190 91534 23196 91598
rect 22984 91528 23196 91534
rect 23392 91734 23604 91740
rect 23392 91670 23534 91734
rect 23598 91670 23604 91734
rect 23392 91598 23604 91670
rect 28288 91664 28636 91876
rect 190128 91664 190340 91876
rect 195840 91800 196052 92148
rect 196150 92142 196460 92148
rect 196112 92078 196118 92142
rect 196182 92078 196460 92142
rect 196150 92072 196460 92078
rect 196248 91876 196460 92072
rect 196656 92142 196868 92148
rect 196656 92078 196662 92142
rect 196726 92078 196868 92142
rect 196656 92006 196868 92078
rect 196656 91942 196798 92006
rect 196862 91942 196868 92006
rect 196656 91936 196868 91942
rect 195976 91740 196052 91800
rect 196112 91800 196460 91876
rect 196112 91740 196188 91800
rect 28424 91604 28500 91664
rect 190264 91604 190340 91664
rect 23392 91534 23534 91598
rect 23598 91534 23604 91598
rect 23392 91528 23604 91534
rect 1632 91252 1844 91332
rect 1632 91196 1702 91252
rect 1758 91196 1844 91252
rect 1224 91190 1844 91196
rect 1224 91126 1230 91190
rect 1294 91126 1844 91190
rect 1224 91120 1844 91126
rect 21760 91326 21972 91332
rect 21760 91262 21902 91326
rect 21966 91262 21972 91326
rect 21760 91190 21972 91262
rect 21760 91126 21766 91190
rect 21830 91126 21972 91190
rect 21760 91120 21972 91126
rect 22168 91196 22380 91332
rect 22576 91326 22788 91332
rect 22576 91262 22718 91326
rect 22782 91262 22788 91326
rect 22576 91196 22788 91262
rect 22168 91190 22788 91196
rect 22168 91126 22174 91190
rect 22238 91126 22582 91190
rect 22646 91126 22788 91190
rect 22168 91120 22788 91126
rect 22984 91326 23196 91332
rect 22984 91262 23126 91326
rect 23190 91262 23196 91326
rect 22984 91190 23196 91262
rect 22984 91126 22990 91190
rect 23054 91126 23196 91190
rect 22984 91120 23196 91126
rect 23392 91326 23604 91332
rect 23392 91262 23534 91326
rect 23598 91262 23604 91326
rect 23392 91190 23604 91262
rect 23392 91126 23534 91190
rect 23598 91126 23604 91190
rect 23392 91120 23604 91126
rect 28288 91120 28636 91604
rect 190128 91120 190340 91604
rect 195024 91734 195236 91740
rect 195024 91670 195166 91734
rect 195230 91670 195236 91734
rect 195024 91598 195236 91670
rect 195024 91534 195030 91598
rect 195094 91534 195236 91598
rect 195024 91528 195236 91534
rect 195432 91734 195644 91740
rect 195432 91670 195438 91734
rect 195502 91670 195644 91734
rect 195432 91598 195644 91670
rect 195432 91534 195438 91598
rect 195502 91534 195644 91598
rect 195432 91528 195644 91534
rect 195840 91664 196188 91740
rect 196248 91740 196324 91800
rect 195840 91528 196052 91664
rect 196248 91598 196460 91740
rect 196248 91534 196254 91598
rect 196318 91534 196460 91598
rect 196248 91528 196460 91534
rect 196656 91734 196868 91740
rect 196656 91670 196798 91734
rect 196862 91670 196868 91734
rect 196656 91598 196868 91670
rect 196656 91534 196662 91598
rect 196726 91534 196868 91598
rect 196656 91528 196868 91534
rect 195024 91326 195236 91332
rect 195024 91262 195030 91326
rect 195094 91262 195236 91326
rect 195024 91190 195236 91262
rect 195024 91126 195166 91190
rect 195230 91126 195236 91190
rect 195024 91120 195236 91126
rect 195432 91326 195644 91332
rect 195432 91262 195438 91326
rect 195502 91262 195644 91326
rect 195432 91190 195644 91262
rect 195432 91126 195574 91190
rect 195638 91126 195644 91190
rect 195432 91120 195644 91126
rect 195840 91326 196460 91332
rect 195840 91262 196254 91326
rect 196318 91262 196460 91326
rect 195840 91256 196460 91262
rect 195840 91190 196052 91256
rect 195840 91126 195846 91190
rect 195910 91126 196052 91190
rect 195840 91120 196052 91126
rect 196248 91120 196460 91256
rect 196656 91326 196868 91332
rect 196656 91262 196662 91326
rect 196726 91262 196868 91326
rect 196656 91190 196868 91262
rect 196656 91126 196662 91190
rect 196726 91126 196868 91190
rect 196656 91120 196868 91126
rect 216784 91326 217540 91332
rect 216784 91262 217470 91326
rect 217534 91262 217540 91326
rect 216784 91256 217540 91262
rect 216784 91252 216996 91256
rect 216784 91196 216908 91252
rect 216964 91196 216996 91252
rect 216784 91120 216996 91196
rect 28288 91060 28364 91120
rect 190128 91060 190204 91120
rect 21760 90918 21972 90924
rect 21760 90854 21766 90918
rect 21830 90854 21972 90918
rect 21760 90782 21972 90854
rect 21760 90718 21902 90782
rect 21966 90718 21972 90782
rect 21760 90712 21972 90718
rect 22168 90918 22380 90924
rect 22168 90854 22174 90918
rect 22238 90854 22380 90918
rect 22168 90712 22380 90854
rect 22576 90918 22788 90924
rect 22576 90854 22582 90918
rect 22646 90854 22788 90918
rect 22576 90782 22788 90854
rect 22576 90718 22718 90782
rect 22782 90718 22788 90782
rect 22576 90712 22788 90718
rect 22984 90918 23196 90924
rect 22984 90854 22990 90918
rect 23054 90854 23196 90918
rect 22984 90782 23196 90854
rect 22984 90718 23126 90782
rect 23190 90718 23196 90782
rect 22984 90712 23196 90718
rect 23392 90918 23604 90924
rect 23392 90854 23534 90918
rect 23598 90854 23604 90918
rect 23392 90782 23604 90854
rect 23392 90718 23398 90782
rect 23462 90718 23604 90782
rect 23392 90712 23604 90718
rect 28288 90848 28636 91060
rect 190128 90848 190340 91060
rect 28288 90788 28364 90848
rect 190264 90788 190340 90848
rect 28288 90576 28636 90788
rect 190128 90576 190340 90788
rect 195024 90918 195236 90924
rect 195024 90854 195166 90918
rect 195230 90854 195236 90918
rect 195024 90782 195236 90854
rect 195024 90718 195030 90782
rect 195094 90718 195236 90782
rect 195024 90712 195236 90718
rect 195432 90918 195644 90924
rect 195432 90854 195574 90918
rect 195638 90854 195644 90918
rect 195432 90782 195644 90854
rect 195432 90718 195574 90782
rect 195638 90718 195644 90782
rect 195432 90712 195644 90718
rect 195840 90918 196460 90924
rect 195840 90854 195846 90918
rect 195910 90854 196460 90918
rect 195840 90848 196460 90854
rect 195840 90712 196052 90848
rect 196248 90788 196460 90848
rect 196150 90782 196460 90788
rect 196112 90718 196118 90782
rect 196182 90718 196460 90782
rect 196150 90712 196460 90718
rect 196656 90918 196868 90924
rect 196656 90854 196662 90918
rect 196726 90854 196868 90918
rect 196656 90782 196868 90854
rect 196656 90718 196798 90782
rect 196862 90718 196868 90782
rect 196656 90712 196868 90718
rect 195976 90652 196052 90712
rect 195976 90576 196324 90652
rect 28560 90516 28636 90576
rect 190264 90516 190340 90576
rect 196248 90516 196324 90576
rect 21760 90510 21972 90516
rect 21760 90446 21902 90510
rect 21966 90446 21972 90510
rect 21760 90374 21972 90446
rect 21760 90310 21902 90374
rect 21966 90310 21972 90374
rect 21760 90304 21972 90310
rect 22168 90380 22380 90516
rect 22576 90510 22788 90516
rect 22576 90446 22718 90510
rect 22782 90446 22788 90510
rect 22576 90380 22788 90446
rect 22168 90374 22788 90380
rect 22168 90310 22310 90374
rect 22374 90310 22788 90374
rect 22168 90304 22788 90310
rect 22984 90510 23196 90516
rect 22984 90446 23126 90510
rect 23190 90446 23196 90510
rect 22984 90374 23196 90446
rect 22984 90310 22990 90374
rect 23054 90310 23196 90374
rect 22984 90304 23196 90310
rect 23392 90510 23604 90516
rect 23392 90446 23398 90510
rect 23462 90446 23604 90510
rect 23392 90374 23604 90446
rect 23392 90310 23534 90374
rect 23598 90310 23604 90374
rect 23392 90304 23604 90310
rect 28288 90304 28636 90516
rect 190128 90304 190340 90516
rect 195024 90510 195236 90516
rect 195024 90446 195030 90510
rect 195094 90446 195236 90510
rect 195024 90374 195236 90446
rect 195024 90310 195030 90374
rect 195094 90310 195236 90374
rect 195024 90304 195236 90310
rect 195432 90510 195644 90516
rect 195432 90446 195574 90510
rect 195638 90446 195644 90510
rect 195432 90374 195644 90446
rect 195432 90310 195574 90374
rect 195638 90310 195644 90374
rect 195432 90304 195644 90310
rect 195840 90510 196188 90516
rect 195840 90446 196118 90510
rect 196182 90446 196188 90510
rect 195840 90440 196188 90446
rect 195840 90374 196052 90440
rect 195840 90310 195846 90374
rect 195910 90310 196052 90374
rect 195840 90304 196052 90310
rect 196248 90304 196460 90516
rect 196656 90510 196868 90516
rect 196656 90446 196798 90510
rect 196862 90446 196868 90510
rect 196656 90374 196868 90446
rect 196656 90310 196798 90374
rect 196862 90310 196868 90374
rect 196656 90304 196868 90310
rect 28424 90244 28500 90304
rect 190264 90244 190340 90304
rect 21760 90102 21972 90108
rect 21760 90038 21902 90102
rect 21966 90038 21972 90102
rect 21760 89896 21972 90038
rect 22168 90102 22380 90108
rect 22168 90038 22310 90102
rect 22374 90038 22380 90102
rect 22168 89966 22380 90038
rect 22168 89902 22174 89966
rect 22238 89902 22380 89966
rect 22168 89896 22380 89902
rect 22576 89966 22788 90108
rect 22576 89902 22718 89966
rect 22782 89902 22788 89966
rect 22576 89896 22788 89902
rect 22984 90102 23196 90108
rect 22984 90038 22990 90102
rect 23054 90038 23196 90102
rect 22984 89966 23196 90038
rect 22984 89902 22990 89966
rect 23054 89902 23196 89966
rect 22984 89896 23196 89902
rect 23392 90102 23604 90108
rect 23392 90038 23534 90102
rect 23598 90038 23604 90102
rect 23392 89966 23604 90038
rect 23392 89902 23534 89966
rect 23598 89902 23604 89966
rect 23392 89896 23604 89902
rect 28288 90032 28636 90244
rect 190128 90032 190340 90244
rect 195024 90102 195236 90108
rect 195024 90038 195030 90102
rect 195094 90038 195236 90102
rect 28288 89972 28364 90032
rect 190128 89972 190204 90032
rect 21760 89836 21836 89896
rect 1632 89572 1844 89700
rect 1632 89564 1702 89572
rect 1224 89558 1702 89564
rect 1224 89494 1230 89558
rect 1294 89516 1702 89558
rect 1758 89516 1844 89572
rect 1294 89494 1844 89516
rect 1224 89488 1844 89494
rect 21760 89488 21972 89836
rect 28288 89830 28636 89972
rect 28288 89766 28566 89830
rect 28630 89766 28636 89830
rect 28288 89760 28636 89766
rect 28560 89700 28636 89760
rect 22168 89694 22380 89700
rect 22168 89630 22174 89694
rect 22238 89630 22380 89694
rect 22168 89564 22380 89630
rect 22576 89694 22788 89700
rect 22576 89630 22718 89694
rect 22782 89630 22788 89694
rect 22576 89564 22788 89630
rect 22168 89488 22788 89564
rect 22984 89694 23196 89700
rect 22984 89630 22990 89694
rect 23054 89630 23196 89694
rect 22984 89558 23196 89630
rect 22984 89494 23126 89558
rect 23190 89494 23196 89558
rect 22984 89488 23196 89494
rect 23392 89694 23604 89700
rect 23392 89630 23534 89694
rect 23598 89630 23604 89694
rect 23392 89558 23604 89630
rect 23392 89494 23398 89558
rect 23462 89494 23604 89558
rect 23392 89488 23604 89494
rect 28288 89558 28636 89700
rect 28288 89494 28566 89558
rect 28630 89494 28636 89558
rect 21760 89428 21836 89488
rect 22304 89428 22380 89488
rect 22712 89428 22788 89488
rect 21760 89080 21972 89428
rect 22168 89150 22380 89428
rect 22168 89086 22174 89150
rect 22238 89086 22380 89150
rect 22168 89080 22380 89086
rect 22576 89080 22788 89428
rect 22984 89286 23196 89292
rect 22984 89222 23126 89286
rect 23190 89222 23196 89286
rect 22984 89150 23196 89222
rect 22984 89086 23126 89150
rect 23190 89086 23196 89150
rect 22984 89080 23196 89086
rect 23392 89286 23604 89292
rect 23392 89222 23398 89286
rect 23462 89222 23604 89286
rect 23392 89150 23604 89222
rect 28288 89216 28636 89494
rect 28560 89156 28636 89216
rect 23392 89086 23534 89150
rect 23598 89086 23604 89150
rect 23392 89080 23604 89086
rect 21896 89020 21972 89080
rect 21760 88878 21972 89020
rect 28288 88944 28636 89156
rect 190128 89760 190340 89972
rect 195024 89966 195236 90038
rect 195024 89902 195030 89966
rect 195094 89902 195236 89966
rect 195024 89896 195236 89902
rect 195432 90102 195644 90108
rect 195432 90038 195574 90102
rect 195638 90038 195644 90102
rect 195432 89966 195644 90038
rect 195432 89902 195438 89966
rect 195502 89902 195644 89966
rect 195432 89896 195644 89902
rect 195840 90102 196052 90108
rect 195840 90038 195846 90102
rect 195910 90038 196052 90102
rect 195840 89966 196052 90038
rect 196248 89972 196460 90108
rect 196150 89966 196460 89972
rect 195840 89902 195982 89966
rect 196046 89902 196052 89966
rect 196112 89902 196118 89966
rect 196182 89902 196460 89966
rect 195840 89896 196052 89902
rect 196150 89896 196460 89902
rect 196656 90102 196868 90108
rect 196656 90038 196798 90102
rect 196862 90038 196868 90102
rect 196656 89896 196868 90038
rect 196656 89836 196732 89896
rect 190128 89700 190204 89760
rect 190128 89216 190340 89700
rect 195024 89694 195236 89700
rect 195024 89630 195030 89694
rect 195094 89630 195236 89694
rect 195024 89558 195236 89630
rect 195024 89494 195030 89558
rect 195094 89494 195236 89558
rect 195024 89488 195236 89494
rect 195432 89694 195644 89700
rect 195432 89630 195438 89694
rect 195502 89630 195644 89694
rect 195432 89558 195644 89630
rect 195432 89494 195438 89558
rect 195502 89494 195644 89558
rect 195432 89488 195644 89494
rect 195840 89694 196188 89700
rect 195840 89630 195982 89694
rect 196046 89630 196118 89694
rect 196182 89630 196188 89694
rect 195840 89624 196188 89630
rect 195840 89564 196052 89624
rect 195840 89488 196188 89564
rect 196248 89488 196460 89700
rect 196656 89488 196868 89836
rect 216784 89694 217540 89700
rect 216784 89630 217470 89694
rect 217534 89630 217540 89694
rect 216784 89624 217540 89630
rect 216784 89572 216996 89624
rect 216784 89516 216908 89572
rect 216964 89516 216996 89572
rect 216784 89488 216996 89516
rect 196112 89428 196188 89488
rect 196384 89428 196460 89488
rect 196792 89428 196868 89488
rect 195024 89286 195236 89292
rect 195024 89222 195030 89286
rect 195094 89222 195236 89286
rect 190128 89156 190204 89216
rect 190128 89014 190340 89156
rect 195024 89150 195236 89222
rect 195024 89086 195166 89150
rect 195230 89086 195236 89150
rect 195024 89080 195236 89086
rect 195432 89286 195644 89292
rect 195432 89222 195438 89286
rect 195502 89222 195644 89286
rect 195432 89150 195644 89222
rect 195432 89086 195438 89150
rect 195502 89086 195644 89150
rect 195432 89080 195644 89086
rect 195840 89150 196052 89428
rect 196112 89352 196460 89428
rect 195840 89086 195982 89150
rect 196046 89086 196052 89150
rect 195840 89080 196052 89086
rect 196248 89150 196460 89352
rect 196248 89086 196254 89150
rect 196318 89086 196460 89150
rect 196248 89080 196460 89086
rect 196656 89080 196868 89428
rect 190128 88950 190134 89014
rect 190198 88950 190340 89014
rect 190128 88944 190340 88950
rect 196656 89020 196732 89080
rect 28424 88884 28500 88944
rect 190128 88884 190204 88944
rect 21760 88814 21902 88878
rect 21966 88814 21972 88878
rect 21760 88808 21972 88814
rect 22168 88878 22380 88884
rect 22168 88814 22174 88878
rect 22238 88814 22380 88878
rect 22168 88672 22380 88814
rect 22576 88672 22788 88884
rect 22984 88878 23196 88884
rect 22984 88814 23126 88878
rect 23190 88814 23196 88878
rect 22984 88672 23196 88814
rect 23392 88878 23604 88884
rect 23392 88814 23534 88878
rect 23598 88814 23604 88878
rect 23392 88672 23604 88814
rect 22304 88612 22380 88672
rect 22712 88612 22788 88672
rect 23120 88612 23196 88672
rect 23528 88612 23604 88672
rect 21760 88606 21972 88612
rect 21760 88542 21902 88606
rect 21966 88542 21972 88606
rect 21760 88470 21972 88542
rect 21760 88406 21902 88470
rect 21966 88406 21972 88470
rect 21760 88400 21972 88406
rect 22168 88470 22380 88612
rect 22576 88476 22788 88612
rect 22478 88470 22788 88476
rect 22168 88406 22174 88470
rect 22238 88406 22380 88470
rect 22440 88406 22446 88470
rect 22510 88406 22788 88470
rect 22168 88400 22380 88406
rect 22478 88400 22788 88406
rect 22984 88264 23196 88612
rect 23392 88264 23604 88612
rect 28288 88606 28636 88884
rect 28288 88542 28430 88606
rect 28494 88542 28636 88606
rect 28288 88536 28636 88542
rect 190128 88742 190340 88884
rect 190128 88678 190134 88742
rect 190198 88678 190270 88742
rect 190334 88678 190340 88742
rect 190128 88536 190340 88678
rect 195024 88878 195236 88884
rect 195024 88814 195166 88878
rect 195230 88814 195236 88878
rect 195024 88672 195236 88814
rect 195432 88878 195644 88884
rect 195432 88814 195438 88878
rect 195502 88814 195644 88878
rect 195432 88672 195644 88814
rect 195840 88878 196052 88884
rect 195840 88814 195982 88878
rect 196046 88814 196052 88878
rect 195840 88672 196052 88814
rect 196248 88878 196460 88884
rect 196248 88814 196254 88878
rect 196318 88814 196460 88878
rect 196248 88672 196460 88814
rect 196656 88878 196868 89020
rect 196656 88814 196662 88878
rect 196726 88814 196868 88878
rect 196656 88808 196868 88814
rect 195024 88612 195100 88672
rect 195432 88612 195508 88672
rect 195840 88612 195916 88672
rect 196248 88612 196324 88672
rect 22984 88204 23060 88264
rect 23528 88204 23604 88264
rect 21760 88198 21972 88204
rect 21760 88134 21902 88198
rect 21966 88134 21972 88198
rect 21760 88062 21972 88134
rect 21760 87998 21766 88062
rect 21830 87998 21972 88062
rect 21760 87992 21972 87998
rect 22168 88198 22516 88204
rect 22168 88134 22174 88198
rect 22238 88134 22446 88198
rect 22510 88134 22516 88198
rect 22168 88128 22516 88134
rect 22168 88068 22380 88128
rect 22576 88068 22788 88204
rect 22168 87992 22788 88068
rect 1224 87926 1844 87932
rect 1224 87862 1230 87926
rect 1294 87892 1844 87926
rect 1294 87862 1702 87892
rect 1224 87856 1702 87862
rect 1632 87836 1702 87856
rect 1758 87836 1844 87892
rect 22168 87856 22380 87992
rect 22576 87856 22788 87992
rect 22984 87856 23196 88204
rect 23392 87856 23604 88204
rect 1632 87720 1844 87836
rect 22576 87796 22652 87856
rect 23120 87796 23196 87856
rect 23528 87796 23604 87856
rect 21760 87790 21972 87796
rect 21760 87726 21766 87790
rect 21830 87726 21972 87790
rect 21760 87654 21972 87726
rect 21760 87590 21766 87654
rect 21830 87590 21972 87654
rect 21760 87584 21972 87590
rect 22168 87654 22380 87796
rect 22576 87660 22788 87796
rect 22478 87654 22788 87660
rect 22168 87590 22310 87654
rect 22374 87590 22380 87654
rect 22440 87590 22446 87654
rect 22510 87590 22582 87654
rect 22646 87590 22788 87654
rect 22168 87584 22380 87590
rect 22478 87584 22788 87590
rect 22984 87654 23196 87796
rect 22984 87590 23126 87654
rect 23190 87590 23196 87654
rect 22984 87584 23196 87590
rect 23392 87654 23604 87796
rect 28288 88334 28636 88340
rect 28288 88270 28430 88334
rect 28494 88270 28636 88334
rect 28288 88198 28636 88270
rect 28288 88134 28566 88198
rect 28630 88134 28636 88198
rect 28288 87926 28636 88134
rect 28288 87862 28566 87926
rect 28630 87862 28636 87926
rect 28288 87720 28636 87862
rect 190128 88334 190340 88340
rect 190128 88270 190270 88334
rect 190334 88270 190340 88334
rect 190128 87926 190340 88270
rect 190128 87862 190134 87926
rect 190198 87862 190340 87926
rect 190128 87720 190340 87862
rect 195024 88264 195236 88612
rect 195432 88264 195644 88612
rect 195840 88536 196460 88612
rect 195840 88476 196052 88536
rect 195840 88470 196188 88476
rect 195840 88406 196118 88470
rect 196182 88406 196188 88470
rect 195840 88400 196188 88406
rect 196248 88400 196460 88536
rect 196656 88606 196868 88612
rect 196656 88542 196662 88606
rect 196726 88542 196868 88606
rect 196656 88470 196868 88542
rect 196656 88406 196798 88470
rect 196862 88406 196868 88470
rect 196656 88400 196868 88406
rect 195024 88204 195100 88264
rect 195568 88204 195644 88264
rect 195024 87856 195236 88204
rect 195432 87856 195644 88204
rect 195160 87796 195236 87856
rect 195568 87796 195644 87856
rect 28424 87660 28500 87720
rect 190128 87660 190204 87720
rect 23392 87590 23534 87654
rect 23598 87590 23604 87654
rect 23392 87584 23604 87590
rect 21760 87382 21972 87388
rect 21760 87318 21766 87382
rect 21830 87318 21972 87382
rect 21760 87246 21972 87318
rect 21760 87182 21766 87246
rect 21830 87182 21972 87246
rect 21760 87176 21972 87182
rect 22168 87382 22516 87388
rect 22168 87318 22310 87382
rect 22374 87318 22446 87382
rect 22510 87318 22516 87382
rect 22168 87312 22516 87318
rect 22576 87382 22788 87388
rect 22576 87318 22582 87382
rect 22646 87318 22788 87382
rect 22168 87252 22380 87312
rect 22168 87246 22516 87252
rect 22168 87182 22174 87246
rect 22238 87182 22446 87246
rect 22510 87182 22516 87246
rect 22168 87176 22516 87182
rect 22576 87176 22788 87318
rect 22984 87382 23196 87388
rect 22984 87318 23126 87382
rect 23190 87318 23196 87382
rect 22984 87246 23196 87318
rect 22984 87182 22990 87246
rect 23054 87182 23196 87246
rect 22984 87176 23196 87182
rect 23392 87382 23604 87388
rect 23392 87318 23534 87382
rect 23598 87318 23604 87382
rect 23392 87246 23604 87318
rect 23392 87182 23398 87246
rect 23462 87182 23604 87246
rect 23392 87176 23604 87182
rect 28288 87382 28636 87660
rect 28288 87318 28430 87382
rect 28494 87318 28636 87382
rect 28288 87176 28636 87318
rect 190128 87654 190340 87660
rect 190128 87590 190134 87654
rect 190198 87590 190340 87654
rect 190128 87382 190340 87590
rect 195024 87654 195236 87796
rect 195024 87590 195030 87654
rect 195094 87590 195236 87654
rect 195024 87584 195236 87590
rect 195432 87654 195644 87796
rect 195432 87590 195574 87654
rect 195638 87590 195644 87654
rect 195432 87584 195644 87590
rect 195840 87856 196052 88204
rect 196150 88198 196460 88204
rect 196112 88134 196118 88198
rect 196182 88134 196460 88198
rect 196150 88128 196460 88134
rect 196248 87856 196460 88128
rect 196656 88198 196868 88204
rect 196656 88134 196798 88198
rect 196862 88134 196868 88198
rect 196656 88062 196868 88134
rect 196656 87998 196662 88062
rect 196726 87998 196868 88062
rect 196656 87992 196868 87998
rect 216784 87892 216996 87932
rect 195840 87796 195916 87856
rect 196248 87796 196324 87856
rect 216784 87836 216908 87892
rect 216964 87836 216996 87892
rect 216784 87796 216996 87836
rect 195840 87654 196052 87796
rect 195840 87590 195982 87654
rect 196046 87590 196052 87654
rect 195840 87584 196052 87590
rect 196248 87654 196460 87796
rect 196248 87590 196390 87654
rect 196454 87590 196460 87654
rect 196248 87584 196460 87590
rect 196656 87790 196868 87796
rect 196656 87726 196662 87790
rect 196726 87726 196868 87790
rect 196656 87654 196868 87726
rect 216784 87790 217540 87796
rect 216784 87726 217470 87790
rect 217534 87726 217540 87790
rect 216784 87720 217540 87726
rect 196656 87590 196662 87654
rect 196726 87590 196868 87654
rect 196656 87584 196868 87590
rect 190128 87318 190270 87382
rect 190334 87318 190340 87382
rect 190128 87176 190340 87318
rect 195024 87382 195236 87388
rect 195024 87318 195030 87382
rect 195094 87318 195236 87382
rect 195024 87246 195236 87318
rect 195024 87182 195030 87246
rect 195094 87182 195236 87246
rect 195024 87176 195236 87182
rect 195432 87382 195644 87388
rect 195432 87318 195574 87382
rect 195638 87318 195644 87382
rect 195432 87246 195644 87318
rect 195432 87182 195438 87246
rect 195502 87182 195644 87246
rect 195432 87176 195644 87182
rect 195840 87382 196460 87388
rect 195840 87318 195982 87382
rect 196046 87318 196390 87382
rect 196454 87318 196460 87382
rect 195840 87312 196460 87318
rect 195840 87176 196052 87312
rect 196248 87246 196460 87312
rect 196248 87182 196254 87246
rect 196318 87182 196460 87246
rect 196248 87176 196460 87182
rect 196656 87382 196868 87388
rect 196656 87318 196662 87382
rect 196726 87318 196868 87382
rect 196656 87246 196868 87318
rect 196656 87182 196662 87246
rect 196726 87182 196868 87246
rect 196656 87176 196868 87182
rect 28424 87116 28500 87176
rect 190264 87116 190340 87176
rect 28288 87110 28636 87116
rect 28288 87046 28430 87110
rect 28494 87046 28636 87110
rect 21760 86974 21972 86980
rect 21760 86910 21766 86974
rect 21830 86910 21972 86974
rect 21760 86838 21972 86910
rect 21760 86774 21766 86838
rect 21830 86774 21972 86838
rect 21760 86768 21972 86774
rect 22168 86974 22380 86980
rect 22478 86974 22788 86980
rect 22168 86910 22174 86974
rect 22238 86910 22380 86974
rect 22440 86910 22446 86974
rect 22510 86910 22788 86974
rect 22168 86768 22380 86910
rect 22478 86904 22788 86910
rect 22576 86838 22788 86904
rect 22576 86774 22582 86838
rect 22646 86774 22788 86838
rect 22576 86768 22788 86774
rect 22984 86974 23196 86980
rect 22984 86910 22990 86974
rect 23054 86910 23196 86974
rect 22984 86838 23196 86910
rect 22984 86774 23126 86838
rect 23190 86774 23196 86838
rect 22984 86768 23196 86774
rect 23392 86974 23604 86980
rect 23392 86910 23398 86974
rect 23462 86910 23604 86974
rect 23392 86838 23604 86910
rect 28288 86904 28636 87046
rect 190128 87110 190340 87116
rect 190128 87046 190270 87110
rect 190334 87046 190340 87110
rect 190128 86904 190340 87046
rect 195024 86974 195236 86980
rect 195024 86910 195030 86974
rect 195094 86910 195236 86974
rect 28424 86844 28500 86904
rect 190128 86844 190204 86904
rect 23392 86774 23534 86838
rect 23598 86774 23604 86838
rect 23392 86768 23604 86774
rect 28288 86632 28636 86844
rect 190128 86632 190340 86844
rect 195024 86838 195236 86910
rect 195024 86774 195166 86838
rect 195230 86774 195236 86838
rect 195024 86768 195236 86774
rect 195432 86974 195644 86980
rect 195432 86910 195438 86974
rect 195502 86910 195644 86974
rect 195432 86838 195644 86910
rect 195432 86774 195574 86838
rect 195638 86774 195644 86838
rect 195432 86768 195644 86774
rect 195840 86838 196052 86980
rect 196248 86974 196460 86980
rect 196248 86910 196254 86974
rect 196318 86910 196460 86974
rect 196248 86844 196460 86910
rect 196150 86838 196460 86844
rect 195840 86774 195846 86838
rect 195910 86774 196052 86838
rect 196112 86774 196118 86838
rect 196182 86774 196460 86838
rect 195840 86768 196052 86774
rect 196150 86768 196460 86774
rect 196656 86974 196868 86980
rect 196656 86910 196662 86974
rect 196726 86910 196868 86974
rect 196656 86838 196868 86910
rect 196656 86774 196662 86838
rect 196726 86774 196868 86838
rect 196656 86768 196868 86774
rect 28288 86572 28364 86632
rect 190128 86572 190204 86632
rect 21760 86566 21972 86572
rect 21760 86502 21766 86566
rect 21830 86502 21972 86566
rect 21760 86430 21972 86502
rect 21760 86366 21902 86430
rect 21966 86366 21972 86430
rect 21760 86360 21972 86366
rect 22168 86436 22380 86572
rect 22576 86566 22788 86572
rect 22576 86502 22582 86566
rect 22646 86502 22788 86566
rect 22576 86436 22788 86502
rect 22168 86430 22788 86436
rect 22168 86366 22310 86430
rect 22374 86366 22788 86430
rect 22168 86360 22788 86366
rect 22984 86566 23196 86572
rect 22984 86502 23126 86566
rect 23190 86502 23196 86566
rect 22984 86430 23196 86502
rect 22984 86366 23126 86430
rect 23190 86366 23196 86430
rect 22984 86360 23196 86366
rect 23392 86566 23604 86572
rect 23392 86502 23534 86566
rect 23598 86502 23604 86566
rect 23392 86430 23604 86502
rect 23392 86366 23398 86430
rect 23462 86366 23604 86430
rect 23392 86360 23604 86366
rect 28288 86360 28636 86572
rect 190128 86360 190340 86572
rect 195024 86566 195236 86572
rect 195024 86502 195166 86566
rect 195230 86502 195236 86566
rect 195024 86430 195236 86502
rect 195024 86366 195030 86430
rect 195094 86366 195236 86430
rect 195024 86360 195236 86366
rect 195432 86566 195644 86572
rect 195432 86502 195574 86566
rect 195638 86502 195644 86566
rect 195432 86430 195644 86502
rect 195432 86366 195438 86430
rect 195502 86366 195644 86430
rect 195432 86360 195644 86366
rect 195840 86566 196188 86572
rect 195840 86502 195846 86566
rect 195910 86502 196118 86566
rect 196182 86502 196188 86566
rect 195840 86496 196188 86502
rect 195840 86436 196052 86496
rect 195840 86430 196188 86436
rect 195840 86366 195982 86430
rect 196046 86366 196118 86430
rect 196182 86366 196188 86430
rect 195840 86360 196188 86366
rect 196248 86360 196460 86572
rect 196656 86566 196868 86572
rect 196656 86502 196662 86566
rect 196726 86502 196868 86566
rect 196656 86430 196868 86502
rect 196656 86366 196798 86430
rect 196862 86366 196868 86430
rect 196656 86360 196868 86366
rect 28288 86300 28364 86360
rect 190264 86300 190340 86360
rect 1224 86294 1844 86300
rect 1224 86230 1230 86294
rect 1294 86230 1844 86294
rect 1224 86224 1844 86230
rect 1632 86212 1844 86224
rect 1632 86156 1702 86212
rect 1758 86156 1844 86212
rect 1632 86088 1844 86156
rect 21760 86158 21972 86164
rect 21760 86094 21902 86158
rect 21966 86094 21972 86158
rect 21760 85952 21972 86094
rect 22168 86158 22380 86164
rect 22168 86094 22310 86158
rect 22374 86094 22380 86158
rect 22168 86028 22380 86094
rect 22576 86028 22788 86164
rect 22168 85952 22788 86028
rect 22984 86158 23196 86164
rect 22984 86094 23126 86158
rect 23190 86094 23196 86158
rect 22984 86022 23196 86094
rect 22984 85958 23126 86022
rect 23190 85958 23196 86022
rect 22984 85952 23196 85958
rect 23392 86158 23604 86164
rect 23392 86094 23398 86158
rect 23462 86094 23604 86158
rect 23392 86022 23604 86094
rect 23392 85958 23398 86022
rect 23462 85958 23604 86022
rect 23392 85952 23604 85958
rect 28288 86088 28636 86300
rect 190128 86088 190340 86300
rect 195976 86300 196052 86360
rect 196248 86300 196324 86360
rect 195976 86224 196324 86300
rect 216784 86212 216996 86300
rect 28288 86028 28364 86088
rect 190264 86028 190340 86088
rect 21896 85892 21972 85952
rect 21760 85614 21972 85892
rect 22304 85892 22380 85952
rect 22304 85816 22652 85892
rect 28288 85816 28636 86028
rect 190128 85816 190340 86028
rect 195024 86158 195236 86164
rect 195024 86094 195030 86158
rect 195094 86094 195236 86158
rect 195024 86022 195236 86094
rect 195024 85958 195030 86022
rect 195094 85958 195236 86022
rect 195024 85952 195236 85958
rect 195432 86158 195644 86164
rect 195432 86094 195438 86158
rect 195502 86094 195644 86158
rect 195432 86022 195644 86094
rect 195432 85958 195574 86022
rect 195638 85958 195644 86022
rect 195432 85952 195644 85958
rect 195840 86158 196052 86164
rect 196150 86158 196460 86164
rect 195840 86094 195982 86158
rect 196046 86094 196052 86158
rect 196112 86094 196118 86158
rect 196182 86094 196460 86158
rect 195840 86022 196052 86094
rect 196150 86088 196460 86094
rect 195840 85958 195846 86022
rect 195910 85958 196052 86022
rect 195840 85952 196052 85958
rect 196248 85952 196460 86088
rect 196656 86158 196868 86164
rect 196656 86094 196798 86158
rect 196862 86094 196868 86158
rect 196656 85952 196868 86094
rect 216784 86156 216908 86212
rect 216964 86164 216996 86212
rect 216964 86158 217540 86164
rect 216964 86156 217470 86158
rect 216784 86094 217470 86156
rect 217534 86094 217540 86158
rect 216784 86088 217540 86094
rect 196792 85892 196868 85952
rect 22576 85756 22652 85816
rect 28424 85756 28500 85816
rect 190128 85756 190204 85816
rect 21760 85550 21902 85614
rect 21966 85550 21972 85614
rect 21760 85544 21972 85550
rect 22168 85614 22380 85756
rect 22168 85550 22174 85614
rect 22238 85550 22380 85614
rect 22168 85544 22380 85550
rect 22576 85614 22788 85756
rect 22576 85550 22582 85614
rect 22646 85550 22788 85614
rect 22576 85544 22788 85550
rect 22984 85750 23196 85756
rect 22984 85686 23126 85750
rect 23190 85686 23196 85750
rect 22984 85614 23196 85686
rect 22984 85550 23126 85614
rect 23190 85550 23196 85614
rect 22984 85544 23196 85550
rect 23392 85750 23604 85756
rect 23392 85686 23398 85750
rect 23462 85686 23604 85750
rect 23392 85614 23604 85686
rect 23392 85550 23398 85614
rect 23462 85550 23604 85614
rect 23392 85544 23604 85550
rect 28288 85544 28636 85756
rect 190128 85544 190340 85756
rect 195024 85750 195236 85756
rect 195024 85686 195030 85750
rect 195094 85686 195236 85750
rect 195024 85614 195236 85686
rect 195024 85550 195030 85614
rect 195094 85550 195236 85614
rect 195024 85544 195236 85550
rect 195432 85750 195644 85756
rect 195432 85686 195574 85750
rect 195638 85686 195644 85750
rect 195432 85614 195644 85686
rect 195432 85550 195438 85614
rect 195502 85550 195644 85614
rect 195432 85544 195644 85550
rect 195840 85750 196052 85756
rect 195840 85686 195846 85750
rect 195910 85686 196052 85750
rect 195840 85614 196052 85686
rect 195840 85550 195982 85614
rect 196046 85550 196052 85614
rect 195840 85544 196052 85550
rect 196248 85544 196460 85756
rect 196656 85614 196868 85892
rect 196656 85550 196798 85614
rect 196862 85550 196868 85614
rect 196656 85544 196868 85550
rect 28288 85484 28364 85544
rect 190128 85484 190204 85544
rect 196248 85484 196324 85544
rect 21760 85342 21972 85348
rect 21760 85278 21902 85342
rect 21966 85278 21972 85342
rect 21760 85136 21972 85278
rect 22168 85342 22380 85348
rect 22168 85278 22174 85342
rect 22238 85278 22380 85342
rect 22168 85212 22380 85278
rect 22576 85342 22788 85348
rect 22576 85278 22582 85342
rect 22646 85278 22788 85342
rect 22576 85212 22788 85278
rect 22168 85206 22788 85212
rect 22168 85142 22310 85206
rect 22374 85142 22788 85206
rect 22168 85136 22788 85142
rect 22984 85342 23196 85348
rect 22984 85278 23126 85342
rect 23190 85278 23196 85342
rect 22984 85206 23196 85278
rect 22984 85142 23126 85206
rect 23190 85142 23196 85206
rect 22984 85136 23196 85142
rect 23392 85342 23604 85348
rect 23392 85278 23398 85342
rect 23462 85278 23604 85342
rect 23392 85206 23604 85278
rect 28288 85272 28636 85484
rect 190128 85272 190340 85484
rect 195976 85408 196324 85484
rect 195976 85348 196052 85408
rect 28424 85212 28500 85272
rect 190264 85212 190340 85272
rect 23392 85142 23398 85206
rect 23462 85142 23604 85206
rect 23392 85136 23604 85142
rect 21896 85076 21972 85136
rect 21760 84934 21972 85076
rect 28288 85070 28636 85212
rect 28288 85006 28294 85070
rect 28358 85006 28636 85070
rect 28288 85000 28636 85006
rect 190128 85000 190340 85212
rect 195024 85342 195236 85348
rect 195024 85278 195030 85342
rect 195094 85278 195236 85342
rect 195024 85206 195236 85278
rect 195024 85142 195030 85206
rect 195094 85142 195236 85206
rect 195024 85136 195236 85142
rect 195432 85342 195644 85348
rect 195432 85278 195438 85342
rect 195502 85278 195644 85342
rect 195432 85206 195644 85278
rect 195432 85142 195574 85206
rect 195638 85142 195644 85206
rect 195432 85136 195644 85142
rect 195840 85342 196460 85348
rect 195840 85278 195982 85342
rect 196046 85278 196460 85342
rect 195840 85272 196460 85278
rect 195840 85136 196052 85272
rect 196248 85206 196460 85272
rect 196248 85142 196390 85206
rect 196454 85142 196460 85206
rect 196248 85136 196460 85142
rect 196656 85342 196868 85348
rect 196656 85278 196798 85342
rect 196862 85278 196868 85342
rect 196656 85136 196868 85278
rect 196792 85076 196868 85136
rect 28560 84940 28636 85000
rect 190264 84940 190340 85000
rect 21760 84870 21902 84934
rect 21966 84870 21972 84934
rect 21760 84864 21972 84870
rect 22168 84934 22788 84940
rect 22168 84870 22310 84934
rect 22374 84870 22788 84934
rect 22168 84864 22788 84870
rect 22168 84728 22380 84864
rect 22576 84728 22788 84864
rect 22984 84934 23196 84940
rect 22984 84870 23126 84934
rect 23190 84870 23196 84934
rect 22984 84798 23196 84870
rect 22984 84734 23126 84798
rect 23190 84734 23196 84798
rect 22984 84728 23196 84734
rect 23392 84934 23604 84940
rect 23392 84870 23398 84934
rect 23462 84870 23604 84934
rect 23392 84798 23604 84870
rect 23392 84734 23534 84798
rect 23598 84734 23604 84798
rect 23392 84728 23604 84734
rect 28288 84798 28636 84940
rect 28288 84734 28294 84798
rect 28358 84734 28636 84798
rect 22304 84668 22380 84728
rect 1632 84532 1844 84668
rect 1224 84526 1702 84532
rect 1224 84462 1230 84526
rect 1294 84476 1702 84526
rect 1758 84476 1844 84532
rect 1294 84462 1844 84476
rect 1224 84456 1844 84462
rect 1632 84320 1844 84456
rect 21760 84662 21972 84668
rect 21760 84598 21902 84662
rect 21966 84598 21972 84662
rect 21760 84320 21972 84598
rect 22168 84390 22380 84668
rect 22576 84592 22788 84668
rect 22688 84396 22788 84592
rect 22478 84390 22788 84396
rect 22168 84326 22310 84390
rect 22374 84326 22380 84390
rect 22440 84326 22446 84390
rect 22510 84326 22788 84390
rect 22168 84320 22380 84326
rect 22478 84320 22788 84326
rect 22984 84526 23196 84532
rect 22984 84462 23126 84526
rect 23190 84462 23196 84526
rect 22984 84320 23196 84462
rect 21896 84260 21972 84320
rect 23120 84260 23196 84320
rect 21760 84118 21972 84260
rect 21760 84054 21902 84118
rect 21966 84054 21972 84118
rect 21760 84048 21972 84054
rect 22168 84118 22516 84124
rect 22168 84054 22310 84118
rect 22374 84054 22446 84118
rect 22510 84054 22516 84118
rect 22168 84048 22516 84054
rect 22168 83988 22380 84048
rect 22168 83912 22516 83988
rect 22576 83912 22788 84124
rect 22984 83912 23196 84260
rect 22440 83852 22516 83912
rect 22712 83852 22788 83912
rect 23120 83852 23196 83912
rect 21760 83846 21972 83852
rect 21760 83782 21902 83846
rect 21966 83782 21972 83846
rect 21760 83710 21972 83782
rect 21760 83646 21766 83710
rect 21830 83646 21972 83710
rect 21760 83640 21972 83646
rect 22168 83716 22380 83852
rect 22440 83776 22788 83852
rect 22576 83716 22788 83776
rect 22168 83710 22788 83716
rect 22168 83646 22310 83710
rect 22374 83646 22582 83710
rect 22646 83646 22788 83710
rect 22168 83640 22788 83646
rect 22984 83710 23196 83852
rect 22984 83646 23126 83710
rect 23190 83646 23196 83710
rect 22984 83640 23196 83646
rect 23392 84526 23604 84532
rect 23392 84462 23534 84526
rect 23598 84462 23604 84526
rect 23392 84320 23604 84462
rect 28288 84526 28636 84734
rect 28288 84462 28430 84526
rect 28494 84462 28636 84526
rect 28288 84456 28636 84462
rect 190128 84456 190340 84940
rect 195024 84934 195236 84940
rect 195024 84870 195030 84934
rect 195094 84870 195236 84934
rect 195024 84798 195236 84870
rect 195024 84734 195166 84798
rect 195230 84734 195236 84798
rect 195024 84728 195236 84734
rect 195432 84934 195644 84940
rect 195432 84870 195574 84934
rect 195638 84870 195644 84934
rect 195432 84798 195644 84870
rect 195432 84734 195438 84798
rect 195502 84734 195644 84798
rect 195432 84728 195644 84734
rect 195840 84728 196052 84940
rect 196248 84934 196460 84940
rect 196248 84870 196390 84934
rect 196454 84870 196460 84934
rect 196248 84728 196460 84870
rect 196656 84934 196868 85076
rect 196656 84870 196798 84934
rect 196862 84870 196868 84934
rect 196656 84864 196868 84870
rect 195976 84668 196052 84728
rect 196384 84668 196460 84728
rect 195024 84526 195236 84532
rect 195024 84462 195166 84526
rect 195230 84462 195236 84526
rect 28424 84396 28500 84456
rect 190128 84396 190204 84456
rect 23392 84260 23468 84320
rect 23392 83912 23604 84260
rect 28288 84254 28636 84396
rect 28288 84190 28430 84254
rect 28494 84190 28566 84254
rect 28630 84190 28636 84254
rect 28288 83982 28636 84190
rect 28288 83918 28566 83982
rect 28630 83918 28636 83982
rect 23392 83852 23468 83912
rect 23392 83710 23604 83852
rect 28288 83846 28636 83918
rect 28288 83782 28566 83846
rect 28630 83782 28636 83846
rect 28288 83776 28636 83782
rect 190128 84254 190340 84396
rect 190128 84190 190270 84254
rect 190334 84190 190340 84254
rect 190128 83982 190340 84190
rect 190128 83918 190270 83982
rect 190334 83918 190340 83982
rect 190128 83776 190340 83918
rect 190264 83716 190340 83776
rect 23392 83646 23534 83710
rect 23598 83646 23604 83710
rect 23392 83640 23604 83646
rect 21760 83438 21972 83444
rect 21760 83374 21766 83438
rect 21830 83374 21972 83438
rect 21760 83302 21972 83374
rect 21760 83238 21766 83302
rect 21830 83238 21972 83302
rect 21760 83232 21972 83238
rect 22168 83438 22380 83444
rect 22168 83374 22310 83438
rect 22374 83374 22380 83438
rect 22168 83232 22380 83374
rect 22576 83438 22788 83444
rect 22576 83374 22582 83438
rect 22646 83374 22788 83438
rect 22576 83232 22788 83374
rect 22984 83438 23196 83444
rect 22984 83374 23126 83438
rect 23190 83374 23196 83438
rect 22984 83302 23196 83374
rect 22984 83238 23126 83302
rect 23190 83238 23196 83302
rect 22984 83232 23196 83238
rect 23392 83438 23604 83444
rect 23392 83374 23534 83438
rect 23598 83374 23604 83438
rect 23392 83302 23604 83374
rect 23392 83238 23534 83302
rect 23598 83238 23604 83302
rect 23392 83232 23604 83238
rect 28288 83438 28636 83716
rect 28288 83374 28430 83438
rect 28494 83374 28566 83438
rect 28630 83374 28636 83438
rect 28288 83232 28636 83374
rect 22576 83172 22652 83232
rect 28560 83172 28636 83232
rect 22304 83096 22652 83172
rect 28288 83166 28636 83172
rect 28288 83102 28430 83166
rect 28494 83102 28636 83166
rect 22304 83036 22380 83096
rect 21760 83030 21972 83036
rect 21760 82966 21766 83030
rect 21830 82966 21972 83030
rect 1632 82852 1844 82900
rect 1632 82796 1702 82852
rect 1758 82796 1844 82852
rect 21760 82894 21972 82966
rect 21760 82830 21766 82894
rect 21830 82830 21972 82894
rect 21760 82824 21972 82830
rect 22168 82960 22788 83036
rect 22168 82824 22380 82960
rect 22576 82894 22788 82960
rect 22576 82830 22718 82894
rect 22782 82830 22788 82894
rect 22576 82824 22788 82830
rect 22984 83030 23196 83036
rect 22984 82966 23126 83030
rect 23190 82966 23196 83030
rect 22984 82894 23196 82966
rect 22984 82830 23126 82894
rect 23190 82830 23196 82894
rect 22984 82824 23196 82830
rect 23392 83030 23604 83036
rect 23392 82966 23534 83030
rect 23598 82966 23604 83030
rect 23392 82894 23604 82966
rect 28288 82960 28636 83102
rect 190128 83232 190340 83716
rect 195024 84320 195236 84462
rect 195432 84526 195644 84532
rect 195432 84462 195438 84526
rect 195502 84462 195644 84526
rect 195432 84320 195644 84462
rect 195840 84390 196052 84668
rect 196248 84396 196460 84668
rect 196150 84390 196460 84396
rect 195840 84326 195846 84390
rect 195910 84326 196052 84390
rect 196112 84326 196118 84390
rect 196182 84326 196460 84390
rect 195840 84320 196052 84326
rect 196150 84320 196460 84326
rect 196656 84662 196868 84668
rect 196656 84598 196798 84662
rect 196862 84598 196868 84662
rect 196656 84320 196868 84598
rect 216784 84532 216996 84668
rect 216784 84476 216908 84532
rect 216964 84476 216996 84532
rect 216784 84396 216996 84476
rect 216784 84390 217540 84396
rect 216784 84326 217470 84390
rect 217534 84326 217540 84390
rect 216784 84320 217540 84326
rect 195024 84260 195100 84320
rect 195432 84260 195508 84320
rect 196792 84260 196868 84320
rect 195024 83912 195236 84260
rect 195432 83912 195644 84260
rect 195840 84118 196188 84124
rect 195840 84054 195846 84118
rect 195910 84054 196118 84118
rect 196182 84054 196188 84118
rect 195840 84048 196188 84054
rect 195840 83988 196052 84048
rect 196248 83988 196460 84124
rect 196656 84118 196868 84260
rect 196656 84054 196798 84118
rect 196862 84054 196868 84118
rect 196656 84048 196868 84054
rect 195840 83912 196460 83988
rect 195024 83852 195100 83912
rect 195568 83852 195644 83912
rect 195976 83852 196052 83912
rect 196384 83852 196460 83912
rect 195024 83710 195236 83852
rect 195024 83646 195166 83710
rect 195230 83646 195236 83710
rect 195024 83640 195236 83646
rect 195432 83710 195644 83852
rect 195432 83646 195438 83710
rect 195502 83646 195644 83710
rect 195432 83640 195644 83646
rect 195840 83710 196052 83852
rect 195840 83646 195846 83710
rect 195910 83646 196052 83710
rect 195840 83640 196052 83646
rect 196248 83640 196460 83852
rect 196656 83846 196868 83852
rect 196656 83782 196798 83846
rect 196862 83782 196868 83846
rect 196656 83710 196868 83782
rect 196656 83646 196662 83710
rect 196726 83646 196868 83710
rect 196656 83640 196868 83646
rect 195024 83438 195236 83444
rect 195024 83374 195166 83438
rect 195230 83374 195236 83438
rect 195024 83302 195236 83374
rect 195024 83238 195166 83302
rect 195230 83238 195236 83302
rect 195024 83232 195236 83238
rect 195432 83438 195644 83444
rect 195432 83374 195438 83438
rect 195502 83374 195644 83438
rect 195432 83302 195644 83374
rect 195432 83238 195574 83302
rect 195638 83238 195644 83302
rect 195432 83232 195644 83238
rect 195840 83438 196052 83444
rect 195840 83374 195846 83438
rect 195910 83374 196052 83438
rect 195840 83302 196052 83374
rect 195840 83238 195982 83302
rect 196046 83238 196052 83302
rect 195840 83232 196052 83238
rect 196248 83302 196460 83444
rect 196248 83238 196390 83302
rect 196454 83238 196460 83302
rect 196248 83232 196460 83238
rect 196656 83438 196868 83444
rect 196656 83374 196662 83438
rect 196726 83374 196868 83438
rect 196656 83302 196868 83374
rect 196656 83238 196662 83302
rect 196726 83238 196868 83302
rect 196656 83232 196868 83238
rect 190128 83172 190204 83232
rect 190128 82960 190340 83172
rect 28560 82900 28636 82960
rect 190264 82900 190340 82960
rect 23392 82830 23534 82894
rect 23598 82830 23604 82894
rect 23392 82824 23604 82830
rect 1632 82764 1844 82796
rect 1224 82758 1844 82764
rect 1224 82694 1230 82758
rect 1294 82694 1844 82758
rect 1224 82688 1844 82694
rect 28288 82688 28636 82900
rect 190128 82688 190340 82900
rect 195024 83030 195236 83036
rect 195024 82966 195166 83030
rect 195230 82966 195236 83030
rect 195024 82894 195236 82966
rect 195024 82830 195166 82894
rect 195230 82830 195236 82894
rect 195024 82824 195236 82830
rect 195432 83030 195644 83036
rect 195432 82966 195574 83030
rect 195638 82966 195644 83030
rect 195432 82894 195644 82966
rect 195432 82830 195438 82894
rect 195502 82830 195644 82894
rect 195432 82824 195644 82830
rect 195840 83030 196460 83036
rect 195840 82966 195982 83030
rect 196046 82966 196390 83030
rect 196454 82966 196460 83030
rect 195840 82960 196460 82966
rect 195840 82824 196052 82960
rect 196248 82894 196460 82960
rect 196248 82830 196254 82894
rect 196318 82830 196460 82894
rect 196248 82824 196460 82830
rect 196656 83030 196868 83036
rect 196656 82966 196662 83030
rect 196726 82966 196868 83030
rect 196656 82894 196868 82966
rect 196656 82830 196798 82894
rect 196862 82830 196868 82894
rect 196656 82824 196868 82830
rect 216784 82894 217540 82900
rect 216784 82852 217470 82894
rect 216784 82796 216908 82852
rect 216964 82830 217470 82852
rect 217534 82830 217540 82894
rect 216964 82824 217540 82830
rect 216964 82796 216996 82824
rect 216784 82688 216996 82796
rect 28424 82628 28500 82688
rect 190128 82628 190204 82688
rect 21760 82622 21972 82628
rect 21760 82558 21766 82622
rect 21830 82558 21972 82622
rect 21760 82486 21972 82558
rect 21760 82422 21766 82486
rect 21830 82422 21972 82486
rect 21760 82416 21972 82422
rect 22168 82492 22380 82628
rect 22576 82622 22788 82628
rect 22576 82558 22718 82622
rect 22782 82558 22788 82622
rect 22576 82492 22788 82558
rect 22168 82486 22788 82492
rect 22168 82422 22174 82486
rect 22238 82422 22582 82486
rect 22646 82422 22788 82486
rect 22168 82416 22788 82422
rect 22984 82622 23196 82628
rect 22984 82558 23126 82622
rect 23190 82558 23196 82622
rect 22984 82486 23196 82558
rect 22984 82422 23126 82486
rect 23190 82422 23196 82486
rect 22984 82416 23196 82422
rect 23392 82622 23604 82628
rect 23392 82558 23534 82622
rect 23598 82558 23604 82622
rect 23392 82486 23604 82558
rect 23392 82422 23534 82486
rect 23598 82422 23604 82486
rect 23392 82416 23604 82422
rect 28288 82416 28636 82628
rect 190128 82416 190340 82628
rect 195024 82622 195236 82628
rect 195024 82558 195166 82622
rect 195230 82558 195236 82622
rect 195024 82486 195236 82558
rect 195024 82422 195166 82486
rect 195230 82422 195236 82486
rect 195024 82416 195236 82422
rect 195432 82622 195644 82628
rect 195432 82558 195438 82622
rect 195502 82558 195644 82622
rect 195432 82486 195644 82558
rect 195432 82422 195438 82486
rect 195502 82422 195644 82486
rect 195432 82416 195644 82422
rect 195840 82486 196052 82628
rect 195840 82422 195846 82486
rect 195910 82422 196052 82486
rect 195840 82416 196052 82422
rect 196248 82622 196460 82628
rect 196248 82558 196254 82622
rect 196318 82558 196460 82622
rect 196248 82486 196460 82558
rect 196248 82422 196254 82486
rect 196318 82422 196460 82486
rect 196248 82416 196460 82422
rect 196656 82622 196868 82628
rect 196656 82558 196798 82622
rect 196862 82558 196868 82622
rect 196656 82486 196868 82558
rect 196656 82422 196662 82486
rect 196726 82422 196868 82486
rect 196656 82416 196868 82422
rect 28288 82356 28364 82416
rect 190128 82356 190204 82416
rect 21760 82214 21972 82220
rect 21760 82150 21766 82214
rect 21830 82150 21972 82214
rect 21760 82078 21972 82150
rect 21760 82014 21902 82078
rect 21966 82014 21972 82078
rect 21760 82008 21972 82014
rect 22168 82214 22380 82220
rect 22168 82150 22174 82214
rect 22238 82150 22380 82214
rect 22168 82008 22380 82150
rect 22576 82214 22788 82220
rect 22576 82150 22582 82214
rect 22646 82150 22788 82214
rect 22576 82078 22788 82150
rect 22576 82014 22718 82078
rect 22782 82014 22788 82078
rect 22576 82008 22788 82014
rect 22984 82214 23196 82220
rect 22984 82150 23126 82214
rect 23190 82150 23196 82214
rect 22984 82078 23196 82150
rect 22984 82014 23126 82078
rect 23190 82014 23196 82078
rect 22984 82008 23196 82014
rect 23392 82214 23604 82220
rect 23392 82150 23534 82214
rect 23598 82150 23604 82214
rect 23392 82078 23604 82150
rect 23392 82014 23398 82078
rect 23462 82014 23604 82078
rect 23392 82008 23604 82014
rect 28288 82144 28636 82356
rect 190128 82144 190340 82356
rect 195024 82214 195236 82220
rect 195024 82150 195166 82214
rect 195230 82150 195236 82214
rect 28288 82084 28364 82144
rect 190128 82084 190204 82144
rect 28288 81872 28636 82084
rect 190128 81872 190340 82084
rect 195024 82078 195236 82150
rect 195024 82014 195030 82078
rect 195094 82014 195236 82078
rect 195024 82008 195236 82014
rect 195432 82214 195644 82220
rect 195432 82150 195438 82214
rect 195502 82150 195644 82214
rect 195432 82078 195644 82150
rect 195432 82014 195438 82078
rect 195502 82014 195644 82078
rect 195432 82008 195644 82014
rect 195840 82214 196052 82220
rect 195840 82150 195846 82214
rect 195910 82150 196052 82214
rect 195840 82084 196052 82150
rect 196248 82214 196460 82220
rect 196248 82150 196254 82214
rect 196318 82150 196460 82214
rect 196248 82084 196460 82150
rect 195840 82078 196460 82084
rect 195840 82014 195982 82078
rect 196046 82014 196460 82078
rect 195840 82008 196460 82014
rect 196656 82214 196868 82220
rect 196656 82150 196662 82214
rect 196726 82150 196868 82214
rect 196656 82078 196868 82150
rect 196656 82014 196798 82078
rect 196862 82014 196868 82078
rect 196656 82008 196868 82014
rect 195976 81948 196052 82008
rect 195976 81872 196324 81948
rect 28424 81812 28500 81872
rect 190264 81812 190340 81872
rect 196248 81812 196324 81872
rect 21760 81806 21972 81812
rect 21760 81742 21902 81806
rect 21966 81742 21972 81806
rect 21760 81670 21972 81742
rect 21760 81606 21766 81670
rect 21830 81606 21972 81670
rect 21760 81600 21972 81606
rect 22168 81806 22788 81812
rect 22168 81742 22718 81806
rect 22782 81742 22788 81806
rect 22168 81736 22788 81742
rect 22168 81676 22380 81736
rect 22168 81670 22516 81676
rect 22168 81606 22310 81670
rect 22374 81606 22446 81670
rect 22510 81606 22516 81670
rect 22168 81600 22516 81606
rect 22576 81600 22788 81736
rect 22984 81806 23196 81812
rect 22984 81742 23126 81806
rect 23190 81742 23196 81806
rect 22984 81670 23196 81742
rect 22984 81606 23126 81670
rect 23190 81606 23196 81670
rect 22984 81600 23196 81606
rect 23392 81806 23604 81812
rect 23392 81742 23398 81806
rect 23462 81742 23604 81806
rect 23392 81670 23604 81742
rect 23392 81606 23534 81670
rect 23598 81606 23604 81670
rect 23392 81600 23604 81606
rect 28288 81600 28636 81812
rect 190128 81600 190340 81812
rect 195024 81806 195236 81812
rect 195024 81742 195030 81806
rect 195094 81742 195236 81806
rect 195024 81670 195236 81742
rect 195024 81606 195166 81670
rect 195230 81606 195236 81670
rect 195024 81600 195236 81606
rect 195432 81806 195644 81812
rect 195432 81742 195438 81806
rect 195502 81742 195644 81806
rect 195432 81670 195644 81742
rect 195432 81606 195438 81670
rect 195502 81606 195644 81670
rect 195432 81600 195644 81606
rect 195840 81806 196052 81812
rect 195840 81742 195982 81806
rect 196046 81742 196052 81806
rect 195840 81676 196052 81742
rect 195840 81670 196188 81676
rect 195840 81606 196118 81670
rect 196182 81606 196188 81670
rect 195840 81600 196188 81606
rect 196248 81600 196460 81812
rect 196656 81806 196868 81812
rect 196656 81742 196798 81806
rect 196862 81742 196868 81806
rect 196656 81670 196868 81742
rect 196656 81606 196662 81670
rect 196726 81606 196868 81670
rect 196656 81600 196868 81606
rect 28288 81540 28364 81600
rect 190128 81540 190204 81600
rect 21760 81398 21972 81404
rect 21760 81334 21766 81398
rect 21830 81334 21972 81398
rect 1632 81172 1844 81268
rect 1632 81132 1702 81172
rect 1224 81126 1702 81132
rect 1224 81062 1230 81126
rect 1294 81116 1702 81126
rect 1758 81116 1844 81172
rect 1294 81062 1844 81116
rect 1224 81056 1844 81062
rect 21760 81192 21972 81334
rect 22168 81398 22380 81404
rect 22478 81398 22788 81404
rect 22168 81334 22310 81398
rect 22374 81334 22380 81398
rect 22440 81334 22446 81398
rect 22510 81334 22788 81398
rect 22168 81192 22380 81334
rect 22478 81328 22788 81334
rect 22576 81262 22788 81328
rect 22576 81198 22582 81262
rect 22646 81198 22788 81262
rect 22576 81192 22788 81198
rect 22984 81398 23196 81404
rect 22984 81334 23126 81398
rect 23190 81334 23196 81398
rect 22984 81262 23196 81334
rect 22984 81198 22990 81262
rect 23054 81198 23196 81262
rect 22984 81192 23196 81198
rect 23392 81398 23604 81404
rect 23392 81334 23534 81398
rect 23598 81334 23604 81398
rect 23392 81262 23604 81334
rect 23392 81198 23534 81262
rect 23598 81198 23604 81262
rect 23392 81192 23604 81198
rect 28288 81328 28636 81540
rect 190128 81328 190340 81540
rect 195024 81398 195236 81404
rect 195024 81334 195166 81398
rect 195230 81334 195236 81398
rect 28288 81268 28364 81328
rect 190128 81268 190204 81328
rect 21760 81132 21836 81192
rect 21760 80990 21972 81132
rect 28288 81126 28636 81268
rect 28288 81062 28566 81126
rect 28630 81062 28636 81126
rect 28288 81056 28636 81062
rect 190128 81056 190340 81268
rect 195024 81262 195236 81334
rect 195024 81198 195166 81262
rect 195230 81198 195236 81262
rect 195024 81192 195236 81198
rect 195432 81398 195644 81404
rect 195432 81334 195438 81398
rect 195502 81334 195644 81398
rect 195432 81262 195644 81334
rect 195432 81198 195438 81262
rect 195502 81198 195644 81262
rect 195432 81192 195644 81198
rect 195840 81262 196052 81404
rect 196150 81398 196460 81404
rect 196112 81334 196118 81398
rect 196182 81334 196460 81398
rect 196150 81328 196460 81334
rect 196248 81268 196460 81328
rect 196150 81262 196460 81268
rect 195840 81198 195982 81262
rect 196046 81198 196052 81262
rect 196112 81198 196118 81262
rect 196182 81198 196460 81262
rect 195840 81192 196052 81198
rect 196150 81192 196460 81198
rect 196656 81398 196868 81404
rect 196656 81334 196662 81398
rect 196726 81334 196868 81398
rect 196656 81192 196868 81334
rect 216784 81262 217540 81268
rect 216784 81198 217470 81262
rect 217534 81198 217540 81262
rect 216784 81192 217540 81198
rect 28424 80996 28500 81056
rect 190264 80996 190340 81056
rect 196656 81132 196732 81192
rect 216784 81172 216996 81192
rect 21760 80926 21902 80990
rect 21966 80926 21972 80990
rect 21760 80920 21972 80926
rect 22168 80990 22516 80996
rect 22168 80926 22446 80990
rect 22510 80926 22516 80990
rect 22168 80920 22516 80926
rect 22576 80990 22788 80996
rect 22576 80926 22582 80990
rect 22646 80926 22788 80990
rect 22168 80860 22380 80920
rect 22576 80860 22788 80926
rect 22168 80784 22788 80860
rect 22984 80990 23196 80996
rect 22984 80926 22990 80990
rect 23054 80926 23196 80990
rect 22984 80854 23196 80926
rect 22984 80790 22990 80854
rect 23054 80790 23196 80854
rect 22984 80784 23196 80790
rect 23392 80990 23604 80996
rect 23392 80926 23534 80990
rect 23598 80926 23604 80990
rect 23392 80854 23604 80926
rect 23392 80790 23398 80854
rect 23462 80790 23604 80854
rect 23392 80784 23604 80790
rect 28288 80854 28636 80996
rect 28288 80790 28430 80854
rect 28494 80790 28566 80854
rect 28630 80790 28636 80854
rect 22168 80724 22244 80784
rect 21760 80718 21972 80724
rect 21760 80654 21902 80718
rect 21966 80654 21972 80718
rect 21760 80376 21972 80654
rect 22168 80376 22380 80724
rect 22478 80718 22788 80724
rect 22440 80654 22446 80718
rect 22510 80654 22788 80718
rect 22478 80648 22788 80654
rect 22576 80452 22788 80648
rect 22478 80446 22788 80452
rect 22440 80382 22446 80446
rect 22510 80382 22788 80446
rect 22478 80376 22788 80382
rect 22984 80582 23196 80588
rect 22984 80518 22990 80582
rect 23054 80518 23196 80582
rect 22984 80376 23196 80518
rect 23392 80582 23604 80588
rect 23392 80518 23398 80582
rect 23462 80518 23604 80582
rect 23392 80376 23604 80518
rect 28288 80512 28636 80790
rect 190128 80512 190340 80996
rect 195024 80990 195236 80996
rect 195024 80926 195166 80990
rect 195230 80926 195236 80990
rect 195024 80854 195236 80926
rect 195024 80790 195030 80854
rect 195094 80790 195236 80854
rect 195024 80784 195236 80790
rect 195432 80990 195644 80996
rect 195432 80926 195438 80990
rect 195502 80926 195644 80990
rect 195432 80854 195644 80926
rect 195432 80790 195574 80854
rect 195638 80790 195644 80854
rect 195432 80784 195644 80790
rect 195840 80990 196188 80996
rect 195840 80926 195982 80990
rect 196046 80926 196118 80990
rect 196182 80926 196188 80990
rect 195840 80920 196188 80926
rect 195840 80860 196052 80920
rect 196248 80860 196460 80996
rect 196656 80990 196868 81132
rect 216784 81116 216908 81172
rect 216964 81116 216996 81172
rect 216784 81056 216996 81116
rect 196656 80926 196662 80990
rect 196726 80926 196868 80990
rect 196656 80920 196868 80926
rect 195840 80784 196460 80860
rect 195976 80724 196052 80784
rect 196384 80724 196460 80784
rect 190264 80452 190340 80512
rect 21760 80316 21836 80376
rect 22984 80316 23060 80376
rect 23528 80316 23604 80376
rect 21760 80174 21972 80316
rect 21760 80110 21766 80174
rect 21830 80110 21972 80174
rect 21760 80104 21972 80110
rect 22168 80174 22516 80180
rect 22168 80110 22446 80174
rect 22510 80110 22516 80174
rect 22168 80104 22516 80110
rect 22168 79968 22380 80104
rect 22576 80044 22788 80180
rect 22304 79908 22380 79968
rect 22440 79968 22788 80044
rect 22984 79968 23196 80316
rect 23392 79968 23604 80316
rect 22440 79908 22516 79968
rect 22712 79908 22788 79968
rect 23120 79908 23196 79968
rect 23528 79908 23604 79968
rect 21760 79902 21972 79908
rect 21760 79838 21766 79902
rect 21830 79838 21972 79902
rect 21760 79766 21972 79838
rect 21760 79702 21902 79766
rect 21966 79702 21972 79766
rect 21760 79696 21972 79702
rect 22168 79832 22516 79908
rect 22168 79772 22380 79832
rect 22168 79766 22516 79772
rect 22168 79702 22310 79766
rect 22374 79702 22446 79766
rect 22510 79702 22516 79766
rect 22168 79696 22516 79702
rect 22576 79696 22788 79908
rect 1224 79630 1844 79636
rect 1224 79566 1230 79630
rect 1294 79566 1844 79630
rect 1224 79560 1844 79566
rect 1632 79492 1844 79560
rect 22984 79560 23196 79908
rect 23392 79560 23604 79908
rect 28288 80446 28636 80452
rect 28288 80382 28430 80446
rect 28494 80382 28636 80446
rect 28288 80310 28636 80382
rect 28288 80246 28294 80310
rect 28358 80246 28636 80310
rect 28288 80038 28636 80246
rect 28288 79974 28294 80038
rect 28358 79974 28430 80038
rect 28494 79974 28636 80038
rect 28288 79832 28636 79974
rect 190128 80310 190340 80452
rect 195024 80582 195236 80588
rect 195024 80518 195030 80582
rect 195094 80518 195236 80582
rect 195024 80376 195236 80518
rect 195432 80582 195644 80588
rect 195432 80518 195574 80582
rect 195638 80518 195644 80582
rect 195432 80376 195644 80518
rect 195840 80446 196052 80724
rect 195840 80382 195982 80446
rect 196046 80382 196052 80446
rect 195840 80376 196052 80382
rect 196248 80376 196460 80724
rect 196656 80718 196868 80724
rect 196656 80654 196662 80718
rect 196726 80654 196868 80718
rect 196656 80376 196868 80654
rect 195160 80316 195236 80376
rect 195568 80316 195644 80376
rect 190128 80246 190134 80310
rect 190198 80246 190340 80310
rect 190128 80038 190340 80246
rect 190128 79974 190134 80038
rect 190198 79974 190340 80038
rect 190128 79902 190340 79974
rect 195024 79968 195236 80316
rect 195432 79968 195644 80316
rect 196656 80316 196732 80376
rect 195840 80174 196052 80180
rect 195840 80110 195982 80174
rect 196046 80110 196052 80174
rect 195840 79968 196052 80110
rect 196248 80044 196460 80180
rect 196656 80174 196868 80316
rect 196656 80110 196798 80174
rect 196862 80110 196868 80174
rect 196656 80104 196868 80110
rect 195160 79908 195236 79968
rect 195568 79908 195644 79968
rect 195976 79908 196052 79968
rect 196112 79968 196460 80044
rect 196112 79908 196188 79968
rect 196384 79908 196460 79968
rect 190128 79838 190270 79902
rect 190334 79838 190340 79902
rect 190128 79832 190340 79838
rect 28288 79630 28636 79636
rect 28288 79566 28430 79630
rect 28494 79566 28636 79630
rect 22984 79500 23060 79560
rect 23392 79500 23468 79560
rect 1632 79436 1702 79492
rect 1758 79436 1844 79492
rect 1632 79288 1844 79436
rect 21760 79494 21972 79500
rect 21760 79430 21902 79494
rect 21966 79430 21972 79494
rect 21760 79358 21972 79430
rect 21760 79294 21766 79358
rect 21830 79294 21972 79358
rect 21760 79288 21972 79294
rect 22168 79494 22380 79500
rect 22478 79494 22788 79500
rect 22168 79430 22310 79494
rect 22374 79430 22380 79494
rect 22440 79430 22446 79494
rect 22510 79430 22788 79494
rect 22168 79152 22380 79430
rect 22478 79424 22788 79430
rect 22576 79152 22788 79424
rect 22984 79358 23196 79500
rect 22984 79294 23126 79358
rect 23190 79294 23196 79358
rect 22984 79288 23196 79294
rect 23392 79358 23604 79500
rect 23392 79294 23534 79358
rect 23598 79294 23604 79358
rect 23392 79288 23604 79294
rect 28288 79494 28636 79566
rect 28288 79430 28566 79494
rect 28630 79430 28636 79494
rect 28288 79288 28636 79430
rect 28560 79228 28636 79288
rect 28288 79222 28636 79228
rect 28288 79158 28566 79222
rect 28630 79158 28636 79222
rect 22168 79092 22244 79152
rect 22576 79092 22652 79152
rect 21760 79086 21972 79092
rect 21760 79022 21766 79086
rect 21830 79022 21972 79086
rect 21760 78950 21972 79022
rect 21760 78886 21902 78950
rect 21966 78886 21972 78950
rect 21760 78880 21972 78886
rect 22168 78880 22380 79092
rect 22576 78950 22788 79092
rect 22576 78886 22582 78950
rect 22646 78886 22788 78950
rect 22576 78880 22788 78886
rect 22984 79086 23196 79092
rect 22984 79022 23126 79086
rect 23190 79022 23196 79086
rect 22984 78950 23196 79022
rect 22984 78886 22990 78950
rect 23054 78886 23196 78950
rect 22984 78880 23196 78886
rect 23392 79086 23604 79092
rect 23392 79022 23534 79086
rect 23598 79022 23604 79086
rect 23392 78950 23604 79022
rect 23392 78886 23398 78950
rect 23462 78886 23604 78950
rect 23392 78880 23604 78886
rect 28288 79016 28636 79158
rect 190128 79630 190340 79636
rect 190128 79566 190270 79630
rect 190334 79566 190340 79630
rect 190128 79494 190340 79566
rect 190128 79430 190270 79494
rect 190334 79430 190340 79494
rect 190128 79288 190340 79430
rect 195024 79560 195236 79908
rect 195432 79560 195644 79908
rect 195840 79832 196188 79908
rect 195840 79696 196052 79832
rect 196248 79766 196460 79908
rect 196248 79702 196390 79766
rect 196454 79702 196460 79766
rect 196248 79696 196460 79702
rect 196656 79902 196868 79908
rect 196656 79838 196798 79902
rect 196862 79838 196868 79902
rect 196656 79766 196868 79838
rect 196656 79702 196798 79766
rect 196862 79702 196868 79766
rect 196656 79696 196868 79702
rect 195024 79500 195100 79560
rect 195568 79500 195644 79560
rect 195024 79358 195236 79500
rect 195024 79294 195166 79358
rect 195230 79294 195236 79358
rect 195024 79288 195236 79294
rect 195432 79358 195644 79500
rect 195432 79294 195574 79358
rect 195638 79294 195644 79358
rect 195432 79288 195644 79294
rect 190128 79228 190204 79288
rect 190128 79222 190340 79228
rect 190128 79158 190270 79222
rect 190334 79158 190340 79222
rect 190128 79016 190340 79158
rect 195840 79152 196052 79500
rect 196248 79494 196460 79500
rect 196248 79430 196390 79494
rect 196454 79430 196460 79494
rect 196248 79152 196460 79430
rect 196656 79494 196868 79500
rect 196656 79430 196798 79494
rect 196862 79430 196868 79494
rect 196656 79358 196868 79430
rect 196656 79294 196662 79358
rect 196726 79294 196868 79358
rect 196656 79288 196868 79294
rect 216784 79492 216996 79636
rect 216784 79436 216908 79492
rect 216964 79436 216996 79492
rect 216784 79364 216996 79436
rect 216784 79358 217540 79364
rect 216784 79294 217470 79358
rect 217534 79294 217540 79358
rect 216784 79288 217540 79294
rect 195840 79092 195916 79152
rect 196248 79092 196324 79152
rect 195024 79086 195236 79092
rect 195024 79022 195166 79086
rect 195230 79022 195236 79086
rect 28288 78956 28364 79016
rect 190128 78956 190204 79016
rect 28288 78744 28636 78956
rect 190128 78744 190340 78956
rect 195024 78950 195236 79022
rect 195024 78886 195166 78950
rect 195230 78886 195236 78950
rect 195024 78880 195236 78886
rect 195432 79086 195644 79092
rect 195432 79022 195574 79086
rect 195638 79022 195644 79086
rect 195432 78950 195644 79022
rect 195432 78886 195438 78950
rect 195502 78886 195644 78950
rect 195432 78880 195644 78886
rect 195840 78950 196052 79092
rect 196248 78956 196460 79092
rect 196150 78950 196460 78956
rect 195840 78886 195846 78950
rect 195910 78886 196052 78950
rect 196112 78886 196118 78950
rect 196182 78886 196460 78950
rect 195840 78880 196052 78886
rect 196150 78880 196460 78886
rect 196656 79086 196868 79092
rect 196656 79022 196662 79086
rect 196726 79022 196868 79086
rect 196656 78950 196868 79022
rect 196656 78886 196798 78950
rect 196862 78886 196868 78950
rect 196656 78880 196868 78886
rect 28560 78684 28636 78744
rect 190264 78684 190340 78744
rect 21760 78678 21972 78684
rect 21760 78614 21902 78678
rect 21966 78614 21972 78678
rect 21760 78542 21972 78614
rect 21760 78478 21902 78542
rect 21966 78478 21972 78542
rect 21760 78472 21972 78478
rect 22168 78678 22788 78684
rect 22168 78614 22582 78678
rect 22646 78614 22788 78678
rect 22168 78608 22788 78614
rect 22168 78542 22380 78608
rect 22168 78478 22174 78542
rect 22238 78478 22380 78542
rect 22168 78472 22380 78478
rect 22576 78542 22788 78608
rect 22576 78478 22718 78542
rect 22782 78478 22788 78542
rect 22576 78472 22788 78478
rect 22984 78678 23196 78684
rect 22984 78614 22990 78678
rect 23054 78614 23196 78678
rect 22984 78542 23196 78614
rect 22984 78478 22990 78542
rect 23054 78478 23196 78542
rect 22984 78472 23196 78478
rect 23392 78678 23604 78684
rect 23392 78614 23398 78678
rect 23462 78614 23604 78678
rect 23392 78542 23604 78614
rect 23392 78478 23398 78542
rect 23462 78478 23604 78542
rect 23392 78472 23604 78478
rect 28288 78472 28636 78684
rect 190128 78472 190340 78684
rect 195024 78678 195236 78684
rect 195024 78614 195166 78678
rect 195230 78614 195236 78678
rect 195024 78542 195236 78614
rect 195024 78478 195166 78542
rect 195230 78478 195236 78542
rect 195024 78472 195236 78478
rect 195432 78678 195644 78684
rect 195432 78614 195438 78678
rect 195502 78614 195644 78678
rect 195432 78542 195644 78614
rect 195432 78478 195574 78542
rect 195638 78478 195644 78542
rect 195432 78472 195644 78478
rect 195840 78678 196188 78684
rect 195840 78614 195846 78678
rect 195910 78614 196118 78678
rect 196182 78614 196188 78678
rect 195840 78608 196188 78614
rect 195840 78548 196052 78608
rect 196248 78548 196460 78684
rect 195840 78542 196460 78548
rect 195840 78478 195846 78542
rect 195910 78478 196460 78542
rect 195840 78472 196460 78478
rect 196656 78678 196868 78684
rect 196656 78614 196798 78678
rect 196862 78614 196868 78678
rect 196656 78542 196868 78614
rect 196656 78478 196798 78542
rect 196862 78478 196868 78542
rect 196656 78472 196868 78478
rect 28424 78412 28500 78472
rect 190264 78412 190340 78472
rect 21760 78270 21972 78276
rect 21760 78206 21902 78270
rect 21966 78206 21972 78270
rect 21760 78134 21972 78206
rect 21760 78070 21766 78134
rect 21830 78070 21972 78134
rect 21760 78064 21972 78070
rect 22168 78270 22380 78276
rect 22168 78206 22174 78270
rect 22238 78206 22380 78270
rect 22168 78064 22380 78206
rect 22576 78270 22788 78276
rect 22576 78206 22718 78270
rect 22782 78206 22788 78270
rect 22576 78134 22788 78206
rect 22576 78070 22582 78134
rect 22646 78070 22788 78134
rect 22576 78064 22788 78070
rect 22984 78270 23196 78276
rect 22984 78206 22990 78270
rect 23054 78206 23196 78270
rect 22984 78134 23196 78206
rect 22984 78070 22990 78134
rect 23054 78070 23196 78134
rect 22984 78064 23196 78070
rect 23392 78270 23604 78276
rect 23392 78206 23398 78270
rect 23462 78206 23604 78270
rect 23392 78134 23604 78206
rect 28288 78200 28636 78412
rect 190128 78200 190340 78412
rect 195024 78270 195236 78276
rect 195024 78206 195166 78270
rect 195230 78206 195236 78270
rect 28424 78140 28500 78200
rect 190128 78140 190204 78200
rect 23392 78070 23534 78134
rect 23598 78070 23604 78134
rect 23392 78064 23604 78070
rect 28288 77928 28636 78140
rect 190128 77928 190340 78140
rect 195024 78134 195236 78206
rect 195024 78070 195166 78134
rect 195230 78070 195236 78134
rect 195024 78064 195236 78070
rect 195432 78270 195644 78276
rect 195432 78206 195574 78270
rect 195638 78206 195644 78270
rect 195432 78134 195644 78206
rect 195432 78070 195438 78134
rect 195502 78070 195644 78134
rect 195432 78064 195644 78070
rect 195840 78270 196460 78276
rect 195840 78206 195846 78270
rect 195910 78206 196460 78270
rect 195840 78200 196460 78206
rect 195840 78134 196052 78200
rect 195840 78070 195846 78134
rect 195910 78070 196052 78134
rect 195840 78064 196052 78070
rect 196248 78064 196460 78200
rect 196656 78270 196868 78276
rect 196656 78206 196798 78270
rect 196862 78206 196868 78270
rect 196656 78134 196868 78206
rect 196656 78070 196662 78134
rect 196726 78070 196868 78134
rect 196656 78064 196868 78070
rect 28288 77868 28364 77928
rect 190128 77868 190204 77928
rect 1632 77812 1844 77868
rect 1632 77756 1702 77812
rect 1758 77756 1844 77812
rect 1632 77732 1844 77756
rect 1224 77726 1844 77732
rect 1224 77662 1230 77726
rect 1294 77662 1844 77726
rect 1224 77656 1844 77662
rect 21760 77862 21972 77868
rect 21760 77798 21766 77862
rect 21830 77798 21972 77862
rect 21760 77726 21972 77798
rect 21760 77662 21902 77726
rect 21966 77662 21972 77726
rect 21760 77656 21972 77662
rect 22168 77862 22788 77868
rect 22168 77798 22582 77862
rect 22646 77798 22788 77862
rect 22168 77792 22788 77798
rect 22168 77732 22380 77792
rect 22168 77726 22516 77732
rect 22168 77662 22446 77726
rect 22510 77662 22516 77726
rect 22168 77656 22516 77662
rect 22576 77656 22788 77792
rect 22984 77862 23196 77868
rect 22984 77798 22990 77862
rect 23054 77798 23196 77862
rect 22984 77726 23196 77798
rect 22984 77662 22990 77726
rect 23054 77662 23196 77726
rect 22984 77656 23196 77662
rect 23392 77862 23604 77868
rect 23392 77798 23534 77862
rect 23598 77798 23604 77862
rect 23392 77726 23604 77798
rect 23392 77662 23398 77726
rect 23462 77662 23604 77726
rect 23392 77656 23604 77662
rect 28288 77656 28636 77868
rect 190128 77656 190340 77868
rect 195024 77862 195236 77868
rect 195024 77798 195166 77862
rect 195230 77798 195236 77862
rect 195024 77726 195236 77798
rect 195024 77662 195030 77726
rect 195094 77662 195236 77726
rect 195024 77656 195236 77662
rect 195432 77862 195644 77868
rect 195432 77798 195438 77862
rect 195502 77798 195644 77862
rect 195432 77726 195644 77798
rect 195432 77662 195438 77726
rect 195502 77662 195644 77726
rect 195432 77656 195644 77662
rect 195840 77862 196052 77868
rect 195840 77798 195846 77862
rect 195910 77798 196052 77862
rect 195840 77726 196052 77798
rect 195840 77662 195982 77726
rect 196046 77662 196052 77726
rect 195840 77656 196052 77662
rect 196248 77726 196460 77868
rect 196248 77662 196390 77726
rect 196454 77662 196460 77726
rect 196248 77656 196460 77662
rect 196656 77862 196868 77868
rect 196656 77798 196662 77862
rect 196726 77798 196868 77862
rect 196656 77726 196868 77798
rect 196656 77662 196798 77726
rect 196862 77662 196868 77726
rect 196656 77656 196868 77662
rect 216784 77862 217540 77868
rect 216784 77812 217470 77862
rect 216784 77756 216908 77812
rect 216964 77798 217470 77812
rect 217534 77798 217540 77862
rect 216964 77792 217540 77798
rect 216964 77756 216996 77792
rect 216784 77656 216996 77756
rect 28560 77596 28636 77656
rect 190264 77596 190340 77656
rect 21760 77454 21972 77460
rect 21760 77390 21902 77454
rect 21966 77390 21972 77454
rect 21760 77248 21972 77390
rect 22168 77324 22380 77460
rect 22478 77454 22788 77460
rect 22440 77390 22446 77454
rect 22510 77390 22788 77454
rect 22478 77384 22788 77390
rect 22576 77324 22788 77384
rect 22168 77318 22788 77324
rect 22168 77254 22310 77318
rect 22374 77254 22788 77318
rect 22168 77248 22788 77254
rect 22984 77454 23196 77460
rect 22984 77390 22990 77454
rect 23054 77390 23196 77454
rect 22984 77318 23196 77390
rect 22984 77254 22990 77318
rect 23054 77254 23196 77318
rect 22984 77248 23196 77254
rect 23392 77454 23604 77460
rect 23392 77390 23398 77454
rect 23462 77390 23604 77454
rect 23392 77318 23604 77390
rect 28288 77384 28636 77596
rect 190128 77384 190340 77596
rect 28424 77324 28500 77384
rect 190264 77324 190340 77384
rect 23392 77254 23534 77318
rect 23598 77254 23604 77318
rect 23392 77248 23604 77254
rect 21760 77188 21836 77248
rect 22304 77188 22380 77248
rect 21760 76840 21972 77188
rect 22304 77112 22652 77188
rect 22576 77052 22652 77112
rect 28288 77112 28636 77324
rect 190128 77182 190340 77324
rect 195024 77454 195236 77460
rect 195024 77390 195030 77454
rect 195094 77390 195236 77454
rect 195024 77318 195236 77390
rect 195024 77254 195166 77318
rect 195230 77254 195236 77318
rect 195024 77248 195236 77254
rect 195432 77454 195644 77460
rect 195432 77390 195438 77454
rect 195502 77390 195644 77454
rect 195432 77318 195644 77390
rect 195432 77254 195438 77318
rect 195502 77254 195644 77318
rect 195432 77248 195644 77254
rect 195840 77454 196460 77460
rect 195840 77390 195982 77454
rect 196046 77390 196390 77454
rect 196454 77390 196460 77454
rect 195840 77384 196460 77390
rect 195840 77318 196052 77384
rect 195840 77254 195846 77318
rect 195910 77254 196052 77318
rect 195840 77248 196052 77254
rect 196248 77318 196460 77384
rect 196248 77254 196390 77318
rect 196454 77254 196460 77318
rect 196248 77248 196460 77254
rect 196656 77454 196868 77460
rect 196656 77390 196798 77454
rect 196862 77390 196868 77454
rect 196656 77248 196868 77390
rect 196792 77188 196868 77248
rect 190128 77118 190134 77182
rect 190198 77118 190340 77182
rect 190128 77112 190340 77118
rect 28288 77052 28364 77112
rect 190128 77052 190204 77112
rect 21896 76780 21972 76840
rect 21760 76432 21972 76780
rect 22168 77046 22380 77052
rect 22168 76982 22310 77046
rect 22374 76982 22380 77046
rect 22168 76840 22380 76982
rect 22576 76840 22788 77052
rect 22984 77046 23196 77052
rect 22984 76982 22990 77046
rect 23054 76982 23196 77046
rect 22984 76910 23196 76982
rect 22984 76846 22990 76910
rect 23054 76846 23196 76910
rect 22984 76840 23196 76846
rect 23392 77046 23604 77052
rect 23392 76982 23534 77046
rect 23598 76982 23604 77046
rect 23392 76910 23604 76982
rect 23392 76846 23534 76910
rect 23598 76846 23604 76910
rect 23392 76840 23604 76846
rect 22168 76780 22244 76840
rect 22576 76780 22652 76840
rect 22168 76508 22380 76780
rect 22168 76502 22516 76508
rect 22168 76438 22310 76502
rect 22374 76438 22446 76502
rect 22510 76438 22516 76502
rect 22168 76432 22516 76438
rect 22576 76432 22788 76780
rect 22984 76638 23196 76644
rect 22984 76574 22990 76638
rect 23054 76574 23196 76638
rect 22984 76432 23196 76574
rect 23392 76638 23604 76644
rect 23392 76574 23534 76638
rect 23598 76574 23604 76638
rect 23392 76432 23604 76574
rect 28288 76568 28636 77052
rect 190128 76910 190340 77052
rect 190128 76846 190134 76910
rect 190198 76846 190340 76910
rect 190128 76568 190340 76846
rect 195024 77046 195236 77052
rect 195024 76982 195166 77046
rect 195230 76982 195236 77046
rect 195024 76910 195236 76982
rect 195024 76846 195166 76910
rect 195230 76846 195236 76910
rect 195024 76840 195236 76846
rect 195432 77046 195644 77052
rect 195432 76982 195438 77046
rect 195502 76982 195644 77046
rect 195432 76910 195644 76982
rect 195432 76846 195438 76910
rect 195502 76846 195644 76910
rect 195432 76840 195644 76846
rect 195840 77046 196052 77052
rect 195840 76982 195846 77046
rect 195910 76982 196052 77046
rect 195840 76840 196052 76982
rect 196248 77046 196460 77052
rect 196248 76982 196390 77046
rect 196454 76982 196460 77046
rect 196248 76840 196460 76982
rect 196656 76840 196868 77188
rect 196248 76780 196324 76840
rect 196792 76780 196868 76840
rect 195840 76644 196052 76780
rect 196248 76644 196460 76780
rect 28424 76508 28500 76568
rect 190264 76508 190340 76568
rect 21760 76372 21836 76432
rect 22984 76372 23060 76432
rect 23392 76372 23468 76432
rect 1224 76230 1844 76236
rect 1224 76166 1230 76230
rect 1294 76166 1844 76230
rect 1224 76160 1844 76166
rect 21760 76230 21972 76372
rect 21760 76166 21766 76230
rect 21830 76166 21972 76230
rect 21760 76160 21972 76166
rect 22168 76230 22380 76236
rect 22478 76230 22788 76236
rect 22168 76166 22310 76230
rect 22374 76166 22380 76230
rect 22440 76166 22446 76230
rect 22510 76166 22788 76230
rect 1632 76132 1844 76160
rect 1632 76076 1702 76132
rect 1758 76076 1844 76132
rect 1632 76024 1844 76076
rect 22168 76024 22380 76166
rect 22478 76160 22788 76166
rect 22576 76024 22788 76160
rect 22984 76024 23196 76372
rect 23392 76024 23604 76372
rect 28288 76366 28636 76508
rect 28288 76302 28566 76366
rect 28630 76302 28636 76366
rect 28288 76296 28636 76302
rect 190128 76366 190340 76508
rect 190128 76302 190270 76366
rect 190334 76302 190340 76366
rect 28404 76100 28502 76296
rect 22168 75964 22244 76024
rect 23120 75964 23196 76024
rect 23528 75964 23604 76024
rect 21760 75958 21972 75964
rect 21760 75894 21766 75958
rect 21830 75894 21972 75958
rect 21760 75822 21972 75894
rect 21760 75758 21766 75822
rect 21830 75758 21972 75822
rect 21760 75752 21972 75758
rect 22168 75822 22380 75964
rect 22576 75828 22788 75964
rect 22478 75822 22788 75828
rect 22168 75758 22174 75822
rect 22238 75758 22380 75822
rect 22440 75758 22446 75822
rect 22510 75758 22788 75822
rect 22168 75752 22380 75758
rect 22478 75752 22788 75758
rect 22984 75692 23196 75964
rect 23392 75692 23604 75964
rect 28288 76094 28636 76100
rect 28288 76030 28566 76094
rect 28630 76030 28636 76094
rect 28288 75958 28636 76030
rect 28288 75894 28430 75958
rect 28494 75894 28636 75958
rect 28288 75888 28636 75894
rect 190128 76094 190340 76302
rect 190128 76030 190270 76094
rect 190334 76030 190340 76094
rect 190128 75958 190340 76030
rect 195024 76638 195236 76644
rect 195024 76574 195166 76638
rect 195230 76574 195236 76638
rect 195024 76432 195236 76574
rect 195432 76638 195644 76644
rect 195432 76574 195438 76638
rect 195502 76574 195644 76638
rect 195432 76432 195644 76574
rect 195840 76568 196460 76644
rect 195840 76508 196052 76568
rect 195840 76502 196188 76508
rect 195840 76438 195846 76502
rect 195910 76438 196118 76502
rect 196182 76438 196188 76502
rect 195840 76432 196188 76438
rect 196248 76432 196460 76568
rect 196656 76432 196868 76780
rect 195024 76372 195100 76432
rect 195432 76372 195508 76432
rect 196792 76372 196868 76432
rect 195024 76024 195236 76372
rect 195160 75964 195236 76024
rect 190128 75894 190134 75958
rect 190198 75894 190340 75958
rect 190128 75888 190340 75894
rect 22984 75686 23332 75692
rect 22984 75622 23262 75686
rect 23326 75622 23332 75686
rect 22984 75616 23332 75622
rect 23392 75616 24284 75692
rect 23120 75556 23196 75616
rect 21760 75550 21972 75556
rect 21760 75486 21766 75550
rect 21830 75486 21972 75550
rect 21760 75414 21972 75486
rect 21760 75350 21902 75414
rect 21966 75350 21972 75414
rect 21760 75344 21972 75350
rect 22168 75550 22516 75556
rect 22168 75486 22174 75550
rect 22238 75486 22446 75550
rect 22510 75486 22516 75550
rect 22168 75480 22516 75486
rect 22168 75284 22380 75480
rect 22576 75284 22788 75556
rect 22984 75414 23196 75556
rect 22984 75350 23126 75414
rect 23190 75350 23196 75414
rect 22984 75344 23196 75350
rect 23392 75556 23468 75616
rect 24208 75556 24284 75616
rect 26792 75686 28636 75692
rect 26792 75622 28430 75686
rect 28494 75622 28636 75686
rect 26792 75616 28636 75622
rect 26792 75556 26868 75616
rect 23392 75414 23604 75556
rect 23392 75350 23398 75414
rect 23462 75350 23604 75414
rect 23392 75344 23604 75350
rect 23800 75284 24012 75556
rect 24208 75284 24556 75556
rect 25296 75480 26868 75556
rect 25296 75414 25508 75480
rect 25296 75350 25302 75414
rect 25366 75350 25508 75414
rect 25296 75344 25508 75350
rect 26928 75344 27140 75556
rect 28288 75550 28636 75616
rect 28288 75486 28430 75550
rect 28494 75486 28636 75550
rect 28288 75344 28636 75486
rect 190128 75686 190340 75692
rect 190128 75622 190134 75686
rect 190198 75622 190340 75686
rect 190128 75550 190340 75622
rect 194072 75616 194692 75692
rect 195024 75616 195236 75964
rect 195432 76024 195644 76372
rect 195840 76230 196052 76236
rect 196150 76230 196460 76236
rect 195840 76166 195846 76230
rect 195910 76166 196052 76230
rect 196112 76166 196118 76230
rect 196182 76166 196460 76230
rect 195840 76024 196052 76166
rect 196150 76160 196460 76166
rect 196656 76230 196868 76372
rect 196656 76166 196798 76230
rect 196862 76166 196868 76230
rect 196656 76160 196868 76166
rect 196248 76024 196460 76160
rect 216784 76132 216996 76236
rect 216784 76076 216908 76132
rect 216964 76100 216996 76132
rect 216964 76094 217540 76100
rect 216964 76076 217470 76094
rect 216784 76030 217470 76076
rect 217534 76030 217540 76094
rect 216784 76024 217540 76030
rect 195432 75964 195508 76024
rect 195840 75964 195916 76024
rect 196248 75964 196324 76024
rect 195432 75616 195644 75964
rect 195840 75752 196052 75964
rect 196248 75828 196460 75964
rect 196150 75822 196460 75828
rect 196112 75758 196118 75822
rect 196182 75758 196390 75822
rect 196454 75758 196460 75822
rect 196150 75752 196460 75758
rect 196656 75958 196868 75964
rect 196656 75894 196798 75958
rect 196862 75894 196868 75958
rect 196656 75822 196868 75894
rect 196656 75758 196662 75822
rect 196726 75758 196868 75822
rect 196656 75752 196868 75758
rect 194072 75556 194148 75616
rect 194616 75556 194692 75616
rect 195160 75556 195236 75616
rect 195568 75556 195644 75616
rect 190128 75486 190270 75550
rect 190334 75486 190340 75550
rect 190128 75344 190340 75486
rect 191488 75420 191700 75556
rect 193120 75480 194148 75556
rect 191488 75344 193060 75420
rect 193120 75414 193332 75480
rect 193120 75350 193126 75414
rect 193190 75350 193332 75414
rect 193120 75344 193332 75350
rect 26928 75284 27004 75344
rect 22168 75208 22788 75284
rect 23294 75278 24148 75284
rect 23256 75214 23262 75278
rect 23326 75214 24148 75278
rect 23294 75208 24148 75214
rect 24208 75208 27004 75284
rect 28288 75284 28364 75344
rect 190264 75284 190340 75344
rect 28288 75278 28636 75284
rect 28288 75214 28430 75278
rect 28494 75214 28636 75278
rect 22712 75148 22788 75208
rect 24072 75148 24148 75208
rect 21760 75142 21972 75148
rect 21760 75078 21902 75142
rect 21966 75078 21972 75142
rect 21760 75006 21972 75078
rect 21760 74942 21766 75006
rect 21830 74942 21972 75006
rect 21760 74936 21972 74942
rect 22168 75012 22380 75148
rect 22576 75012 22788 75148
rect 22168 75006 22788 75012
rect 22168 74942 22174 75006
rect 22238 74942 22788 75006
rect 22168 74936 22788 74942
rect 22984 75142 23196 75148
rect 22984 75078 23126 75142
rect 23190 75078 23196 75142
rect 22984 75006 23196 75078
rect 22984 74942 22990 75006
rect 23054 74942 23196 75006
rect 22984 74936 23196 74942
rect 23392 75142 23604 75148
rect 23392 75078 23398 75142
rect 23462 75078 23604 75142
rect 23392 75006 23604 75078
rect 24072 75142 25372 75148
rect 24072 75078 25302 75142
rect 25366 75078 25372 75142
rect 24072 75072 25372 75078
rect 28288 75072 28636 75214
rect 190128 75278 190340 75284
rect 190128 75214 190270 75278
rect 190334 75214 190340 75278
rect 190128 75148 190340 75214
rect 192984 75284 193060 75344
rect 194208 75284 194420 75556
rect 194616 75284 194828 75556
rect 195024 75414 195236 75556
rect 195024 75350 195030 75414
rect 195094 75350 195236 75414
rect 195024 75344 195236 75350
rect 195432 75414 195644 75556
rect 195432 75350 195438 75414
rect 195502 75350 195644 75414
rect 195432 75344 195644 75350
rect 195840 75550 196188 75556
rect 195840 75486 196118 75550
rect 196182 75486 196188 75550
rect 195840 75480 196188 75486
rect 196248 75550 196460 75556
rect 196248 75486 196390 75550
rect 196454 75486 196460 75550
rect 192984 75208 194556 75284
rect 194616 75208 195508 75284
rect 195840 75208 196052 75480
rect 196248 75284 196460 75486
rect 196656 75550 196868 75556
rect 196656 75486 196662 75550
rect 196726 75486 196868 75550
rect 196656 75414 196868 75486
rect 196656 75350 196798 75414
rect 196862 75350 196868 75414
rect 196656 75344 196868 75350
rect 196112 75208 196460 75284
rect 194480 75148 194556 75208
rect 195432 75148 195508 75208
rect 196112 75148 196188 75208
rect 190128 75142 193196 75148
rect 190128 75078 193126 75142
rect 193190 75078 193196 75142
rect 190128 75072 193196 75078
rect 194480 75142 195236 75148
rect 194480 75078 195030 75142
rect 195094 75078 195236 75142
rect 194480 75072 195236 75078
rect 23392 74942 23534 75006
rect 23598 74942 23604 75006
rect 23392 74936 23604 74942
rect 28288 75012 28364 75072
rect 190264 75012 190340 75072
rect 22304 74876 22380 74936
rect 22304 74800 22652 74876
rect 22576 74740 22652 74800
rect 21760 74734 21972 74740
rect 21760 74670 21766 74734
rect 21830 74670 21972 74734
rect 1224 74598 1844 74604
rect 1224 74534 1230 74598
rect 1294 74534 1844 74598
rect 1224 74528 1844 74534
rect 21760 74598 21972 74670
rect 21760 74534 21766 74598
rect 21830 74534 21972 74598
rect 21760 74528 21972 74534
rect 22168 74734 22380 74740
rect 22168 74670 22174 74734
rect 22238 74670 22380 74734
rect 22168 74528 22380 74670
rect 22576 74528 22788 74740
rect 22984 74734 23196 74740
rect 22984 74670 22990 74734
rect 23054 74670 23196 74734
rect 22984 74598 23196 74670
rect 22984 74534 22990 74598
rect 23054 74534 23196 74598
rect 22984 74528 23196 74534
rect 23392 74734 23604 74740
rect 23392 74670 23534 74734
rect 23598 74670 23604 74734
rect 23392 74598 23604 74670
rect 23392 74534 23534 74598
rect 23598 74534 23604 74598
rect 23392 74528 23604 74534
rect 28288 74528 28636 75012
rect 190128 74528 190340 75012
rect 195024 75006 195236 75072
rect 195024 74942 195166 75006
rect 195230 74942 195236 75006
rect 195024 74936 195236 74942
rect 195432 75142 195644 75148
rect 195432 75078 195438 75142
rect 195502 75078 195644 75142
rect 195432 75006 195644 75078
rect 195432 74942 195438 75006
rect 195502 74942 195644 75006
rect 195432 74936 195644 74942
rect 195840 75072 196188 75148
rect 195840 75012 196052 75072
rect 196248 75012 196460 75148
rect 195840 75006 196460 75012
rect 195840 74942 196254 75006
rect 196318 74942 196460 75006
rect 195840 74936 196460 74942
rect 196656 75142 196868 75148
rect 196656 75078 196798 75142
rect 196862 75078 196868 75142
rect 196656 75006 196868 75078
rect 196656 74942 196662 75006
rect 196726 74942 196868 75006
rect 196656 74936 196868 74942
rect 195024 74734 195236 74740
rect 195024 74670 195166 74734
rect 195230 74670 195236 74734
rect 195024 74598 195236 74670
rect 195024 74534 195166 74598
rect 195230 74534 195236 74598
rect 195024 74528 195236 74534
rect 195432 74734 195644 74740
rect 195432 74670 195438 74734
rect 195502 74670 195644 74734
rect 195432 74598 195644 74670
rect 195432 74534 195438 74598
rect 195502 74534 195644 74598
rect 195432 74528 195644 74534
rect 195840 74598 196052 74740
rect 195840 74534 195846 74598
rect 195910 74534 196052 74598
rect 195840 74528 196052 74534
rect 196248 74734 196460 74740
rect 196248 74670 196254 74734
rect 196318 74670 196460 74734
rect 196248 74598 196460 74670
rect 196248 74534 196390 74598
rect 196454 74534 196460 74598
rect 196248 74528 196460 74534
rect 196656 74734 196868 74740
rect 196656 74670 196662 74734
rect 196726 74670 196868 74734
rect 196656 74598 196868 74670
rect 196656 74534 196798 74598
rect 196862 74534 196868 74598
rect 196656 74528 196868 74534
rect 216784 74598 217540 74604
rect 216784 74534 217470 74598
rect 217534 74534 217540 74598
rect 216784 74528 217540 74534
rect 1632 74452 1844 74528
rect 22576 74468 22652 74528
rect 28560 74468 28636 74528
rect 190264 74468 190340 74528
rect 1632 74396 1702 74452
rect 1758 74396 1844 74452
rect 1632 74256 1844 74396
rect 22304 74392 22652 74468
rect 22304 74332 22380 74392
rect 21760 74326 21972 74332
rect 21760 74262 21766 74326
rect 21830 74262 21972 74326
rect 21760 74190 21972 74262
rect 21760 74126 21766 74190
rect 21830 74126 21972 74190
rect 21760 74120 21972 74126
rect 22168 74256 22788 74332
rect 22168 74190 22380 74256
rect 22168 74126 22174 74190
rect 22238 74126 22380 74190
rect 22168 74120 22380 74126
rect 22576 74190 22788 74256
rect 22576 74126 22718 74190
rect 22782 74126 22788 74190
rect 22576 74120 22788 74126
rect 22984 74326 23196 74332
rect 22984 74262 22990 74326
rect 23054 74262 23196 74326
rect 22984 74190 23196 74262
rect 22984 74126 22990 74190
rect 23054 74126 23196 74190
rect 22984 74120 23196 74126
rect 23392 74326 23604 74332
rect 23392 74262 23534 74326
rect 23598 74262 23604 74326
rect 23392 74190 23604 74262
rect 28288 74256 28636 74468
rect 190128 74256 190340 74468
rect 216784 74452 216996 74528
rect 216784 74396 216908 74452
rect 216964 74396 216996 74452
rect 28560 74196 28636 74256
rect 190264 74196 190340 74256
rect 23392 74126 23534 74190
rect 23598 74126 23604 74190
rect 23392 74120 23604 74126
rect 28288 73984 28636 74196
rect 190128 73984 190340 74196
rect 195024 74326 195236 74332
rect 195024 74262 195166 74326
rect 195230 74262 195236 74326
rect 195024 74190 195236 74262
rect 195024 74126 195166 74190
rect 195230 74126 195236 74190
rect 195024 74120 195236 74126
rect 195432 74326 195644 74332
rect 195432 74262 195438 74326
rect 195502 74262 195644 74326
rect 195432 74190 195644 74262
rect 195432 74126 195438 74190
rect 195502 74126 195644 74190
rect 195432 74120 195644 74126
rect 195840 74326 196460 74332
rect 195840 74262 195846 74326
rect 195910 74262 196390 74326
rect 196454 74262 196460 74326
rect 195840 74256 196460 74262
rect 195840 74196 196052 74256
rect 195840 74190 196188 74196
rect 195840 74126 196118 74190
rect 196182 74126 196188 74190
rect 195840 74120 196188 74126
rect 196248 74120 196460 74256
rect 196656 74326 196868 74332
rect 196656 74262 196798 74326
rect 196862 74262 196868 74326
rect 196656 74190 196868 74262
rect 216784 74256 216996 74396
rect 196656 74126 196662 74190
rect 196726 74126 196868 74190
rect 196656 74120 196868 74126
rect 28424 73924 28500 73984
rect 190264 73924 190340 73984
rect 21760 73918 21972 73924
rect 21760 73854 21766 73918
rect 21830 73854 21972 73918
rect 21760 73782 21972 73854
rect 21760 73718 21766 73782
rect 21830 73718 21972 73782
rect 21760 73712 21972 73718
rect 22168 73918 22380 73924
rect 22168 73854 22174 73918
rect 22238 73854 22380 73918
rect 22168 73712 22380 73854
rect 22576 73918 22788 73924
rect 22576 73854 22718 73918
rect 22782 73854 22788 73918
rect 22576 73782 22788 73854
rect 22576 73718 22582 73782
rect 22646 73718 22788 73782
rect 22576 73712 22788 73718
rect 22984 73918 23196 73924
rect 22984 73854 22990 73918
rect 23054 73854 23196 73918
rect 22984 73782 23196 73854
rect 22984 73718 23126 73782
rect 23190 73718 23196 73782
rect 22984 73712 23196 73718
rect 23392 73918 23604 73924
rect 23392 73854 23534 73918
rect 23598 73854 23604 73918
rect 23392 73782 23604 73854
rect 23392 73718 23534 73782
rect 23598 73718 23604 73782
rect 23392 73712 23604 73718
rect 28288 73712 28636 73924
rect 190128 73712 190340 73924
rect 195024 73918 195236 73924
rect 195024 73854 195166 73918
rect 195230 73854 195236 73918
rect 195024 73782 195236 73854
rect 195024 73718 195166 73782
rect 195230 73718 195236 73782
rect 195024 73712 195236 73718
rect 195432 73918 195644 73924
rect 195432 73854 195438 73918
rect 195502 73854 195644 73918
rect 195432 73782 195644 73854
rect 195432 73718 195574 73782
rect 195638 73718 195644 73782
rect 195432 73712 195644 73718
rect 195840 73782 196052 73924
rect 196150 73918 196460 73924
rect 196112 73854 196118 73918
rect 196182 73854 196460 73918
rect 196150 73848 196460 73854
rect 195840 73718 195846 73782
rect 195910 73718 196052 73782
rect 195840 73712 196052 73718
rect 196248 73782 196460 73848
rect 196248 73718 196254 73782
rect 196318 73718 196460 73782
rect 196248 73712 196460 73718
rect 196656 73918 196868 73924
rect 196656 73854 196662 73918
rect 196726 73854 196868 73918
rect 196656 73782 196868 73854
rect 196656 73718 196662 73782
rect 196726 73718 196868 73782
rect 196656 73712 196868 73718
rect 28424 73652 28500 73712
rect 190128 73652 190204 73712
rect 21760 73510 21972 73516
rect 21760 73446 21766 73510
rect 21830 73446 21972 73510
rect 21760 73304 21972 73446
rect 22168 73374 22380 73516
rect 22168 73310 22174 73374
rect 22238 73310 22380 73374
rect 22168 73304 22380 73310
rect 22576 73510 22788 73516
rect 22576 73446 22582 73510
rect 22646 73446 22788 73510
rect 22576 73374 22788 73446
rect 22576 73310 22718 73374
rect 22782 73310 22788 73374
rect 22576 73304 22788 73310
rect 22984 73510 23196 73516
rect 22984 73446 23126 73510
rect 23190 73446 23196 73510
rect 22984 73374 23196 73446
rect 22984 73310 23126 73374
rect 23190 73310 23196 73374
rect 22984 73304 23196 73310
rect 23392 73510 23604 73516
rect 23392 73446 23534 73510
rect 23598 73446 23604 73510
rect 23392 73374 23604 73446
rect 23392 73310 23398 73374
rect 23462 73310 23604 73374
rect 23392 73304 23604 73310
rect 28288 73440 28636 73652
rect 190128 73440 190340 73652
rect 28288 73380 28364 73440
rect 190264 73380 190340 73440
rect 21760 73244 21836 73304
rect 21760 72896 21972 73244
rect 28288 73168 28636 73380
rect 190128 73168 190340 73380
rect 195024 73510 195236 73516
rect 195024 73446 195166 73510
rect 195230 73446 195236 73510
rect 195024 73374 195236 73446
rect 195024 73310 195030 73374
rect 195094 73310 195236 73374
rect 195024 73304 195236 73310
rect 195432 73510 195644 73516
rect 195432 73446 195574 73510
rect 195638 73446 195644 73510
rect 195432 73374 195644 73446
rect 195432 73310 195438 73374
rect 195502 73310 195644 73374
rect 195432 73304 195644 73310
rect 195840 73510 196052 73516
rect 195840 73446 195846 73510
rect 195910 73446 196052 73510
rect 195840 73374 196052 73446
rect 196248 73510 196460 73516
rect 196248 73446 196254 73510
rect 196318 73446 196460 73510
rect 196248 73380 196460 73446
rect 196150 73374 196460 73380
rect 195840 73310 195982 73374
rect 196046 73310 196052 73374
rect 196112 73310 196118 73374
rect 196182 73310 196460 73374
rect 195840 73304 196052 73310
rect 196150 73304 196460 73310
rect 196656 73510 196868 73516
rect 196656 73446 196662 73510
rect 196726 73446 196868 73510
rect 196656 73304 196868 73446
rect 196792 73244 196868 73304
rect 28424 73108 28500 73168
rect 190264 73108 190340 73168
rect 195976 73168 196324 73244
rect 195976 73108 196052 73168
rect 196248 73108 196324 73168
rect 22168 73102 22380 73108
rect 22168 73038 22174 73102
rect 22238 73038 22380 73102
rect 22168 72972 22380 73038
rect 22576 73102 22788 73108
rect 22576 73038 22718 73102
rect 22782 73038 22788 73102
rect 22168 72896 22516 72972
rect 22576 72896 22788 73038
rect 22984 73102 23196 73108
rect 22984 73038 23126 73102
rect 23190 73038 23196 73102
rect 22984 72966 23196 73038
rect 22984 72902 23126 72966
rect 23190 72902 23196 72966
rect 22984 72896 23196 72902
rect 23392 73102 23604 73108
rect 23392 73038 23398 73102
rect 23462 73038 23604 73102
rect 23392 72966 23604 73038
rect 23392 72902 23534 72966
rect 23598 72902 23604 72966
rect 23392 72896 23604 72902
rect 28288 72966 28636 73108
rect 28288 72902 28294 72966
rect 28358 72902 28636 72966
rect 21896 72836 21972 72896
rect 22304 72836 22380 72896
rect 1632 72772 1844 72836
rect 1632 72716 1702 72772
rect 1758 72716 1844 72772
rect 1632 72700 1844 72716
rect 1224 72694 1844 72700
rect 1224 72630 1230 72694
rect 1294 72630 1844 72694
rect 1224 72624 1844 72630
rect 21760 72488 21972 72836
rect 22168 72488 22380 72836
rect 22440 72836 22516 72896
rect 22712 72836 22788 72896
rect 22440 72760 22788 72836
rect 22576 72558 22788 72760
rect 22576 72494 22718 72558
rect 22782 72494 22788 72558
rect 22576 72488 22788 72494
rect 22984 72694 23196 72700
rect 22984 72630 23126 72694
rect 23190 72630 23196 72694
rect 22984 72558 23196 72630
rect 22984 72494 22990 72558
rect 23054 72494 23196 72558
rect 22984 72488 23196 72494
rect 23392 72694 23604 72700
rect 23392 72630 23534 72694
rect 23598 72630 23604 72694
rect 23392 72558 23604 72630
rect 23392 72494 23398 72558
rect 23462 72494 23604 72558
rect 23392 72488 23604 72494
rect 28288 72624 28636 72902
rect 190128 72624 190340 73108
rect 195024 73102 195236 73108
rect 195024 73038 195030 73102
rect 195094 73038 195236 73102
rect 195024 72966 195236 73038
rect 195024 72902 195030 72966
rect 195094 72902 195236 72966
rect 195024 72896 195236 72902
rect 195432 73102 195644 73108
rect 195432 73038 195438 73102
rect 195502 73038 195644 73102
rect 195432 72966 195644 73038
rect 195432 72902 195574 72966
rect 195638 72902 195644 72966
rect 195432 72896 195644 72902
rect 195840 73102 196188 73108
rect 195840 73038 195982 73102
rect 196046 73038 196118 73102
rect 196182 73038 196188 73102
rect 195840 73032 196188 73038
rect 195840 72972 196052 73032
rect 195840 72896 196188 72972
rect 196248 72896 196460 73108
rect 196656 72896 196868 73244
rect 195840 72836 195916 72896
rect 196112 72836 196188 72896
rect 196792 72836 196868 72896
rect 195024 72694 195236 72700
rect 195024 72630 195030 72694
rect 195094 72630 195236 72694
rect 28288 72564 28364 72624
rect 190128 72564 190204 72624
rect 28288 72558 28636 72564
rect 28288 72494 28294 72558
rect 28358 72494 28636 72558
rect 21760 72428 21836 72488
rect 21760 72286 21972 72428
rect 28288 72422 28636 72494
rect 28288 72358 28566 72422
rect 28630 72358 28636 72422
rect 28288 72352 28636 72358
rect 190128 72352 190340 72564
rect 195024 72558 195236 72630
rect 195024 72494 195030 72558
rect 195094 72494 195236 72558
rect 195024 72488 195236 72494
rect 195432 72694 195644 72700
rect 195432 72630 195574 72694
rect 195638 72630 195644 72694
rect 195432 72558 195644 72630
rect 195432 72494 195438 72558
rect 195502 72494 195644 72558
rect 195432 72488 195644 72494
rect 195840 72488 196052 72836
rect 196112 72760 196460 72836
rect 196248 72564 196460 72760
rect 196150 72558 196460 72564
rect 196112 72494 196118 72558
rect 196182 72494 196460 72558
rect 196150 72488 196460 72494
rect 196656 72488 196868 72836
rect 216784 72830 217540 72836
rect 216784 72772 217470 72830
rect 216784 72716 216908 72772
rect 216964 72766 217470 72772
rect 217534 72766 217540 72830
rect 216964 72760 217540 72766
rect 216964 72716 216996 72760
rect 216784 72624 216996 72716
rect 196792 72428 196868 72488
rect 28424 72292 28500 72352
rect 190264 72292 190340 72352
rect 21760 72222 21902 72286
rect 21966 72222 21972 72286
rect 21760 72216 21972 72222
rect 22168 72156 22380 72292
rect 22576 72286 22788 72292
rect 22576 72222 22718 72286
rect 22782 72222 22788 72286
rect 22576 72156 22788 72222
rect 22168 72080 22788 72156
rect 22304 72020 22380 72080
rect 22712 72020 22788 72080
rect 21760 72014 21972 72020
rect 21760 71950 21902 72014
rect 21966 71950 21972 72014
rect 21760 71878 21972 71950
rect 21760 71814 21902 71878
rect 21966 71814 21972 71878
rect 21760 71808 21972 71814
rect 22168 71884 22380 72020
rect 22168 71878 22516 71884
rect 22168 71814 22310 71878
rect 22374 71814 22446 71878
rect 22510 71814 22516 71878
rect 22168 71808 22516 71814
rect 22576 71808 22788 72020
rect 22984 72286 23196 72292
rect 22984 72222 22990 72286
rect 23054 72222 23196 72286
rect 22984 72080 23196 72222
rect 23392 72286 23604 72292
rect 23392 72222 23398 72286
rect 23462 72222 23604 72286
rect 23392 72080 23604 72222
rect 28288 72150 28636 72292
rect 28288 72086 28566 72150
rect 28630 72086 28636 72150
rect 22984 72020 23060 72080
rect 23392 72020 23468 72080
rect 22984 71672 23196 72020
rect 23392 71672 23604 72020
rect 28288 72014 28636 72086
rect 28288 71950 28566 72014
rect 28630 71950 28636 72014
rect 28288 71944 28636 71950
rect 190128 72014 190340 72292
rect 190128 71950 190134 72014
rect 190198 71950 190340 72014
rect 190128 71944 190340 71950
rect 195024 72286 195236 72292
rect 195024 72222 195030 72286
rect 195094 72222 195236 72286
rect 195024 72080 195236 72222
rect 195432 72286 195644 72292
rect 195432 72222 195438 72286
rect 195502 72222 195644 72286
rect 195432 72080 195644 72222
rect 195840 72286 196188 72292
rect 195840 72222 196118 72286
rect 196182 72222 196188 72286
rect 195840 72216 196188 72222
rect 195840 72080 196052 72216
rect 196248 72080 196460 72292
rect 196656 72286 196868 72428
rect 196656 72222 196798 72286
rect 196862 72222 196868 72286
rect 196656 72216 196868 72222
rect 195024 72020 195100 72080
rect 195432 72020 195508 72080
rect 195976 72020 196052 72080
rect 196384 72020 196460 72080
rect 22984 71612 23060 71672
rect 23528 71612 23604 71672
rect 21760 71606 21972 71612
rect 21760 71542 21902 71606
rect 21966 71542 21972 71606
rect 21760 71470 21972 71542
rect 21760 71406 21902 71470
rect 21966 71406 21972 71470
rect 21760 71400 21972 71406
rect 22168 71606 22380 71612
rect 22478 71606 22788 71612
rect 22168 71542 22310 71606
rect 22374 71542 22380 71606
rect 22440 71542 22446 71606
rect 22510 71542 22788 71606
rect 22168 71264 22380 71542
rect 22478 71536 22788 71542
rect 22576 71264 22788 71536
rect 22304 71204 22380 71264
rect 22712 71204 22788 71264
rect 1632 71092 1844 71204
rect 1632 71068 1702 71092
rect 1224 71062 1702 71068
rect 1224 70998 1230 71062
rect 1294 71036 1702 71062
rect 1758 71036 1844 71092
rect 1294 70998 1844 71036
rect 1224 70992 1844 70998
rect 21760 71198 21972 71204
rect 21760 71134 21902 71198
rect 21966 71134 21972 71198
rect 21760 71062 21972 71134
rect 21760 70998 21902 71062
rect 21966 70998 21972 71062
rect 21760 70992 21972 70998
rect 22168 71068 22380 71204
rect 22168 70992 22516 71068
rect 22576 70992 22788 71204
rect 22984 71264 23196 71612
rect 23392 71264 23604 71612
rect 22984 71204 23060 71264
rect 23528 71204 23604 71264
rect 22984 71062 23196 71204
rect 22984 70998 22990 71062
rect 23054 70998 23196 71062
rect 22984 70992 23196 70998
rect 23392 71062 23604 71204
rect 28288 71742 28636 71748
rect 28288 71678 28566 71742
rect 28630 71678 28636 71742
rect 28288 71334 28636 71678
rect 28288 71270 28430 71334
rect 28494 71270 28636 71334
rect 28288 71198 28636 71270
rect 28288 71134 28294 71198
rect 28358 71134 28636 71198
rect 28288 71128 28636 71134
rect 190128 71742 190340 71748
rect 190128 71678 190134 71742
rect 190198 71678 190340 71742
rect 190128 71606 190340 71678
rect 195024 71672 195236 72020
rect 195160 71612 195236 71672
rect 190128 71542 190134 71606
rect 190198 71542 190340 71606
rect 190128 71334 190340 71542
rect 190128 71270 190134 71334
rect 190198 71270 190270 71334
rect 190334 71270 190340 71334
rect 190128 71128 190340 71270
rect 195024 71264 195236 71612
rect 195432 71672 195644 72020
rect 195840 71944 196460 72020
rect 195840 71808 196052 71944
rect 196248 71878 196460 71944
rect 196248 71814 196390 71878
rect 196454 71814 196460 71878
rect 196248 71808 196460 71814
rect 196656 72014 196868 72020
rect 196656 71950 196798 72014
rect 196862 71950 196868 72014
rect 196656 71878 196868 71950
rect 196656 71814 196798 71878
rect 196862 71814 196868 71878
rect 196656 71808 196868 71814
rect 195432 71612 195508 71672
rect 195432 71264 195644 71612
rect 195160 71204 195236 71264
rect 195568 71204 195644 71264
rect 190264 71068 190340 71128
rect 23392 70998 23398 71062
rect 23462 70998 23604 71062
rect 23392 70992 23604 70998
rect 28288 71062 28636 71068
rect 28288 70998 28430 71062
rect 28494 70998 28636 71062
rect 22440 70932 22516 70992
rect 22440 70856 22652 70932
rect 22576 70796 22652 70856
rect 21760 70790 21972 70796
rect 21760 70726 21902 70790
rect 21966 70726 21972 70790
rect 21760 70654 21972 70726
rect 21760 70590 21766 70654
rect 21830 70590 21972 70654
rect 21760 70584 21972 70590
rect 22168 70720 22788 70796
rect 22168 70584 22380 70720
rect 22576 70660 22788 70720
rect 22478 70654 22788 70660
rect 22440 70590 22446 70654
rect 22510 70590 22788 70654
rect 22478 70584 22788 70590
rect 22984 70790 23196 70796
rect 22984 70726 22990 70790
rect 23054 70726 23196 70790
rect 22984 70654 23196 70726
rect 22984 70590 22990 70654
rect 23054 70590 23196 70654
rect 22984 70584 23196 70590
rect 23392 70790 23604 70796
rect 23392 70726 23398 70790
rect 23462 70726 23604 70790
rect 23392 70654 23604 70726
rect 23392 70590 23534 70654
rect 23598 70590 23604 70654
rect 23392 70584 23604 70590
rect 28288 70790 28636 70998
rect 28288 70726 28294 70790
rect 28358 70726 28566 70790
rect 28630 70726 28636 70790
rect 28288 70584 28636 70726
rect 28560 70524 28636 70584
rect 28288 70518 28636 70524
rect 28288 70454 28566 70518
rect 28630 70454 28636 70518
rect 21760 70382 21972 70388
rect 21760 70318 21766 70382
rect 21830 70318 21972 70382
rect 21760 70246 21972 70318
rect 21760 70182 21902 70246
rect 21966 70182 21972 70246
rect 21760 70176 21972 70182
rect 22168 70382 22516 70388
rect 22168 70318 22446 70382
rect 22510 70318 22516 70382
rect 22168 70312 22516 70318
rect 22168 70246 22380 70312
rect 22168 70182 22310 70246
rect 22374 70182 22380 70246
rect 22168 70176 22380 70182
rect 22576 70246 22788 70388
rect 22576 70182 22582 70246
rect 22646 70182 22788 70246
rect 22576 70176 22788 70182
rect 22984 70382 23196 70388
rect 22984 70318 22990 70382
rect 23054 70318 23196 70382
rect 22984 70246 23196 70318
rect 22984 70182 22990 70246
rect 23054 70182 23196 70246
rect 22984 70176 23196 70182
rect 23392 70382 23604 70388
rect 23392 70318 23534 70382
rect 23598 70318 23604 70382
rect 23392 70246 23604 70318
rect 23392 70182 23534 70246
rect 23598 70182 23604 70246
rect 23392 70176 23604 70182
rect 28288 70312 28636 70454
rect 190128 71062 190340 71068
rect 190128 70998 190270 71062
rect 190334 70998 190340 71062
rect 190128 70790 190340 70998
rect 195024 71062 195236 71204
rect 195024 70998 195030 71062
rect 195094 70998 195236 71062
rect 195024 70992 195236 70998
rect 195432 71062 195644 71204
rect 195432 70998 195574 71062
rect 195638 70998 195644 71062
rect 195432 70992 195644 70998
rect 195840 71264 196052 71612
rect 196248 71606 196460 71612
rect 196248 71542 196390 71606
rect 196454 71542 196460 71606
rect 196248 71340 196460 71542
rect 196656 71606 196868 71612
rect 196656 71542 196798 71606
rect 196862 71542 196868 71606
rect 196656 71470 196868 71542
rect 196656 71406 196662 71470
rect 196726 71406 196868 71470
rect 196656 71400 196868 71406
rect 196112 71264 196460 71340
rect 195840 71204 195916 71264
rect 196112 71204 196188 71264
rect 196384 71204 196460 71264
rect 195840 71128 196188 71204
rect 195840 70992 196052 71128
rect 196248 71062 196460 71204
rect 196248 70998 196390 71062
rect 196454 70998 196460 71062
rect 196248 70992 196460 70998
rect 196656 71198 196868 71204
rect 196656 71134 196662 71198
rect 196726 71134 196868 71198
rect 196656 71062 196868 71134
rect 196656 70998 196798 71062
rect 196862 70998 196868 71062
rect 196656 70992 196868 70998
rect 216784 71198 217540 71204
rect 216784 71134 217470 71198
rect 217534 71134 217540 71198
rect 216784 71128 217540 71134
rect 216784 71092 216996 71128
rect 216784 71036 216908 71092
rect 216964 71036 216996 71092
rect 216784 70992 216996 71036
rect 190128 70726 190134 70790
rect 190198 70726 190340 70790
rect 190128 70584 190340 70726
rect 195024 70790 195236 70796
rect 195024 70726 195030 70790
rect 195094 70726 195236 70790
rect 195024 70654 195236 70726
rect 195024 70590 195166 70654
rect 195230 70590 195236 70654
rect 195024 70584 195236 70590
rect 195432 70790 195644 70796
rect 195432 70726 195574 70790
rect 195638 70726 195644 70790
rect 195432 70654 195644 70726
rect 195432 70590 195438 70654
rect 195502 70590 195644 70654
rect 195432 70584 195644 70590
rect 195840 70660 196052 70796
rect 196248 70790 196460 70796
rect 196248 70726 196390 70790
rect 196454 70726 196460 70790
rect 195840 70654 196188 70660
rect 195840 70590 196118 70654
rect 196182 70590 196188 70654
rect 195840 70584 196188 70590
rect 196248 70654 196460 70726
rect 196248 70590 196254 70654
rect 196318 70590 196460 70654
rect 196248 70584 196460 70590
rect 196656 70790 196868 70796
rect 196656 70726 196798 70790
rect 196862 70726 196868 70790
rect 196656 70654 196868 70726
rect 196656 70590 196662 70654
rect 196726 70590 196868 70654
rect 196656 70584 196868 70590
rect 190128 70524 190204 70584
rect 190128 70518 190340 70524
rect 190128 70454 190134 70518
rect 190198 70454 190340 70518
rect 190128 70312 190340 70454
rect 195024 70382 195236 70388
rect 195024 70318 195166 70382
rect 195230 70318 195236 70382
rect 28288 70252 28364 70312
rect 190128 70252 190204 70312
rect 28288 70040 28636 70252
rect 190128 70040 190340 70252
rect 195024 70246 195236 70318
rect 195024 70182 195030 70246
rect 195094 70182 195236 70246
rect 195024 70176 195236 70182
rect 195432 70382 195644 70388
rect 195432 70318 195438 70382
rect 195502 70318 195644 70382
rect 195432 70246 195644 70318
rect 195432 70182 195438 70246
rect 195502 70182 195644 70246
rect 195432 70176 195644 70182
rect 195840 70246 196052 70388
rect 196150 70382 196460 70388
rect 196112 70318 196118 70382
rect 196182 70318 196254 70382
rect 196318 70318 196460 70382
rect 196150 70312 196460 70318
rect 196248 70252 196460 70312
rect 196150 70246 196460 70252
rect 195840 70182 195982 70246
rect 196046 70182 196052 70246
rect 196112 70182 196118 70246
rect 196182 70182 196460 70246
rect 195840 70176 196052 70182
rect 196150 70176 196460 70182
rect 196656 70382 196868 70388
rect 196656 70318 196662 70382
rect 196726 70318 196868 70382
rect 196656 70246 196868 70318
rect 196656 70182 196662 70246
rect 196726 70182 196868 70246
rect 196656 70176 196868 70182
rect 28560 69980 28636 70040
rect 190264 69980 190340 70040
rect 21760 69974 21972 69980
rect 21760 69910 21902 69974
rect 21966 69910 21972 69974
rect 21760 69838 21972 69910
rect 21760 69774 21766 69838
rect 21830 69774 21972 69838
rect 21760 69768 21972 69774
rect 22168 69974 22788 69980
rect 22168 69910 22310 69974
rect 22374 69910 22582 69974
rect 22646 69910 22788 69974
rect 22168 69904 22788 69910
rect 22168 69838 22380 69904
rect 22168 69774 22310 69838
rect 22374 69774 22380 69838
rect 22168 69768 22380 69774
rect 22576 69838 22788 69904
rect 22576 69774 22582 69838
rect 22646 69774 22788 69838
rect 22576 69768 22788 69774
rect 22984 69974 23196 69980
rect 22984 69910 22990 69974
rect 23054 69910 23196 69974
rect 22984 69838 23196 69910
rect 22984 69774 22990 69838
rect 23054 69774 23196 69838
rect 22984 69768 23196 69774
rect 23392 69974 23604 69980
rect 23392 69910 23534 69974
rect 23598 69910 23604 69974
rect 23392 69838 23604 69910
rect 23392 69774 23534 69838
rect 23598 69774 23604 69838
rect 23392 69768 23604 69774
rect 28288 69768 28636 69980
rect 190128 69768 190340 69980
rect 195024 69974 195236 69980
rect 195024 69910 195030 69974
rect 195094 69910 195236 69974
rect 195024 69838 195236 69910
rect 195024 69774 195030 69838
rect 195094 69774 195236 69838
rect 195024 69768 195236 69774
rect 195432 69974 195644 69980
rect 195432 69910 195438 69974
rect 195502 69910 195644 69974
rect 195432 69838 195644 69910
rect 195432 69774 195438 69838
rect 195502 69774 195644 69838
rect 195432 69768 195644 69774
rect 195840 69974 196188 69980
rect 195840 69910 195982 69974
rect 196046 69910 196118 69974
rect 196182 69910 196188 69974
rect 195840 69904 196188 69910
rect 195840 69844 196052 69904
rect 196248 69844 196460 69980
rect 195840 69838 196460 69844
rect 195840 69774 196254 69838
rect 196318 69774 196460 69838
rect 195840 69768 196460 69774
rect 196656 69974 196868 69980
rect 196656 69910 196662 69974
rect 196726 69910 196868 69974
rect 196656 69838 196868 69910
rect 196656 69774 196798 69838
rect 196862 69774 196868 69838
rect 196656 69768 196868 69774
rect 28424 69708 28500 69768
rect 190264 69708 190340 69768
rect 21760 69566 21972 69572
rect 21760 69502 21766 69566
rect 21830 69502 21972 69566
rect 1224 69430 1844 69436
rect 1224 69366 1230 69430
rect 1294 69412 1844 69430
rect 1294 69366 1702 69412
rect 1224 69360 1702 69366
rect 1632 69356 1702 69360
rect 1758 69356 1844 69412
rect 1632 69224 1844 69356
rect 21760 69360 21972 69502
rect 22168 69566 22380 69572
rect 22168 69502 22310 69566
rect 22374 69502 22380 69566
rect 22168 69360 22380 69502
rect 22576 69566 22788 69572
rect 22576 69502 22582 69566
rect 22646 69502 22788 69566
rect 22576 69430 22788 69502
rect 22576 69366 22582 69430
rect 22646 69366 22788 69430
rect 22576 69360 22788 69366
rect 22984 69566 23196 69572
rect 22984 69502 22990 69566
rect 23054 69502 23196 69566
rect 22984 69430 23196 69502
rect 22984 69366 22990 69430
rect 23054 69366 23196 69430
rect 22984 69360 23196 69366
rect 23392 69566 23604 69572
rect 23392 69502 23534 69566
rect 23598 69502 23604 69566
rect 23392 69430 23604 69502
rect 28288 69496 28636 69708
rect 190128 69496 190340 69708
rect 195024 69566 195236 69572
rect 195024 69502 195030 69566
rect 195094 69502 195236 69566
rect 28424 69436 28500 69496
rect 190128 69436 190204 69496
rect 23392 69366 23534 69430
rect 23598 69366 23604 69430
rect 23392 69360 23604 69366
rect 21760 69300 21836 69360
rect 21760 69022 21972 69300
rect 28288 69224 28636 69436
rect 190128 69224 190340 69436
rect 195024 69430 195236 69502
rect 195024 69366 195166 69430
rect 195230 69366 195236 69430
rect 195024 69360 195236 69366
rect 195432 69566 195644 69572
rect 195432 69502 195438 69566
rect 195502 69502 195644 69566
rect 195432 69430 195644 69502
rect 195432 69366 195574 69430
rect 195638 69366 195644 69430
rect 195432 69360 195644 69366
rect 195840 69430 196052 69572
rect 196248 69566 196460 69572
rect 196248 69502 196254 69566
rect 196318 69502 196460 69566
rect 196248 69436 196460 69502
rect 196150 69430 196460 69436
rect 195840 69366 195846 69430
rect 195910 69366 196052 69430
rect 196112 69366 196118 69430
rect 196182 69366 196460 69430
rect 195840 69360 196052 69366
rect 196150 69360 196460 69366
rect 196656 69566 196868 69572
rect 196656 69502 196798 69566
rect 196862 69502 196868 69566
rect 196656 69360 196868 69502
rect 216784 69412 216996 69436
rect 196656 69300 196732 69360
rect 216784 69356 216908 69412
rect 216964 69356 216996 69412
rect 216784 69300 216996 69356
rect 28424 69164 28500 69224
rect 190128 69164 190204 69224
rect 21760 68958 21902 69022
rect 21966 68958 21972 69022
rect 21760 68952 21972 68958
rect 22168 69028 22380 69164
rect 22576 69158 22788 69164
rect 22576 69094 22582 69158
rect 22646 69094 22788 69158
rect 22576 69028 22788 69094
rect 22168 69022 22788 69028
rect 22168 68958 22718 69022
rect 22782 68958 22788 69022
rect 22168 68952 22788 68958
rect 22984 69158 23196 69164
rect 22984 69094 22990 69158
rect 23054 69094 23196 69158
rect 22984 69022 23196 69094
rect 22984 68958 23126 69022
rect 23190 68958 23196 69022
rect 22984 68952 23196 68958
rect 23392 69158 23604 69164
rect 23392 69094 23534 69158
rect 23598 69094 23604 69158
rect 23392 69022 23604 69094
rect 23392 68958 23398 69022
rect 23462 68958 23604 69022
rect 23392 68952 23604 68958
rect 28288 68952 28636 69164
rect 190128 68952 190340 69164
rect 195024 69158 195236 69164
rect 195024 69094 195166 69158
rect 195230 69094 195236 69158
rect 195024 69022 195236 69094
rect 195024 68958 195030 69022
rect 195094 68958 195236 69022
rect 195024 68952 195236 68958
rect 195432 69158 195644 69164
rect 195432 69094 195574 69158
rect 195638 69094 195644 69158
rect 195432 69022 195644 69094
rect 195432 68958 195438 69022
rect 195502 68958 195644 69022
rect 195432 68952 195644 68958
rect 195840 69158 196188 69164
rect 195840 69094 195846 69158
rect 195910 69094 196118 69158
rect 196182 69094 196188 69158
rect 195840 69088 196188 69094
rect 195840 69028 196052 69088
rect 196248 69028 196460 69164
rect 195840 68952 196460 69028
rect 196656 69022 196868 69300
rect 216784 69294 217540 69300
rect 216784 69230 217470 69294
rect 217534 69230 217540 69294
rect 216784 69224 217540 69230
rect 196656 68958 196798 69022
rect 196862 68958 196868 69022
rect 196656 68952 196868 68958
rect 28560 68892 28636 68952
rect 190264 68892 190340 68952
rect 196248 68892 196324 68952
rect 21760 68750 21972 68756
rect 21760 68686 21902 68750
rect 21966 68686 21972 68750
rect 21760 68544 21972 68686
rect 22168 68620 22380 68756
rect 22576 68750 22788 68756
rect 22576 68686 22718 68750
rect 22782 68686 22788 68750
rect 22576 68620 22788 68686
rect 22168 68614 22788 68620
rect 22168 68550 22310 68614
rect 22374 68550 22788 68614
rect 22168 68544 22788 68550
rect 22984 68750 23196 68756
rect 22984 68686 23126 68750
rect 23190 68686 23196 68750
rect 22984 68614 23196 68686
rect 22984 68550 22990 68614
rect 23054 68550 23196 68614
rect 22984 68544 23196 68550
rect 23392 68750 23604 68756
rect 23392 68686 23398 68750
rect 23462 68686 23604 68750
rect 23392 68614 23604 68686
rect 28288 68680 28636 68892
rect 190128 68680 190340 68892
rect 196112 68816 196324 68892
rect 196112 68756 196188 68816
rect 28424 68620 28500 68680
rect 190264 68620 190340 68680
rect 23392 68550 23534 68614
rect 23598 68550 23604 68614
rect 23392 68544 23604 68550
rect 21896 68484 21972 68544
rect 21760 68342 21972 68484
rect 22304 68484 22380 68544
rect 22304 68408 22652 68484
rect 28288 68408 28636 68620
rect 190128 68478 190340 68620
rect 195024 68750 195236 68756
rect 195024 68686 195030 68750
rect 195094 68686 195236 68750
rect 195024 68614 195236 68686
rect 195024 68550 195030 68614
rect 195094 68550 195236 68614
rect 195024 68544 195236 68550
rect 195432 68750 195644 68756
rect 195432 68686 195438 68750
rect 195502 68686 195644 68750
rect 195432 68614 195644 68686
rect 195432 68550 195574 68614
rect 195638 68550 195644 68614
rect 195432 68544 195644 68550
rect 195840 68680 196188 68756
rect 195840 68620 196052 68680
rect 196248 68620 196460 68756
rect 195840 68614 196460 68620
rect 195840 68550 195846 68614
rect 195910 68550 196460 68614
rect 195840 68544 196460 68550
rect 196656 68750 196868 68756
rect 196656 68686 196798 68750
rect 196862 68686 196868 68750
rect 196656 68544 196868 68686
rect 196792 68484 196868 68544
rect 190128 68414 190134 68478
rect 190198 68414 190340 68478
rect 190128 68408 190340 68414
rect 22576 68348 22652 68408
rect 28424 68348 28500 68408
rect 190128 68348 190204 68408
rect 21760 68278 21766 68342
rect 21830 68278 21972 68342
rect 21760 68272 21972 68278
rect 22168 68342 22380 68348
rect 22168 68278 22310 68342
rect 22374 68278 22380 68342
rect 22168 68136 22380 68278
rect 22576 68136 22788 68348
rect 22984 68342 23196 68348
rect 22984 68278 22990 68342
rect 23054 68278 23196 68342
rect 22984 68136 23196 68278
rect 23392 68342 23604 68348
rect 23392 68278 23534 68342
rect 23598 68278 23604 68342
rect 23392 68136 23604 68278
rect 22168 68076 22244 68136
rect 22576 68076 22652 68136
rect 23120 68076 23196 68136
rect 23528 68076 23604 68136
rect 21760 68070 21972 68076
rect 21760 68006 21766 68070
rect 21830 68006 21972 68070
rect 21760 67934 21972 68006
rect 21760 67870 21902 67934
rect 21966 67870 21972 67934
rect 21760 67864 21972 67870
rect 22168 67864 22380 68076
rect 22576 67940 22788 68076
rect 22478 67934 22788 67940
rect 22440 67870 22446 67934
rect 22510 67870 22788 67934
rect 22478 67864 22788 67870
rect 1224 67798 1844 67804
rect 1224 67734 1230 67798
rect 1294 67734 1844 67798
rect 1224 67732 1844 67734
rect 1224 67728 1702 67732
rect 1632 67676 1702 67728
rect 1758 67676 1844 67732
rect 1632 67592 1844 67676
rect 22984 67728 23196 68076
rect 23392 67728 23604 68076
rect 28288 68070 28636 68348
rect 28288 68006 28430 68070
rect 28494 68006 28636 68070
rect 28288 68000 28636 68006
rect 190128 68206 190340 68348
rect 190128 68142 190134 68206
rect 190198 68142 190340 68206
rect 190128 68070 190340 68142
rect 195024 68342 195236 68348
rect 195024 68278 195030 68342
rect 195094 68278 195236 68342
rect 195024 68136 195236 68278
rect 195160 68076 195236 68136
rect 190128 68006 190134 68070
rect 190198 68006 190340 68070
rect 190128 68000 190340 68006
rect 28288 67798 28636 67804
rect 28288 67734 28430 67798
rect 28494 67734 28636 67798
rect 22984 67668 23060 67728
rect 23392 67668 23468 67728
rect 21760 67662 21972 67668
rect 21760 67598 21902 67662
rect 21966 67598 21972 67662
rect 21760 67526 21972 67598
rect 21760 67462 21902 67526
rect 21966 67462 21972 67526
rect 21760 67456 21972 67462
rect 22168 67662 22516 67668
rect 22168 67598 22446 67662
rect 22510 67598 22516 67662
rect 22168 67592 22516 67598
rect 22576 67592 22788 67668
rect 22168 67396 22380 67592
rect 22688 67396 22788 67592
rect 22168 67320 22516 67396
rect 22168 67260 22244 67320
rect 22440 67260 22516 67320
rect 22576 67320 22788 67396
rect 22984 67320 23196 67668
rect 23392 67320 23604 67668
rect 22576 67260 22652 67320
rect 22984 67260 23060 67320
rect 23528 67260 23604 67320
rect 21760 67254 21972 67260
rect 21760 67190 21902 67254
rect 21966 67190 21972 67254
rect 21760 67118 21972 67190
rect 21760 67054 21902 67118
rect 21966 67054 21972 67118
rect 21760 67048 21972 67054
rect 22168 67048 22380 67260
rect 22440 67184 22788 67260
rect 22576 67118 22788 67184
rect 22576 67054 22582 67118
rect 22646 67054 22788 67118
rect 22576 67048 22788 67054
rect 22984 67118 23196 67260
rect 22984 67054 23126 67118
rect 23190 67054 23196 67118
rect 22984 67048 23196 67054
rect 23392 67118 23604 67260
rect 23392 67054 23398 67118
rect 23462 67054 23604 67118
rect 23392 67048 23604 67054
rect 28288 67662 28636 67734
rect 28288 67598 28294 67662
rect 28358 67598 28636 67662
rect 28288 67390 28636 67598
rect 28288 67326 28294 67390
rect 28358 67326 28636 67390
rect 28288 67184 28636 67326
rect 190128 67798 190340 67804
rect 190128 67734 190134 67798
rect 190198 67734 190340 67798
rect 190128 67184 190340 67734
rect 195024 67728 195236 68076
rect 195432 68342 195644 68348
rect 195432 68278 195574 68342
rect 195638 68278 195644 68342
rect 195432 68136 195644 68278
rect 195840 68342 196052 68348
rect 195840 68278 195846 68342
rect 195910 68278 196052 68342
rect 195840 68136 196052 68278
rect 196248 68136 196460 68348
rect 196656 68342 196868 68484
rect 196656 68278 196662 68342
rect 196726 68278 196868 68342
rect 196656 68272 196868 68278
rect 195432 68076 195508 68136
rect 195840 68076 195916 68136
rect 196248 68076 196324 68136
rect 195432 67728 195644 68076
rect 195840 67940 196052 68076
rect 196248 67940 196460 68076
rect 195840 67864 196460 67940
rect 196656 68070 196868 68076
rect 196656 68006 196662 68070
rect 196726 68006 196868 68070
rect 196656 67934 196868 68006
rect 196656 67870 196798 67934
rect 196862 67870 196868 67934
rect 196656 67864 196868 67870
rect 195976 67804 196052 67864
rect 195976 67728 196324 67804
rect 195024 67668 195100 67728
rect 195568 67668 195644 67728
rect 196248 67668 196324 67728
rect 216784 67732 216996 67804
rect 216784 67676 216908 67732
rect 216964 67676 216996 67732
rect 216784 67668 216996 67676
rect 195024 67320 195236 67668
rect 195432 67320 195644 67668
rect 195840 67320 196052 67668
rect 196248 67396 196460 67668
rect 196656 67662 196868 67668
rect 196656 67598 196798 67662
rect 196862 67598 196868 67662
rect 196656 67526 196868 67598
rect 216784 67662 217540 67668
rect 216784 67598 217470 67662
rect 217534 67598 217540 67662
rect 216784 67592 217540 67598
rect 196656 67462 196662 67526
rect 196726 67462 196868 67526
rect 196656 67456 196868 67462
rect 196112 67320 196460 67396
rect 195024 67260 195100 67320
rect 195432 67260 195508 67320
rect 195840 67260 195916 67320
rect 196112 67260 196188 67320
rect 28288 67124 28364 67184
rect 190128 67124 190204 67184
rect 21760 66846 21972 66852
rect 21760 66782 21902 66846
rect 21966 66782 21972 66846
rect 21760 66710 21972 66782
rect 21760 66646 21902 66710
rect 21966 66646 21972 66710
rect 21760 66640 21972 66646
rect 22168 66716 22380 66852
rect 22576 66846 22788 66852
rect 22576 66782 22582 66846
rect 22646 66782 22788 66846
rect 22576 66716 22788 66782
rect 22168 66710 22788 66716
rect 22168 66646 22310 66710
rect 22374 66646 22718 66710
rect 22782 66646 22788 66710
rect 22168 66640 22788 66646
rect 22984 66846 23196 66852
rect 22984 66782 23126 66846
rect 23190 66782 23196 66846
rect 22984 66710 23196 66782
rect 22984 66646 22990 66710
rect 23054 66646 23196 66710
rect 22984 66640 23196 66646
rect 23392 66846 23604 66852
rect 23392 66782 23398 66846
rect 23462 66782 23604 66846
rect 23392 66710 23604 66782
rect 23392 66646 23398 66710
rect 23462 66646 23604 66710
rect 23392 66640 23604 66646
rect 28288 66846 28636 67124
rect 28288 66782 28294 66846
rect 28358 66782 28636 66846
rect 28288 66640 28636 66782
rect 190128 66846 190340 67124
rect 195024 67118 195236 67260
rect 195024 67054 195030 67118
rect 195094 67054 195236 67118
rect 195024 67048 195236 67054
rect 195432 67118 195644 67260
rect 195432 67054 195438 67118
rect 195502 67054 195644 67118
rect 195432 67048 195644 67054
rect 195840 67184 196188 67260
rect 196248 67260 196324 67320
rect 195840 67048 196052 67184
rect 196248 67048 196460 67260
rect 196656 67254 196868 67260
rect 196656 67190 196662 67254
rect 196726 67190 196868 67254
rect 196656 67118 196868 67190
rect 196656 67054 196798 67118
rect 196862 67054 196868 67118
rect 196656 67048 196868 67054
rect 196248 66988 196324 67048
rect 195976 66912 196324 66988
rect 195976 66852 196052 66912
rect 190128 66782 190270 66846
rect 190334 66782 190340 66846
rect 190128 66640 190340 66782
rect 195024 66846 195236 66852
rect 195024 66782 195030 66846
rect 195094 66782 195236 66846
rect 195024 66710 195236 66782
rect 195024 66646 195030 66710
rect 195094 66646 195236 66710
rect 195024 66640 195236 66646
rect 195432 66846 195644 66852
rect 195432 66782 195438 66846
rect 195502 66782 195644 66846
rect 195432 66710 195644 66782
rect 195432 66646 195438 66710
rect 195502 66646 195644 66710
rect 195432 66640 195644 66646
rect 195840 66776 196460 66852
rect 195840 66640 196052 66776
rect 196248 66710 196460 66776
rect 196248 66646 196390 66710
rect 196454 66646 196460 66710
rect 196248 66640 196460 66646
rect 196656 66846 196868 66852
rect 196656 66782 196798 66846
rect 196862 66782 196868 66846
rect 196656 66710 196868 66782
rect 196656 66646 196798 66710
rect 196862 66646 196868 66710
rect 196656 66640 196868 66646
rect 28288 66580 28364 66640
rect 190264 66580 190340 66640
rect 28288 66574 28636 66580
rect 28288 66510 28294 66574
rect 28358 66510 28636 66574
rect 21760 66438 21972 66444
rect 21760 66374 21902 66438
rect 21966 66374 21972 66438
rect 21760 66302 21972 66374
rect 21760 66238 21766 66302
rect 21830 66238 21972 66302
rect 21760 66232 21972 66238
rect 22168 66438 22380 66444
rect 22168 66374 22310 66438
rect 22374 66374 22380 66438
rect 22168 66308 22380 66374
rect 22576 66438 22788 66444
rect 22576 66374 22718 66438
rect 22782 66374 22788 66438
rect 22168 66302 22516 66308
rect 22168 66238 22174 66302
rect 22238 66238 22446 66302
rect 22510 66238 22516 66302
rect 22168 66232 22516 66238
rect 22576 66232 22788 66374
rect 22984 66438 23196 66444
rect 22984 66374 22990 66438
rect 23054 66374 23196 66438
rect 22984 66302 23196 66374
rect 22984 66238 23126 66302
rect 23190 66238 23196 66302
rect 22984 66232 23196 66238
rect 23392 66438 23604 66444
rect 23392 66374 23398 66438
rect 23462 66374 23604 66438
rect 23392 66302 23604 66374
rect 28288 66368 28636 66510
rect 190128 66574 190340 66580
rect 190128 66510 190270 66574
rect 190334 66510 190340 66574
rect 190128 66368 190340 66510
rect 28560 66308 28636 66368
rect 190264 66308 190340 66368
rect 23392 66238 23534 66302
rect 23598 66238 23604 66302
rect 23392 66232 23604 66238
rect 1224 66166 1844 66172
rect 1224 66102 1230 66166
rect 1294 66102 1844 66166
rect 1224 66096 1844 66102
rect 28288 66096 28636 66308
rect 190128 66096 190340 66308
rect 195024 66438 195236 66444
rect 195024 66374 195030 66438
rect 195094 66374 195236 66438
rect 195024 66302 195236 66374
rect 195024 66238 195166 66302
rect 195230 66238 195236 66302
rect 195024 66232 195236 66238
rect 195432 66438 195644 66444
rect 195432 66374 195438 66438
rect 195502 66374 195644 66438
rect 195432 66302 195644 66374
rect 195432 66238 195438 66302
rect 195502 66238 195644 66302
rect 195432 66232 195644 66238
rect 195840 66302 196052 66444
rect 195840 66238 195846 66302
rect 195910 66238 196052 66302
rect 195840 66232 196052 66238
rect 196248 66438 196460 66444
rect 196248 66374 196390 66438
rect 196454 66374 196460 66438
rect 196248 66302 196460 66374
rect 196248 66238 196254 66302
rect 196318 66238 196460 66302
rect 196248 66232 196460 66238
rect 196656 66438 196868 66444
rect 196656 66374 196798 66438
rect 196862 66374 196868 66438
rect 196656 66302 196868 66374
rect 196656 66238 196662 66302
rect 196726 66238 196868 66302
rect 196656 66232 196868 66238
rect 1632 66052 1844 66096
rect 1632 65996 1702 66052
rect 1758 65996 1844 66052
rect 28424 66036 28500 66096
rect 190128 66036 190204 66096
rect 216784 66052 216996 66172
rect 1632 65960 1844 65996
rect 21760 66030 21972 66036
rect 21760 65966 21766 66030
rect 21830 65966 21972 66030
rect 21760 65894 21972 65966
rect 21760 65830 21766 65894
rect 21830 65830 21972 65894
rect 21760 65824 21972 65830
rect 22168 66030 22380 66036
rect 22478 66030 22788 66036
rect 22168 65966 22174 66030
rect 22238 65966 22380 66030
rect 22440 65966 22446 66030
rect 22510 65966 22788 66030
rect 22168 65824 22380 65966
rect 22478 65960 22788 65966
rect 22576 65894 22788 65960
rect 22576 65830 22582 65894
rect 22646 65830 22788 65894
rect 22576 65824 22788 65830
rect 22984 66030 23196 66036
rect 22984 65966 23126 66030
rect 23190 65966 23196 66030
rect 22984 65894 23196 65966
rect 22984 65830 23126 65894
rect 23190 65830 23196 65894
rect 22984 65824 23196 65830
rect 23392 66030 23604 66036
rect 23392 65966 23534 66030
rect 23598 65966 23604 66030
rect 23392 65894 23604 65966
rect 23392 65830 23398 65894
rect 23462 65830 23604 65894
rect 23392 65824 23604 65830
rect 28288 65824 28636 66036
rect 28560 65764 28636 65824
rect 21760 65622 21972 65628
rect 21760 65558 21766 65622
rect 21830 65558 21972 65622
rect 21760 65416 21972 65558
rect 22168 65622 22788 65628
rect 22168 65558 22582 65622
rect 22646 65558 22788 65622
rect 22168 65552 22788 65558
rect 22168 65492 22380 65552
rect 22168 65486 22516 65492
rect 22168 65422 22174 65486
rect 22238 65422 22446 65486
rect 22510 65422 22516 65486
rect 22168 65416 22516 65422
rect 22576 65416 22788 65552
rect 22984 65622 23196 65628
rect 22984 65558 23126 65622
rect 23190 65558 23196 65622
rect 22984 65486 23196 65558
rect 22984 65422 22990 65486
rect 23054 65422 23196 65486
rect 22984 65416 23196 65422
rect 23392 65622 23604 65628
rect 23392 65558 23398 65622
rect 23462 65558 23604 65622
rect 23392 65486 23604 65558
rect 28288 65552 28636 65764
rect 190128 65824 190340 66036
rect 195024 66030 195236 66036
rect 195024 65966 195166 66030
rect 195230 65966 195236 66030
rect 195024 65894 195236 65966
rect 195024 65830 195166 65894
rect 195230 65830 195236 65894
rect 195024 65824 195236 65830
rect 195432 66030 195644 66036
rect 195432 65966 195438 66030
rect 195502 65966 195644 66030
rect 195432 65894 195644 65966
rect 195432 65830 195574 65894
rect 195638 65830 195644 65894
rect 195432 65824 195644 65830
rect 195840 66030 196052 66036
rect 195840 65966 195846 66030
rect 195910 65966 196052 66030
rect 195840 65894 196052 65966
rect 196248 66030 196460 66036
rect 196248 65966 196254 66030
rect 196318 65966 196460 66030
rect 196248 65900 196460 65966
rect 196150 65894 196460 65900
rect 195840 65830 195982 65894
rect 196046 65830 196052 65894
rect 196112 65830 196118 65894
rect 196182 65830 196460 65894
rect 195840 65824 196052 65830
rect 196150 65824 196460 65830
rect 196656 66030 196868 66036
rect 196656 65966 196662 66030
rect 196726 65966 196868 66030
rect 196656 65894 196868 65966
rect 216784 65996 216908 66052
rect 216964 66036 216996 66052
rect 216964 66030 217540 66036
rect 216964 65996 217470 66030
rect 216784 65966 217470 65996
rect 217534 65966 217540 66030
rect 216784 65960 217540 65966
rect 196656 65830 196662 65894
rect 196726 65830 196868 65894
rect 196656 65824 196868 65830
rect 190128 65764 190204 65824
rect 190128 65552 190340 65764
rect 28560 65492 28636 65552
rect 190264 65492 190340 65552
rect 23392 65422 23398 65486
rect 23462 65422 23604 65486
rect 23392 65416 23604 65422
rect 21760 65356 21836 65416
rect 21760 65078 21972 65356
rect 28288 65280 28636 65492
rect 190128 65280 190340 65492
rect 195024 65622 195236 65628
rect 195024 65558 195166 65622
rect 195230 65558 195236 65622
rect 195024 65486 195236 65558
rect 195024 65422 195030 65486
rect 195094 65422 195236 65486
rect 195024 65416 195236 65422
rect 195432 65622 195644 65628
rect 195432 65558 195574 65622
rect 195638 65558 195644 65622
rect 195432 65486 195644 65558
rect 195432 65422 195438 65486
rect 195502 65422 195644 65486
rect 195432 65416 195644 65422
rect 195840 65622 196188 65628
rect 195840 65558 195982 65622
rect 196046 65558 196118 65622
rect 196182 65558 196188 65622
rect 195840 65552 196188 65558
rect 195840 65492 196052 65552
rect 196248 65492 196460 65628
rect 195840 65486 196460 65492
rect 195840 65422 196254 65486
rect 196318 65422 196460 65486
rect 195840 65416 196460 65422
rect 196656 65622 196868 65628
rect 196656 65558 196662 65622
rect 196726 65558 196868 65622
rect 196656 65416 196868 65558
rect 196792 65356 196868 65416
rect 28424 65220 28500 65280
rect 190264 65220 190340 65280
rect 21760 65014 21766 65078
rect 21830 65014 21972 65078
rect 21760 65008 21972 65014
rect 22168 65214 22380 65220
rect 22478 65214 22788 65220
rect 22168 65150 22174 65214
rect 22238 65150 22380 65214
rect 22440 65150 22446 65214
rect 22510 65150 22788 65214
rect 22168 65008 22380 65150
rect 22478 65144 22788 65150
rect 22576 65078 22788 65144
rect 22576 65014 22582 65078
rect 22646 65014 22788 65078
rect 22576 65008 22788 65014
rect 22984 65214 23196 65220
rect 22984 65150 22990 65214
rect 23054 65150 23196 65214
rect 22984 65078 23196 65150
rect 22984 65014 23126 65078
rect 23190 65014 23196 65078
rect 22984 65008 23196 65014
rect 23392 65214 23604 65220
rect 23392 65150 23398 65214
rect 23462 65150 23604 65214
rect 23392 65078 23604 65150
rect 23392 65014 23534 65078
rect 23598 65014 23604 65078
rect 23392 65008 23604 65014
rect 28288 65008 28636 65220
rect 190128 65008 190340 65220
rect 195024 65214 195236 65220
rect 195024 65150 195030 65214
rect 195094 65150 195236 65214
rect 195024 65078 195236 65150
rect 195024 65014 195166 65078
rect 195230 65014 195236 65078
rect 195024 65008 195236 65014
rect 195432 65214 195644 65220
rect 195432 65150 195438 65214
rect 195502 65150 195644 65214
rect 195432 65078 195644 65150
rect 195432 65014 195574 65078
rect 195638 65014 195644 65078
rect 195432 65008 195644 65014
rect 195840 65078 196052 65220
rect 196248 65214 196460 65220
rect 196248 65150 196254 65214
rect 196318 65150 196460 65214
rect 196248 65084 196460 65150
rect 196150 65078 196460 65084
rect 195840 65014 195846 65078
rect 195910 65014 196052 65078
rect 196112 65014 196118 65078
rect 196182 65014 196460 65078
rect 195840 65008 196052 65014
rect 196150 65008 196460 65014
rect 196656 65078 196868 65356
rect 196656 65014 196662 65078
rect 196726 65014 196868 65078
rect 196656 65008 196868 65014
rect 28288 64948 28364 65008
rect 190128 64948 190204 65008
rect 21760 64806 21972 64812
rect 21760 64742 21766 64806
rect 21830 64742 21972 64806
rect 21760 64600 21972 64742
rect 22168 64676 22380 64812
rect 22576 64806 22788 64812
rect 22576 64742 22582 64806
rect 22646 64742 22788 64806
rect 22168 64670 22516 64676
rect 22168 64606 22446 64670
rect 22510 64606 22516 64670
rect 22168 64600 22516 64606
rect 22576 64670 22788 64742
rect 22576 64606 22718 64670
rect 22782 64606 22788 64670
rect 22576 64600 22788 64606
rect 22984 64806 23196 64812
rect 22984 64742 23126 64806
rect 23190 64742 23196 64806
rect 22984 64670 23196 64742
rect 22984 64606 23126 64670
rect 23190 64606 23196 64670
rect 22984 64600 23196 64606
rect 23392 64806 23604 64812
rect 23392 64742 23534 64806
rect 23598 64742 23604 64806
rect 23392 64670 23604 64742
rect 23392 64606 23398 64670
rect 23462 64606 23604 64670
rect 23392 64600 23604 64606
rect 28288 64736 28636 64948
rect 190128 64736 190340 64948
rect 28288 64676 28364 64736
rect 190264 64676 190340 64736
rect 21896 64540 21972 64600
rect 1632 64372 1844 64404
rect 1632 64316 1702 64372
rect 1758 64316 1844 64372
rect 21760 64398 21972 64540
rect 28288 64534 28636 64676
rect 28288 64470 28566 64534
rect 28630 64470 28636 64534
rect 28288 64464 28636 64470
rect 190128 64464 190340 64676
rect 195024 64806 195236 64812
rect 195024 64742 195166 64806
rect 195230 64742 195236 64806
rect 195024 64670 195236 64742
rect 195024 64606 195030 64670
rect 195094 64606 195236 64670
rect 195024 64600 195236 64606
rect 195432 64806 195644 64812
rect 195432 64742 195574 64806
rect 195638 64742 195644 64806
rect 195432 64670 195644 64742
rect 195432 64606 195574 64670
rect 195638 64606 195644 64670
rect 195432 64600 195644 64606
rect 195840 64806 196188 64812
rect 195840 64742 195846 64806
rect 195910 64742 196118 64806
rect 196182 64742 196188 64806
rect 195840 64736 196188 64742
rect 195840 64670 196052 64736
rect 195840 64606 195982 64670
rect 196046 64606 196052 64670
rect 195840 64600 196052 64606
rect 196248 64600 196460 64812
rect 196656 64806 196868 64812
rect 196656 64742 196662 64806
rect 196726 64742 196868 64806
rect 196656 64600 196868 64742
rect 196248 64540 196324 64600
rect 196792 64540 196868 64600
rect 28424 64404 28500 64464
rect 190264 64404 190340 64464
rect 195976 64464 196324 64540
rect 195976 64404 196052 64464
rect 21760 64334 21902 64398
rect 21966 64334 21972 64398
rect 21760 64328 21972 64334
rect 1632 64268 1844 64316
rect 1224 64262 1844 64268
rect 1224 64198 1230 64262
rect 1294 64198 1844 64262
rect 1224 64192 1844 64198
rect 22168 64268 22380 64404
rect 22478 64398 22788 64404
rect 22440 64334 22446 64398
rect 22510 64334 22718 64398
rect 22782 64334 22788 64398
rect 22478 64328 22788 64334
rect 22576 64268 22788 64328
rect 22168 64192 22788 64268
rect 22984 64398 23196 64404
rect 22984 64334 23126 64398
rect 23190 64334 23196 64398
rect 22984 64262 23196 64334
rect 22984 64198 23126 64262
rect 23190 64198 23196 64262
rect 22984 64192 23196 64198
rect 23392 64398 23604 64404
rect 23392 64334 23398 64398
rect 23462 64334 23604 64398
rect 23392 64262 23604 64334
rect 23392 64198 23398 64262
rect 23462 64198 23604 64262
rect 23392 64192 23604 64198
rect 28288 64262 28636 64404
rect 28288 64198 28566 64262
rect 28630 64198 28636 64262
rect 22304 64132 22380 64192
rect 22712 64132 22788 64192
rect 21760 64126 21972 64132
rect 21760 64062 21902 64126
rect 21966 64062 21972 64126
rect 21760 63784 21972 64062
rect 22168 63784 22380 64132
rect 22576 63854 22788 64132
rect 22576 63790 22718 63854
rect 22782 63790 22788 63854
rect 22576 63784 22788 63790
rect 22984 63990 23196 63996
rect 22984 63926 23126 63990
rect 23190 63926 23196 63990
rect 22984 63784 23196 63926
rect 23392 63990 23604 63996
rect 23392 63926 23398 63990
rect 23462 63926 23604 63990
rect 23392 63784 23604 63926
rect 21896 63724 21972 63784
rect 23120 63724 23196 63784
rect 23528 63724 23604 63784
rect 21760 63582 21972 63724
rect 21760 63518 21902 63582
rect 21966 63518 21972 63582
rect 21760 63512 21972 63518
rect 22168 63452 22380 63588
rect 22576 63582 22788 63588
rect 22576 63518 22718 63582
rect 22782 63518 22788 63582
rect 22168 63376 22516 63452
rect 22576 63376 22788 63518
rect 22984 63376 23196 63724
rect 22304 63316 22380 63376
rect 21760 63310 21972 63316
rect 21760 63246 21902 63310
rect 21966 63246 21972 63310
rect 21760 63174 21972 63246
rect 21760 63110 21902 63174
rect 21966 63110 21972 63174
rect 21760 63104 21972 63110
rect 22168 63180 22380 63316
rect 22440 63316 22516 63376
rect 22712 63316 22788 63376
rect 23120 63316 23196 63376
rect 22440 63240 22788 63316
rect 22168 63174 22516 63180
rect 22168 63110 22310 63174
rect 22374 63110 22446 63174
rect 22510 63110 22516 63174
rect 22168 63104 22516 63110
rect 22576 63104 22788 63240
rect 22984 62968 23196 63316
rect 23392 63376 23604 63724
rect 28288 63920 28636 64198
rect 190128 63920 190340 64404
rect 195024 64398 195236 64404
rect 195024 64334 195030 64398
rect 195094 64334 195236 64398
rect 195024 64262 195236 64334
rect 195024 64198 195166 64262
rect 195230 64198 195236 64262
rect 195024 64192 195236 64198
rect 195432 64398 195644 64404
rect 195432 64334 195574 64398
rect 195638 64334 195644 64398
rect 195432 64262 195644 64334
rect 195432 64198 195574 64262
rect 195638 64198 195644 64262
rect 195432 64192 195644 64198
rect 195840 64398 196460 64404
rect 195840 64334 195982 64398
rect 196046 64334 196460 64398
rect 195840 64328 196460 64334
rect 196656 64398 196868 64540
rect 196656 64334 196798 64398
rect 196862 64334 196868 64398
rect 196656 64328 196868 64334
rect 216784 64398 217540 64404
rect 216784 64372 217470 64398
rect 195840 64192 196052 64328
rect 196248 64192 196460 64328
rect 216784 64316 216908 64372
rect 216964 64334 217470 64372
rect 217534 64334 217540 64398
rect 216964 64328 217540 64334
rect 216964 64316 216996 64328
rect 216784 64192 216996 64316
rect 195840 64132 195916 64192
rect 196384 64132 196460 64192
rect 195024 63990 195236 63996
rect 195024 63926 195166 63990
rect 195230 63926 195236 63990
rect 28288 63860 28364 63920
rect 190128 63860 190204 63920
rect 28288 63718 28636 63860
rect 28288 63654 28430 63718
rect 28494 63654 28636 63718
rect 28288 63446 28636 63654
rect 28288 63382 28294 63446
rect 28358 63382 28430 63446
rect 28494 63382 28636 63446
rect 23392 63316 23468 63376
rect 23392 62968 23604 63316
rect 28288 63240 28636 63382
rect 190128 63718 190340 63860
rect 195024 63784 195236 63926
rect 195432 63990 195644 63996
rect 195432 63926 195574 63990
rect 195638 63926 195644 63990
rect 195432 63784 195644 63926
rect 195840 63854 196052 64132
rect 195840 63790 195982 63854
rect 196046 63790 196052 63854
rect 195840 63784 196052 63790
rect 196248 63784 196460 64132
rect 196656 64126 196868 64132
rect 196656 64062 196798 64126
rect 196862 64062 196868 64126
rect 196656 63784 196868 64062
rect 195160 63724 195236 63784
rect 195568 63724 195644 63784
rect 190128 63654 190134 63718
rect 190198 63654 190340 63718
rect 190128 63446 190340 63654
rect 190128 63382 190134 63446
rect 190198 63382 190340 63446
rect 190128 63310 190340 63382
rect 195024 63376 195236 63724
rect 195160 63316 195236 63376
rect 190128 63246 190134 63310
rect 190198 63246 190340 63310
rect 190128 63240 190340 63246
rect 22984 62908 23060 62968
rect 23528 62908 23604 62968
rect 21760 62902 21972 62908
rect 21760 62838 21902 62902
rect 21966 62838 21972 62902
rect 1632 62692 1844 62772
rect 21760 62766 21972 62838
rect 21760 62702 21766 62766
rect 21830 62702 21972 62766
rect 21760 62696 21972 62702
rect 22168 62902 22380 62908
rect 22478 62902 22788 62908
rect 22168 62838 22310 62902
rect 22374 62838 22380 62902
rect 22440 62838 22446 62902
rect 22510 62838 22788 62902
rect 1632 62636 1702 62692
rect 1758 62636 1844 62692
rect 1224 62630 1844 62636
rect 1224 62566 1230 62630
rect 1294 62566 1844 62630
rect 1224 62560 1844 62566
rect 22168 62560 22380 62838
rect 22478 62832 22788 62838
rect 22576 62560 22788 62832
rect 22984 62766 23196 62908
rect 22984 62702 22990 62766
rect 23054 62702 23196 62766
rect 22984 62696 23196 62702
rect 23392 62766 23604 62908
rect 23392 62702 23398 62766
rect 23462 62702 23604 62766
rect 23392 62696 23604 62702
rect 28288 63038 28636 63044
rect 28288 62974 28294 63038
rect 28358 62974 28636 63038
rect 28288 62696 28636 62974
rect 190128 63038 190340 63044
rect 190128 62974 190134 63038
rect 190198 62974 190340 63038
rect 190128 62902 190340 62974
rect 190128 62838 190134 62902
rect 190198 62838 190340 62902
rect 190128 62696 190340 62838
rect 195024 62968 195236 63316
rect 195432 63376 195644 63724
rect 196656 63724 196732 63784
rect 195840 63582 196052 63588
rect 195840 63518 195982 63582
rect 196046 63518 196052 63582
rect 195840 63376 196052 63518
rect 196248 63376 196460 63588
rect 196656 63582 196868 63724
rect 196656 63518 196798 63582
rect 196862 63518 196868 63582
rect 196656 63512 196868 63518
rect 195432 63316 195508 63376
rect 195976 63316 196052 63376
rect 196384 63316 196460 63376
rect 195432 62968 195644 63316
rect 195840 63240 196460 63316
rect 195840 63180 196052 63240
rect 195840 63174 196188 63180
rect 195840 63110 196118 63174
rect 196182 63110 196188 63174
rect 195840 63104 196188 63110
rect 196248 63104 196460 63240
rect 196656 63310 196868 63316
rect 196656 63246 196798 63310
rect 196862 63246 196868 63310
rect 196656 63174 196868 63246
rect 196656 63110 196662 63174
rect 196726 63110 196868 63174
rect 196656 63104 196868 63110
rect 195024 62908 195100 62968
rect 195432 62908 195508 62968
rect 195024 62766 195236 62908
rect 195024 62702 195030 62766
rect 195094 62702 195236 62766
rect 195024 62696 195236 62702
rect 195432 62766 195644 62908
rect 195432 62702 195438 62766
rect 195502 62702 195644 62766
rect 195432 62696 195644 62702
rect 28424 62636 28500 62696
rect 190128 62636 190204 62696
rect 22304 62500 22380 62560
rect 22712 62500 22788 62560
rect 21760 62494 21972 62500
rect 21760 62430 21766 62494
rect 21830 62430 21972 62494
rect 21760 62358 21972 62430
rect 21760 62294 21902 62358
rect 21966 62294 21972 62358
rect 21760 62288 21972 62294
rect 22168 62288 22380 62500
rect 22576 62358 22788 62500
rect 22576 62294 22718 62358
rect 22782 62294 22788 62358
rect 22576 62288 22788 62294
rect 22984 62494 23196 62500
rect 22984 62430 22990 62494
rect 23054 62430 23196 62494
rect 22984 62358 23196 62430
rect 22984 62294 23126 62358
rect 23190 62294 23196 62358
rect 22984 62288 23196 62294
rect 23392 62494 23604 62500
rect 23392 62430 23398 62494
rect 23462 62430 23604 62494
rect 23392 62358 23604 62430
rect 23392 62294 23398 62358
rect 23462 62294 23604 62358
rect 23392 62288 23604 62294
rect 28288 62424 28636 62636
rect 190128 62630 190340 62636
rect 190128 62566 190134 62630
rect 190198 62566 190340 62630
rect 190128 62424 190340 62566
rect 195840 62560 196052 62908
rect 196150 62902 196460 62908
rect 196112 62838 196118 62902
rect 196182 62838 196460 62902
rect 196150 62832 196460 62838
rect 196248 62636 196460 62832
rect 196656 62902 196868 62908
rect 196656 62838 196662 62902
rect 196726 62838 196868 62902
rect 196656 62766 196868 62838
rect 196656 62702 196798 62766
rect 196862 62702 196868 62766
rect 196656 62696 196868 62702
rect 216784 62766 217540 62772
rect 216784 62702 217470 62766
rect 217534 62702 217540 62766
rect 216784 62696 217540 62702
rect 196112 62560 196460 62636
rect 216784 62692 216996 62696
rect 216784 62636 216908 62692
rect 216964 62636 216996 62692
rect 216784 62560 216996 62636
rect 195840 62500 195916 62560
rect 196112 62500 196188 62560
rect 28288 62364 28364 62424
rect 190264 62364 190340 62424
rect 28288 62152 28636 62364
rect 190128 62152 190340 62364
rect 195024 62494 195236 62500
rect 195024 62430 195030 62494
rect 195094 62430 195236 62494
rect 195024 62358 195236 62430
rect 195024 62294 195030 62358
rect 195094 62294 195236 62358
rect 195024 62288 195236 62294
rect 195432 62494 195644 62500
rect 195432 62430 195438 62494
rect 195502 62430 195644 62494
rect 195432 62358 195644 62430
rect 195432 62294 195438 62358
rect 195502 62294 195644 62358
rect 195432 62288 195644 62294
rect 195840 62424 196188 62500
rect 195840 62364 196052 62424
rect 196248 62364 196460 62500
rect 195840 62358 196460 62364
rect 195840 62294 195982 62358
rect 196046 62294 196460 62358
rect 195840 62288 196460 62294
rect 196656 62494 196868 62500
rect 196656 62430 196798 62494
rect 196862 62430 196868 62494
rect 196656 62358 196868 62430
rect 196656 62294 196798 62358
rect 196862 62294 196868 62358
rect 196656 62288 196868 62294
rect 28288 62092 28364 62152
rect 190264 62092 190340 62152
rect 21760 62086 21972 62092
rect 21760 62022 21902 62086
rect 21966 62022 21972 62086
rect 21760 61950 21972 62022
rect 21760 61886 21766 61950
rect 21830 61886 21972 61950
rect 21760 61880 21972 61886
rect 22168 61950 22380 62092
rect 22168 61886 22174 61950
rect 22238 61886 22380 61950
rect 22168 61880 22380 61886
rect 22576 62086 22788 62092
rect 22576 62022 22718 62086
rect 22782 62022 22788 62086
rect 22576 61950 22788 62022
rect 22576 61886 22582 61950
rect 22646 61886 22788 61950
rect 22576 61880 22788 61886
rect 22984 62086 23196 62092
rect 22984 62022 23126 62086
rect 23190 62022 23196 62086
rect 22984 61950 23196 62022
rect 22984 61886 22990 61950
rect 23054 61886 23196 61950
rect 22984 61880 23196 61886
rect 23392 62086 23604 62092
rect 23392 62022 23398 62086
rect 23462 62022 23604 62086
rect 23392 61950 23604 62022
rect 23392 61886 23534 61950
rect 23598 61886 23604 61950
rect 23392 61880 23604 61886
rect 28288 61880 28636 62092
rect 190128 61880 190340 62092
rect 195024 62086 195236 62092
rect 195024 62022 195030 62086
rect 195094 62022 195236 62086
rect 195024 61950 195236 62022
rect 195024 61886 195166 61950
rect 195230 61886 195236 61950
rect 195024 61880 195236 61886
rect 195432 62086 195644 62092
rect 195432 62022 195438 62086
rect 195502 62022 195644 62086
rect 195432 61950 195644 62022
rect 195432 61886 195574 61950
rect 195638 61886 195644 61950
rect 195432 61880 195644 61886
rect 195840 62086 196052 62092
rect 195840 62022 195982 62086
rect 196046 62022 196052 62086
rect 195840 61956 196052 62022
rect 195840 61950 196188 61956
rect 195840 61886 196118 61950
rect 196182 61886 196188 61950
rect 195840 61880 196188 61886
rect 196248 61950 196460 62092
rect 196248 61886 196254 61950
rect 196318 61886 196460 61950
rect 196248 61880 196460 61886
rect 196656 62086 196868 62092
rect 196656 62022 196798 62086
rect 196862 62022 196868 62086
rect 196656 61950 196868 62022
rect 196656 61886 196662 61950
rect 196726 61886 196868 61950
rect 196656 61880 196868 61886
rect 28288 61820 28364 61880
rect 190128 61820 190204 61880
rect 21760 61678 21972 61684
rect 21760 61614 21766 61678
rect 21830 61614 21972 61678
rect 21760 61542 21972 61614
rect 21760 61478 21902 61542
rect 21966 61478 21972 61542
rect 21760 61472 21972 61478
rect 22168 61678 22380 61684
rect 22168 61614 22174 61678
rect 22238 61614 22380 61678
rect 22168 61548 22380 61614
rect 22576 61678 22788 61684
rect 22576 61614 22582 61678
rect 22646 61614 22788 61678
rect 22576 61548 22788 61614
rect 22168 61472 22788 61548
rect 22984 61678 23196 61684
rect 22984 61614 22990 61678
rect 23054 61614 23196 61678
rect 22984 61542 23196 61614
rect 22984 61478 23126 61542
rect 23190 61478 23196 61542
rect 22984 61472 23196 61478
rect 23392 61678 23604 61684
rect 23392 61614 23534 61678
rect 23598 61614 23604 61678
rect 23392 61542 23604 61614
rect 28288 61608 28636 61820
rect 190128 61608 190340 61820
rect 195024 61678 195236 61684
rect 195024 61614 195166 61678
rect 195230 61614 195236 61678
rect 28424 61548 28500 61608
rect 190128 61548 190204 61608
rect 23392 61478 23534 61542
rect 23598 61478 23604 61542
rect 23392 61472 23604 61478
rect 22576 61412 22652 61472
rect 22304 61336 22652 61412
rect 28288 61336 28636 61548
rect 190128 61336 190340 61548
rect 195024 61542 195236 61614
rect 195024 61478 195166 61542
rect 195230 61478 195236 61542
rect 195024 61472 195236 61478
rect 195432 61678 195644 61684
rect 195432 61614 195574 61678
rect 195638 61614 195644 61678
rect 195432 61542 195644 61614
rect 195432 61478 195574 61542
rect 195638 61478 195644 61542
rect 195432 61472 195644 61478
rect 195840 61542 196052 61684
rect 196150 61678 196460 61684
rect 196112 61614 196118 61678
rect 196182 61614 196254 61678
rect 196318 61614 196460 61678
rect 196150 61608 196460 61614
rect 195840 61478 195982 61542
rect 196046 61478 196052 61542
rect 195840 61472 196052 61478
rect 196248 61472 196460 61608
rect 196656 61678 196868 61684
rect 196656 61614 196662 61678
rect 196726 61614 196868 61678
rect 196656 61542 196868 61614
rect 196656 61478 196662 61542
rect 196726 61478 196868 61542
rect 196656 61472 196868 61478
rect 196248 61412 196324 61472
rect 22304 61276 22380 61336
rect 28560 61276 28636 61336
rect 190264 61276 190340 61336
rect 195976 61336 196324 61412
rect 195976 61276 196052 61336
rect 21760 61270 21972 61276
rect 21760 61206 21902 61270
rect 21966 61206 21972 61270
rect 1632 61012 1844 61140
rect 21760 61134 21972 61206
rect 21760 61070 21902 61134
rect 21966 61070 21972 61134
rect 21760 61064 21972 61070
rect 22168 61200 22788 61276
rect 22168 61134 22380 61200
rect 22168 61070 22174 61134
rect 22238 61070 22380 61134
rect 22168 61064 22380 61070
rect 22576 61140 22788 61200
rect 22984 61270 23196 61276
rect 22984 61206 23126 61270
rect 23190 61206 23196 61270
rect 22576 61134 22924 61140
rect 22576 61070 22718 61134
rect 22782 61070 22924 61134
rect 22576 61064 22924 61070
rect 22984 61134 23196 61206
rect 22984 61070 22990 61134
rect 23054 61070 23196 61134
rect 22984 61064 23196 61070
rect 23392 61270 23604 61276
rect 23392 61206 23534 61270
rect 23598 61206 23604 61270
rect 23392 61134 23604 61206
rect 23392 61070 23534 61134
rect 23598 61070 23604 61134
rect 23392 61064 23604 61070
rect 28288 61064 28636 61276
rect 190128 61064 190340 61276
rect 195024 61270 195236 61276
rect 195024 61206 195166 61270
rect 195230 61206 195236 61270
rect 195024 61134 195236 61206
rect 195024 61070 195030 61134
rect 195094 61070 195236 61134
rect 195024 61064 195236 61070
rect 195432 61270 195644 61276
rect 195432 61206 195574 61270
rect 195638 61206 195644 61270
rect 195432 61134 195644 61206
rect 195432 61070 195438 61134
rect 195502 61070 195644 61134
rect 195432 61064 195644 61070
rect 195840 61270 196460 61276
rect 195840 61206 195982 61270
rect 196046 61206 196460 61270
rect 195840 61200 196460 61206
rect 195840 61140 196052 61200
rect 195840 61134 196188 61140
rect 195840 61070 196118 61134
rect 196182 61070 196188 61134
rect 195840 61064 196188 61070
rect 196248 61064 196460 61200
rect 196656 61270 196868 61276
rect 196656 61206 196662 61270
rect 196726 61206 196868 61270
rect 196656 61134 196868 61206
rect 196656 61070 196662 61134
rect 196726 61070 196868 61134
rect 196656 61064 196868 61070
rect 216784 61134 217540 61140
rect 216784 61070 217470 61134
rect 217534 61070 217540 61134
rect 216784 61064 217540 61070
rect 1632 61004 1702 61012
rect 1224 60998 1702 61004
rect 1224 60934 1230 60998
rect 1294 60956 1702 60998
rect 1758 60956 1844 61012
rect 1294 60934 1844 60956
rect 1224 60928 1844 60934
rect 22848 61004 22924 61064
rect 28424 61004 28500 61064
rect 190264 61004 190340 61064
rect 22848 60928 23468 61004
rect 23392 60868 23468 60928
rect 21760 60862 21972 60868
rect 21760 60798 21902 60862
rect 21966 60798 21972 60862
rect 21760 60656 21972 60798
rect 22168 60862 22380 60868
rect 22168 60798 22174 60862
rect 22238 60798 22380 60862
rect 22168 60656 22380 60798
rect 22576 60862 22788 60868
rect 22576 60798 22718 60862
rect 22782 60798 22788 60862
rect 22576 60726 22788 60798
rect 22576 60662 22582 60726
rect 22646 60662 22788 60726
rect 22576 60656 22788 60662
rect 22984 60862 23196 60868
rect 22984 60798 22990 60862
rect 23054 60798 23196 60862
rect 22984 60726 23196 60798
rect 22984 60662 22990 60726
rect 23054 60662 23196 60726
rect 22984 60656 23196 60662
rect 23392 60862 23604 60868
rect 23392 60798 23534 60862
rect 23598 60798 23604 60862
rect 23392 60726 23604 60798
rect 28288 60792 28636 61004
rect 190128 60792 190340 61004
rect 216784 61012 216996 61064
rect 216784 60956 216908 61012
rect 216964 60956 216996 61012
rect 216784 60928 216996 60956
rect 195024 60862 195236 60868
rect 195024 60798 195030 60862
rect 195094 60798 195236 60862
rect 28424 60732 28500 60792
rect 190128 60732 190204 60792
rect 23392 60662 23534 60726
rect 23598 60662 23604 60726
rect 23392 60656 23604 60662
rect 21760 60596 21836 60656
rect 21760 60248 21972 60596
rect 28288 60520 28636 60732
rect 190128 60520 190340 60732
rect 195024 60726 195236 60798
rect 195024 60662 195166 60726
rect 195230 60662 195236 60726
rect 195024 60656 195236 60662
rect 195432 60862 195644 60868
rect 195432 60798 195438 60862
rect 195502 60798 195644 60862
rect 195432 60726 195644 60798
rect 195432 60662 195438 60726
rect 195502 60662 195644 60726
rect 195432 60656 195644 60662
rect 195840 60726 196052 60868
rect 196150 60862 196460 60868
rect 196112 60798 196118 60862
rect 196182 60798 196460 60862
rect 196150 60792 196460 60798
rect 195840 60662 195846 60726
rect 195910 60662 196052 60726
rect 195840 60656 196052 60662
rect 196248 60726 196460 60792
rect 196248 60662 196254 60726
rect 196318 60662 196460 60726
rect 196248 60656 196460 60662
rect 196656 60862 196868 60868
rect 196656 60798 196662 60862
rect 196726 60798 196868 60862
rect 196656 60656 196868 60798
rect 196656 60596 196732 60656
rect 28288 60460 28364 60520
rect 190128 60460 190204 60520
rect 22168 60248 22380 60460
rect 22576 60454 22788 60460
rect 22576 60390 22582 60454
rect 22646 60390 22788 60454
rect 22576 60248 22788 60390
rect 22984 60454 23196 60460
rect 22984 60390 22990 60454
rect 23054 60390 23196 60454
rect 22984 60318 23196 60390
rect 22984 60254 23126 60318
rect 23190 60254 23196 60318
rect 22984 60248 23196 60254
rect 23392 60454 23604 60460
rect 23392 60390 23534 60454
rect 23598 60390 23604 60454
rect 23392 60318 23604 60390
rect 23392 60254 23398 60318
rect 23462 60254 23604 60318
rect 23392 60248 23604 60254
rect 28288 60318 28636 60460
rect 28288 60254 28294 60318
rect 28358 60254 28636 60318
rect 21760 60188 21836 60248
rect 22168 60188 22244 60248
rect 22576 60188 22652 60248
rect 21760 59840 21972 60188
rect 22168 60112 22788 60188
rect 22168 59840 22380 60112
rect 22576 59910 22788 60112
rect 22576 59846 22582 59910
rect 22646 59846 22788 59910
rect 22576 59840 22788 59846
rect 22984 60046 23196 60052
rect 22984 59982 23126 60046
rect 23190 59982 23196 60046
rect 22984 59840 23196 59982
rect 23392 60046 23604 60052
rect 23392 59982 23398 60046
rect 23462 59982 23604 60046
rect 23392 59840 23604 59982
rect 28288 59976 28636 60254
rect 190128 59976 190340 60460
rect 195024 60454 195236 60460
rect 195024 60390 195166 60454
rect 195230 60390 195236 60454
rect 195024 60318 195236 60390
rect 195024 60254 195030 60318
rect 195094 60254 195236 60318
rect 195024 60248 195236 60254
rect 195432 60454 195644 60460
rect 195432 60390 195438 60454
rect 195502 60390 195644 60454
rect 195432 60318 195644 60390
rect 195432 60254 195438 60318
rect 195502 60254 195644 60318
rect 195432 60248 195644 60254
rect 195840 60454 196052 60460
rect 195840 60390 195846 60454
rect 195910 60390 196052 60454
rect 195840 60248 196052 60390
rect 196248 60454 196460 60460
rect 196248 60390 196254 60454
rect 196318 60390 196460 60454
rect 196248 60324 196460 60390
rect 196112 60248 196460 60324
rect 196656 60248 196868 60596
rect 195840 60188 195916 60248
rect 196112 60188 196188 60248
rect 196792 60188 196868 60248
rect 195840 60112 196188 60188
rect 28424 59916 28500 59976
rect 190264 59916 190340 59976
rect 21760 59780 21836 59840
rect 22984 59780 23060 59840
rect 23528 59780 23604 59840
rect 21760 59638 21972 59780
rect 21760 59574 21766 59638
rect 21830 59574 21972 59638
rect 21760 59568 21972 59574
rect 22168 59432 22380 59644
rect 22576 59638 22788 59644
rect 22576 59574 22582 59638
rect 22646 59574 22788 59638
rect 22576 59432 22788 59574
rect 22984 59432 23196 59780
rect 22168 59372 22244 59432
rect 22576 59372 22652 59432
rect 23120 59372 23196 59432
rect 1632 59332 1844 59372
rect 1632 59276 1702 59332
rect 1758 59276 1844 59332
rect 1632 59236 1844 59276
rect 1224 59230 1844 59236
rect 1224 59166 1230 59230
rect 1294 59166 1844 59230
rect 1224 59160 1844 59166
rect 21760 59366 21972 59372
rect 21760 59302 21766 59366
rect 21830 59302 21972 59366
rect 21760 59230 21972 59302
rect 21760 59166 21902 59230
rect 21966 59166 21972 59230
rect 21760 59160 21972 59166
rect 22168 59236 22380 59372
rect 22576 59236 22788 59372
rect 22168 59230 22788 59236
rect 22168 59166 22582 59230
rect 22646 59166 22788 59230
rect 22168 59160 22788 59166
rect 22984 59024 23196 59372
rect 23120 58964 23196 59024
rect 21760 58958 21972 58964
rect 21760 58894 21902 58958
rect 21966 58894 21972 58958
rect 21760 58822 21972 58894
rect 21760 58758 21766 58822
rect 21830 58758 21972 58822
rect 21760 58752 21972 58758
rect 22168 58828 22380 58964
rect 22576 58958 22788 58964
rect 22576 58894 22582 58958
rect 22646 58894 22788 58958
rect 22576 58828 22788 58894
rect 22168 58752 22788 58828
rect 22984 58822 23196 58964
rect 22984 58758 22990 58822
rect 23054 58758 23196 58822
rect 22984 58752 23196 58758
rect 23392 59432 23604 59780
rect 28288 59910 28636 59916
rect 28288 59846 28294 59910
rect 28358 59846 28636 59910
rect 23392 59372 23468 59432
rect 23392 59024 23604 59372
rect 28288 59366 28636 59846
rect 28288 59302 28566 59366
rect 28630 59302 28636 59366
rect 28288 59296 28636 59302
rect 190128 59366 190340 59916
rect 195024 60046 195236 60052
rect 195024 59982 195030 60046
rect 195094 59982 195236 60046
rect 195024 59840 195236 59982
rect 195432 60046 195644 60052
rect 195432 59982 195438 60046
rect 195502 59982 195644 60046
rect 195432 59840 195644 59982
rect 195840 59916 196052 60112
rect 196248 59916 196460 60188
rect 195840 59840 196460 59916
rect 196656 59840 196868 60188
rect 195024 59780 195100 59840
rect 195568 59780 195644 59840
rect 196248 59780 196324 59840
rect 195024 59432 195236 59780
rect 195160 59372 195236 59432
rect 190128 59302 190270 59366
rect 190334 59302 190340 59366
rect 190128 59296 190340 59302
rect 28288 59094 28636 59100
rect 28288 59030 28566 59094
rect 28630 59030 28636 59094
rect 23392 58964 23468 59024
rect 23392 58822 23604 58964
rect 23392 58758 23534 58822
rect 23598 58758 23604 58822
rect 23392 58752 23604 58758
rect 28288 58958 28636 59030
rect 28288 58894 28566 58958
rect 28630 58894 28636 58958
rect 28288 58752 28636 58894
rect 22168 58616 22380 58752
rect 22576 58616 22788 58752
rect 28560 58692 28636 58752
rect 28288 58686 28636 58692
rect 28288 58622 28566 58686
rect 28630 58622 28636 58686
rect 22168 58556 22244 58616
rect 22576 58556 22652 58616
rect 21760 58550 21972 58556
rect 21760 58486 21766 58550
rect 21830 58486 21972 58550
rect 21760 58414 21972 58486
rect 21760 58350 21902 58414
rect 21966 58350 21972 58414
rect 21760 58344 21972 58350
rect 22168 58344 22380 58556
rect 22576 58414 22788 58556
rect 22576 58350 22582 58414
rect 22646 58350 22788 58414
rect 22576 58344 22788 58350
rect 22984 58550 23196 58556
rect 22984 58486 22990 58550
rect 23054 58486 23196 58550
rect 22984 58414 23196 58486
rect 22984 58350 22990 58414
rect 23054 58350 23196 58414
rect 22984 58344 23196 58350
rect 23392 58550 23604 58556
rect 23392 58486 23534 58550
rect 23598 58486 23604 58550
rect 23392 58414 23604 58486
rect 28288 58480 28636 58622
rect 190128 59094 190340 59100
rect 190128 59030 190270 59094
rect 190334 59030 190340 59094
rect 190128 58958 190340 59030
rect 195024 59024 195236 59372
rect 195432 59432 195644 59780
rect 196112 59704 196324 59780
rect 196656 59780 196732 59840
rect 196112 59644 196188 59704
rect 195840 59568 196188 59644
rect 195840 59432 196052 59568
rect 196248 59432 196460 59644
rect 196656 59638 196868 59780
rect 196656 59574 196662 59638
rect 196726 59574 196868 59638
rect 196656 59568 196868 59574
rect 195432 59372 195508 59432
rect 195840 59372 195916 59432
rect 196248 59372 196324 59432
rect 195432 59024 195644 59372
rect 195840 59236 196052 59372
rect 196248 59236 196460 59372
rect 195840 59230 196460 59236
rect 195840 59166 195982 59230
rect 196046 59166 196460 59230
rect 195840 59160 196460 59166
rect 196656 59366 196868 59372
rect 196656 59302 196662 59366
rect 196726 59302 196868 59366
rect 196656 59230 196868 59302
rect 196656 59166 196798 59230
rect 196862 59166 196868 59230
rect 196656 59160 196868 59166
rect 216784 59366 217540 59372
rect 216784 59332 217470 59366
rect 216784 59276 216908 59332
rect 216964 59302 217470 59332
rect 217534 59302 217540 59366
rect 216964 59296 217540 59302
rect 216964 59276 216996 59296
rect 216784 59160 216996 59276
rect 195976 59100 196052 59160
rect 195976 59024 196324 59100
rect 195160 58964 195236 59024
rect 195568 58964 195644 59024
rect 196248 58964 196324 59024
rect 190128 58894 190134 58958
rect 190198 58894 190340 58958
rect 190128 58752 190340 58894
rect 195024 58822 195236 58964
rect 195024 58758 195166 58822
rect 195230 58758 195236 58822
rect 195024 58752 195236 58758
rect 195432 58822 195644 58964
rect 195432 58758 195438 58822
rect 195502 58758 195644 58822
rect 195432 58752 195644 58758
rect 195840 58958 196052 58964
rect 195840 58894 195982 58958
rect 196046 58894 196052 58958
rect 190128 58692 190204 58752
rect 190128 58686 190340 58692
rect 190128 58622 190134 58686
rect 190198 58622 190340 58686
rect 190128 58480 190340 58622
rect 195840 58616 196052 58894
rect 196248 58616 196460 58964
rect 196656 58958 196868 58964
rect 196656 58894 196798 58958
rect 196862 58894 196868 58958
rect 196656 58822 196868 58894
rect 196656 58758 196798 58822
rect 196862 58758 196868 58822
rect 196656 58752 196868 58758
rect 195840 58556 195916 58616
rect 195024 58550 195236 58556
rect 195024 58486 195166 58550
rect 195230 58486 195236 58550
rect 28424 58420 28500 58480
rect 190128 58420 190204 58480
rect 23392 58350 23534 58414
rect 23598 58350 23604 58414
rect 23392 58344 23604 58350
rect 21760 58142 21972 58148
rect 21760 58078 21902 58142
rect 21966 58078 21972 58142
rect 21760 58006 21972 58078
rect 21760 57942 21902 58006
rect 21966 57942 21972 58006
rect 21760 57936 21972 57942
rect 22168 58012 22380 58148
rect 22576 58142 22788 58148
rect 22576 58078 22582 58142
rect 22646 58078 22788 58142
rect 22576 58012 22788 58078
rect 22168 57936 22788 58012
rect 22984 58142 23196 58148
rect 22984 58078 22990 58142
rect 23054 58078 23196 58142
rect 22984 58006 23196 58078
rect 22984 57942 22990 58006
rect 23054 57942 23196 58006
rect 22984 57936 23196 57942
rect 23392 58142 23604 58148
rect 23392 58078 23534 58142
rect 23598 58078 23604 58142
rect 23392 58006 23604 58078
rect 23392 57942 23398 58006
rect 23462 57942 23604 58006
rect 23392 57936 23604 57942
rect 28288 58142 28636 58420
rect 28288 58078 28430 58142
rect 28494 58078 28636 58142
rect 28288 57936 28636 58078
rect 190128 57936 190340 58420
rect 195024 58414 195236 58486
rect 195024 58350 195030 58414
rect 195094 58350 195236 58414
rect 195024 58344 195236 58350
rect 195432 58550 195644 58556
rect 195432 58486 195438 58550
rect 195502 58486 195644 58550
rect 195432 58414 195644 58486
rect 195432 58350 195438 58414
rect 195502 58350 195644 58414
rect 195432 58344 195644 58350
rect 195840 58414 196052 58556
rect 196248 58420 196460 58556
rect 196150 58414 196460 58420
rect 195840 58350 195982 58414
rect 196046 58350 196052 58414
rect 196112 58350 196118 58414
rect 196182 58350 196460 58414
rect 195840 58344 196052 58350
rect 196150 58344 196460 58350
rect 196656 58550 196868 58556
rect 196656 58486 196798 58550
rect 196862 58486 196868 58550
rect 196656 58414 196868 58486
rect 196656 58350 196662 58414
rect 196726 58350 196868 58414
rect 196656 58344 196868 58350
rect 195024 58142 195236 58148
rect 195024 58078 195030 58142
rect 195094 58078 195236 58142
rect 195024 58006 195236 58078
rect 195024 57942 195030 58006
rect 195094 57942 195236 58006
rect 195024 57936 195236 57942
rect 195432 58142 195644 58148
rect 195432 58078 195438 58142
rect 195502 58078 195644 58142
rect 195432 58006 195644 58078
rect 195432 57942 195574 58006
rect 195638 57942 195644 58006
rect 195432 57936 195644 57942
rect 195840 58142 196188 58148
rect 195840 58078 195982 58142
rect 196046 58078 196118 58142
rect 196182 58078 196188 58142
rect 195840 58072 196188 58078
rect 195840 58012 196052 58072
rect 196248 58012 196460 58148
rect 195840 58006 196460 58012
rect 195840 57942 196390 58006
rect 196454 57942 196460 58006
rect 195840 57936 196460 57942
rect 196656 58142 196868 58148
rect 196656 58078 196662 58142
rect 196726 58078 196868 58142
rect 196656 58006 196868 58078
rect 196656 57942 196798 58006
rect 196862 57942 196868 58006
rect 196656 57936 196868 57942
rect 22304 57876 22380 57936
rect 28288 57876 28364 57936
rect 190264 57876 190340 57936
rect 22304 57800 22652 57876
rect 22576 57740 22652 57800
rect 28288 57870 28636 57876
rect 28288 57806 28430 57870
rect 28494 57806 28636 57870
rect 1224 57734 1844 57740
rect 1224 57670 1230 57734
rect 1294 57670 1844 57734
rect 1224 57664 1844 57670
rect 1632 57652 1844 57664
rect 1632 57596 1702 57652
rect 1758 57596 1844 57652
rect 1632 57528 1844 57596
rect 21760 57734 21972 57740
rect 21760 57670 21902 57734
rect 21966 57670 21972 57734
rect 21760 57598 21972 57670
rect 21760 57534 21766 57598
rect 21830 57534 21972 57598
rect 21760 57528 21972 57534
rect 22168 57664 22788 57740
rect 22168 57598 22380 57664
rect 22168 57534 22174 57598
rect 22238 57534 22380 57598
rect 22168 57528 22380 57534
rect 22576 57598 22788 57664
rect 22576 57534 22582 57598
rect 22646 57534 22788 57598
rect 22576 57528 22788 57534
rect 22984 57734 23196 57740
rect 22984 57670 22990 57734
rect 23054 57670 23196 57734
rect 22984 57598 23196 57670
rect 22984 57534 22990 57598
rect 23054 57534 23196 57598
rect 22984 57528 23196 57534
rect 23392 57734 23604 57740
rect 23392 57670 23398 57734
rect 23462 57670 23604 57734
rect 23392 57598 23604 57670
rect 28288 57664 28636 57806
rect 28560 57604 28636 57664
rect 23392 57534 23534 57598
rect 23598 57534 23604 57598
rect 23392 57528 23604 57534
rect 28288 57392 28636 57604
rect 190128 57664 190340 57876
rect 195024 57734 195236 57740
rect 195024 57670 195030 57734
rect 195094 57670 195236 57734
rect 190128 57604 190204 57664
rect 190128 57392 190340 57604
rect 195024 57598 195236 57670
rect 195024 57534 195166 57598
rect 195230 57534 195236 57598
rect 195024 57528 195236 57534
rect 195432 57734 195644 57740
rect 195432 57670 195574 57734
rect 195638 57670 195644 57734
rect 195432 57598 195644 57670
rect 195432 57534 195438 57598
rect 195502 57534 195644 57598
rect 195432 57528 195644 57534
rect 195840 57604 196052 57740
rect 196248 57734 196460 57740
rect 196248 57670 196390 57734
rect 196454 57670 196460 57734
rect 195840 57598 196188 57604
rect 195840 57534 196118 57598
rect 196182 57534 196188 57598
rect 195840 57528 196188 57534
rect 196248 57598 196460 57670
rect 196248 57534 196254 57598
rect 196318 57534 196460 57598
rect 196248 57528 196460 57534
rect 196656 57734 196868 57740
rect 196656 57670 196798 57734
rect 196862 57670 196868 57734
rect 196656 57598 196868 57670
rect 196656 57534 196662 57598
rect 196726 57534 196868 57598
rect 196656 57528 196868 57534
rect 216784 57652 216996 57740
rect 216784 57596 216908 57652
rect 216964 57604 216996 57652
rect 216964 57598 217540 57604
rect 216964 57596 217470 57598
rect 216784 57534 217470 57596
rect 217534 57534 217540 57598
rect 216784 57528 217540 57534
rect 28424 57332 28500 57392
rect 190128 57332 190204 57392
rect 21760 57326 21972 57332
rect 21760 57262 21766 57326
rect 21830 57262 21972 57326
rect 21760 57190 21972 57262
rect 21760 57126 21766 57190
rect 21830 57126 21972 57190
rect 21760 57120 21972 57126
rect 22168 57326 22380 57332
rect 22168 57262 22174 57326
rect 22238 57262 22380 57326
rect 22168 57120 22380 57262
rect 22576 57326 22788 57332
rect 22576 57262 22582 57326
rect 22646 57262 22788 57326
rect 22576 57120 22788 57262
rect 22984 57326 23196 57332
rect 22984 57262 22990 57326
rect 23054 57262 23196 57326
rect 22984 57190 23196 57262
rect 22984 57126 23126 57190
rect 23190 57126 23196 57190
rect 22984 57120 23196 57126
rect 23392 57326 23604 57332
rect 23392 57262 23534 57326
rect 23598 57262 23604 57326
rect 23392 57190 23604 57262
rect 23392 57126 23534 57190
rect 23598 57126 23604 57190
rect 23392 57120 23604 57126
rect 28288 57120 28636 57332
rect 190128 57120 190340 57332
rect 195024 57326 195236 57332
rect 195024 57262 195166 57326
rect 195230 57262 195236 57326
rect 195024 57190 195236 57262
rect 195024 57126 195166 57190
rect 195230 57126 195236 57190
rect 195024 57120 195236 57126
rect 195432 57326 195644 57332
rect 195432 57262 195438 57326
rect 195502 57262 195644 57326
rect 195432 57190 195644 57262
rect 195432 57126 195438 57190
rect 195502 57126 195644 57190
rect 195432 57120 195644 57126
rect 195840 57190 196052 57332
rect 196150 57326 196460 57332
rect 196112 57262 196118 57326
rect 196182 57262 196254 57326
rect 196318 57262 196460 57326
rect 196150 57256 196460 57262
rect 196248 57196 196460 57256
rect 196150 57190 196460 57196
rect 195840 57126 195846 57190
rect 195910 57126 196052 57190
rect 196112 57126 196118 57190
rect 196182 57126 196460 57190
rect 195840 57120 196052 57126
rect 196150 57120 196460 57126
rect 196656 57326 196868 57332
rect 196656 57262 196662 57326
rect 196726 57262 196868 57326
rect 196656 57190 196868 57262
rect 196656 57126 196798 57190
rect 196862 57126 196868 57190
rect 196656 57120 196868 57126
rect 22576 57060 22652 57120
rect 22304 56984 22652 57060
rect 28288 57060 28364 57120
rect 190264 57060 190340 57120
rect 22304 56924 22380 56984
rect 21760 56918 21972 56924
rect 21760 56854 21766 56918
rect 21830 56854 21972 56918
rect 21760 56788 21972 56854
rect 22168 56848 22788 56924
rect 21760 56712 22108 56788
rect 22168 56782 22380 56848
rect 22168 56718 22174 56782
rect 22238 56718 22380 56782
rect 22168 56712 22380 56718
rect 22576 56782 22788 56848
rect 22576 56718 22718 56782
rect 22782 56718 22788 56782
rect 22576 56712 22788 56718
rect 22984 56918 23196 56924
rect 22984 56854 23126 56918
rect 23190 56854 23196 56918
rect 22984 56782 23196 56854
rect 22984 56718 22990 56782
rect 23054 56718 23196 56782
rect 22984 56712 23196 56718
rect 23392 56918 23604 56924
rect 23392 56854 23534 56918
rect 23598 56854 23604 56918
rect 23392 56782 23604 56854
rect 28288 56848 28636 57060
rect 190128 56848 190340 57060
rect 28424 56788 28500 56848
rect 190264 56788 190340 56848
rect 23392 56718 23534 56782
rect 23598 56718 23604 56782
rect 23392 56712 23604 56718
rect 21896 56652 21972 56712
rect 21760 56304 21972 56652
rect 22032 56652 22108 56712
rect 22032 56576 23060 56652
rect 28288 56576 28636 56788
rect 190128 56646 190340 56788
rect 195024 56918 195236 56924
rect 195024 56854 195166 56918
rect 195230 56854 195236 56918
rect 195024 56782 195236 56854
rect 195024 56718 195166 56782
rect 195230 56718 195236 56782
rect 195024 56712 195236 56718
rect 195432 56918 195644 56924
rect 195432 56854 195438 56918
rect 195502 56854 195644 56918
rect 195432 56782 195644 56854
rect 195432 56718 195438 56782
rect 195502 56718 195644 56782
rect 195432 56712 195644 56718
rect 195840 56918 196188 56924
rect 195840 56854 195846 56918
rect 195910 56854 196118 56918
rect 196182 56854 196188 56918
rect 195840 56848 196188 56854
rect 195840 56788 196052 56848
rect 196248 56788 196460 56924
rect 195840 56782 196460 56788
rect 195840 56718 196254 56782
rect 196318 56718 196460 56782
rect 195840 56712 196460 56718
rect 196656 56918 196868 56924
rect 196656 56854 196798 56918
rect 196862 56854 196868 56918
rect 196656 56712 196868 56854
rect 196792 56652 196868 56712
rect 190128 56582 190270 56646
rect 190334 56582 190340 56646
rect 190128 56576 190340 56582
rect 22984 56516 23060 56576
rect 28424 56516 28500 56576
rect 190128 56516 190204 56576
rect 21896 56244 21972 56304
rect 1632 55972 1844 56108
rect 1224 55966 1702 55972
rect 1224 55902 1230 55966
rect 1294 55916 1702 55966
rect 1758 55916 1844 55972
rect 1294 55902 1844 55916
rect 1224 55896 1844 55902
rect 21760 55896 21972 56244
rect 22168 56510 22380 56516
rect 22168 56446 22174 56510
rect 22238 56446 22380 56510
rect 22168 56304 22380 56446
rect 22576 56510 22788 56516
rect 22576 56446 22718 56510
rect 22782 56446 22788 56510
rect 22576 56304 22788 56446
rect 22984 56510 23196 56516
rect 22984 56446 22990 56510
rect 23054 56446 23196 56510
rect 22984 56374 23196 56446
rect 22984 56310 22990 56374
rect 23054 56310 23196 56374
rect 22984 56304 23196 56310
rect 23392 56510 23604 56516
rect 23392 56446 23534 56510
rect 23598 56446 23604 56510
rect 23392 56374 23604 56446
rect 23392 56310 23534 56374
rect 23598 56310 23604 56374
rect 23392 56304 23604 56310
rect 22168 56244 22244 56304
rect 22576 56244 22652 56304
rect 22168 55896 22380 56244
rect 22576 55966 22788 56244
rect 22576 55902 22718 55966
rect 22782 55902 22788 55966
rect 22576 55896 22788 55902
rect 22984 56102 23196 56108
rect 22984 56038 22990 56102
rect 23054 56038 23196 56102
rect 22984 55966 23196 56038
rect 22984 55902 22990 55966
rect 23054 55902 23196 55966
rect 22984 55896 23196 55902
rect 23392 56102 23604 56108
rect 23392 56038 23534 56102
rect 23598 56038 23604 56102
rect 23392 55966 23604 56038
rect 23392 55902 23398 55966
rect 23462 55902 23604 55966
rect 23392 55896 23604 55902
rect 28288 56032 28636 56516
rect 190128 56374 190340 56516
rect 190128 56310 190270 56374
rect 190334 56310 190340 56374
rect 190128 56032 190340 56310
rect 195024 56510 195236 56516
rect 195024 56446 195166 56510
rect 195230 56446 195236 56510
rect 195024 56374 195236 56446
rect 195024 56310 195166 56374
rect 195230 56310 195236 56374
rect 195024 56304 195236 56310
rect 195432 56510 195644 56516
rect 195432 56446 195438 56510
rect 195502 56446 195644 56510
rect 195432 56374 195644 56446
rect 195432 56310 195574 56374
rect 195638 56310 195644 56374
rect 195432 56304 195644 56310
rect 195840 56510 196460 56516
rect 195840 56446 196254 56510
rect 196318 56446 196460 56510
rect 195840 56440 196460 56446
rect 195840 56304 196052 56440
rect 196248 56304 196460 56440
rect 196656 56304 196868 56652
rect 196248 56244 196324 56304
rect 196792 56244 196868 56304
rect 195840 56108 196052 56244
rect 196248 56108 196460 56244
rect 28288 55972 28364 56032
rect 190264 55972 190340 56032
rect 1632 55760 1844 55896
rect 21896 55836 21972 55896
rect 21760 55694 21972 55836
rect 28288 55830 28636 55972
rect 28288 55766 28294 55830
rect 28358 55766 28636 55830
rect 28288 55760 28636 55766
rect 190128 55760 190340 55972
rect 195024 56102 195236 56108
rect 195024 56038 195166 56102
rect 195230 56038 195236 56102
rect 195024 55966 195236 56038
rect 195024 55902 195030 55966
rect 195094 55902 195236 55966
rect 195024 55896 195236 55902
rect 195432 56102 195644 56108
rect 195432 56038 195574 56102
rect 195638 56038 195644 56102
rect 195432 55966 195644 56038
rect 195432 55902 195438 55966
rect 195502 55902 195644 55966
rect 195432 55896 195644 55902
rect 195840 56032 196460 56108
rect 195840 55972 196052 56032
rect 195840 55966 196188 55972
rect 195840 55902 195982 55966
rect 196046 55902 196118 55966
rect 196182 55902 196188 55966
rect 195840 55896 196188 55902
rect 196248 55896 196460 56032
rect 196656 55896 196868 56244
rect 196792 55836 196868 55896
rect 28560 55700 28636 55760
rect 190264 55700 190340 55760
rect 21760 55630 21766 55694
rect 21830 55630 21972 55694
rect 21760 55624 21972 55630
rect 22168 55564 22380 55700
rect 22576 55694 22788 55700
rect 22576 55630 22718 55694
rect 22782 55630 22788 55694
rect 22576 55564 22788 55630
rect 22168 55488 22788 55564
rect 22304 55428 22380 55488
rect 22712 55428 22788 55488
rect 21760 55422 21972 55428
rect 21760 55358 21766 55422
rect 21830 55358 21972 55422
rect 21760 55286 21972 55358
rect 21760 55222 21766 55286
rect 21830 55222 21972 55286
rect 21760 55216 21972 55222
rect 22168 55216 22380 55428
rect 22576 55286 22788 55428
rect 22576 55222 22582 55286
rect 22646 55222 22788 55286
rect 22576 55216 22788 55222
rect 22984 55694 23196 55700
rect 22984 55630 22990 55694
rect 23054 55630 23196 55694
rect 22984 55488 23196 55630
rect 23392 55694 23604 55700
rect 23392 55630 23398 55694
rect 23462 55630 23604 55694
rect 23392 55488 23604 55630
rect 22984 55428 23060 55488
rect 23528 55428 23604 55488
rect 22984 55080 23196 55428
rect 23120 55020 23196 55080
rect 21760 55014 21972 55020
rect 21760 54950 21766 55014
rect 21830 54950 21972 55014
rect 21760 54878 21972 54950
rect 21760 54814 21902 54878
rect 21966 54814 21972 54878
rect 21760 54808 21972 54814
rect 22168 54884 22380 55020
rect 22576 55014 22788 55020
rect 22576 54950 22582 55014
rect 22646 54950 22788 55014
rect 22576 54884 22788 54950
rect 22168 54808 22788 54884
rect 22168 54748 22380 54808
rect 22168 54672 22516 54748
rect 22576 54672 22788 54808
rect 22984 54672 23196 55020
rect 22304 54612 22380 54672
rect 21760 54606 21972 54612
rect 21760 54542 21902 54606
rect 21966 54542 21972 54606
rect 21760 54470 21972 54542
rect 21760 54406 21766 54470
rect 21830 54406 21972 54470
rect 21760 54400 21972 54406
rect 22168 54476 22380 54612
rect 22440 54612 22516 54672
rect 23120 54612 23196 54672
rect 22440 54536 22788 54612
rect 22168 54470 22516 54476
rect 22168 54406 22446 54470
rect 22510 54406 22516 54470
rect 22168 54400 22516 54406
rect 22576 54400 22788 54536
rect 22984 54470 23196 54612
rect 22984 54406 23126 54470
rect 23190 54406 23196 54470
rect 22984 54400 23196 54406
rect 23392 55080 23604 55428
rect 28288 55558 28636 55700
rect 28288 55494 28294 55558
rect 28358 55494 28636 55558
rect 28288 55422 28636 55494
rect 28288 55358 28294 55422
rect 28358 55358 28636 55422
rect 28288 55352 28636 55358
rect 190128 55422 190340 55700
rect 190128 55358 190134 55422
rect 190198 55358 190340 55422
rect 190128 55352 190340 55358
rect 195024 55694 195236 55700
rect 195024 55630 195030 55694
rect 195094 55630 195236 55694
rect 195024 55488 195236 55630
rect 195432 55694 195644 55700
rect 195432 55630 195438 55694
rect 195502 55630 195644 55694
rect 195432 55488 195644 55630
rect 195840 55694 196052 55700
rect 196150 55694 196460 55700
rect 195840 55630 195982 55694
rect 196046 55630 196052 55694
rect 196112 55630 196118 55694
rect 196182 55630 196460 55694
rect 195840 55488 196052 55630
rect 196150 55624 196460 55630
rect 196656 55694 196868 55836
rect 216784 55972 216996 56108
rect 216784 55916 216908 55972
rect 216964 55966 217540 55972
rect 216964 55916 217470 55966
rect 216784 55902 217470 55916
rect 217534 55902 217540 55966
rect 216784 55896 217540 55902
rect 216784 55760 216996 55896
rect 196656 55630 196662 55694
rect 196726 55630 196868 55694
rect 196656 55624 196868 55630
rect 196248 55488 196460 55624
rect 195024 55428 195100 55488
rect 195568 55428 195644 55488
rect 195976 55428 196052 55488
rect 196384 55428 196460 55488
rect 28288 55150 28636 55156
rect 28288 55086 28294 55150
rect 28358 55086 28636 55150
rect 23392 55020 23468 55080
rect 23392 54672 23604 55020
rect 28288 55014 28636 55086
rect 28288 54950 28566 55014
rect 28630 54950 28636 55014
rect 28288 54944 28636 54950
rect 190128 55150 190340 55156
rect 190128 55086 190134 55150
rect 190198 55086 190340 55150
rect 190128 55014 190340 55086
rect 195024 55080 195236 55428
rect 195160 55020 195236 55080
rect 190128 54950 190270 55014
rect 190334 54950 190340 55014
rect 28404 54748 28502 54944
rect 28288 54742 28636 54748
rect 28288 54678 28294 54742
rect 28358 54678 28566 54742
rect 28630 54678 28636 54742
rect 23392 54612 23468 54672
rect 23392 54470 23604 54612
rect 28288 54536 28636 54678
rect 190128 54742 190340 54950
rect 190128 54678 190270 54742
rect 190334 54678 190340 54742
rect 190128 54536 190340 54678
rect 28560 54476 28636 54536
rect 190264 54476 190340 54536
rect 23392 54406 23398 54470
rect 23462 54406 23604 54470
rect 23392 54400 23604 54406
rect 28288 54470 28636 54476
rect 28288 54406 28294 54470
rect 28358 54406 28636 54470
rect 1632 54292 1844 54340
rect 1632 54236 1702 54292
rect 1758 54236 1844 54292
rect 1632 54204 1844 54236
rect 1224 54198 1844 54204
rect 1224 54134 1230 54198
rect 1294 54134 1844 54198
rect 1224 54128 1844 54134
rect 21760 54198 21972 54204
rect 21760 54134 21766 54198
rect 21830 54134 21972 54198
rect 21760 54062 21972 54134
rect 21760 53998 21902 54062
rect 21966 53998 21972 54062
rect 21760 53992 21972 53998
rect 22168 54062 22380 54204
rect 22478 54198 22788 54204
rect 22440 54134 22446 54198
rect 22510 54134 22788 54198
rect 22478 54128 22788 54134
rect 22168 53998 22310 54062
rect 22374 53998 22380 54062
rect 22168 53992 22380 53998
rect 22576 54062 22788 54128
rect 22576 53998 22718 54062
rect 22782 53998 22788 54062
rect 22576 53992 22788 53998
rect 22984 54198 23196 54204
rect 22984 54134 23126 54198
rect 23190 54134 23196 54198
rect 22984 54062 23196 54134
rect 22984 53998 22990 54062
rect 23054 53998 23196 54062
rect 22984 53992 23196 53998
rect 23392 54198 23604 54204
rect 23392 54134 23398 54198
rect 23462 54134 23604 54198
rect 23392 54062 23604 54134
rect 23392 53998 23398 54062
rect 23462 53998 23604 54062
rect 23392 53992 23604 53998
rect 28288 53992 28636 54406
rect 190128 53992 190340 54476
rect 195024 54672 195236 55020
rect 195432 55080 195644 55428
rect 195840 55292 196052 55428
rect 195840 55286 196188 55292
rect 195840 55222 196118 55286
rect 196182 55222 196188 55286
rect 195840 55216 196188 55222
rect 196248 55216 196460 55428
rect 196656 55422 196868 55428
rect 196656 55358 196662 55422
rect 196726 55358 196868 55422
rect 196656 55286 196868 55358
rect 196656 55222 196662 55286
rect 196726 55222 196868 55286
rect 196656 55216 196868 55222
rect 195432 55020 195508 55080
rect 195432 54672 195644 55020
rect 195024 54612 195100 54672
rect 195568 54612 195644 54672
rect 195024 54470 195236 54612
rect 195024 54406 195166 54470
rect 195230 54406 195236 54470
rect 195024 54400 195236 54406
rect 195432 54470 195644 54612
rect 195432 54406 195574 54470
rect 195638 54406 195644 54470
rect 195432 54400 195644 54406
rect 195840 54672 196052 55020
rect 196150 55014 196460 55020
rect 196112 54950 196118 55014
rect 196182 54950 196460 55014
rect 196150 54944 196460 54950
rect 196248 54748 196460 54944
rect 196656 55014 196868 55020
rect 196656 54950 196662 55014
rect 196726 54950 196868 55014
rect 196656 54878 196868 54950
rect 196656 54814 196798 54878
rect 196862 54814 196868 54878
rect 196656 54808 196868 54814
rect 196112 54672 196460 54748
rect 195840 54612 195916 54672
rect 196112 54612 196188 54672
rect 196384 54612 196460 54672
rect 195840 54536 196188 54612
rect 195840 54470 196052 54536
rect 195840 54406 195846 54470
rect 195910 54406 196052 54470
rect 195840 54400 196052 54406
rect 196248 54470 196460 54612
rect 196248 54406 196390 54470
rect 196454 54406 196460 54470
rect 196248 54400 196460 54406
rect 196656 54606 196868 54612
rect 196656 54542 196798 54606
rect 196862 54542 196868 54606
rect 196656 54470 196868 54542
rect 196656 54406 196798 54470
rect 196862 54406 196868 54470
rect 196656 54400 196868 54406
rect 216784 54334 217540 54340
rect 216784 54292 217470 54334
rect 216784 54236 216908 54292
rect 216964 54270 217470 54292
rect 217534 54270 217540 54334
rect 216964 54264 217540 54270
rect 216964 54236 216996 54264
rect 195024 54198 195236 54204
rect 195024 54134 195166 54198
rect 195230 54134 195236 54198
rect 195024 54062 195236 54134
rect 195024 53998 195166 54062
rect 195230 53998 195236 54062
rect 195024 53992 195236 53998
rect 195432 54198 195644 54204
rect 195432 54134 195574 54198
rect 195638 54134 195644 54198
rect 195432 54062 195644 54134
rect 195432 53998 195574 54062
rect 195638 53998 195644 54062
rect 195432 53992 195644 53998
rect 195840 54198 196052 54204
rect 195840 54134 195846 54198
rect 195910 54134 196052 54198
rect 195840 53992 196052 54134
rect 196248 54198 196460 54204
rect 196248 54134 196390 54198
rect 196454 54134 196460 54198
rect 196248 53992 196460 54134
rect 196656 54198 196868 54204
rect 196656 54134 196798 54198
rect 196862 54134 196868 54198
rect 196656 54062 196868 54134
rect 216784 54128 216996 54236
rect 196656 53998 196798 54062
rect 196862 53998 196868 54062
rect 196656 53992 196868 53998
rect 28424 53932 28500 53992
rect 190128 53932 190204 53992
rect 196248 53932 196324 53992
rect 21760 53790 21972 53796
rect 21760 53726 21902 53790
rect 21966 53726 21972 53790
rect 21760 53654 21972 53726
rect 21760 53590 21902 53654
rect 21966 53590 21972 53654
rect 21760 53584 21972 53590
rect 22168 53790 22788 53796
rect 22168 53726 22310 53790
rect 22374 53726 22718 53790
rect 22782 53726 22788 53790
rect 22168 53720 22788 53726
rect 22168 53660 22380 53720
rect 22168 53584 22516 53660
rect 22576 53584 22788 53720
rect 22984 53790 23196 53796
rect 22984 53726 22990 53790
rect 23054 53726 23196 53790
rect 22984 53654 23196 53726
rect 22984 53590 23126 53654
rect 23190 53590 23196 53654
rect 22984 53584 23196 53590
rect 23392 53790 23604 53796
rect 23392 53726 23398 53790
rect 23462 53726 23604 53790
rect 23392 53654 23604 53726
rect 28288 53720 28636 53932
rect 190128 53720 190340 53932
rect 195976 53856 196324 53932
rect 195976 53796 196052 53856
rect 28424 53660 28500 53720
rect 190264 53660 190340 53720
rect 23392 53590 23398 53654
rect 23462 53590 23604 53654
rect 23392 53584 23604 53590
rect 22440 53524 22516 53584
rect 22440 53448 22652 53524
rect 28288 53448 28636 53660
rect 190128 53448 190340 53660
rect 195024 53790 195236 53796
rect 195024 53726 195166 53790
rect 195230 53726 195236 53790
rect 195024 53654 195236 53726
rect 195024 53590 195030 53654
rect 195094 53590 195236 53654
rect 195024 53584 195236 53590
rect 195432 53790 195644 53796
rect 195432 53726 195574 53790
rect 195638 53726 195644 53790
rect 195432 53654 195644 53726
rect 195432 53590 195574 53654
rect 195638 53590 195644 53654
rect 195432 53584 195644 53590
rect 195840 53720 196460 53796
rect 195840 53584 196052 53720
rect 196248 53654 196460 53720
rect 196248 53590 196390 53654
rect 196454 53590 196460 53654
rect 196248 53584 196460 53590
rect 196656 53790 196868 53796
rect 196656 53726 196798 53790
rect 196862 53726 196868 53790
rect 196656 53654 196868 53726
rect 196656 53590 196798 53654
rect 196862 53590 196868 53654
rect 196656 53584 196868 53590
rect 22576 53388 22652 53448
rect 28560 53388 28636 53448
rect 190264 53388 190340 53448
rect 21760 53382 21972 53388
rect 21760 53318 21902 53382
rect 21966 53318 21972 53382
rect 21760 53246 21972 53318
rect 21760 53182 21766 53246
rect 21830 53182 21972 53246
rect 21760 53176 21972 53182
rect 22168 53312 22788 53388
rect 22168 53252 22380 53312
rect 22168 53246 22516 53252
rect 22168 53182 22446 53246
rect 22510 53182 22516 53246
rect 22168 53176 22516 53182
rect 22576 53176 22788 53312
rect 22984 53382 23196 53388
rect 22984 53318 23126 53382
rect 23190 53318 23196 53382
rect 22984 53246 23196 53318
rect 22984 53182 22990 53246
rect 23054 53182 23196 53246
rect 22984 53176 23196 53182
rect 23392 53382 23604 53388
rect 23392 53318 23398 53382
rect 23462 53318 23604 53382
rect 23392 53246 23604 53318
rect 23392 53182 23534 53246
rect 23598 53182 23604 53246
rect 23392 53176 23604 53182
rect 28288 53176 28636 53388
rect 28560 53116 28636 53176
rect 21760 52974 21972 52980
rect 21760 52910 21766 52974
rect 21830 52910 21972 52974
rect 21760 52768 21972 52910
rect 22168 52838 22380 52980
rect 22478 52974 22788 52980
rect 22440 52910 22446 52974
rect 22510 52910 22788 52974
rect 22478 52904 22788 52910
rect 22168 52774 22310 52838
rect 22374 52774 22380 52838
rect 22168 52768 22380 52774
rect 22576 52768 22788 52904
rect 22984 52974 23196 52980
rect 22984 52910 22990 52974
rect 23054 52910 23196 52974
rect 22984 52838 23196 52910
rect 22984 52774 22990 52838
rect 23054 52774 23196 52838
rect 22984 52768 23196 52774
rect 23392 52974 23604 52980
rect 23392 52910 23534 52974
rect 23598 52910 23604 52974
rect 23392 52838 23604 52910
rect 28288 52904 28636 53116
rect 190128 53176 190340 53388
rect 195024 53382 195236 53388
rect 195024 53318 195030 53382
rect 195094 53318 195236 53382
rect 195024 53246 195236 53318
rect 195024 53182 195166 53246
rect 195230 53182 195236 53246
rect 195024 53176 195236 53182
rect 195432 53382 195644 53388
rect 195432 53318 195574 53382
rect 195638 53318 195644 53382
rect 195432 53246 195644 53318
rect 195432 53182 195438 53246
rect 195502 53182 195644 53246
rect 195432 53176 195644 53182
rect 195840 53246 196052 53388
rect 195840 53182 195846 53246
rect 195910 53182 196052 53246
rect 195840 53176 196052 53182
rect 196248 53382 196460 53388
rect 196248 53318 196390 53382
rect 196454 53318 196460 53382
rect 196248 53246 196460 53318
rect 196248 53182 196390 53246
rect 196454 53182 196460 53246
rect 196248 53176 196460 53182
rect 196656 53382 196868 53388
rect 196656 53318 196798 53382
rect 196862 53318 196868 53382
rect 196656 53246 196868 53318
rect 196656 53182 196662 53246
rect 196726 53182 196868 53246
rect 196656 53176 196868 53182
rect 190128 53116 190204 53176
rect 190128 52904 190340 53116
rect 195024 52974 195236 52980
rect 195024 52910 195166 52974
rect 195230 52910 195236 52974
rect 28424 52844 28500 52904
rect 190128 52844 190204 52904
rect 23392 52774 23398 52838
rect 23462 52774 23604 52838
rect 23392 52768 23604 52774
rect 21760 52708 21836 52768
rect 22576 52708 22652 52768
rect 1632 52612 1844 52708
rect 1632 52572 1702 52612
rect 1224 52566 1702 52572
rect 1224 52502 1230 52566
rect 1294 52556 1702 52566
rect 1758 52556 1844 52612
rect 1294 52502 1844 52556
rect 1224 52496 1844 52502
rect 21760 52360 21972 52708
rect 22304 52632 22652 52708
rect 28288 52632 28636 52844
rect 190128 52632 190340 52844
rect 195024 52838 195236 52910
rect 195024 52774 195166 52838
rect 195230 52774 195236 52838
rect 195024 52768 195236 52774
rect 195432 52974 195644 52980
rect 195432 52910 195438 52974
rect 195502 52910 195644 52974
rect 195432 52838 195644 52910
rect 195432 52774 195438 52838
rect 195502 52774 195644 52838
rect 195432 52768 195644 52774
rect 195840 52974 196052 52980
rect 195840 52910 195846 52974
rect 195910 52910 196052 52974
rect 195840 52838 196052 52910
rect 196248 52974 196460 52980
rect 196248 52910 196390 52974
rect 196454 52910 196460 52974
rect 196248 52844 196460 52910
rect 196150 52838 196460 52844
rect 195840 52774 195982 52838
rect 196046 52774 196052 52838
rect 196112 52774 196118 52838
rect 196182 52774 196390 52838
rect 196454 52774 196460 52838
rect 195840 52768 196052 52774
rect 196150 52768 196460 52774
rect 196656 52974 196868 52980
rect 196656 52910 196662 52974
rect 196726 52910 196868 52974
rect 196656 52768 196868 52910
rect 22304 52572 22380 52632
rect 28560 52572 28636 52632
rect 190264 52572 190340 52632
rect 196656 52708 196732 52768
rect 22168 52566 22788 52572
rect 22168 52502 22310 52566
rect 22374 52502 22788 52566
rect 22168 52496 22788 52502
rect 22168 52360 22380 52496
rect 22576 52360 22788 52496
rect 22984 52566 23196 52572
rect 22984 52502 22990 52566
rect 23054 52502 23196 52566
rect 22984 52430 23196 52502
rect 22984 52366 22990 52430
rect 23054 52366 23196 52430
rect 22984 52360 23196 52366
rect 23392 52566 23604 52572
rect 23392 52502 23398 52566
rect 23462 52502 23604 52566
rect 23392 52430 23604 52502
rect 23392 52366 23398 52430
rect 23462 52366 23604 52430
rect 23392 52360 23604 52366
rect 28288 52360 28636 52572
rect 190128 52360 190340 52572
rect 195024 52566 195236 52572
rect 195024 52502 195166 52566
rect 195230 52502 195236 52566
rect 195024 52430 195236 52502
rect 195024 52366 195166 52430
rect 195230 52366 195236 52430
rect 195024 52360 195236 52366
rect 195432 52566 195644 52572
rect 195432 52502 195438 52566
rect 195502 52502 195644 52566
rect 195432 52430 195644 52502
rect 195432 52366 195438 52430
rect 195502 52366 195644 52430
rect 195432 52360 195644 52366
rect 195840 52566 196188 52572
rect 195840 52502 195982 52566
rect 196046 52502 196118 52566
rect 196182 52502 196188 52566
rect 195840 52496 196188 52502
rect 196248 52566 196460 52572
rect 196248 52502 196390 52566
rect 196454 52502 196460 52566
rect 195840 52360 196052 52496
rect 196248 52360 196460 52502
rect 21760 52300 21836 52360
rect 22304 52300 22380 52360
rect 22712 52300 22788 52360
rect 28424 52300 28500 52360
rect 190264 52300 190340 52360
rect 195976 52300 196052 52360
rect 196384 52300 196460 52360
rect 21760 51952 21972 52300
rect 22168 51952 22380 52300
rect 22576 52224 22788 52300
rect 22688 52028 22788 52224
rect 22478 52022 22788 52028
rect 22440 51958 22446 52022
rect 22510 51958 22788 52022
rect 22478 51952 22788 51958
rect 22984 52158 23196 52164
rect 22984 52094 22990 52158
rect 23054 52094 23196 52158
rect 22984 52022 23196 52094
rect 22984 51958 23126 52022
rect 23190 51958 23196 52022
rect 22984 51952 23196 51958
rect 23392 52158 23604 52164
rect 23392 52094 23398 52158
rect 23462 52094 23604 52158
rect 23392 52022 23604 52094
rect 28288 52088 28636 52300
rect 190128 52088 190340 52300
rect 195024 52158 195236 52164
rect 195024 52094 195166 52158
rect 195230 52094 195236 52158
rect 28424 52028 28500 52088
rect 190128 52028 190204 52088
rect 23392 51958 23534 52022
rect 23598 51958 23604 52022
rect 23392 51952 23604 51958
rect 21760 51892 21836 51952
rect 21760 51750 21972 51892
rect 28288 51886 28636 52028
rect 28288 51822 28294 51886
rect 28358 51822 28636 51886
rect 28288 51816 28636 51822
rect 190128 51816 190340 52028
rect 195024 52022 195236 52094
rect 195024 51958 195166 52022
rect 195230 51958 195236 52022
rect 195024 51952 195236 51958
rect 195432 52158 195644 52164
rect 195432 52094 195438 52158
rect 195502 52094 195644 52158
rect 195432 52022 195644 52094
rect 195432 51958 195438 52022
rect 195502 51958 195644 52022
rect 195432 51952 195644 51958
rect 195840 52022 196052 52300
rect 195840 51958 195846 52022
rect 195910 51958 196052 52022
rect 195840 51952 196052 51958
rect 196248 51952 196460 52300
rect 196656 52360 196868 52708
rect 216784 52702 217540 52708
rect 216784 52638 217470 52702
rect 217534 52638 217540 52702
rect 216784 52632 217540 52638
rect 216784 52612 216996 52632
rect 216784 52556 216908 52612
rect 216964 52556 216996 52612
rect 216784 52496 216996 52556
rect 196656 52300 196732 52360
rect 196656 51952 196868 52300
rect 196656 51892 196732 51952
rect 28288 51756 28364 51816
rect 190128 51756 190204 51816
rect 21760 51686 21902 51750
rect 21966 51686 21972 51750
rect 21760 51680 21972 51686
rect 22168 51750 22516 51756
rect 22168 51686 22446 51750
rect 22510 51686 22516 51750
rect 22168 51680 22516 51686
rect 22168 51544 22380 51680
rect 22576 51620 22788 51756
rect 22304 51484 22380 51544
rect 22440 51544 22788 51620
rect 22440 51484 22516 51544
rect 22712 51484 22788 51544
rect 21760 51478 21972 51484
rect 21760 51414 21902 51478
rect 21966 51414 21972 51478
rect 21760 51342 21972 51414
rect 21760 51278 21766 51342
rect 21830 51278 21972 51342
rect 21760 51272 21972 51278
rect 22168 51408 22516 51484
rect 22168 51272 22380 51408
rect 22576 51342 22788 51484
rect 22576 51278 22718 51342
rect 22782 51278 22788 51342
rect 22576 51272 22788 51278
rect 22984 51750 23196 51756
rect 22984 51686 23126 51750
rect 23190 51686 23196 51750
rect 22984 51544 23196 51686
rect 23392 51750 23604 51756
rect 23392 51686 23534 51750
rect 23598 51686 23604 51750
rect 23392 51544 23604 51686
rect 28288 51614 28636 51756
rect 28288 51550 28294 51614
rect 28358 51550 28636 51614
rect 22984 51484 23060 51544
rect 23392 51484 23468 51544
rect 22984 51136 23196 51484
rect 23392 51136 23604 51484
rect 28288 51478 28636 51550
rect 28288 51414 28294 51478
rect 28358 51414 28636 51478
rect 28288 51408 28636 51414
rect 190128 51478 190340 51756
rect 190128 51414 190270 51478
rect 190334 51414 190340 51478
rect 190128 51408 190340 51414
rect 195024 51750 195236 51756
rect 195024 51686 195166 51750
rect 195230 51686 195236 51750
rect 195024 51544 195236 51686
rect 195432 51750 195644 51756
rect 195432 51686 195438 51750
rect 195502 51686 195644 51750
rect 195432 51544 195644 51686
rect 195840 51750 196052 51756
rect 195840 51686 195846 51750
rect 195910 51686 196052 51750
rect 195840 51620 196052 51686
rect 195840 51544 196188 51620
rect 196248 51544 196460 51756
rect 196656 51750 196868 51892
rect 196656 51686 196662 51750
rect 196726 51686 196868 51750
rect 196656 51680 196868 51686
rect 195024 51484 195100 51544
rect 195568 51484 195644 51544
rect 195976 51484 196052 51544
rect 22984 51076 23060 51136
rect 23528 51076 23604 51136
rect 1632 50940 1844 51076
rect 1224 50934 1844 50940
rect 1224 50870 1230 50934
rect 1294 50932 1844 50934
rect 1294 50876 1702 50932
rect 1758 50876 1844 50932
rect 1294 50870 1844 50876
rect 1224 50864 1844 50870
rect 21760 51070 21972 51076
rect 21760 51006 21766 51070
rect 21830 51006 21972 51070
rect 21760 50934 21972 51006
rect 21760 50870 21766 50934
rect 21830 50870 21972 50934
rect 21760 50864 21972 50870
rect 1632 50728 1844 50864
rect 22168 50728 22380 51076
rect 22576 51070 22788 51076
rect 22576 51006 22718 51070
rect 22782 51006 22788 51070
rect 22576 50804 22788 51006
rect 22304 50668 22380 50728
rect 22440 50728 22788 50804
rect 22984 50728 23196 51076
rect 22440 50668 22516 50728
rect 22712 50668 22788 50728
rect 23120 50668 23196 50728
rect 21760 50662 21972 50668
rect 21760 50598 21766 50662
rect 21830 50598 21972 50662
rect 21760 50526 21972 50598
rect 21760 50462 21902 50526
rect 21966 50462 21972 50526
rect 21760 50456 21972 50462
rect 22168 50592 22516 50668
rect 22168 50456 22380 50592
rect 22576 50526 22788 50668
rect 22576 50462 22718 50526
rect 22782 50462 22788 50526
rect 22576 50456 22788 50462
rect 22984 50526 23196 50668
rect 22984 50462 22990 50526
rect 23054 50462 23196 50526
rect 22984 50456 23196 50462
rect 23392 50728 23604 51076
rect 28288 51206 28636 51212
rect 28288 51142 28294 51206
rect 28358 51142 28636 51206
rect 23392 50668 23468 50728
rect 23392 50526 23604 50668
rect 28288 50592 28636 51142
rect 28560 50532 28636 50592
rect 23392 50462 23398 50526
rect 23462 50462 23604 50526
rect 23392 50456 23604 50462
rect 21760 50254 21972 50260
rect 21760 50190 21902 50254
rect 21966 50190 21972 50254
rect 21760 50118 21972 50190
rect 21760 50054 21766 50118
rect 21830 50054 21972 50118
rect 21760 50048 21972 50054
rect 22168 50124 22380 50260
rect 22576 50254 22788 50260
rect 22576 50190 22718 50254
rect 22782 50190 22788 50254
rect 22576 50124 22788 50190
rect 22168 50118 22788 50124
rect 22168 50054 22310 50118
rect 22374 50054 22788 50118
rect 22168 50048 22788 50054
rect 22984 50254 23196 50260
rect 22984 50190 22990 50254
rect 23054 50190 23196 50254
rect 22984 50118 23196 50190
rect 22984 50054 22990 50118
rect 23054 50054 23196 50118
rect 22984 50048 23196 50054
rect 23392 50254 23604 50260
rect 23392 50190 23398 50254
rect 23462 50190 23604 50254
rect 23392 50118 23604 50190
rect 23392 50054 23398 50118
rect 23462 50054 23604 50118
rect 23392 50048 23604 50054
rect 28288 50254 28636 50532
rect 28288 50190 28294 50254
rect 28358 50190 28636 50254
rect 28288 50048 28636 50190
rect 28560 49988 28636 50048
rect 28288 49982 28636 49988
rect 28288 49918 28294 49982
rect 28358 49918 28636 49982
rect 21760 49846 21972 49852
rect 21760 49782 21766 49846
rect 21830 49782 21972 49846
rect 21760 49710 21972 49782
rect 21760 49646 21766 49710
rect 21830 49646 21972 49710
rect 21760 49640 21972 49646
rect 22168 49846 22380 49852
rect 22168 49782 22310 49846
rect 22374 49782 22380 49846
rect 22168 49710 22380 49782
rect 22168 49646 22174 49710
rect 22238 49646 22380 49710
rect 22168 49640 22380 49646
rect 22576 49710 22788 49852
rect 22576 49646 22718 49710
rect 22782 49646 22788 49710
rect 22576 49640 22788 49646
rect 22984 49846 23196 49852
rect 22984 49782 22990 49846
rect 23054 49782 23196 49846
rect 22984 49710 23196 49782
rect 22984 49646 22990 49710
rect 23054 49646 23196 49710
rect 22984 49640 23196 49646
rect 23392 49846 23604 49852
rect 23392 49782 23398 49846
rect 23462 49782 23604 49846
rect 23392 49710 23604 49782
rect 23392 49646 23398 49710
rect 23462 49646 23604 49710
rect 23392 49640 23604 49646
rect 28288 49776 28636 49918
rect 190128 51206 190340 51212
rect 190128 51142 190270 51206
rect 190334 51142 190340 51206
rect 190128 50592 190340 51142
rect 195024 51136 195236 51484
rect 195160 51076 195236 51136
rect 195024 50728 195236 51076
rect 195432 51136 195644 51484
rect 195840 51342 196052 51484
rect 196112 51484 196188 51544
rect 196384 51484 196460 51544
rect 196112 51408 196460 51484
rect 195840 51278 195982 51342
rect 196046 51278 196052 51342
rect 195840 51272 196052 51278
rect 196248 51272 196460 51408
rect 196656 51478 196868 51484
rect 196656 51414 196662 51478
rect 196726 51414 196868 51478
rect 196656 51342 196868 51414
rect 196656 51278 196662 51342
rect 196726 51278 196868 51342
rect 196656 51272 196868 51278
rect 195432 51076 195508 51136
rect 195432 50728 195644 51076
rect 195160 50668 195236 50728
rect 195568 50668 195644 50728
rect 190128 50532 190204 50592
rect 190128 50048 190340 50532
rect 195024 50526 195236 50668
rect 195024 50462 195030 50526
rect 195094 50462 195236 50526
rect 195024 50456 195236 50462
rect 195432 50526 195644 50668
rect 195432 50462 195438 50526
rect 195502 50462 195644 50526
rect 195432 50456 195644 50462
rect 195840 51070 196052 51076
rect 195840 51006 195982 51070
rect 196046 51006 196052 51070
rect 195840 50728 196052 51006
rect 196248 50728 196460 51076
rect 196656 51070 196868 51076
rect 196656 51006 196662 51070
rect 196726 51006 196868 51070
rect 196656 50934 196868 51006
rect 196656 50870 196662 50934
rect 196726 50870 196868 50934
rect 196656 50864 196868 50870
rect 216784 50932 216996 51076
rect 216784 50876 216908 50932
rect 216964 50876 216996 50932
rect 216784 50804 216996 50876
rect 216784 50798 217540 50804
rect 216784 50734 217470 50798
rect 217534 50734 217540 50798
rect 216784 50728 217540 50734
rect 195840 50668 195916 50728
rect 196248 50668 196324 50728
rect 195840 50526 196052 50668
rect 195840 50462 195982 50526
rect 196046 50462 196052 50526
rect 195840 50456 196052 50462
rect 196248 50456 196460 50668
rect 196656 50662 196868 50668
rect 196656 50598 196662 50662
rect 196726 50598 196868 50662
rect 196656 50526 196868 50598
rect 196656 50462 196798 50526
rect 196862 50462 196868 50526
rect 196656 50456 196868 50462
rect 196248 50396 196324 50456
rect 195976 50320 196324 50396
rect 195976 50260 196052 50320
rect 195024 50254 195236 50260
rect 195024 50190 195030 50254
rect 195094 50190 195236 50254
rect 195024 50118 195236 50190
rect 195024 50054 195030 50118
rect 195094 50054 195236 50118
rect 195024 50048 195236 50054
rect 195432 50254 195644 50260
rect 195432 50190 195438 50254
rect 195502 50190 195644 50254
rect 195432 50118 195644 50190
rect 195432 50054 195438 50118
rect 195502 50054 195644 50118
rect 195432 50048 195644 50054
rect 195840 50254 196460 50260
rect 195840 50190 195982 50254
rect 196046 50190 196460 50254
rect 195840 50184 196460 50190
rect 195840 50048 196052 50184
rect 196248 50118 196460 50184
rect 196248 50054 196390 50118
rect 196454 50054 196460 50118
rect 196248 50048 196460 50054
rect 196656 50254 196868 50260
rect 196656 50190 196798 50254
rect 196862 50190 196868 50254
rect 196656 50118 196868 50190
rect 196656 50054 196798 50118
rect 196862 50054 196868 50118
rect 196656 50048 196868 50054
rect 190128 49988 190204 50048
rect 190128 49776 190340 49988
rect 195024 49846 195236 49852
rect 195024 49782 195030 49846
rect 195094 49782 195236 49846
rect 28288 49716 28364 49776
rect 190128 49716 190204 49776
rect 195024 49716 195236 49782
rect 195432 49846 195644 49852
rect 195432 49782 195438 49846
rect 195502 49782 195644 49846
rect 28288 49504 28636 49716
rect 190128 49504 190340 49716
rect 195024 49710 195372 49716
rect 195024 49646 195030 49710
rect 195094 49646 195372 49710
rect 195024 49640 195372 49646
rect 195432 49710 195644 49782
rect 195432 49646 195438 49710
rect 195502 49646 195644 49710
rect 195432 49640 195644 49646
rect 195840 49710 196052 49852
rect 195840 49646 195846 49710
rect 195910 49646 196052 49710
rect 195840 49640 196052 49646
rect 196248 49846 196460 49852
rect 196248 49782 196390 49846
rect 196454 49782 196460 49846
rect 196248 49640 196460 49782
rect 196656 49846 196868 49852
rect 196656 49782 196798 49846
rect 196862 49782 196868 49846
rect 196656 49710 196868 49782
rect 196656 49646 196662 49710
rect 196726 49646 196868 49710
rect 196656 49640 196868 49646
rect 195296 49580 195372 49640
rect 195840 49580 195916 49640
rect 196248 49580 196324 49640
rect 195296 49504 195916 49580
rect 195976 49504 196324 49580
rect 28424 49444 28500 49504
rect 190264 49444 190340 49504
rect 195976 49444 196052 49504
rect 21760 49438 21972 49444
rect 21760 49374 21766 49438
rect 21830 49374 21972 49438
rect 1224 49302 1844 49308
rect 1224 49238 1230 49302
rect 1294 49252 1844 49302
rect 1294 49238 1702 49252
rect 1224 49232 1702 49238
rect 1632 49196 1702 49232
rect 1758 49196 1844 49252
rect 21760 49302 21972 49374
rect 21760 49238 21902 49302
rect 21966 49238 21972 49302
rect 21760 49232 21972 49238
rect 22168 49438 22380 49444
rect 22168 49374 22174 49438
rect 22238 49374 22380 49438
rect 22168 49308 22380 49374
rect 22576 49438 22788 49444
rect 22576 49374 22718 49438
rect 22782 49374 22788 49438
rect 22576 49308 22788 49374
rect 22168 49302 22788 49308
rect 22168 49238 22310 49302
rect 22374 49238 22788 49302
rect 22168 49232 22788 49238
rect 22984 49438 23196 49444
rect 22984 49374 22990 49438
rect 23054 49374 23196 49438
rect 22984 49302 23196 49374
rect 22984 49238 23126 49302
rect 23190 49238 23196 49302
rect 22984 49232 23196 49238
rect 23392 49438 23604 49444
rect 23392 49374 23398 49438
rect 23462 49374 23604 49438
rect 23392 49302 23604 49374
rect 23392 49238 23398 49302
rect 23462 49238 23604 49302
rect 23392 49232 23604 49238
rect 28288 49232 28636 49444
rect 190128 49232 190340 49444
rect 195024 49438 195236 49444
rect 195024 49374 195030 49438
rect 195094 49374 195236 49438
rect 195024 49302 195236 49374
rect 195024 49238 195030 49302
rect 195094 49238 195236 49302
rect 195024 49232 195236 49238
rect 195432 49438 195644 49444
rect 195432 49374 195438 49438
rect 195502 49374 195644 49438
rect 195432 49302 195644 49374
rect 195432 49238 195574 49302
rect 195638 49238 195644 49302
rect 195432 49232 195644 49238
rect 195840 49438 196460 49444
rect 195840 49374 195846 49438
rect 195910 49374 196460 49438
rect 195840 49368 196460 49374
rect 195840 49232 196052 49368
rect 196248 49302 196460 49368
rect 196248 49238 196390 49302
rect 196454 49238 196460 49302
rect 196248 49232 196460 49238
rect 196656 49438 196868 49444
rect 196656 49374 196662 49438
rect 196726 49374 196868 49438
rect 196656 49302 196868 49374
rect 196656 49238 196798 49302
rect 196862 49238 196868 49302
rect 196656 49232 196868 49238
rect 216784 49252 216996 49308
rect 1632 49096 1844 49196
rect 22304 49172 22380 49232
rect 28288 49172 28364 49232
rect 190264 49172 190340 49232
rect 22304 49096 22652 49172
rect 22576 49036 22652 49096
rect 21760 49030 21972 49036
rect 21760 48966 21902 49030
rect 21966 48966 21972 49030
rect 21760 48824 21972 48966
rect 22168 49030 22380 49036
rect 22168 48966 22310 49030
rect 22374 48966 22380 49030
rect 22168 48894 22380 48966
rect 22168 48830 22174 48894
rect 22238 48830 22380 48894
rect 22168 48824 22380 48830
rect 22576 48824 22788 49036
rect 22984 49030 23196 49036
rect 22984 48966 23126 49030
rect 23190 48966 23196 49030
rect 22984 48894 23196 48966
rect 22984 48830 22990 48894
rect 23054 48830 23196 48894
rect 22984 48824 23196 48830
rect 23392 49030 23604 49036
rect 23392 48966 23398 49030
rect 23462 48966 23604 49030
rect 23392 48894 23604 48966
rect 28288 48960 28636 49172
rect 28560 48900 28636 48960
rect 23392 48830 23534 48894
rect 23598 48830 23604 48894
rect 23392 48824 23604 48830
rect 21760 48764 21836 48824
rect 21760 48486 21972 48764
rect 28288 48688 28636 48900
rect 190128 48960 190340 49172
rect 216784 49196 216908 49252
rect 216964 49196 216996 49252
rect 216784 49172 216996 49196
rect 216784 49166 217540 49172
rect 216784 49102 217470 49166
rect 217534 49102 217540 49166
rect 216784 49096 217540 49102
rect 195024 49030 195236 49036
rect 195024 48966 195030 49030
rect 195094 48966 195236 49030
rect 190128 48900 190204 48960
rect 190128 48688 190340 48900
rect 195024 48894 195236 48966
rect 195024 48830 195166 48894
rect 195230 48830 195236 48894
rect 195024 48824 195236 48830
rect 195432 49030 195644 49036
rect 195432 48966 195574 49030
rect 195638 48966 195644 49030
rect 195432 48894 195644 48966
rect 195432 48830 195438 48894
rect 195502 48830 195644 48894
rect 195432 48824 195644 48830
rect 195840 48894 196052 49036
rect 195840 48830 195846 48894
rect 195910 48830 196052 48894
rect 195840 48824 196052 48830
rect 196248 49030 196460 49036
rect 196248 48966 196390 49030
rect 196454 48966 196460 49030
rect 196248 48894 196460 48966
rect 196248 48830 196254 48894
rect 196318 48830 196460 48894
rect 196248 48824 196460 48830
rect 196656 49030 196868 49036
rect 196656 48966 196798 49030
rect 196862 48966 196868 49030
rect 196656 48824 196868 48966
rect 196656 48764 196732 48824
rect 28424 48628 28500 48688
rect 190128 48628 190204 48688
rect 21760 48422 21902 48486
rect 21966 48422 21972 48486
rect 21760 48416 21972 48422
rect 22168 48622 22380 48628
rect 22168 48558 22174 48622
rect 22238 48558 22380 48622
rect 22168 48486 22380 48558
rect 22168 48422 22310 48486
rect 22374 48422 22380 48486
rect 22168 48416 22380 48422
rect 22576 48486 22788 48628
rect 22576 48422 22582 48486
rect 22646 48422 22788 48486
rect 22576 48416 22788 48422
rect 22984 48622 23196 48628
rect 22984 48558 22990 48622
rect 23054 48558 23196 48622
rect 22984 48486 23196 48558
rect 22984 48422 23126 48486
rect 23190 48422 23196 48486
rect 22984 48416 23196 48422
rect 23392 48622 23604 48628
rect 23392 48558 23534 48622
rect 23598 48558 23604 48622
rect 23392 48486 23604 48558
rect 23392 48422 23534 48486
rect 23598 48422 23604 48486
rect 23392 48416 23604 48422
rect 28288 48416 28636 48628
rect 28560 48356 28636 48416
rect 21760 48214 21972 48220
rect 21760 48150 21902 48214
rect 21966 48150 21972 48214
rect 21760 48008 21972 48150
rect 22168 48214 22788 48220
rect 22168 48150 22310 48214
rect 22374 48150 22582 48214
rect 22646 48150 22788 48214
rect 22168 48144 22788 48150
rect 22168 48008 22380 48144
rect 22576 48078 22788 48144
rect 22576 48014 22718 48078
rect 22782 48014 22788 48078
rect 22576 48008 22788 48014
rect 22984 48214 23196 48220
rect 22984 48150 23126 48214
rect 23190 48150 23196 48214
rect 22984 48078 23196 48150
rect 22984 48014 22990 48078
rect 23054 48014 23196 48078
rect 22984 48008 23196 48014
rect 23392 48214 23604 48220
rect 23392 48150 23534 48214
rect 23598 48150 23604 48214
rect 23392 48078 23604 48150
rect 28288 48144 28636 48356
rect 190128 48416 190340 48628
rect 195024 48622 195236 48628
rect 195024 48558 195166 48622
rect 195230 48558 195236 48622
rect 195024 48486 195236 48558
rect 195024 48422 195030 48486
rect 195094 48422 195236 48486
rect 195024 48416 195236 48422
rect 195432 48622 195644 48628
rect 195432 48558 195438 48622
rect 195502 48558 195644 48622
rect 195432 48486 195644 48558
rect 195432 48422 195574 48486
rect 195638 48422 195644 48486
rect 195432 48416 195644 48422
rect 195840 48622 196052 48628
rect 195840 48558 195846 48622
rect 195910 48558 196052 48622
rect 195840 48486 196052 48558
rect 196248 48622 196460 48628
rect 196248 48558 196254 48622
rect 196318 48558 196460 48622
rect 196248 48492 196460 48558
rect 196150 48486 196460 48492
rect 195840 48422 195846 48486
rect 195910 48422 196052 48486
rect 196112 48422 196118 48486
rect 196182 48422 196460 48486
rect 195840 48416 196052 48422
rect 196150 48416 196460 48422
rect 196656 48486 196868 48764
rect 196656 48422 196798 48486
rect 196862 48422 196868 48486
rect 196656 48416 196868 48422
rect 190128 48356 190204 48416
rect 190128 48144 190340 48356
rect 28560 48084 28636 48144
rect 190264 48084 190340 48144
rect 23392 48014 23534 48078
rect 23598 48014 23604 48078
rect 23392 48008 23604 48014
rect 21896 47948 21972 48008
rect 21760 47806 21972 47948
rect 28288 47872 28636 48084
rect 190128 47872 190340 48084
rect 195024 48214 195236 48220
rect 195024 48150 195030 48214
rect 195094 48150 195236 48214
rect 195024 48078 195236 48150
rect 195024 48014 195166 48078
rect 195230 48014 195236 48078
rect 195024 48008 195236 48014
rect 195432 48214 195644 48220
rect 195432 48150 195574 48214
rect 195638 48150 195644 48214
rect 195432 48078 195644 48150
rect 195432 48014 195438 48078
rect 195502 48014 195644 48078
rect 195432 48008 195644 48014
rect 195840 48214 196188 48220
rect 195840 48150 195846 48214
rect 195910 48150 196118 48214
rect 196182 48150 196188 48214
rect 195840 48144 196188 48150
rect 195840 48084 196052 48144
rect 196248 48084 196460 48220
rect 195840 48078 196460 48084
rect 195840 48014 196254 48078
rect 196318 48014 196460 48078
rect 195840 48008 196460 48014
rect 196656 48214 196868 48220
rect 196656 48150 196798 48214
rect 196862 48150 196868 48214
rect 196656 48008 196868 48150
rect 196792 47948 196868 48008
rect 28424 47812 28500 47872
rect 190264 47812 190340 47872
rect 21760 47742 21902 47806
rect 21966 47742 21972 47806
rect 21760 47736 21972 47742
rect 22168 47676 22380 47812
rect 22576 47806 22788 47812
rect 22576 47742 22718 47806
rect 22782 47742 22788 47806
rect 1224 47670 1844 47676
rect 1224 47606 1230 47670
rect 1294 47606 1844 47670
rect 1224 47600 1844 47606
rect 1632 47572 1844 47600
rect 1632 47516 1702 47572
rect 1758 47516 1844 47572
rect 22168 47600 22516 47676
rect 22168 47540 22244 47600
rect 22440 47540 22516 47600
rect 22576 47600 22788 47742
rect 22984 47806 23196 47812
rect 22984 47742 22990 47806
rect 23054 47742 23196 47806
rect 22984 47670 23196 47742
rect 22984 47606 22990 47670
rect 23054 47606 23196 47670
rect 22984 47600 23196 47606
rect 23392 47806 23604 47812
rect 23392 47742 23534 47806
rect 23598 47742 23604 47806
rect 23392 47670 23604 47742
rect 23392 47606 23534 47670
rect 23598 47606 23604 47670
rect 23392 47600 23604 47606
rect 22576 47540 22652 47600
rect 1632 47464 1844 47516
rect 21760 47534 21972 47540
rect 21760 47470 21902 47534
rect 21966 47470 21972 47534
rect 21760 47192 21972 47470
rect 22168 47192 22380 47540
rect 22440 47464 22788 47540
rect 22576 47268 22788 47464
rect 22478 47262 22788 47268
rect 22440 47198 22446 47262
rect 22510 47198 22788 47262
rect 22478 47192 22788 47198
rect 22984 47398 23196 47404
rect 22984 47334 22990 47398
rect 23054 47334 23196 47398
rect 22984 47192 23196 47334
rect 23392 47398 23604 47404
rect 23392 47334 23534 47398
rect 23598 47334 23604 47398
rect 23392 47192 23604 47334
rect 28288 47328 28636 47812
rect 190128 47328 190340 47812
rect 195024 47806 195236 47812
rect 195024 47742 195166 47806
rect 195230 47742 195236 47806
rect 195024 47670 195236 47742
rect 195024 47606 195166 47670
rect 195230 47606 195236 47670
rect 195024 47600 195236 47606
rect 195432 47806 195644 47812
rect 195432 47742 195438 47806
rect 195502 47742 195644 47806
rect 195432 47670 195644 47742
rect 195432 47606 195438 47670
rect 195502 47606 195644 47670
rect 195432 47600 195644 47606
rect 195840 47600 196052 47812
rect 195976 47540 196052 47600
rect 28288 47268 28364 47328
rect 190264 47268 190340 47328
rect 21896 47132 21972 47192
rect 21760 46990 21972 47132
rect 22984 47132 23060 47192
rect 23392 47132 23468 47192
rect 21760 46926 21902 46990
rect 21966 46926 21972 46990
rect 21760 46920 21972 46926
rect 22168 46990 22516 46996
rect 22168 46926 22446 46990
rect 22510 46926 22516 46990
rect 22168 46920 22516 46926
rect 22168 46860 22380 46920
rect 22576 46860 22788 46996
rect 22168 46854 22788 46860
rect 22168 46790 22310 46854
rect 22374 46790 22788 46854
rect 22168 46784 22788 46790
rect 22984 46784 23196 47132
rect 23392 46784 23604 47132
rect 28288 47126 28636 47268
rect 28288 47062 28294 47126
rect 28358 47062 28636 47126
rect 28288 46854 28636 47062
rect 28288 46790 28294 46854
rect 28358 46790 28636 46854
rect 22168 46724 22244 46784
rect 22984 46724 23060 46784
rect 23392 46724 23468 46784
rect 21760 46718 21972 46724
rect 21760 46654 21902 46718
rect 21966 46654 21972 46718
rect 21760 46582 21972 46654
rect 21760 46518 21766 46582
rect 21830 46518 21972 46582
rect 21760 46512 21972 46518
rect 22168 46512 22380 46724
rect 22478 46718 22788 46724
rect 22440 46654 22446 46718
rect 22510 46654 22788 46718
rect 22478 46648 22788 46654
rect 22576 46582 22788 46648
rect 22576 46518 22582 46582
rect 22646 46518 22788 46582
rect 22576 46512 22788 46518
rect 22984 46582 23196 46724
rect 22984 46518 22990 46582
rect 23054 46518 23196 46582
rect 22984 46512 23196 46518
rect 23392 46582 23604 46724
rect 28288 46648 28636 46790
rect 190128 46648 190340 47268
rect 195024 47398 195236 47404
rect 195024 47334 195166 47398
rect 195230 47334 195236 47398
rect 195024 47192 195236 47334
rect 195432 47398 195644 47404
rect 195432 47334 195438 47398
rect 195502 47334 195644 47398
rect 195432 47192 195644 47334
rect 195840 47268 196052 47540
rect 196248 47806 196460 47812
rect 196248 47742 196254 47806
rect 196318 47742 196460 47806
rect 196248 47600 196460 47742
rect 196656 47806 196868 47948
rect 196656 47742 196662 47806
rect 196726 47742 196868 47806
rect 196656 47736 196868 47742
rect 196248 47540 196324 47600
rect 216784 47572 216996 47676
rect 196248 47268 196460 47540
rect 195840 47192 196460 47268
rect 196656 47534 196868 47540
rect 196656 47470 196662 47534
rect 196726 47470 196868 47534
rect 196656 47192 196868 47470
rect 216784 47516 216908 47572
rect 216964 47540 216996 47572
rect 216964 47534 217540 47540
rect 216964 47516 217470 47534
rect 216784 47470 217470 47516
rect 217534 47470 217540 47534
rect 216784 47464 217540 47470
rect 195024 47132 195100 47192
rect 195432 47132 195508 47192
rect 196248 47132 196324 47192
rect 196792 47132 196868 47192
rect 195024 46784 195236 47132
rect 195160 46724 195236 46784
rect 28424 46588 28500 46648
rect 190128 46588 190204 46648
rect 23392 46518 23534 46582
rect 23598 46518 23604 46582
rect 23392 46512 23604 46518
rect 21760 46310 21972 46316
rect 21760 46246 21766 46310
rect 21830 46246 21972 46310
rect 21760 46174 21972 46246
rect 21760 46110 21902 46174
rect 21966 46110 21972 46174
rect 21760 46104 21972 46110
rect 1224 46038 1844 46044
rect 1224 45974 1230 46038
rect 1294 45974 1844 46038
rect 1224 45968 1844 45974
rect 22168 45968 22380 46316
rect 22576 46310 22788 46316
rect 22576 46246 22582 46310
rect 22646 46246 22788 46310
rect 22576 46240 22788 46246
rect 22688 46044 22788 46240
rect 22984 46310 23196 46316
rect 22984 46246 22990 46310
rect 23054 46246 23196 46310
rect 22984 46174 23196 46246
rect 22984 46110 23126 46174
rect 23190 46110 23196 46174
rect 22984 46104 23196 46110
rect 23392 46310 23604 46316
rect 23392 46246 23534 46310
rect 23598 46246 23604 46310
rect 23392 46174 23604 46246
rect 23392 46110 23398 46174
rect 23462 46110 23604 46174
rect 23392 46104 23604 46110
rect 28288 46104 28636 46588
rect 190128 46310 190340 46588
rect 195024 46582 195236 46724
rect 195024 46518 195166 46582
rect 195230 46518 195236 46582
rect 195024 46512 195236 46518
rect 195432 46784 195644 47132
rect 195976 47056 196324 47132
rect 195976 46996 196052 47056
rect 195840 46920 196460 46996
rect 196656 46990 196868 47132
rect 196656 46926 196798 46990
rect 196862 46926 196868 46990
rect 196656 46920 196868 46926
rect 195840 46784 196052 46920
rect 196248 46784 196460 46920
rect 195432 46724 195508 46784
rect 195840 46724 195916 46784
rect 196248 46724 196324 46784
rect 195432 46582 195644 46724
rect 195432 46518 195438 46582
rect 195502 46518 195644 46582
rect 195432 46512 195644 46518
rect 195840 46512 196052 46724
rect 196248 46582 196460 46724
rect 196248 46518 196254 46582
rect 196318 46518 196460 46582
rect 196248 46512 196460 46518
rect 196656 46718 196868 46724
rect 196656 46654 196798 46718
rect 196862 46654 196868 46718
rect 196656 46582 196868 46654
rect 196656 46518 196662 46582
rect 196726 46518 196868 46582
rect 196656 46512 196868 46518
rect 190128 46246 190134 46310
rect 190198 46246 190340 46310
rect 190128 46104 190340 46246
rect 195024 46310 195236 46316
rect 195024 46246 195166 46310
rect 195230 46246 195236 46310
rect 195024 46174 195236 46246
rect 195024 46110 195030 46174
rect 195094 46110 195236 46174
rect 195024 46104 195236 46110
rect 195432 46310 195644 46316
rect 195432 46246 195438 46310
rect 195502 46246 195644 46310
rect 195432 46174 195644 46246
rect 195432 46110 195574 46174
rect 195638 46110 195644 46174
rect 195432 46104 195644 46110
rect 28424 46044 28500 46104
rect 190264 46044 190340 46104
rect 1632 45892 1844 45968
rect 22304 45908 22380 45968
rect 22440 45968 22788 46044
rect 22440 45908 22516 45968
rect 1632 45836 1702 45892
rect 1758 45836 1844 45892
rect 1632 45696 1844 45836
rect 21760 45902 21972 45908
rect 21760 45838 21902 45902
rect 21966 45838 21972 45902
rect 14552 45630 14764 45772
rect 21760 45766 21972 45838
rect 21760 45702 21902 45766
rect 21966 45702 21972 45766
rect 21760 45696 21972 45702
rect 22168 45832 22516 45908
rect 22168 45772 22380 45832
rect 22576 45772 22788 45908
rect 22168 45766 22788 45772
rect 22168 45702 22174 45766
rect 22238 45702 22788 45766
rect 22168 45696 22788 45702
rect 22984 45902 23196 45908
rect 22984 45838 23126 45902
rect 23190 45838 23196 45902
rect 22984 45766 23196 45838
rect 22984 45702 23126 45766
rect 23190 45702 23196 45766
rect 22984 45696 23196 45702
rect 23392 45902 23604 45908
rect 23392 45838 23398 45902
rect 23462 45838 23604 45902
rect 23392 45766 23604 45838
rect 28288 45832 28636 46044
rect 190128 46038 190340 46044
rect 190128 45974 190134 46038
rect 190198 45974 190340 46038
rect 190128 45832 190340 45974
rect 195840 45968 196052 46316
rect 196248 46310 196460 46316
rect 196248 46246 196254 46310
rect 196318 46246 196460 46310
rect 196248 46044 196460 46246
rect 196656 46310 196868 46316
rect 196656 46246 196662 46310
rect 196726 46246 196868 46310
rect 196656 46174 196868 46246
rect 196656 46110 196798 46174
rect 196862 46110 196868 46174
rect 196656 46104 196868 46110
rect 196112 45968 196460 46044
rect 195840 45908 195916 45968
rect 196112 45908 196188 45968
rect 196384 45908 196460 45968
rect 216784 46038 217540 46044
rect 216784 45974 217470 46038
rect 217534 45974 217540 46038
rect 216784 45968 217540 45974
rect 28560 45772 28636 45832
rect 190264 45772 190340 45832
rect 23392 45702 23534 45766
rect 23598 45702 23604 45766
rect 23392 45696 23604 45702
rect 14552 45566 14694 45630
rect 14758 45566 14764 45630
rect 14552 45560 14764 45566
rect 22304 45636 22380 45696
rect 22304 45560 22652 45636
rect 22576 45500 22652 45560
rect 28288 45560 28636 45772
rect 190128 45560 190340 45772
rect 195024 45902 195236 45908
rect 195024 45838 195030 45902
rect 195094 45838 195236 45902
rect 195024 45766 195236 45838
rect 195024 45702 195166 45766
rect 195230 45702 195236 45766
rect 195024 45696 195236 45702
rect 195432 45902 195644 45908
rect 195432 45838 195574 45902
rect 195638 45838 195644 45902
rect 195432 45766 195644 45838
rect 195432 45702 195574 45766
rect 195638 45702 195644 45766
rect 195432 45696 195644 45702
rect 195840 45832 196188 45908
rect 195840 45766 196052 45832
rect 195840 45702 195846 45766
rect 195910 45702 196052 45766
rect 195840 45696 196052 45702
rect 196248 45696 196460 45908
rect 196656 45902 196868 45908
rect 196656 45838 196798 45902
rect 196862 45838 196868 45902
rect 196656 45766 196868 45838
rect 196656 45702 196662 45766
rect 196726 45702 196868 45766
rect 196656 45696 196868 45702
rect 216784 45892 216996 45968
rect 216784 45836 216908 45892
rect 216964 45836 216996 45892
rect 216784 45696 216996 45836
rect 28288 45500 28364 45560
rect 190128 45500 190204 45560
rect 21760 45494 21972 45500
rect 21760 45430 21902 45494
rect 21966 45430 21972 45494
rect 21760 45358 21972 45430
rect 21760 45294 21902 45358
rect 21966 45294 21972 45358
rect 21760 45288 21972 45294
rect 22168 45494 22380 45500
rect 22168 45430 22174 45494
rect 22238 45430 22380 45494
rect 22168 45288 22380 45430
rect 22576 45358 22788 45500
rect 22576 45294 22718 45358
rect 22782 45294 22788 45358
rect 22576 45288 22788 45294
rect 22984 45494 23196 45500
rect 22984 45430 23126 45494
rect 23190 45430 23196 45494
rect 22984 45358 23196 45430
rect 22984 45294 22990 45358
rect 23054 45294 23196 45358
rect 22984 45288 23196 45294
rect 23392 45494 23604 45500
rect 23392 45430 23534 45494
rect 23598 45430 23604 45494
rect 23392 45358 23604 45430
rect 23392 45294 23534 45358
rect 23598 45294 23604 45358
rect 23392 45288 23604 45294
rect 28288 45288 28636 45500
rect 190128 45288 190340 45500
rect 195024 45494 195236 45500
rect 195024 45430 195166 45494
rect 195230 45430 195236 45494
rect 195024 45358 195236 45430
rect 195024 45294 195166 45358
rect 195230 45294 195236 45358
rect 195024 45288 195236 45294
rect 195432 45494 195644 45500
rect 195432 45430 195574 45494
rect 195638 45430 195644 45494
rect 195432 45358 195644 45430
rect 195432 45294 195438 45358
rect 195502 45294 195644 45358
rect 195432 45288 195644 45294
rect 195840 45494 196052 45500
rect 195840 45430 195846 45494
rect 195910 45430 196052 45494
rect 195840 45358 196052 45430
rect 196248 45364 196460 45500
rect 196150 45358 196460 45364
rect 195840 45294 195846 45358
rect 195910 45294 196052 45358
rect 196112 45294 196118 45358
rect 196182 45294 196460 45358
rect 195840 45288 196052 45294
rect 196150 45288 196460 45294
rect 196656 45494 196868 45500
rect 196656 45430 196662 45494
rect 196726 45430 196868 45494
rect 196656 45358 196868 45430
rect 196656 45294 196662 45358
rect 196726 45294 196868 45358
rect 196656 45288 196868 45294
rect 28424 45228 28500 45288
rect 190128 45228 190204 45288
rect 0 45152 14356 45228
rect 14144 45093 14356 45152
rect 14144 45037 14212 45093
rect 14268 45037 14356 45093
rect 14144 44880 14356 45037
rect 21760 45086 21972 45092
rect 15152 45024 15218 45027
rect 15966 45024 16032 45027
rect 15152 45022 16032 45024
rect 15152 44966 15157 45022
rect 15213 44966 15971 45022
rect 16027 44966 16032 45022
rect 15152 44964 16032 44966
rect 15152 44961 15218 44964
rect 15966 44961 16032 44964
rect 21760 45022 21902 45086
rect 21966 45022 21972 45086
rect 21760 44950 21972 45022
rect 21760 44886 21902 44950
rect 21966 44886 21972 44950
rect 21760 44880 21972 44886
rect 22168 44956 22380 45092
rect 22576 45086 22788 45092
rect 22576 45022 22718 45086
rect 22782 45022 22788 45086
rect 22576 44956 22788 45022
rect 22168 44950 22788 44956
rect 22168 44886 22310 44950
rect 22374 44886 22788 44950
rect 22168 44880 22788 44886
rect 22984 45086 23196 45092
rect 22984 45022 22990 45086
rect 23054 45022 23196 45086
rect 22984 44950 23196 45022
rect 22984 44886 23126 44950
rect 23190 44886 23196 44950
rect 22984 44880 23196 44886
rect 23392 45086 23604 45092
rect 23392 45022 23534 45086
rect 23598 45022 23604 45086
rect 23392 44950 23604 45022
rect 28288 45016 28636 45228
rect 190128 45016 190340 45228
rect 28424 44956 28500 45016
rect 190264 44956 190340 45016
rect 23392 44886 23398 44950
rect 23462 44886 23604 44950
rect 23392 44880 23604 44886
rect 22304 44820 22380 44880
rect 22304 44744 22652 44820
rect 28288 44744 28636 44956
rect 190128 44744 190340 44956
rect 195024 45086 195236 45092
rect 195024 45022 195166 45086
rect 195230 45022 195236 45086
rect 195024 44950 195236 45022
rect 195024 44886 195030 44950
rect 195094 44886 195236 44950
rect 195024 44880 195236 44886
rect 195432 45086 195644 45092
rect 195432 45022 195438 45086
rect 195502 45022 195644 45086
rect 195432 44950 195644 45022
rect 195432 44886 195438 44950
rect 195502 44886 195644 44950
rect 195432 44880 195644 44886
rect 195840 45086 196188 45092
rect 195840 45022 195846 45086
rect 195910 45022 196118 45086
rect 196182 45022 196188 45086
rect 195840 45016 196188 45022
rect 195840 44956 196052 45016
rect 196248 44956 196460 45092
rect 195840 44950 196460 44956
rect 195840 44886 196390 44950
rect 196454 44886 196460 44950
rect 195840 44880 196460 44886
rect 196656 45086 196868 45092
rect 196656 45022 196662 45086
rect 196726 45022 196868 45086
rect 196656 44950 196868 45022
rect 196656 44886 196798 44950
rect 196862 44886 196868 44950
rect 196656 44880 196868 44886
rect 22576 44684 22652 44744
rect 28560 44684 28636 44744
rect 190264 44684 190340 44744
rect 21760 44678 21972 44684
rect 21760 44614 21902 44678
rect 21966 44614 21972 44678
rect 21760 44542 21972 44614
rect 21760 44478 21766 44542
rect 21830 44478 21972 44542
rect 21760 44472 21972 44478
rect 22168 44678 22380 44684
rect 22168 44614 22310 44678
rect 22374 44614 22380 44678
rect 22168 44542 22380 44614
rect 22168 44478 22174 44542
rect 22238 44478 22380 44542
rect 22168 44472 22380 44478
rect 22576 44542 22788 44684
rect 22576 44478 22582 44542
rect 22646 44478 22788 44542
rect 22576 44472 22788 44478
rect 22984 44678 23196 44684
rect 22984 44614 23126 44678
rect 23190 44614 23196 44678
rect 22984 44542 23196 44614
rect 22984 44478 22990 44542
rect 23054 44478 23196 44542
rect 22984 44472 23196 44478
rect 23392 44678 23604 44684
rect 23392 44614 23398 44678
rect 23462 44614 23604 44678
rect 23392 44542 23604 44614
rect 23392 44478 23534 44542
rect 23598 44478 23604 44542
rect 23392 44472 23604 44478
rect 28288 44472 28636 44684
rect 28560 44412 28636 44472
rect 1632 44212 1844 44276
rect 1632 44156 1702 44212
rect 1758 44156 1844 44212
rect 1632 44140 1844 44156
rect 1224 44134 1844 44140
rect 1224 44070 1230 44134
rect 1294 44070 1844 44134
rect 1224 44064 1844 44070
rect 14552 44134 14764 44276
rect 14552 44070 14558 44134
rect 14622 44070 14764 44134
rect 14552 44064 14764 44070
rect 21760 44270 21972 44276
rect 21760 44206 21766 44270
rect 21830 44206 21972 44270
rect 21760 44064 21972 44206
rect 22168 44270 22380 44276
rect 22168 44206 22174 44270
rect 22238 44206 22380 44270
rect 22168 44064 22380 44206
rect 22576 44270 22788 44276
rect 22576 44206 22582 44270
rect 22646 44206 22788 44270
rect 22576 44140 22788 44206
rect 22478 44134 22788 44140
rect 22440 44070 22446 44134
rect 22510 44070 22788 44134
rect 22478 44064 22788 44070
rect 22984 44270 23196 44276
rect 22984 44206 22990 44270
rect 23054 44206 23196 44270
rect 22984 44134 23196 44206
rect 22984 44070 23126 44134
rect 23190 44070 23196 44134
rect 22984 44064 23196 44070
rect 23392 44270 23604 44276
rect 23392 44206 23534 44270
rect 23598 44206 23604 44270
rect 23392 44134 23604 44206
rect 28288 44200 28636 44412
rect 190128 44472 190340 44684
rect 195024 44678 195236 44684
rect 195024 44614 195030 44678
rect 195094 44614 195236 44678
rect 195024 44542 195236 44614
rect 195024 44478 195166 44542
rect 195230 44478 195236 44542
rect 195024 44472 195236 44478
rect 195432 44678 195644 44684
rect 195432 44614 195438 44678
rect 195502 44614 195644 44678
rect 195432 44542 195644 44614
rect 195432 44478 195574 44542
rect 195638 44478 195644 44542
rect 195432 44472 195644 44478
rect 195840 44678 196460 44684
rect 195840 44614 196390 44678
rect 196454 44614 196460 44678
rect 195840 44608 196460 44614
rect 195840 44472 196052 44608
rect 196248 44542 196460 44608
rect 196248 44478 196254 44542
rect 196318 44478 196460 44542
rect 196248 44472 196460 44478
rect 196656 44678 196868 44684
rect 196656 44614 196798 44678
rect 196862 44614 196868 44678
rect 196656 44542 196868 44614
rect 196656 44478 196662 44542
rect 196726 44478 196868 44542
rect 196656 44472 196868 44478
rect 190128 44412 190204 44472
rect 190128 44200 190340 44412
rect 195024 44270 195236 44276
rect 195024 44206 195166 44270
rect 195230 44206 195236 44270
rect 28424 44140 28500 44200
rect 190128 44140 190204 44200
rect 23392 44070 23534 44134
rect 23598 44070 23604 44134
rect 23392 44064 23604 44070
rect 21896 44004 21972 44064
rect 21760 43656 21972 44004
rect 28288 43928 28636 44140
rect 190128 43928 190340 44140
rect 195024 44134 195236 44206
rect 195024 44070 195030 44134
rect 195094 44070 195236 44134
rect 195024 44064 195236 44070
rect 195432 44270 195644 44276
rect 195432 44206 195574 44270
rect 195638 44206 195644 44270
rect 195432 44134 195644 44206
rect 195432 44070 195574 44134
rect 195638 44070 195644 44134
rect 195432 44064 195644 44070
rect 195840 44134 196052 44276
rect 195840 44070 195982 44134
rect 196046 44070 196052 44134
rect 195840 44064 196052 44070
rect 196248 44270 196460 44276
rect 196248 44206 196254 44270
rect 196318 44206 196460 44270
rect 196248 44134 196460 44206
rect 196248 44070 196390 44134
rect 196454 44070 196460 44134
rect 196248 44064 196460 44070
rect 196656 44270 196868 44276
rect 196656 44206 196662 44270
rect 196726 44206 196868 44270
rect 196656 44064 196868 44206
rect 216784 44270 217540 44276
rect 216784 44212 217470 44270
rect 216784 44156 216908 44212
rect 216964 44206 217470 44212
rect 217534 44206 217540 44270
rect 216964 44200 217540 44206
rect 216964 44156 216996 44200
rect 216784 44064 216996 44156
rect 28560 43868 28636 43928
rect 190264 43868 190340 43928
rect 196656 44004 196732 44064
rect 22168 43862 22516 43868
rect 22168 43798 22446 43862
rect 22510 43798 22516 43862
rect 22168 43792 22516 43798
rect 22168 43732 22380 43792
rect 22168 43656 22516 43732
rect 22576 43656 22788 43868
rect 22984 43862 23196 43868
rect 22984 43798 23126 43862
rect 23190 43798 23196 43862
rect 22984 43726 23196 43798
rect 22984 43662 22990 43726
rect 23054 43662 23196 43726
rect 22984 43656 23196 43662
rect 23392 43862 23604 43868
rect 23392 43798 23534 43862
rect 23598 43798 23604 43862
rect 23392 43726 23604 43798
rect 23392 43662 23398 43726
rect 23462 43662 23604 43726
rect 23392 43656 23604 43662
rect 21760 43596 21836 43656
rect 22304 43596 22380 43656
rect 15152 43466 15218 43469
rect 15886 43466 15952 43469
rect 15152 43464 15952 43466
rect 14144 43393 14356 43460
rect 15152 43408 15157 43464
rect 15213 43408 15891 43464
rect 15947 43408 15952 43464
rect 15152 43406 15952 43408
rect 15152 43403 15218 43406
rect 15886 43403 15952 43406
rect 14144 43337 14212 43393
rect 14268 43337 14356 43393
rect 14144 43324 14356 43337
rect 0 43248 14356 43324
rect 21760 43248 21972 43596
rect 22168 43248 22380 43596
rect 22440 43596 22516 43656
rect 22712 43596 22788 43656
rect 22440 43520 22788 43596
rect 22576 43324 22788 43520
rect 22478 43318 22788 43324
rect 22440 43254 22446 43318
rect 22510 43254 22788 43318
rect 22478 43248 22788 43254
rect 22984 43454 23196 43460
rect 22984 43390 22990 43454
rect 23054 43390 23196 43454
rect 22984 43248 23196 43390
rect 23392 43454 23604 43460
rect 23392 43390 23398 43454
rect 23462 43390 23604 43454
rect 23392 43248 23604 43390
rect 28288 43384 28636 43868
rect 190128 43454 190340 43868
rect 195024 43862 195236 43868
rect 195024 43798 195030 43862
rect 195094 43798 195236 43862
rect 195024 43726 195236 43798
rect 195024 43662 195030 43726
rect 195094 43662 195236 43726
rect 195024 43656 195236 43662
rect 195432 43862 195644 43868
rect 195432 43798 195574 43862
rect 195638 43798 195644 43862
rect 195432 43726 195644 43798
rect 195432 43662 195574 43726
rect 195638 43662 195644 43726
rect 195432 43656 195644 43662
rect 195840 43862 196052 43868
rect 195840 43798 195982 43862
rect 196046 43798 196052 43862
rect 195840 43732 196052 43798
rect 196248 43862 196460 43868
rect 196248 43798 196390 43862
rect 196454 43798 196460 43862
rect 195840 43656 196188 43732
rect 196248 43656 196460 43798
rect 196656 43656 196868 44004
rect 195840 43596 195916 43656
rect 196112 43596 196188 43656
rect 196384 43596 196460 43656
rect 196792 43596 196868 43656
rect 190128 43390 190134 43454
rect 190198 43390 190340 43454
rect 190128 43384 190340 43390
rect 195024 43454 195236 43460
rect 195024 43390 195030 43454
rect 195094 43390 195236 43454
rect 28424 43324 28500 43384
rect 190128 43324 190204 43384
rect 21760 43188 21836 43248
rect 22984 43188 23060 43248
rect 23528 43188 23604 43248
rect 21760 43046 21972 43188
rect 21760 42982 21766 43046
rect 21830 42982 21972 43046
rect 21760 42976 21972 42982
rect 22168 43046 22516 43052
rect 22168 42982 22446 43046
rect 22510 42982 22516 43046
rect 22168 42976 22516 42982
rect 14552 42910 14764 42916
rect 14552 42846 14694 42910
rect 14758 42846 14764 42910
rect 14552 42774 14764 42846
rect 22168 42840 22380 42976
rect 22576 42916 22788 43052
rect 22478 42910 22788 42916
rect 22440 42846 22446 42910
rect 22510 42846 22788 42910
rect 22478 42840 22788 42846
rect 22984 42840 23196 43188
rect 23392 42840 23604 43188
rect 22304 42780 22380 42840
rect 22984 42780 23060 42840
rect 23528 42780 23604 42840
rect 14552 42710 14694 42774
rect 14758 42710 14764 42774
rect 14552 42704 14764 42710
rect 21760 42774 21972 42780
rect 21760 42710 21766 42774
rect 21830 42710 21972 42774
rect 1632 42532 1844 42644
rect 21760 42638 21972 42710
rect 21760 42574 21766 42638
rect 21830 42574 21972 42638
rect 21760 42568 21972 42574
rect 22168 42704 22788 42780
rect 22168 42644 22380 42704
rect 22168 42638 22516 42644
rect 22168 42574 22446 42638
rect 22510 42574 22516 42638
rect 22168 42568 22516 42574
rect 22576 42638 22788 42704
rect 22576 42574 22718 42638
rect 22782 42574 22788 42638
rect 22576 42568 22788 42574
rect 1632 42508 1702 42532
rect 1224 42502 1702 42508
rect 1224 42438 1230 42502
rect 1294 42476 1702 42502
rect 1758 42476 1844 42532
rect 1294 42438 1844 42476
rect 1224 42432 1844 42438
rect 22984 42432 23196 42780
rect 23392 42432 23604 42780
rect 28288 43182 28636 43324
rect 28288 43118 28294 43182
rect 28358 43118 28636 43182
rect 28288 42910 28636 43118
rect 28288 42846 28294 42910
rect 28358 42846 28566 42910
rect 28630 42846 28636 42910
rect 28288 42774 28636 42846
rect 28288 42710 28294 42774
rect 28358 42710 28636 42774
rect 28288 42704 28636 42710
rect 190128 43182 190340 43324
rect 195024 43248 195236 43390
rect 195160 43188 195236 43248
rect 190128 43118 190134 43182
rect 190198 43118 190270 43182
rect 190334 43118 190340 43182
rect 190128 42910 190340 43118
rect 190128 42846 190270 42910
rect 190334 42846 190340 42910
rect 190128 42774 190340 42846
rect 190128 42710 190270 42774
rect 190334 42710 190340 42774
rect 190128 42704 190340 42710
rect 195024 42840 195236 43188
rect 195432 43454 195644 43460
rect 195432 43390 195574 43454
rect 195638 43390 195644 43454
rect 195432 43248 195644 43390
rect 195840 43248 196052 43596
rect 196112 43520 196460 43596
rect 196248 43318 196460 43520
rect 196248 43254 196390 43318
rect 196454 43254 196460 43318
rect 196248 43248 196460 43254
rect 196656 43248 196868 43596
rect 195432 43188 195508 43248
rect 196792 43188 196868 43248
rect 195432 42840 195644 43188
rect 195840 42916 196052 43052
rect 196248 43046 196460 43052
rect 196248 42982 196390 43046
rect 196454 42982 196460 43046
rect 195840 42840 196188 42916
rect 196248 42840 196460 42982
rect 196656 43046 196868 43188
rect 196656 42982 196662 43046
rect 196726 42982 196868 43046
rect 196656 42976 196868 42982
rect 195024 42780 195100 42840
rect 195568 42780 195644 42840
rect 195976 42780 196052 42840
rect 23120 42372 23196 42432
rect 23528 42372 23604 42432
rect 14144 42265 14356 42372
rect 14144 42236 14212 42265
rect 0 42209 14212 42236
rect 14268 42209 14356 42265
rect 0 42160 14356 42209
rect 21760 42366 21972 42372
rect 21760 42302 21766 42366
rect 21830 42302 21972 42366
rect 21760 42230 21972 42302
rect 15152 42196 15218 42199
rect 15806 42196 15872 42199
rect 15152 42194 15872 42196
rect 15152 42138 15157 42194
rect 15213 42138 15811 42194
rect 15867 42138 15872 42194
rect 21760 42166 21766 42230
rect 21830 42166 21972 42230
rect 21760 42160 21972 42166
rect 15152 42136 15872 42138
rect 15152 42133 15218 42136
rect 15806 42133 15872 42136
rect 22168 42024 22380 42372
rect 22576 42366 22788 42372
rect 22576 42302 22718 42366
rect 22782 42302 22788 42366
rect 22576 42100 22788 42302
rect 22984 42230 23196 42372
rect 22984 42166 23126 42230
rect 23190 42166 23196 42230
rect 22984 42160 23196 42166
rect 23392 42230 23604 42372
rect 23392 42166 23534 42230
rect 23598 42166 23604 42230
rect 23392 42160 23604 42166
rect 28288 42502 28636 42508
rect 28288 42438 28294 42502
rect 28358 42438 28566 42502
rect 28630 42438 28636 42502
rect 28288 42160 28636 42438
rect 190128 42502 190340 42508
rect 190128 42438 190270 42502
rect 190334 42438 190340 42502
rect 190128 42160 190340 42438
rect 195024 42432 195236 42780
rect 195160 42372 195236 42432
rect 195024 42230 195236 42372
rect 195024 42166 195166 42230
rect 195230 42166 195236 42230
rect 195024 42160 195236 42166
rect 195432 42432 195644 42780
rect 195840 42568 196052 42780
rect 196112 42780 196188 42840
rect 196384 42780 196460 42840
rect 196112 42704 196460 42780
rect 196248 42638 196460 42704
rect 196248 42574 196390 42638
rect 196454 42574 196460 42638
rect 196248 42568 196460 42574
rect 196656 42774 196868 42780
rect 196656 42710 196662 42774
rect 196726 42710 196868 42774
rect 196656 42638 196868 42710
rect 196656 42574 196662 42638
rect 196726 42574 196868 42638
rect 196656 42568 196868 42574
rect 216784 42638 217540 42644
rect 216784 42574 217470 42638
rect 217534 42574 217540 42638
rect 216784 42568 217540 42574
rect 216784 42532 216996 42568
rect 216784 42476 216908 42532
rect 216964 42476 216996 42532
rect 216784 42432 216996 42476
rect 195432 42372 195508 42432
rect 195432 42230 195644 42372
rect 195432 42166 195574 42230
rect 195638 42166 195644 42230
rect 195432 42160 195644 42166
rect 22440 42024 22788 42100
rect 28288 42100 28364 42160
rect 190128 42100 190204 42160
rect 22168 41964 22244 42024
rect 22440 41964 22516 42024
rect 21760 41958 21972 41964
rect 21760 41894 21766 41958
rect 21830 41894 21972 41958
rect 21760 41822 21972 41894
rect 21760 41758 21902 41822
rect 21966 41758 21972 41822
rect 21760 41752 21972 41758
rect 22168 41888 22516 41964
rect 22168 41828 22380 41888
rect 22168 41822 22516 41828
rect 22168 41758 22446 41822
rect 22510 41758 22516 41822
rect 22168 41752 22516 41758
rect 22576 41822 22788 41964
rect 22576 41758 22718 41822
rect 22782 41758 22788 41822
rect 22576 41752 22788 41758
rect 22984 41958 23196 41964
rect 22984 41894 23126 41958
rect 23190 41894 23196 41958
rect 22984 41822 23196 41894
rect 22984 41758 22990 41822
rect 23054 41758 23196 41822
rect 22984 41752 23196 41758
rect 23392 41958 23604 41964
rect 23392 41894 23534 41958
rect 23598 41894 23604 41958
rect 23392 41822 23604 41894
rect 28288 41888 28636 42100
rect 28560 41828 28636 41888
rect 23392 41758 23398 41822
rect 23462 41758 23604 41822
rect 23392 41752 23604 41758
rect 14552 41550 14764 41556
rect 14552 41486 14558 41550
rect 14622 41486 14764 41550
rect 14552 41278 14764 41486
rect 21760 41550 21972 41556
rect 21760 41486 21902 41550
rect 21966 41486 21972 41550
rect 21760 41414 21972 41486
rect 21760 41350 21902 41414
rect 21966 41350 21972 41414
rect 21760 41344 21972 41350
rect 22168 41420 22380 41556
rect 22478 41550 22788 41556
rect 22440 41486 22446 41550
rect 22510 41486 22718 41550
rect 22782 41486 22788 41550
rect 22478 41480 22788 41486
rect 22576 41420 22788 41480
rect 22168 41414 22788 41420
rect 22168 41350 22310 41414
rect 22374 41350 22788 41414
rect 22168 41344 22788 41350
rect 22984 41550 23196 41556
rect 22984 41486 22990 41550
rect 23054 41486 23196 41550
rect 22984 41414 23196 41486
rect 22984 41350 23126 41414
rect 23190 41350 23196 41414
rect 22984 41344 23196 41350
rect 23392 41550 23604 41556
rect 23392 41486 23398 41550
rect 23462 41486 23604 41550
rect 23392 41414 23604 41486
rect 23392 41350 23398 41414
rect 23462 41350 23604 41414
rect 23392 41344 23604 41350
rect 28288 41550 28636 41828
rect 28288 41486 28294 41550
rect 28358 41486 28636 41550
rect 28288 41344 28636 41486
rect 190128 41888 190340 42100
rect 195840 42024 196052 42372
rect 196248 42366 196460 42372
rect 196248 42302 196390 42366
rect 196454 42302 196460 42366
rect 196248 42100 196460 42302
rect 196656 42366 196868 42372
rect 196656 42302 196662 42366
rect 196726 42302 196868 42366
rect 196656 42230 196868 42302
rect 196656 42166 196662 42230
rect 196726 42166 196868 42230
rect 196656 42160 196868 42166
rect 195976 41964 196052 42024
rect 196112 42024 196460 42100
rect 196112 41964 196188 42024
rect 196384 41964 196460 42024
rect 195024 41958 195236 41964
rect 195024 41894 195166 41958
rect 195230 41894 195236 41958
rect 190128 41828 190204 41888
rect 190128 41550 190340 41828
rect 195024 41822 195236 41894
rect 195024 41758 195030 41822
rect 195094 41758 195236 41822
rect 195024 41752 195236 41758
rect 195432 41958 195644 41964
rect 195432 41894 195574 41958
rect 195638 41894 195644 41958
rect 195432 41822 195644 41894
rect 195432 41758 195438 41822
rect 195502 41758 195644 41822
rect 195432 41752 195644 41758
rect 195840 41888 196188 41964
rect 195840 41752 196052 41888
rect 196248 41752 196460 41964
rect 196656 41958 196868 41964
rect 196656 41894 196662 41958
rect 196726 41894 196868 41958
rect 196656 41822 196868 41894
rect 196656 41758 196798 41822
rect 196862 41758 196868 41822
rect 196656 41752 196868 41758
rect 196248 41692 196324 41752
rect 195976 41616 196324 41692
rect 195976 41556 196052 41616
rect 190128 41486 190134 41550
rect 190198 41486 190340 41550
rect 190128 41344 190340 41486
rect 195024 41550 195236 41556
rect 195024 41486 195030 41550
rect 195094 41486 195236 41550
rect 195024 41414 195236 41486
rect 195024 41350 195166 41414
rect 195230 41350 195236 41414
rect 195024 41344 195236 41350
rect 195432 41550 195644 41556
rect 195432 41486 195438 41550
rect 195502 41486 195644 41550
rect 195432 41414 195644 41486
rect 195432 41350 195574 41414
rect 195638 41350 195644 41414
rect 195432 41344 195644 41350
rect 195840 41480 196460 41556
rect 195840 41414 196052 41480
rect 195840 41350 195846 41414
rect 195910 41350 196052 41414
rect 195840 41344 196052 41350
rect 196248 41414 196460 41480
rect 196248 41350 196390 41414
rect 196454 41350 196460 41414
rect 196248 41344 196460 41350
rect 196656 41550 196868 41556
rect 196656 41486 196798 41550
rect 196862 41486 196868 41550
rect 196656 41414 196868 41486
rect 196656 41350 196798 41414
rect 196862 41350 196868 41414
rect 196656 41344 196868 41350
rect 14552 41214 14558 41278
rect 14622 41214 14764 41278
rect 14552 41208 14764 41214
rect 22304 41284 22380 41344
rect 28288 41284 28364 41344
rect 190128 41284 190204 41344
rect 22304 41208 22652 41284
rect 22576 41148 22652 41208
rect 28288 41278 28636 41284
rect 28288 41214 28294 41278
rect 28358 41214 28636 41278
rect 21760 41142 21972 41148
rect 21760 41078 21902 41142
rect 21966 41078 21972 41142
rect 21760 41006 21972 41078
rect 21760 40942 21902 41006
rect 21966 40942 21972 41006
rect 21760 40936 21972 40942
rect 22168 41142 22380 41148
rect 22168 41078 22310 41142
rect 22374 41078 22380 41142
rect 22168 40936 22380 41078
rect 22576 41006 22788 41148
rect 22576 40942 22582 41006
rect 22646 40942 22788 41006
rect 22576 40936 22788 40942
rect 22984 41142 23196 41148
rect 22984 41078 23126 41142
rect 23190 41078 23196 41142
rect 22984 41006 23196 41078
rect 22984 40942 22990 41006
rect 23054 40942 23196 41006
rect 22984 40936 23196 40942
rect 23392 41142 23604 41148
rect 23392 41078 23398 41142
rect 23462 41078 23604 41142
rect 23392 41006 23604 41078
rect 23392 40942 23534 41006
rect 23598 40942 23604 41006
rect 23392 40936 23604 40942
rect 28288 41072 28636 41214
rect 190128 41278 190340 41284
rect 190128 41214 190134 41278
rect 190198 41214 190340 41278
rect 190128 41072 190340 41214
rect 195024 41142 195236 41148
rect 195024 41078 195166 41142
rect 195230 41078 195236 41142
rect 28288 41012 28364 41072
rect 190128 41012 190204 41072
rect 1224 40870 1844 40876
rect 1224 40806 1230 40870
rect 1294 40852 1844 40870
rect 1294 40806 1702 40852
rect 1224 40800 1702 40806
rect 1681 40796 1702 40800
rect 1758 40800 1844 40852
rect 28288 40800 28636 41012
rect 190128 40800 190340 41012
rect 195024 41006 195236 41078
rect 195024 40942 195166 41006
rect 195230 40942 195236 41006
rect 195024 40936 195236 40942
rect 195432 41142 195644 41148
rect 195432 41078 195574 41142
rect 195638 41078 195644 41142
rect 195432 41006 195644 41078
rect 195432 40942 195438 41006
rect 195502 40942 195644 41006
rect 195432 40936 195644 40942
rect 195840 41142 196052 41148
rect 195840 41078 195846 41142
rect 195910 41078 196052 41142
rect 195840 40936 196052 41078
rect 196248 41142 196460 41148
rect 196248 41078 196390 41142
rect 196454 41078 196460 41142
rect 196248 40936 196460 41078
rect 196656 41142 196868 41148
rect 196656 41078 196798 41142
rect 196862 41078 196868 41142
rect 196656 41006 196868 41078
rect 196656 40942 196662 41006
rect 196726 40942 196868 41006
rect 196656 40936 196868 40942
rect 196248 40876 196324 40936
rect 195976 40800 196324 40876
rect 216784 40870 217540 40876
rect 216784 40852 217470 40870
rect 1758 40796 1779 40800
rect 1681 40775 1779 40796
rect 28424 40740 28500 40800
rect 190128 40740 190204 40800
rect 195976 40740 196052 40800
rect 216784 40796 216908 40852
rect 216964 40806 217470 40852
rect 217534 40806 217540 40870
rect 216964 40800 217540 40806
rect 216964 40796 216996 40800
rect 21760 40734 21972 40740
rect 21760 40670 21902 40734
rect 21966 40670 21972 40734
rect 15152 40638 15218 40641
rect 15726 40638 15792 40641
rect 15152 40636 15792 40638
rect 0 40565 14356 40604
rect 15152 40580 15157 40636
rect 15213 40580 15731 40636
rect 15787 40580 15792 40636
rect 15152 40578 15792 40580
rect 15152 40575 15218 40578
rect 15726 40575 15792 40578
rect 21760 40598 21972 40670
rect 0 40528 14212 40565
rect 14144 40509 14212 40528
rect 14268 40509 14356 40565
rect 21760 40534 21902 40598
rect 21966 40534 21972 40598
rect 21760 40528 21972 40534
rect 22168 40604 22380 40740
rect 22576 40734 22788 40740
rect 22576 40670 22582 40734
rect 22646 40670 22788 40734
rect 22576 40604 22788 40670
rect 22168 40598 22788 40604
rect 22168 40534 22310 40598
rect 22374 40534 22788 40598
rect 22168 40528 22788 40534
rect 22984 40734 23196 40740
rect 22984 40670 22990 40734
rect 23054 40670 23196 40734
rect 22984 40598 23196 40670
rect 22984 40534 23126 40598
rect 23190 40534 23196 40598
rect 22984 40528 23196 40534
rect 23392 40734 23604 40740
rect 23392 40670 23534 40734
rect 23598 40670 23604 40734
rect 23392 40598 23604 40670
rect 23392 40534 23398 40598
rect 23462 40534 23604 40598
rect 23392 40528 23604 40534
rect 28288 40528 28636 40740
rect 190128 40528 190340 40740
rect 195024 40734 195236 40740
rect 195024 40670 195166 40734
rect 195230 40670 195236 40734
rect 195024 40598 195236 40670
rect 195024 40534 195030 40598
rect 195094 40534 195236 40598
rect 195024 40528 195236 40534
rect 195432 40734 195644 40740
rect 195432 40670 195438 40734
rect 195502 40670 195644 40734
rect 195432 40598 195644 40670
rect 195432 40534 195438 40598
rect 195502 40534 195644 40598
rect 195432 40528 195644 40534
rect 195840 40664 196460 40740
rect 195840 40528 196052 40664
rect 196248 40598 196460 40664
rect 196248 40534 196390 40598
rect 196454 40534 196460 40598
rect 196248 40528 196460 40534
rect 196656 40734 196868 40740
rect 196656 40670 196662 40734
rect 196726 40670 196868 40734
rect 196656 40598 196868 40670
rect 216784 40664 216996 40796
rect 196656 40534 196798 40598
rect 196862 40534 196868 40598
rect 196656 40528 196868 40534
rect 14144 40392 14356 40509
rect 22304 40468 22380 40528
rect 28288 40468 28364 40528
rect 190264 40468 190340 40528
rect 22304 40392 22652 40468
rect 22576 40332 22652 40392
rect 21760 40326 21972 40332
rect 21760 40262 21902 40326
rect 21966 40262 21972 40326
rect 21760 40120 21972 40262
rect 22168 40326 22380 40332
rect 22168 40262 22310 40326
rect 22374 40262 22380 40326
rect 22168 40196 22380 40262
rect 22168 40190 22516 40196
rect 22168 40126 22174 40190
rect 22238 40126 22446 40190
rect 22510 40126 22516 40190
rect 22168 40120 22516 40126
rect 22576 40120 22788 40332
rect 22984 40326 23196 40332
rect 22984 40262 23126 40326
rect 23190 40262 23196 40326
rect 22984 40190 23196 40262
rect 22984 40126 22990 40190
rect 23054 40126 23196 40190
rect 22984 40120 23196 40126
rect 23392 40326 23604 40332
rect 23392 40262 23398 40326
rect 23462 40262 23604 40326
rect 23392 40190 23604 40262
rect 28288 40256 28636 40468
rect 28560 40196 28636 40256
rect 23392 40126 23534 40190
rect 23598 40126 23604 40190
rect 23392 40120 23604 40126
rect 21760 40060 21836 40120
rect 14552 40054 14764 40060
rect 14552 39990 14694 40054
rect 14758 39990 14764 40054
rect 14552 39918 14764 39990
rect 14552 39854 14694 39918
rect 14758 39854 14764 39918
rect 14552 39848 14764 39854
rect 21760 39712 21972 40060
rect 28288 40054 28636 40196
rect 28288 39990 28294 40054
rect 28358 39990 28636 40054
rect 28288 39984 28636 39990
rect 190128 40256 190340 40468
rect 195024 40326 195236 40332
rect 195024 40262 195030 40326
rect 195094 40262 195236 40326
rect 190128 40196 190204 40256
rect 190128 40054 190340 40196
rect 195024 40190 195236 40262
rect 195024 40126 195166 40190
rect 195230 40126 195236 40190
rect 195024 40120 195236 40126
rect 195432 40326 195644 40332
rect 195432 40262 195438 40326
rect 195502 40262 195644 40326
rect 195432 40190 195644 40262
rect 195432 40126 195574 40190
rect 195638 40126 195644 40190
rect 195432 40120 195644 40126
rect 195840 40190 196052 40332
rect 195840 40126 195846 40190
rect 195910 40126 196052 40190
rect 195840 40120 196052 40126
rect 196248 40326 196460 40332
rect 196248 40262 196390 40326
rect 196454 40262 196460 40326
rect 196248 40190 196460 40262
rect 196248 40126 196254 40190
rect 196318 40126 196460 40190
rect 196248 40120 196460 40126
rect 196656 40326 196868 40332
rect 196656 40262 196798 40326
rect 196862 40262 196868 40326
rect 196656 40120 196868 40262
rect 190128 39990 190134 40054
rect 190198 39990 190340 40054
rect 190128 39984 190340 39990
rect 196656 40060 196732 40120
rect 28424 39924 28500 39984
rect 190128 39924 190204 39984
rect 21896 39652 21972 39712
rect 0 39440 14356 39516
rect 14144 39437 14356 39440
rect 14144 39381 14212 39437
rect 14268 39381 14356 39437
rect 14144 39304 14356 39381
rect 15152 39368 15218 39371
rect 15646 39368 15712 39371
rect 15152 39366 15712 39368
rect 15152 39310 15157 39366
rect 15213 39310 15651 39366
rect 15707 39310 15712 39366
rect 15152 39308 15712 39310
rect 15152 39305 15218 39308
rect 15646 39305 15712 39308
rect 21760 39304 21972 39652
rect 22168 39918 22380 39924
rect 22478 39918 22788 39924
rect 22168 39854 22174 39918
rect 22238 39854 22380 39918
rect 22440 39854 22446 39918
rect 22510 39854 22788 39918
rect 22168 39712 22380 39854
rect 22478 39848 22788 39854
rect 22576 39712 22788 39848
rect 22984 39918 23196 39924
rect 22984 39854 22990 39918
rect 23054 39854 23196 39918
rect 22984 39782 23196 39854
rect 22984 39718 22990 39782
rect 23054 39718 23196 39782
rect 22984 39712 23196 39718
rect 23392 39918 23604 39924
rect 23392 39854 23534 39918
rect 23598 39854 23604 39918
rect 23392 39782 23604 39854
rect 23392 39718 23398 39782
rect 23462 39718 23604 39782
rect 23392 39712 23604 39718
rect 28288 39782 28636 39924
rect 28288 39718 28294 39782
rect 28358 39718 28636 39782
rect 22168 39652 22244 39712
rect 22576 39652 22652 39712
rect 22168 39380 22380 39652
rect 22168 39374 22516 39380
rect 22168 39310 22174 39374
rect 22238 39310 22446 39374
rect 22510 39310 22516 39374
rect 22168 39304 22516 39310
rect 22576 39304 22788 39652
rect 22984 39510 23196 39516
rect 22984 39446 22990 39510
rect 23054 39446 23196 39510
rect 22984 39374 23196 39446
rect 22984 39310 22990 39374
rect 23054 39310 23196 39374
rect 22984 39304 23196 39310
rect 23392 39510 23604 39516
rect 23392 39446 23398 39510
rect 23462 39446 23604 39510
rect 23392 39374 23604 39446
rect 28288 39440 28636 39718
rect 190128 39782 190340 39924
rect 190128 39718 190134 39782
rect 190198 39718 190340 39782
rect 190128 39440 190340 39718
rect 195024 39918 195236 39924
rect 195024 39854 195166 39918
rect 195230 39854 195236 39918
rect 195024 39782 195236 39854
rect 195024 39718 195166 39782
rect 195230 39718 195236 39782
rect 195024 39712 195236 39718
rect 195432 39918 195644 39924
rect 195432 39854 195574 39918
rect 195638 39854 195644 39918
rect 195432 39782 195644 39854
rect 195432 39718 195574 39782
rect 195638 39718 195644 39782
rect 195432 39712 195644 39718
rect 195840 39918 196052 39924
rect 195840 39854 195846 39918
rect 195910 39854 196052 39918
rect 195840 39712 196052 39854
rect 196248 39918 196460 39924
rect 196248 39854 196254 39918
rect 196318 39854 196460 39918
rect 196248 39788 196460 39854
rect 196112 39712 196460 39788
rect 196656 39712 196868 40060
rect 195840 39652 195916 39712
rect 196112 39652 196188 39712
rect 195840 39576 196188 39652
rect 196248 39652 196324 39712
rect 196656 39652 196732 39712
rect 28424 39380 28500 39440
rect 190264 39380 190340 39440
rect 23392 39310 23398 39374
rect 23462 39310 23604 39374
rect 23392 39304 23604 39310
rect 21896 39244 21972 39304
rect 1224 39238 1844 39244
rect 1224 39174 1230 39238
rect 1294 39174 1844 39238
rect 1224 39172 1844 39174
rect 1224 39168 1702 39172
rect 1632 39116 1702 39168
rect 1758 39116 1844 39172
rect 1632 39032 1844 39116
rect 21760 39102 21972 39244
rect 28288 39168 28636 39380
rect 190128 39168 190340 39380
rect 195024 39510 195236 39516
rect 195024 39446 195166 39510
rect 195230 39446 195236 39510
rect 195024 39374 195236 39446
rect 195024 39310 195166 39374
rect 195230 39310 195236 39374
rect 195024 39304 195236 39310
rect 195432 39510 195644 39516
rect 195432 39446 195574 39510
rect 195638 39446 195644 39510
rect 195432 39374 195644 39446
rect 195432 39310 195438 39374
rect 195502 39310 195644 39374
rect 195432 39304 195644 39310
rect 195840 39304 196052 39576
rect 196248 39374 196460 39652
rect 196248 39310 196254 39374
rect 196318 39310 196460 39374
rect 196248 39304 196460 39310
rect 196656 39304 196868 39652
rect 196656 39244 196732 39304
rect 28424 39108 28500 39168
rect 190128 39108 190204 39168
rect 21760 39038 21766 39102
rect 21830 39038 21972 39102
rect 21760 39032 21972 39038
rect 22168 39102 22380 39108
rect 22478 39102 22788 39108
rect 22168 39038 22174 39102
rect 22238 39038 22380 39102
rect 22440 39038 22446 39102
rect 22510 39038 22788 39102
rect 22168 38896 22380 39038
rect 22478 39032 22788 39038
rect 22576 38896 22788 39032
rect 22984 39102 23196 39108
rect 22984 39038 22990 39102
rect 23054 39038 23196 39102
rect 22984 38896 23196 39038
rect 23392 39102 23604 39108
rect 23392 39038 23398 39102
rect 23462 39038 23604 39102
rect 23392 38896 23604 39038
rect 22168 38836 22244 38896
rect 22576 38836 22652 38896
rect 22984 38836 23060 38896
rect 23528 38836 23604 38896
rect 21760 38830 21972 38836
rect 21760 38766 21766 38830
rect 21830 38766 21972 38830
rect 14552 38694 14764 38700
rect 14552 38630 14558 38694
rect 14622 38630 14764 38694
rect 14552 38558 14764 38630
rect 21760 38694 21972 38766
rect 21760 38630 21902 38694
rect 21966 38630 21972 38694
rect 21760 38624 21972 38630
rect 22168 38624 22380 38836
rect 22576 38694 22788 38836
rect 22576 38630 22582 38694
rect 22646 38630 22788 38694
rect 22576 38624 22788 38630
rect 14552 38494 14558 38558
rect 14622 38494 14764 38558
rect 14552 38488 14764 38494
rect 22984 38488 23196 38836
rect 23120 38428 23196 38488
rect 21760 38422 21972 38428
rect 21760 38358 21902 38422
rect 21966 38358 21972 38422
rect 21760 38286 21972 38358
rect 21760 38222 21902 38286
rect 21966 38222 21972 38286
rect 21760 38216 21972 38222
rect 22168 38422 22788 38428
rect 22168 38358 22582 38422
rect 22646 38358 22788 38422
rect 22168 38352 22788 38358
rect 22168 38156 22380 38352
rect 22168 38080 22516 38156
rect 22576 38080 22788 38352
rect 22984 38286 23196 38428
rect 22984 38222 22990 38286
rect 23054 38222 23196 38286
rect 22984 38216 23196 38222
rect 23392 38488 23604 38836
rect 28288 38830 28636 39108
rect 28288 38766 28294 38830
rect 28358 38766 28636 38830
rect 28288 38760 28636 38766
rect 190128 38966 190340 39108
rect 190128 38902 190134 38966
rect 190198 38902 190340 38966
rect 190128 38830 190340 38902
rect 195024 39102 195236 39108
rect 195024 39038 195166 39102
rect 195230 39038 195236 39102
rect 195024 38896 195236 39038
rect 195160 38836 195236 38896
rect 190128 38766 190270 38830
rect 190334 38766 190340 38830
rect 190128 38760 190340 38766
rect 28288 38558 28636 38564
rect 28288 38494 28294 38558
rect 28358 38494 28636 38558
rect 23392 38428 23468 38488
rect 23392 38286 23604 38428
rect 23392 38222 23398 38286
rect 23462 38222 23604 38286
rect 23392 38216 23604 38222
rect 28288 38216 28636 38494
rect 190128 38558 190340 38564
rect 190128 38494 190134 38558
rect 190198 38494 190270 38558
rect 190334 38494 190340 38558
rect 190128 38216 190340 38494
rect 195024 38488 195236 38836
rect 195432 39102 195644 39108
rect 195432 39038 195438 39102
rect 195502 39038 195644 39102
rect 195432 38896 195644 39038
rect 195840 38972 196052 39108
rect 196248 39102 196460 39108
rect 196248 39038 196254 39102
rect 196318 39038 196460 39102
rect 195840 38896 196188 38972
rect 195432 38836 195508 38896
rect 195840 38836 195916 38896
rect 196112 38836 196188 38896
rect 196248 38896 196460 39038
rect 196656 39102 196868 39244
rect 196656 39038 196662 39102
rect 196726 39038 196868 39102
rect 196656 39032 196868 39038
rect 216784 39172 216996 39244
rect 216784 39116 216908 39172
rect 216964 39116 216996 39172
rect 216784 39108 216996 39116
rect 216784 39102 217540 39108
rect 216784 39038 217470 39102
rect 217534 39038 217540 39102
rect 216784 39032 217540 39038
rect 196248 38836 196324 38896
rect 195432 38488 195644 38836
rect 195840 38694 196052 38836
rect 196112 38760 196460 38836
rect 195840 38630 195846 38694
rect 195910 38630 196052 38694
rect 195840 38624 196052 38630
rect 196248 38624 196460 38760
rect 196656 38830 196868 38836
rect 196656 38766 196662 38830
rect 196726 38766 196868 38830
rect 196656 38694 196868 38766
rect 196656 38630 196662 38694
rect 196726 38630 196868 38694
rect 196656 38624 196868 38630
rect 195024 38428 195100 38488
rect 195568 38428 195644 38488
rect 195024 38286 195236 38428
rect 195024 38222 195166 38286
rect 195230 38222 195236 38286
rect 195024 38216 195236 38222
rect 195432 38286 195644 38428
rect 195432 38222 195438 38286
rect 195502 38222 195644 38286
rect 195432 38216 195644 38222
rect 195840 38422 196052 38428
rect 195840 38358 195846 38422
rect 195910 38358 196052 38422
rect 28424 38156 28500 38216
rect 190264 38156 190340 38216
rect 22168 38020 22244 38080
rect 22440 38020 22516 38080
rect 21760 38014 21972 38020
rect 21760 37950 21902 38014
rect 21966 37950 21972 38014
rect 0 37808 14356 37884
rect 21760 37878 21972 37950
rect 21760 37814 21766 37878
rect 21830 37814 21972 37878
rect 14144 37737 14356 37808
rect 15152 37810 15218 37813
rect 15566 37810 15632 37813
rect 15152 37808 15632 37810
rect 21760 37808 21972 37814
rect 22168 37878 22380 38020
rect 22440 37944 22788 38020
rect 22168 37814 22174 37878
rect 22238 37814 22380 37878
rect 22168 37808 22380 37814
rect 22576 37878 22788 37944
rect 22576 37814 22582 37878
rect 22646 37814 22788 37878
rect 22576 37808 22788 37814
rect 22984 38014 23196 38020
rect 22984 37950 22990 38014
rect 23054 37950 23196 38014
rect 22984 37878 23196 37950
rect 22984 37814 22990 37878
rect 23054 37814 23196 37878
rect 22984 37808 23196 37814
rect 23392 38014 23604 38020
rect 23392 37950 23398 38014
rect 23462 37950 23604 38014
rect 23392 37878 23604 37950
rect 23392 37814 23534 37878
rect 23598 37814 23604 37878
rect 23392 37808 23604 37814
rect 28288 37944 28636 38156
rect 190128 37944 190340 38156
rect 195840 38156 196052 38358
rect 196248 38156 196460 38428
rect 196656 38422 196868 38428
rect 196656 38358 196662 38422
rect 196726 38358 196868 38422
rect 196656 38286 196868 38358
rect 196656 38222 196798 38286
rect 196862 38222 196868 38286
rect 196656 38216 196868 38222
rect 195840 38080 196460 38156
rect 195976 38020 196052 38080
rect 195024 38014 195236 38020
rect 195024 37950 195166 38014
rect 195230 37950 195236 38014
rect 28288 37884 28364 37944
rect 190128 37884 190204 37944
rect 15152 37752 15157 37808
rect 15213 37752 15571 37808
rect 15627 37752 15632 37808
rect 15152 37750 15632 37752
rect 15152 37747 15218 37750
rect 15566 37747 15632 37750
rect 14144 37681 14212 37737
rect 14268 37681 14356 37737
rect 1632 37492 1844 37612
rect 14144 37536 14356 37681
rect 21760 37606 21972 37612
rect 21760 37542 21766 37606
rect 21830 37542 21972 37606
rect 1632 37476 1702 37492
rect 1224 37470 1702 37476
rect 1224 37406 1230 37470
rect 1294 37436 1702 37470
rect 1758 37436 1844 37492
rect 1294 37406 1844 37436
rect 1224 37400 1844 37406
rect 21760 37470 21972 37542
rect 21760 37406 21902 37470
rect 21966 37406 21972 37470
rect 21760 37400 21972 37406
rect 22168 37606 22380 37612
rect 22168 37542 22174 37606
rect 22238 37542 22380 37606
rect 22168 37400 22380 37542
rect 22576 37606 22788 37612
rect 22576 37542 22582 37606
rect 22646 37542 22788 37606
rect 22576 37470 22788 37542
rect 22576 37406 22718 37470
rect 22782 37406 22788 37470
rect 22576 37400 22788 37406
rect 22984 37606 23196 37612
rect 22984 37542 22990 37606
rect 23054 37542 23196 37606
rect 22984 37470 23196 37542
rect 22984 37406 22990 37470
rect 23054 37406 23196 37470
rect 22984 37400 23196 37406
rect 23392 37606 23604 37612
rect 23392 37542 23534 37606
rect 23598 37542 23604 37606
rect 23392 37470 23604 37542
rect 23392 37406 23398 37470
rect 23462 37406 23604 37470
rect 23392 37400 23604 37406
rect 28288 37400 28636 37884
rect 190128 37606 190340 37884
rect 195024 37878 195236 37950
rect 195024 37814 195166 37878
rect 195230 37814 195236 37878
rect 195024 37808 195236 37814
rect 195432 38014 195644 38020
rect 195432 37950 195438 38014
rect 195502 37950 195644 38014
rect 195432 37878 195644 37950
rect 195432 37814 195438 37878
rect 195502 37814 195644 37878
rect 195432 37808 195644 37814
rect 195840 37808 196052 38020
rect 196248 38020 196324 38080
rect 196248 37878 196460 38020
rect 196248 37814 196254 37878
rect 196318 37814 196460 37878
rect 196248 37808 196460 37814
rect 196656 38014 196868 38020
rect 196656 37950 196798 38014
rect 196862 37950 196868 38014
rect 196656 37878 196868 37950
rect 196656 37814 196662 37878
rect 196726 37814 196868 37878
rect 196656 37808 196868 37814
rect 190128 37542 190134 37606
rect 190198 37542 190340 37606
rect 190128 37400 190340 37542
rect 195024 37606 195236 37612
rect 195024 37542 195166 37606
rect 195230 37542 195236 37606
rect 195024 37470 195236 37542
rect 195024 37406 195030 37470
rect 195094 37406 195236 37470
rect 195024 37400 195236 37406
rect 195432 37606 195644 37612
rect 195432 37542 195438 37606
rect 195502 37542 195644 37606
rect 195432 37470 195644 37542
rect 195432 37406 195574 37470
rect 195638 37406 195644 37470
rect 195432 37400 195644 37406
rect 195840 37476 196052 37612
rect 196248 37606 196460 37612
rect 196248 37542 196254 37606
rect 196318 37542 196460 37606
rect 196248 37476 196460 37542
rect 195840 37400 196460 37476
rect 196656 37606 196868 37612
rect 196656 37542 196662 37606
rect 196726 37542 196868 37606
rect 196656 37470 196868 37542
rect 196656 37406 196798 37470
rect 196862 37406 196868 37470
rect 196656 37400 196868 37406
rect 216784 37606 217540 37612
rect 216784 37542 217470 37606
rect 217534 37542 217540 37606
rect 216784 37536 217540 37542
rect 216784 37492 216996 37536
rect 216784 37436 216908 37492
rect 216964 37436 216996 37492
rect 216784 37400 216996 37436
rect 28424 37340 28500 37400
rect 190264 37340 190340 37400
rect 14552 37198 14764 37204
rect 14552 37134 14694 37198
rect 14758 37134 14764 37198
rect 14552 37062 14764 37134
rect 14552 36998 14694 37062
rect 14758 36998 14764 37062
rect 14552 36992 14764 36998
rect 21760 37198 21972 37204
rect 21760 37134 21902 37198
rect 21966 37134 21972 37198
rect 21760 37062 21972 37134
rect 21760 36998 21902 37062
rect 21966 36998 21972 37062
rect 21760 36992 21972 36998
rect 22168 37068 22380 37204
rect 22576 37198 22788 37204
rect 22576 37134 22718 37198
rect 22782 37134 22788 37198
rect 22576 37068 22788 37134
rect 22168 37062 22788 37068
rect 22168 36998 22310 37062
rect 22374 36998 22788 37062
rect 22168 36992 22788 36998
rect 22984 37198 23196 37204
rect 22984 37134 22990 37198
rect 23054 37134 23196 37198
rect 22984 37062 23196 37134
rect 22984 36998 22990 37062
rect 23054 36998 23196 37062
rect 22984 36992 23196 36998
rect 23392 37198 23604 37204
rect 23392 37134 23398 37198
rect 23462 37134 23604 37198
rect 23392 37062 23604 37134
rect 28288 37128 28636 37340
rect 190128 37334 190340 37340
rect 190128 37270 190134 37334
rect 190198 37270 190340 37334
rect 190128 37128 190340 37270
rect 195976 37340 196052 37400
rect 195976 37264 196324 37340
rect 196248 37204 196324 37264
rect 28560 37068 28636 37128
rect 190264 37068 190340 37128
rect 23392 36998 23534 37062
rect 23598 36998 23604 37062
rect 23392 36992 23604 36998
rect 22304 36932 22380 36992
rect 22304 36856 22652 36932
rect 22576 36796 22652 36856
rect 28288 36856 28636 37068
rect 190128 36856 190340 37068
rect 195024 37198 195236 37204
rect 195024 37134 195030 37198
rect 195094 37134 195236 37198
rect 195024 37062 195236 37134
rect 195024 36998 195166 37062
rect 195230 36998 195236 37062
rect 195024 36992 195236 36998
rect 195432 37198 195644 37204
rect 195432 37134 195574 37198
rect 195638 37134 195644 37198
rect 195432 37062 195644 37134
rect 195432 36998 195574 37062
rect 195638 36998 195644 37062
rect 195432 36992 195644 36998
rect 195840 37128 196460 37204
rect 195840 36992 196052 37128
rect 196248 36992 196460 37128
rect 196656 37198 196868 37204
rect 196656 37134 196798 37198
rect 196862 37134 196868 37198
rect 196656 37062 196868 37134
rect 196656 36998 196798 37062
rect 196862 36998 196868 37062
rect 196656 36992 196868 36998
rect 196248 36932 196324 36992
rect 195976 36856 196324 36932
rect 28288 36796 28364 36856
rect 190128 36796 190204 36856
rect 195976 36796 196052 36856
rect 21760 36790 21972 36796
rect 21760 36726 21902 36790
rect 21966 36726 21972 36790
rect 14144 36609 14356 36660
rect 14144 36553 14212 36609
rect 14268 36553 14356 36609
rect 21760 36654 21972 36726
rect 21760 36590 21902 36654
rect 21966 36590 21972 36654
rect 21760 36584 21972 36590
rect 22168 36790 22380 36796
rect 22168 36726 22310 36790
rect 22374 36726 22380 36790
rect 22168 36584 22380 36726
rect 22576 36654 22788 36796
rect 22576 36590 22582 36654
rect 22646 36590 22788 36654
rect 22576 36584 22788 36590
rect 22984 36790 23196 36796
rect 22984 36726 22990 36790
rect 23054 36726 23196 36790
rect 22984 36654 23196 36726
rect 22984 36590 22990 36654
rect 23054 36590 23196 36654
rect 22984 36584 23196 36590
rect 23392 36790 23604 36796
rect 23392 36726 23534 36790
rect 23598 36726 23604 36790
rect 23392 36654 23604 36726
rect 23392 36590 23534 36654
rect 23598 36590 23604 36654
rect 23392 36584 23604 36590
rect 28288 36584 28636 36796
rect 190128 36584 190340 36796
rect 195024 36790 195236 36796
rect 195024 36726 195166 36790
rect 195230 36726 195236 36790
rect 195024 36654 195236 36726
rect 195024 36590 195166 36654
rect 195230 36590 195236 36654
rect 195024 36584 195236 36590
rect 195432 36790 195644 36796
rect 195432 36726 195574 36790
rect 195638 36726 195644 36790
rect 195432 36654 195644 36726
rect 195432 36590 195438 36654
rect 195502 36590 195644 36654
rect 195432 36584 195644 36590
rect 195840 36720 196460 36796
rect 195840 36584 196052 36720
rect 196248 36584 196460 36720
rect 196656 36790 196868 36796
rect 196656 36726 196798 36790
rect 196862 36726 196868 36790
rect 196656 36654 196868 36726
rect 196656 36590 196798 36654
rect 196862 36590 196868 36654
rect 196656 36584 196868 36590
rect 14144 36524 14356 36553
rect 0 36448 14356 36524
rect 15152 36540 15218 36543
rect 15486 36540 15552 36543
rect 15152 36538 15552 36540
rect 15152 36482 15157 36538
rect 15213 36482 15491 36538
rect 15547 36482 15552 36538
rect 28424 36524 28500 36584
rect 190128 36524 190204 36584
rect 196248 36524 196324 36584
rect 15152 36480 15552 36482
rect 15152 36477 15218 36480
rect 15486 36477 15552 36480
rect 21760 36382 21972 36388
rect 21760 36318 21902 36382
rect 21966 36318 21972 36382
rect 21760 36176 21972 36318
rect 22168 36252 22380 36388
rect 22576 36382 22788 36388
rect 22576 36318 22582 36382
rect 22646 36318 22788 36382
rect 22168 36246 22516 36252
rect 22168 36182 22446 36246
rect 22510 36182 22516 36246
rect 22168 36176 22516 36182
rect 22576 36246 22788 36318
rect 22576 36182 22718 36246
rect 22782 36182 22788 36246
rect 22576 36176 22788 36182
rect 22984 36382 23196 36388
rect 22984 36318 22990 36382
rect 23054 36318 23196 36382
rect 22984 36246 23196 36318
rect 22984 36182 23126 36246
rect 23190 36182 23196 36246
rect 22984 36176 23196 36182
rect 23392 36382 23604 36388
rect 23392 36318 23534 36382
rect 23598 36318 23604 36382
rect 23392 36246 23604 36318
rect 28288 36312 28636 36524
rect 190128 36312 190340 36524
rect 195976 36448 196324 36524
rect 195976 36388 196052 36448
rect 28424 36252 28500 36312
rect 190264 36252 190340 36312
rect 23392 36182 23398 36246
rect 23462 36182 23604 36246
rect 23392 36176 23604 36182
rect 21896 36116 21972 36176
rect 1632 35812 1844 35844
rect 1632 35756 1702 35812
rect 1758 35756 1844 35812
rect 1632 35708 1844 35756
rect 1224 35702 1844 35708
rect 1224 35638 1230 35702
rect 1294 35638 1844 35702
rect 1224 35632 1844 35638
rect 14552 35838 14764 35844
rect 14552 35774 14558 35838
rect 14622 35774 14764 35838
rect 14552 35708 14764 35774
rect 21760 35768 21972 36116
rect 28288 36110 28636 36252
rect 28288 36046 28294 36110
rect 28358 36046 28636 36110
rect 28288 36040 28636 36046
rect 190128 36040 190340 36252
rect 195024 36382 195236 36388
rect 195024 36318 195166 36382
rect 195230 36318 195236 36382
rect 195024 36246 195236 36318
rect 195024 36182 195030 36246
rect 195094 36182 195236 36246
rect 195024 36176 195236 36182
rect 195432 36382 195644 36388
rect 195432 36318 195438 36382
rect 195502 36318 195644 36382
rect 195432 36246 195644 36318
rect 195432 36182 195438 36246
rect 195502 36182 195644 36246
rect 195432 36176 195644 36182
rect 195840 36312 196460 36388
rect 195840 36176 196052 36312
rect 196248 36246 196460 36312
rect 196248 36182 196390 36246
rect 196454 36182 196460 36246
rect 196248 36176 196460 36182
rect 196656 36382 196868 36388
rect 196656 36318 196798 36382
rect 196862 36318 196868 36382
rect 196656 36176 196868 36318
rect 196792 36116 196868 36176
rect 28288 35980 28364 36040
rect 190264 35980 190340 36040
rect 21896 35708 21972 35768
rect 14552 35702 18572 35708
rect 14552 35638 18502 35702
rect 18566 35638 18572 35702
rect 14552 35632 18572 35638
rect 21760 35360 21972 35708
rect 22168 35768 22380 35980
rect 22478 35974 22788 35980
rect 22440 35910 22446 35974
rect 22510 35910 22718 35974
rect 22782 35910 22788 35974
rect 22478 35904 22788 35910
rect 22576 35768 22788 35904
rect 22984 35974 23196 35980
rect 22984 35910 23126 35974
rect 23190 35910 23196 35974
rect 22984 35838 23196 35910
rect 22984 35774 22990 35838
rect 23054 35774 23196 35838
rect 22984 35768 23196 35774
rect 23392 35974 23604 35980
rect 23392 35910 23398 35974
rect 23462 35910 23604 35974
rect 23392 35838 23604 35910
rect 23392 35774 23534 35838
rect 23598 35774 23604 35838
rect 23392 35768 23604 35774
rect 28288 35838 28636 35980
rect 28288 35774 28294 35838
rect 28358 35774 28636 35838
rect 22168 35708 22244 35768
rect 22576 35708 22652 35768
rect 22168 35430 22380 35708
rect 22576 35436 22788 35708
rect 22478 35430 22788 35436
rect 22168 35366 22310 35430
rect 22374 35366 22380 35430
rect 22440 35366 22446 35430
rect 22510 35366 22788 35430
rect 22168 35360 22380 35366
rect 22478 35360 22788 35366
rect 22984 35566 23196 35572
rect 22984 35502 22990 35566
rect 23054 35502 23196 35566
rect 22984 35430 23196 35502
rect 22984 35366 22990 35430
rect 23054 35366 23196 35430
rect 22984 35360 23196 35366
rect 23392 35566 23604 35572
rect 23392 35502 23534 35566
rect 23598 35502 23604 35566
rect 23392 35430 23604 35502
rect 28288 35496 28636 35774
rect 190128 35496 190340 35980
rect 195024 35974 195236 35980
rect 195024 35910 195030 35974
rect 195094 35910 195236 35974
rect 195024 35838 195236 35910
rect 195024 35774 195166 35838
rect 195230 35774 195236 35838
rect 195024 35768 195236 35774
rect 195432 35974 195644 35980
rect 195432 35910 195438 35974
rect 195502 35910 195644 35974
rect 195432 35838 195644 35910
rect 195432 35774 195438 35838
rect 195502 35774 195644 35838
rect 195432 35768 195644 35774
rect 195840 35768 196052 35980
rect 196248 35974 196460 35980
rect 196248 35910 196390 35974
rect 196454 35910 196460 35974
rect 196248 35844 196460 35910
rect 196112 35768 196460 35844
rect 196656 35768 196868 36116
rect 195840 35708 195916 35768
rect 196112 35708 196188 35768
rect 196792 35708 196868 35768
rect 195840 35632 196188 35708
rect 195024 35566 195236 35572
rect 195024 35502 195166 35566
rect 195230 35502 195236 35566
rect 28424 35436 28500 35496
rect 190128 35436 190204 35496
rect 23392 35366 23398 35430
rect 23462 35366 23604 35430
rect 23392 35360 23604 35366
rect 21896 35300 21972 35360
rect 21760 35158 21972 35300
rect 28288 35224 28636 35436
rect 190128 35294 190340 35436
rect 195024 35430 195236 35502
rect 195024 35366 195166 35430
rect 195230 35366 195236 35430
rect 195024 35360 195236 35366
rect 195432 35566 195644 35572
rect 195432 35502 195438 35566
rect 195502 35502 195644 35566
rect 195432 35430 195644 35502
rect 195432 35366 195438 35430
rect 195502 35366 195644 35430
rect 195432 35360 195644 35366
rect 195840 35430 196052 35632
rect 196248 35436 196460 35708
rect 196150 35430 196460 35436
rect 195840 35366 195982 35430
rect 196046 35366 196052 35430
rect 196112 35366 196118 35430
rect 196182 35366 196460 35430
rect 195840 35360 196052 35366
rect 196150 35360 196460 35366
rect 196656 35360 196868 35708
rect 216784 35838 217540 35844
rect 216784 35812 217470 35838
rect 216784 35756 216908 35812
rect 216964 35774 217470 35812
rect 217534 35774 217540 35838
rect 216964 35768 217540 35774
rect 216964 35756 216996 35768
rect 216784 35632 216996 35756
rect 196792 35300 196868 35360
rect 190128 35230 190270 35294
rect 190334 35230 190340 35294
rect 190128 35224 190340 35230
rect 28560 35164 28636 35224
rect 190264 35164 190340 35224
rect 21760 35094 21902 35158
rect 21966 35094 21972 35158
rect 21760 35088 21972 35094
rect 22168 35158 22516 35164
rect 22168 35094 22310 35158
rect 22374 35094 22446 35158
rect 22510 35094 22516 35158
rect 22168 35088 22516 35094
rect 22168 35028 22380 35088
rect 14144 34909 14356 35028
rect 15152 34982 15218 34985
rect 15406 34982 15472 34985
rect 15152 34980 15472 34982
rect 15152 34924 15157 34980
rect 15213 34924 15411 34980
rect 15467 34924 15472 34980
rect 22168 34952 22516 35028
rect 22576 34952 22788 35164
rect 22984 35158 23196 35164
rect 22984 35094 22990 35158
rect 23054 35094 23196 35158
rect 22984 34952 23196 35094
rect 15152 34922 15472 34924
rect 15152 34919 15218 34922
rect 15406 34919 15472 34922
rect 14144 34892 14212 34909
rect 0 34853 14212 34892
rect 14268 34853 14356 34909
rect 22304 34892 22380 34952
rect 0 34816 14356 34853
rect 21760 34886 21972 34892
rect 21760 34822 21902 34886
rect 21966 34822 21972 34886
rect 21760 34750 21972 34822
rect 21760 34686 21766 34750
rect 21830 34686 21972 34750
rect 21760 34680 21972 34686
rect 22168 34750 22380 34892
rect 22440 34892 22516 34952
rect 22712 34892 22788 34952
rect 23120 34892 23196 34952
rect 22440 34816 22788 34892
rect 22168 34686 22174 34750
rect 22238 34686 22380 34750
rect 22168 34680 22380 34686
rect 22576 34750 22788 34816
rect 22576 34686 22582 34750
rect 22646 34686 22788 34750
rect 22576 34680 22788 34686
rect 15238 34658 15322 34662
rect 15238 34653 15355 34658
rect 15238 34597 15294 34653
rect 15350 34597 15355 34653
rect 15238 34592 15355 34597
rect 15238 34588 15322 34592
rect 22984 34544 23196 34892
rect 23392 35158 23604 35164
rect 23392 35094 23398 35158
rect 23462 35094 23604 35158
rect 23392 34952 23604 35094
rect 23392 34892 23468 34952
rect 23392 34544 23604 34892
rect 28288 34886 28636 35164
rect 28288 34822 28430 34886
rect 28494 34822 28636 34886
rect 28288 34816 28636 34822
rect 190128 35022 190340 35164
rect 190128 34958 190270 35022
rect 190334 34958 190340 35022
rect 190128 34886 190340 34958
rect 190128 34822 190134 34886
rect 190198 34822 190340 34886
rect 190128 34816 190340 34822
rect 195024 35158 195236 35164
rect 195024 35094 195166 35158
rect 195230 35094 195236 35158
rect 195024 34952 195236 35094
rect 195432 35158 195644 35164
rect 195432 35094 195438 35158
rect 195502 35094 195644 35158
rect 195432 34952 195644 35094
rect 195840 35158 196188 35164
rect 195840 35094 195982 35158
rect 196046 35094 196118 35158
rect 196182 35094 196188 35158
rect 195840 35088 196188 35094
rect 195840 35028 196052 35088
rect 195840 34952 196188 35028
rect 196248 34952 196460 35164
rect 196656 35158 196868 35300
rect 196656 35094 196798 35158
rect 196862 35094 196868 35158
rect 196656 35088 196868 35094
rect 195024 34892 195100 34952
rect 195432 34892 195508 34952
rect 195976 34892 196052 34952
rect 23120 34484 23196 34544
rect 23528 34484 23604 34544
rect 14552 34478 14764 34484
rect 14552 34414 14694 34478
rect 14758 34414 14764 34478
rect 14552 34212 14764 34414
rect 21760 34478 21972 34484
rect 21760 34414 21766 34478
rect 21830 34414 21972 34478
rect 21760 34342 21972 34414
rect 21760 34278 21766 34342
rect 21830 34278 21972 34342
rect 21760 34272 21972 34278
rect 22168 34478 22380 34484
rect 22168 34414 22174 34478
rect 22238 34414 22380 34478
rect 1632 34132 1844 34212
rect 14552 34206 16668 34212
rect 14552 34142 16598 34206
rect 16662 34142 16668 34206
rect 14552 34136 16668 34142
rect 19176 34136 19796 34212
rect 22168 34136 22380 34414
rect 22576 34478 22788 34484
rect 22576 34414 22582 34478
rect 22646 34414 22788 34478
rect 22576 34212 22788 34414
rect 22440 34136 22788 34212
rect 1632 34076 1702 34132
rect 1758 34076 1844 34132
rect 19176 34076 19252 34136
rect 19720 34076 19796 34136
rect 22440 34076 22516 34136
rect 22712 34076 22788 34136
rect 1224 34070 1844 34076
rect 1224 34006 1230 34070
rect 1294 34006 1844 34070
rect 1224 34000 1844 34006
rect 18088 33940 18300 34076
rect 18496 34070 19252 34076
rect 18496 34006 18502 34070
rect 18566 34006 19252 34070
rect 18496 34000 19252 34006
rect 18088 33934 18436 33940
rect 18088 33870 18230 33934
rect 18294 33870 18436 33934
rect 18088 33864 18436 33870
rect 18496 33864 18708 34000
rect 18904 33934 19116 34000
rect 18904 33870 18910 33934
rect 18974 33870 19116 33934
rect 18904 33864 19116 33870
rect 19312 33934 19524 34076
rect 19312 33870 19318 33934
rect 19382 33870 19524 33934
rect 19312 33864 19524 33870
rect 19720 33864 19932 34076
rect 21760 34070 21972 34076
rect 21760 34006 21766 34070
rect 21830 34006 21972 34070
rect 21760 33934 21972 34006
rect 21760 33870 21766 33934
rect 21830 33870 21972 33934
rect 21760 33864 21972 33870
rect 22168 34000 22516 34076
rect 22168 33934 22380 34000
rect 22168 33870 22174 33934
rect 22238 33870 22380 33934
rect 22168 33864 22380 33870
rect 22576 33934 22788 34076
rect 22576 33870 22582 33934
rect 22646 33870 22788 33934
rect 22576 33864 22788 33870
rect 22984 34136 23196 34484
rect 23392 34136 23604 34484
rect 28288 34614 28636 34620
rect 28288 34550 28430 34614
rect 28494 34550 28636 34614
rect 28288 34478 28636 34550
rect 28288 34414 28294 34478
rect 28358 34414 28636 34478
rect 28288 34206 28636 34414
rect 28288 34142 28294 34206
rect 28358 34142 28430 34206
rect 28494 34142 28636 34206
rect 22984 34076 23060 34136
rect 23392 34076 23468 34136
rect 22984 33934 23196 34076
rect 22984 33870 22990 33934
rect 23054 33870 23196 33934
rect 22984 33864 23196 33870
rect 23392 33934 23604 34076
rect 28288 34000 28636 34142
rect 190128 34614 190340 34620
rect 190128 34550 190134 34614
rect 190198 34550 190340 34614
rect 190128 34478 190340 34550
rect 190128 34414 190134 34478
rect 190198 34414 190340 34478
rect 190128 34206 190340 34414
rect 190128 34142 190134 34206
rect 190198 34142 190340 34206
rect 190128 34000 190340 34142
rect 28560 33940 28636 34000
rect 190264 33940 190340 34000
rect 23392 33870 23534 33934
rect 23598 33870 23604 33934
rect 23392 33864 23604 33870
rect 28288 33934 28636 33940
rect 28288 33870 28430 33934
rect 28494 33870 28636 33934
rect 18360 33804 18436 33864
rect 19312 33804 19388 33864
rect 18360 33728 19388 33804
rect 21760 33662 21972 33668
rect 21760 33598 21766 33662
rect 21830 33598 21972 33662
rect 21760 33526 21972 33598
rect 21760 33462 21766 33526
rect 21830 33462 21972 33526
rect 21760 33456 21972 33462
rect 22168 33662 22380 33668
rect 22168 33598 22174 33662
rect 22238 33598 22380 33662
rect 22168 33456 22380 33598
rect 22576 33662 22788 33668
rect 22576 33598 22582 33662
rect 22646 33598 22788 33662
rect 22576 33526 22788 33598
rect 22576 33462 22582 33526
rect 22646 33462 22788 33526
rect 22576 33456 22788 33462
rect 22984 33662 23196 33668
rect 22984 33598 22990 33662
rect 23054 33598 23196 33662
rect 22984 33526 23196 33598
rect 22984 33462 23126 33526
rect 23190 33462 23196 33526
rect 22984 33456 23196 33462
rect 23392 33662 23604 33668
rect 23392 33598 23534 33662
rect 23598 33598 23604 33662
rect 23392 33526 23604 33598
rect 23392 33462 23534 33526
rect 23598 33462 23604 33526
rect 23392 33456 23604 33462
rect 28288 33456 28636 33870
rect 190128 33456 190340 33940
rect 195024 34544 195236 34892
rect 195432 34544 195644 34892
rect 195840 34750 196052 34892
rect 196112 34892 196188 34952
rect 196384 34892 196460 34952
rect 196112 34816 196460 34892
rect 195840 34686 195846 34750
rect 195910 34686 196052 34750
rect 195840 34680 196052 34686
rect 196248 34680 196460 34816
rect 196656 34886 196868 34892
rect 196656 34822 196798 34886
rect 196862 34822 196868 34886
rect 196656 34750 196868 34822
rect 196656 34686 196662 34750
rect 196726 34686 196868 34750
rect 196656 34680 196868 34686
rect 195024 34484 195100 34544
rect 195432 34484 195508 34544
rect 195024 34136 195236 34484
rect 195432 34136 195644 34484
rect 195840 34478 196052 34484
rect 195840 34414 195846 34478
rect 195910 34414 196052 34478
rect 195840 34212 196052 34414
rect 195840 34136 196188 34212
rect 196248 34136 196460 34484
rect 196656 34478 196868 34484
rect 196656 34414 196662 34478
rect 196726 34414 196868 34478
rect 196656 34342 196868 34414
rect 196656 34278 196662 34342
rect 196726 34278 196868 34342
rect 196656 34272 196868 34278
rect 195024 34076 195100 34136
rect 195432 34076 195508 34136
rect 195976 34076 196052 34136
rect 195024 33934 195236 34076
rect 195024 33870 195166 33934
rect 195230 33870 195236 33934
rect 195024 33864 195236 33870
rect 195432 33934 195644 34076
rect 195432 33870 195438 33934
rect 195502 33870 195644 33934
rect 195432 33864 195644 33870
rect 195840 33864 196052 34076
rect 196112 34076 196188 34136
rect 196384 34076 196460 34136
rect 199376 34136 200540 34212
rect 199376 34076 199452 34136
rect 200464 34076 200540 34136
rect 216784 34206 217540 34212
rect 216784 34142 217470 34206
rect 217534 34142 217540 34206
rect 216784 34136 217540 34142
rect 216784 34132 216996 34136
rect 216784 34076 216908 34132
rect 216964 34076 216996 34132
rect 196112 34000 196460 34076
rect 196248 33934 196460 34000
rect 196248 33870 196390 33934
rect 196454 33870 196460 33934
rect 196248 33864 196460 33870
rect 196656 34070 196868 34076
rect 196656 34006 196662 34070
rect 196726 34006 196868 34070
rect 196656 33934 196868 34006
rect 196656 33870 196662 33934
rect 196726 33870 196868 33934
rect 196656 33864 196868 33870
rect 198832 33934 199044 34076
rect 198832 33870 198838 33934
rect 198902 33870 199044 33934
rect 198832 33864 199044 33870
rect 199104 33934 199452 34076
rect 199104 33870 199110 33934
rect 199174 33870 199452 33934
rect 199104 33864 199452 33870
rect 199512 34000 200268 34076
rect 199512 33864 199724 34000
rect 199920 33864 200268 34000
rect 200464 33934 200676 34076
rect 216784 34000 216996 34076
rect 200464 33870 200470 33934
rect 200534 33870 200676 33934
rect 200464 33864 200676 33870
rect 198968 33804 199044 33864
rect 199512 33804 199588 33864
rect 198968 33728 199588 33804
rect 195024 33662 195236 33668
rect 195024 33598 195166 33662
rect 195230 33598 195236 33662
rect 195024 33526 195236 33598
rect 195024 33462 195166 33526
rect 195230 33462 195236 33526
rect 195024 33456 195236 33462
rect 195432 33662 195644 33668
rect 195432 33598 195438 33662
rect 195502 33598 195644 33662
rect 195432 33526 195644 33598
rect 195432 33462 195574 33526
rect 195638 33462 195644 33526
rect 195432 33456 195644 33462
rect 195840 33532 196052 33668
rect 196248 33662 196460 33668
rect 196248 33598 196390 33662
rect 196454 33598 196460 33662
rect 195840 33526 196188 33532
rect 195840 33462 196118 33526
rect 196182 33462 196188 33526
rect 195840 33456 196188 33462
rect 196248 33526 196460 33598
rect 196248 33462 196390 33526
rect 196454 33462 196460 33526
rect 196248 33456 196460 33462
rect 196656 33662 196868 33668
rect 196656 33598 196662 33662
rect 196726 33598 196868 33662
rect 196656 33526 196868 33598
rect 196656 33462 196662 33526
rect 196726 33462 196868 33526
rect 196656 33456 196868 33462
rect 28288 33396 28364 33456
rect 190128 33396 190204 33456
rect 18088 33254 18300 33260
rect 18088 33190 18230 33254
rect 18294 33190 18300 33254
rect 18088 33118 18300 33190
rect 18088 33054 18094 33118
rect 18158 33054 18300 33118
rect 18088 33048 18300 33054
rect 18496 33254 19116 33260
rect 18496 33190 18910 33254
rect 18974 33190 19116 33254
rect 18496 33184 19116 33190
rect 18496 33124 18708 33184
rect 18904 33124 19116 33184
rect 19312 33254 19524 33260
rect 19312 33190 19318 33254
rect 19382 33190 19524 33254
rect 18496 33118 18844 33124
rect 18496 33054 18774 33118
rect 18838 33054 18844 33118
rect 18496 33048 18844 33054
rect 18904 33048 19252 33124
rect 19312 33118 19524 33190
rect 19312 33054 19454 33118
rect 19518 33054 19524 33118
rect 19312 33048 19524 33054
rect 19720 33048 19932 33260
rect 21760 33254 21972 33260
rect 21760 33190 21766 33254
rect 21830 33190 21972 33254
rect 21760 33118 21972 33190
rect 21760 33054 21902 33118
rect 21966 33054 21972 33118
rect 21760 33048 21972 33054
rect 22168 33254 22788 33260
rect 22168 33190 22582 33254
rect 22646 33190 22788 33254
rect 22168 33184 22788 33190
rect 22168 33124 22380 33184
rect 22168 33118 22516 33124
rect 22168 33054 22446 33118
rect 22510 33054 22516 33118
rect 22168 33048 22516 33054
rect 22576 33048 22788 33184
rect 22984 33254 23196 33260
rect 22984 33190 23126 33254
rect 23190 33190 23196 33254
rect 22984 33118 23196 33190
rect 22984 33054 22990 33118
rect 23054 33054 23196 33118
rect 22984 33048 23196 33054
rect 23392 33254 23604 33260
rect 23392 33190 23534 33254
rect 23598 33190 23604 33254
rect 23392 33118 23604 33190
rect 28288 33184 28636 33396
rect 190128 33184 190340 33396
rect 28424 33124 28500 33184
rect 190264 33124 190340 33184
rect 23392 33054 23398 33118
rect 23462 33054 23604 33118
rect 23392 33048 23604 33054
rect 19176 32988 19252 33048
rect 19720 32988 19796 33048
rect 19176 32912 19796 32988
rect 28288 32912 28636 33124
rect 190128 32912 190340 33124
rect 195024 33254 195236 33260
rect 195024 33190 195166 33254
rect 195230 33190 195236 33254
rect 195024 33118 195236 33190
rect 195024 33054 195030 33118
rect 195094 33054 195236 33118
rect 195024 33048 195236 33054
rect 195432 33254 195644 33260
rect 195432 33190 195574 33254
rect 195638 33190 195644 33254
rect 195432 33118 195644 33190
rect 195432 33054 195574 33118
rect 195638 33054 195644 33118
rect 195432 33048 195644 33054
rect 195840 33118 196052 33260
rect 196150 33254 196460 33260
rect 196112 33190 196118 33254
rect 196182 33190 196390 33254
rect 196454 33190 196460 33254
rect 196150 33184 196460 33190
rect 196248 33124 196460 33184
rect 196150 33118 196460 33124
rect 195840 33054 195982 33118
rect 196046 33054 196052 33118
rect 196112 33054 196118 33118
rect 196182 33054 196460 33118
rect 195840 33048 196052 33054
rect 196150 33048 196460 33054
rect 196656 33254 196868 33260
rect 196656 33190 196662 33254
rect 196726 33190 196868 33254
rect 196656 33118 196868 33190
rect 196656 33054 196798 33118
rect 196862 33054 196868 33118
rect 196656 33048 196868 33054
rect 198832 33254 199044 33260
rect 198832 33190 198838 33254
rect 198902 33190 199044 33254
rect 198832 33048 199044 33190
rect 199104 33254 199452 33260
rect 199104 33190 199110 33254
rect 199174 33190 199452 33254
rect 199104 33118 199452 33190
rect 199104 33054 199110 33118
rect 199174 33054 199452 33118
rect 199104 33048 199452 33054
rect 199512 33184 200268 33260
rect 199512 33124 199724 33184
rect 199512 33118 199860 33124
rect 199512 33054 199790 33118
rect 199854 33054 199860 33118
rect 199512 33048 199860 33054
rect 199920 33048 200268 33184
rect 200464 33254 200676 33260
rect 200464 33190 200470 33254
rect 200534 33190 200676 33254
rect 200464 33118 200676 33190
rect 200464 33054 200470 33118
rect 200534 33054 200676 33118
rect 200464 33048 200676 33054
rect 198968 32988 199044 33048
rect 199512 32988 199588 33048
rect 198968 32912 199588 32988
rect 28424 32852 28500 32912
rect 190264 32852 190340 32912
rect 21760 32846 21972 32852
rect 21760 32782 21902 32846
rect 21966 32782 21972 32846
rect 21760 32710 21972 32782
rect 21760 32646 21902 32710
rect 21966 32646 21972 32710
rect 21760 32640 21972 32646
rect 22168 32716 22380 32852
rect 22478 32846 22788 32852
rect 22440 32782 22446 32846
rect 22510 32782 22788 32846
rect 22478 32776 22788 32782
rect 22576 32716 22788 32776
rect 22168 32640 22788 32716
rect 22984 32846 23196 32852
rect 22984 32782 22990 32846
rect 23054 32782 23196 32846
rect 22984 32710 23196 32782
rect 22984 32646 23126 32710
rect 23190 32646 23196 32710
rect 22984 32640 23196 32646
rect 23392 32846 23604 32852
rect 23392 32782 23398 32846
rect 23462 32782 23604 32846
rect 23392 32710 23604 32782
rect 23392 32646 23398 32710
rect 23462 32646 23604 32710
rect 23392 32640 23604 32646
rect 28288 32640 28636 32852
rect 190128 32640 190340 32852
rect 195024 32846 195236 32852
rect 195024 32782 195030 32846
rect 195094 32782 195236 32846
rect 195024 32710 195236 32782
rect 195024 32646 195166 32710
rect 195230 32646 195236 32710
rect 195024 32640 195236 32646
rect 195432 32846 195644 32852
rect 195432 32782 195574 32846
rect 195638 32782 195644 32846
rect 195432 32710 195644 32782
rect 195432 32646 195438 32710
rect 195502 32646 195644 32710
rect 195432 32640 195644 32646
rect 195840 32846 196188 32852
rect 195840 32782 195982 32846
rect 196046 32782 196118 32846
rect 196182 32782 196188 32846
rect 195840 32776 196188 32782
rect 195840 32716 196052 32776
rect 196248 32716 196460 32852
rect 195840 32710 196460 32716
rect 195840 32646 195982 32710
rect 196046 32646 196390 32710
rect 196454 32646 196460 32710
rect 195840 32640 196460 32646
rect 196656 32846 196868 32852
rect 196656 32782 196798 32846
rect 196862 32782 196868 32846
rect 196656 32710 196868 32782
rect 196656 32646 196798 32710
rect 196862 32646 196868 32710
rect 196656 32640 196868 32646
rect 22304 32580 22380 32640
rect 28288 32580 28364 32640
rect 190128 32580 190204 32640
rect 1632 32452 1844 32580
rect 22304 32504 22652 32580
rect 1632 32444 1702 32452
rect 1224 32438 1702 32444
rect 1224 32374 1230 32438
rect 1294 32396 1702 32438
rect 1758 32396 1844 32452
rect 22576 32444 22652 32504
rect 1294 32374 1844 32396
rect 1224 32368 1844 32374
rect 18088 32438 18300 32444
rect 18088 32374 18094 32438
rect 18158 32374 18300 32438
rect 18088 32302 18300 32374
rect 18088 32238 18094 32302
rect 18158 32238 18300 32302
rect 18088 32232 18300 32238
rect 18496 32438 19116 32444
rect 18496 32374 18910 32438
rect 18974 32374 19116 32438
rect 18496 32368 19116 32374
rect 18496 32232 18708 32368
rect 18904 32302 19116 32368
rect 18904 32238 18910 32302
rect 18974 32238 19116 32302
rect 18904 32232 19116 32238
rect 19312 32438 19524 32444
rect 19312 32374 19454 32438
rect 19518 32374 19524 32438
rect 19312 32302 19524 32374
rect 19312 32238 19454 32302
rect 19518 32238 19524 32302
rect 19312 32232 19524 32238
rect 19720 32302 19932 32444
rect 19720 32238 19862 32302
rect 19926 32238 19932 32302
rect 19720 32232 19932 32238
rect 21760 32438 21972 32444
rect 21760 32374 21902 32438
rect 21966 32374 21972 32438
rect 21760 32232 21972 32374
rect 22168 32302 22380 32444
rect 22168 32238 22174 32302
rect 22238 32238 22380 32302
rect 22168 32232 22380 32238
rect 22576 32302 22788 32444
rect 22576 32238 22718 32302
rect 22782 32238 22788 32302
rect 22576 32232 22788 32238
rect 22984 32438 23196 32444
rect 22984 32374 23126 32438
rect 23190 32374 23196 32438
rect 22984 32302 23196 32374
rect 22984 32238 22990 32302
rect 23054 32238 23196 32302
rect 22984 32232 23196 32238
rect 23392 32438 23604 32444
rect 23392 32374 23398 32438
rect 23462 32374 23604 32438
rect 23392 32302 23604 32374
rect 23392 32238 23534 32302
rect 23598 32238 23604 32302
rect 23392 32232 23604 32238
rect 28288 32368 28636 32580
rect 190128 32368 190340 32580
rect 216784 32574 217540 32580
rect 216784 32510 217470 32574
rect 217534 32510 217540 32574
rect 216784 32504 217540 32510
rect 216784 32452 216996 32504
rect 195024 32438 195236 32444
rect 195024 32374 195166 32438
rect 195230 32374 195236 32438
rect 28288 32308 28364 32368
rect 190128 32308 190204 32368
rect 21760 32172 21836 32232
rect 21760 31894 21972 32172
rect 28288 32096 28636 32308
rect 190128 32096 190340 32308
rect 195024 32302 195236 32374
rect 195024 32238 195166 32302
rect 195230 32238 195236 32302
rect 195024 32232 195236 32238
rect 195432 32438 195644 32444
rect 195432 32374 195438 32438
rect 195502 32374 195644 32438
rect 195432 32302 195644 32374
rect 195432 32238 195438 32302
rect 195502 32238 195644 32302
rect 195432 32232 195644 32238
rect 195840 32438 196052 32444
rect 195840 32374 195982 32438
rect 196046 32374 196052 32438
rect 195840 32232 196052 32374
rect 196248 32438 196460 32444
rect 196248 32374 196390 32438
rect 196454 32374 196460 32438
rect 196248 32308 196460 32374
rect 196150 32302 196460 32308
rect 196112 32238 196118 32302
rect 196182 32238 196460 32302
rect 196150 32232 196460 32238
rect 196656 32438 196868 32444
rect 196656 32374 196798 32438
rect 196862 32374 196868 32438
rect 196656 32232 196868 32374
rect 198832 32302 199044 32444
rect 198832 32238 198974 32302
rect 199038 32238 199044 32302
rect 198832 32232 199044 32238
rect 199104 32438 199452 32444
rect 199104 32374 199110 32438
rect 199174 32374 199452 32438
rect 199104 32302 199452 32374
rect 199104 32238 199246 32302
rect 199310 32238 199452 32302
rect 199104 32232 199452 32238
rect 199512 32438 200268 32444
rect 199512 32374 199926 32438
rect 199990 32374 200268 32438
rect 199512 32368 200268 32374
rect 199512 32232 199724 32368
rect 199920 32232 200268 32368
rect 200464 32438 200676 32444
rect 200464 32374 200470 32438
rect 200534 32374 200676 32438
rect 200464 32308 200676 32374
rect 216784 32396 216908 32452
rect 216964 32396 216996 32452
rect 216784 32368 216996 32396
rect 200464 32302 201900 32308
rect 200464 32238 200470 32302
rect 200534 32238 201830 32302
rect 201894 32238 201900 32302
rect 200464 32232 201900 32238
rect 196792 32172 196868 32232
rect 28424 32036 28500 32096
rect 190264 32036 190340 32096
rect 21760 31830 21902 31894
rect 21966 31830 21972 31894
rect 21760 31824 21972 31830
rect 22168 32030 22380 32036
rect 22168 31966 22174 32030
rect 22238 31966 22380 32030
rect 22168 31894 22380 31966
rect 22576 32030 22788 32036
rect 22576 31966 22718 32030
rect 22782 31966 22788 32030
rect 22576 31900 22788 31966
rect 22478 31894 22788 31900
rect 22168 31830 22310 31894
rect 22374 31830 22380 31894
rect 22440 31830 22446 31894
rect 22510 31830 22788 31894
rect 22168 31824 22380 31830
rect 22478 31824 22788 31830
rect 22984 32030 23196 32036
rect 22984 31966 22990 32030
rect 23054 31966 23196 32030
rect 22984 31894 23196 31966
rect 22984 31830 23126 31894
rect 23190 31830 23196 31894
rect 22984 31824 23196 31830
rect 23392 32030 23604 32036
rect 23392 31966 23534 32030
rect 23598 31966 23604 32030
rect 23392 31894 23604 31966
rect 23392 31830 23398 31894
rect 23462 31830 23604 31894
rect 23392 31824 23604 31830
rect 28288 31824 28636 32036
rect 190128 31824 190340 32036
rect 195024 32030 195236 32036
rect 195024 31966 195166 32030
rect 195230 31966 195236 32030
rect 195024 31894 195236 31966
rect 195024 31830 195030 31894
rect 195094 31830 195236 31894
rect 195024 31824 195236 31830
rect 195432 32030 195644 32036
rect 195432 31966 195438 32030
rect 195502 31966 195644 32030
rect 195432 31894 195644 31966
rect 195432 31830 195438 31894
rect 195502 31830 195644 31894
rect 195432 31824 195644 31830
rect 195840 32030 196188 32036
rect 195840 31966 196118 32030
rect 196182 31966 196188 32030
rect 195840 31960 196188 31966
rect 195840 31900 196052 31960
rect 196248 31900 196460 32036
rect 195840 31894 196460 31900
rect 195840 31830 196390 31894
rect 196454 31830 196460 31894
rect 195840 31824 196460 31830
rect 196656 31894 196868 32172
rect 198968 32172 199044 32232
rect 199512 32172 199588 32232
rect 198968 32096 199588 32172
rect 196656 31830 196662 31894
rect 196726 31830 196868 31894
rect 196656 31824 196868 31830
rect 28288 31764 28364 31824
rect 190264 31764 190340 31824
rect 16864 31688 18164 31764
rect 16864 31628 16940 31688
rect 18088 31628 18164 31688
rect 19176 31688 19796 31764
rect 19176 31628 19252 31688
rect 19720 31628 19796 31688
rect 16592 31622 16940 31628
rect 16592 31558 16598 31622
rect 16662 31558 16940 31622
rect 16592 31552 16940 31558
rect 16592 31416 16804 31552
rect 17000 31492 17212 31628
rect 18088 31622 18300 31628
rect 18088 31558 18094 31622
rect 18158 31558 18300 31622
rect 17000 31416 18028 31492
rect 18088 31416 18300 31558
rect 18496 31622 19252 31628
rect 18496 31558 18910 31622
rect 18974 31558 19252 31622
rect 18496 31552 19252 31558
rect 19312 31622 19524 31628
rect 19312 31558 19454 31622
rect 19518 31558 19524 31622
rect 18496 31416 18708 31552
rect 18904 31486 19116 31552
rect 18904 31422 18910 31486
rect 18974 31422 19116 31486
rect 18904 31416 19116 31422
rect 19312 31486 19524 31558
rect 19312 31422 19318 31486
rect 19382 31422 19524 31486
rect 19312 31416 19524 31422
rect 19720 31622 19932 31628
rect 19720 31558 19862 31622
rect 19926 31558 19932 31622
rect 19720 31416 19932 31558
rect 21760 31622 21972 31628
rect 21760 31558 21902 31622
rect 21966 31558 21972 31622
rect 21760 31416 21972 31558
rect 22168 31622 22516 31628
rect 22168 31558 22310 31622
rect 22374 31558 22446 31622
rect 22510 31558 22516 31622
rect 22168 31552 22516 31558
rect 22168 31492 22380 31552
rect 22576 31492 22788 31628
rect 22168 31486 22788 31492
rect 22168 31422 22582 31486
rect 22646 31422 22788 31486
rect 22168 31416 22788 31422
rect 22984 31622 23196 31628
rect 22984 31558 23126 31622
rect 23190 31558 23196 31622
rect 22984 31486 23196 31558
rect 22984 31422 22990 31486
rect 23054 31422 23196 31486
rect 22984 31416 23196 31422
rect 23392 31622 23604 31628
rect 23392 31558 23398 31622
rect 23462 31558 23604 31622
rect 23392 31486 23604 31558
rect 23392 31422 23534 31486
rect 23598 31422 23604 31486
rect 23392 31416 23604 31422
rect 28288 31552 28636 31764
rect 190128 31552 190340 31764
rect 198968 31688 199588 31764
rect 198968 31628 199044 31688
rect 199512 31628 199588 31688
rect 200328 31688 201492 31764
rect 200328 31628 200404 31688
rect 201416 31628 201492 31688
rect 195024 31622 195236 31628
rect 195024 31558 195030 31622
rect 195094 31558 195236 31622
rect 28288 31492 28364 31552
rect 190128 31492 190204 31552
rect 17952 31356 18028 31416
rect 18496 31356 18572 31416
rect 17952 31280 18572 31356
rect 21760 31356 21836 31416
rect 21760 31214 21972 31356
rect 28288 31350 28636 31492
rect 28288 31286 28566 31350
rect 28630 31286 28636 31350
rect 28288 31280 28636 31286
rect 28560 31220 28636 31280
rect 21760 31150 21766 31214
rect 21830 31150 21972 31214
rect 21760 31144 21972 31150
rect 2720 31008 3748 31084
rect 2720 30872 2932 31008
rect 3400 30872 3748 31008
rect 22168 31008 22380 31220
rect 22576 31214 22788 31220
rect 22576 31150 22582 31214
rect 22646 31150 22788 31214
rect 22576 31084 22788 31150
rect 22440 31008 22788 31084
rect 22984 31214 23196 31220
rect 22984 31150 22990 31214
rect 23054 31150 23196 31214
rect 22984 31078 23196 31150
rect 22984 31014 22990 31078
rect 23054 31014 23196 31078
rect 22984 31008 23196 31014
rect 23392 31214 23604 31220
rect 23392 31150 23534 31214
rect 23598 31150 23604 31214
rect 23392 31078 23604 31150
rect 23392 31014 23534 31078
rect 23598 31014 23604 31078
rect 23392 31008 23604 31014
rect 28288 31078 28636 31220
rect 28288 31014 28566 31078
rect 28630 31014 28636 31078
rect 22168 30948 22244 31008
rect 22440 30948 22516 31008
rect 21760 30942 21972 30948
rect 21760 30878 21766 30942
rect 21830 30878 21972 30942
rect 2720 30812 2796 30872
rect 1224 30806 2796 30812
rect 1224 30742 1230 30806
rect 1294 30772 2796 30806
rect 1294 30742 1702 30772
rect 1224 30736 1702 30742
rect 1632 30716 1702 30736
rect 1758 30736 2796 30772
rect 1758 30716 1844 30736
rect 1632 30600 1844 30716
rect 21760 30600 21972 30878
rect 22168 30872 22516 30948
rect 22576 30948 22652 31008
rect 22576 30872 22788 30948
rect 22168 30676 22380 30872
rect 22688 30676 22788 30872
rect 22070 30670 22380 30676
rect 22032 30606 22038 30670
rect 22102 30606 22174 30670
rect 22238 30606 22380 30670
rect 22070 30600 22380 30606
rect 22576 30670 22788 30676
rect 22576 30606 22582 30670
rect 22646 30606 22788 30670
rect 22576 30600 22788 30606
rect 22984 30806 23196 30812
rect 22984 30742 22990 30806
rect 23054 30742 23196 30806
rect 22984 30600 23196 30742
rect 21896 30540 21972 30600
rect 23120 30540 23196 30600
rect 21760 30398 21972 30540
rect 2108 30356 2174 30357
rect 2066 30292 2109 30356
rect 2173 30292 2216 30356
rect 21760 30334 21766 30398
rect 21830 30334 21972 30398
rect 21760 30328 21972 30334
rect 22168 30398 22380 30404
rect 22168 30334 22174 30398
rect 22238 30334 22380 30398
rect 2108 30291 2174 30292
rect 21624 30262 22108 30268
rect 21624 30198 22038 30262
rect 22102 30198 22108 30262
rect 21624 30192 22108 30198
rect 22168 30192 22380 30334
rect 22576 30398 22788 30404
rect 22576 30334 22582 30398
rect 22646 30334 22788 30398
rect 22576 30192 22788 30334
rect 22984 30192 23196 30540
rect 23392 30806 23604 30812
rect 23392 30742 23534 30806
rect 23598 30742 23604 30806
rect 23392 30600 23604 30742
rect 28288 30736 28636 31014
rect 190128 31350 190340 31492
rect 195024 31486 195236 31558
rect 195024 31422 195166 31486
rect 195230 31422 195236 31486
rect 195024 31416 195236 31422
rect 195432 31622 195644 31628
rect 195432 31558 195438 31622
rect 195502 31558 195644 31622
rect 195432 31486 195644 31558
rect 195432 31422 195438 31486
rect 195502 31422 195644 31486
rect 195432 31416 195644 31422
rect 195840 31486 196052 31628
rect 195840 31422 195846 31486
rect 195910 31422 196052 31486
rect 195840 31416 196052 31422
rect 196248 31622 196460 31628
rect 196248 31558 196390 31622
rect 196454 31558 196460 31622
rect 196248 31486 196460 31558
rect 196248 31422 196254 31486
rect 196318 31422 196460 31486
rect 196248 31416 196460 31422
rect 196656 31622 196868 31628
rect 196656 31558 196662 31622
rect 196726 31558 196868 31622
rect 196656 31416 196868 31558
rect 198832 31622 199044 31628
rect 198832 31558 198974 31622
rect 199038 31558 199044 31622
rect 198832 31486 199044 31558
rect 198832 31422 198838 31486
rect 198902 31422 199044 31486
rect 198832 31416 199044 31422
rect 199104 31622 199452 31628
rect 199104 31558 199246 31622
rect 199310 31558 199452 31622
rect 199104 31486 199452 31558
rect 199104 31422 199110 31486
rect 199174 31422 199452 31486
rect 199104 31416 199452 31422
rect 199512 31552 200404 31628
rect 200464 31622 200676 31628
rect 200464 31558 200470 31622
rect 200534 31558 200676 31622
rect 199512 31416 199724 31552
rect 199920 31492 200268 31552
rect 199822 31486 200268 31492
rect 199784 31422 199790 31486
rect 199854 31422 200268 31486
rect 199822 31416 200268 31422
rect 200464 31416 200676 31558
rect 201416 31416 201764 31628
rect 201824 31622 202036 31628
rect 201824 31558 201830 31622
rect 201894 31558 202036 31622
rect 201824 31416 202036 31558
rect 190128 31286 190134 31350
rect 190198 31286 190340 31350
rect 190128 31280 190340 31286
rect 196656 31356 196732 31416
rect 190128 31220 190204 31280
rect 190128 31078 190340 31220
rect 190128 31014 190134 31078
rect 190198 31014 190340 31078
rect 190128 30736 190340 31014
rect 195024 31214 195236 31220
rect 195024 31150 195166 31214
rect 195230 31150 195236 31214
rect 195024 31078 195236 31150
rect 195024 31014 195030 31078
rect 195094 31014 195236 31078
rect 195024 31008 195236 31014
rect 195432 31214 195644 31220
rect 195432 31150 195438 31214
rect 195502 31150 195644 31214
rect 195432 31078 195644 31150
rect 195432 31014 195574 31078
rect 195638 31014 195644 31078
rect 195432 31008 195644 31014
rect 195840 31214 196052 31220
rect 195840 31150 195846 31214
rect 195910 31150 196052 31214
rect 195840 31008 196052 31150
rect 196248 31214 196460 31220
rect 196248 31150 196254 31214
rect 196318 31150 196460 31214
rect 196248 31084 196460 31150
rect 196656 31214 196868 31356
rect 196656 31150 196662 31214
rect 196726 31150 196868 31214
rect 196656 31144 196868 31150
rect 196112 31008 196460 31084
rect 196520 31078 198908 31084
rect 196520 31014 198838 31078
rect 198902 31014 198908 31078
rect 196520 31008 198908 31014
rect 195840 30948 195916 31008
rect 196112 30948 196188 31008
rect 195840 30872 196188 30948
rect 196248 30948 196324 31008
rect 196520 30948 196596 31008
rect 196248 30872 196596 30948
rect 196656 30942 196868 30948
rect 196656 30878 196662 30942
rect 196726 30878 196868 30942
rect 28424 30676 28500 30736
rect 190264 30676 190340 30736
rect 23392 30540 23468 30600
rect 23392 30192 23604 30540
rect 21624 30132 21700 30192
rect 22168 30132 22244 30192
rect 22576 30132 22652 30192
rect 23120 30132 23196 30192
rect 23528 30132 23604 30192
rect 18088 29990 18300 30132
rect 18088 29926 18230 29990
rect 18294 29926 18300 29990
rect 18088 29920 18300 29926
rect 18496 30126 19116 30132
rect 18496 30062 18910 30126
rect 18974 30062 19116 30126
rect 18496 30056 19116 30062
rect 18496 29996 18708 30056
rect 18496 29990 18844 29996
rect 18496 29926 18774 29990
rect 18838 29926 18844 29990
rect 18496 29920 18844 29926
rect 18904 29920 19116 30056
rect 19312 30126 19524 30132
rect 19312 30062 19318 30126
rect 19382 30062 19524 30126
rect 19312 29990 19524 30062
rect 19312 29926 19318 29990
rect 19382 29926 19524 29990
rect 19312 29920 19524 29926
rect 19720 30056 21700 30132
rect 21760 30126 21972 30132
rect 21760 30062 21766 30126
rect 21830 30062 21972 30126
rect 19720 29990 19932 30056
rect 19720 29926 19862 29990
rect 19926 29926 19932 29990
rect 19720 29920 19932 29926
rect 21760 29990 21972 30062
rect 21760 29926 21902 29990
rect 21966 29926 21972 29990
rect 21760 29920 21972 29926
rect 22168 29920 22380 30132
rect 22576 29996 22788 30132
rect 22478 29990 22788 29996
rect 22440 29926 22446 29990
rect 22510 29926 22788 29990
rect 22478 29920 22788 29926
rect 22984 29990 23196 30132
rect 22984 29926 23126 29990
rect 23190 29926 23196 29990
rect 22984 29920 23196 29926
rect 23392 29990 23604 30132
rect 23392 29926 23398 29990
rect 23462 29926 23604 29990
rect 23392 29920 23604 29926
rect 28288 30056 28636 30676
rect 190128 30534 190340 30676
rect 190128 30470 190134 30534
rect 190198 30470 190340 30534
rect 190128 30262 190340 30470
rect 190128 30198 190134 30262
rect 190198 30198 190340 30262
rect 190128 30056 190340 30198
rect 195024 30806 195236 30812
rect 195024 30742 195030 30806
rect 195094 30742 195236 30806
rect 195024 30600 195236 30742
rect 195432 30806 195644 30812
rect 195432 30742 195574 30806
rect 195638 30742 195644 30806
rect 195432 30600 195644 30742
rect 195840 30600 196052 30872
rect 196248 30670 196460 30872
rect 196248 30606 196254 30670
rect 196318 30606 196460 30670
rect 196248 30600 196460 30606
rect 196656 30600 196868 30878
rect 216784 30772 216996 30812
rect 216784 30716 216908 30772
rect 216964 30716 216996 30772
rect 216784 30676 216996 30716
rect 216784 30670 217540 30676
rect 216784 30606 217470 30670
rect 217534 30606 217540 30670
rect 216784 30600 217540 30606
rect 195024 30540 195100 30600
rect 195432 30540 195508 30600
rect 196656 30540 196732 30600
rect 195024 30192 195236 30540
rect 195432 30192 195644 30540
rect 195160 30132 195236 30192
rect 195568 30132 195644 30192
rect 28288 29996 28364 30056
rect 190264 29996 190340 30056
rect 544 29718 3748 29724
rect 544 29654 550 29718
rect 614 29654 3748 29718
rect 544 29648 3748 29654
rect 2720 29512 2932 29648
rect 3400 29512 3748 29648
rect 21760 29718 21972 29724
rect 21760 29654 21902 29718
rect 21966 29654 21972 29718
rect 21760 29582 21972 29654
rect 21760 29518 21902 29582
rect 21966 29518 21972 29582
rect 21760 29512 21972 29518
rect 22168 29718 22516 29724
rect 22168 29654 22446 29718
rect 22510 29654 22516 29718
rect 22168 29648 22516 29654
rect 22168 29588 22380 29648
rect 22576 29588 22788 29724
rect 22168 29582 22788 29588
rect 22168 29518 22310 29582
rect 22374 29518 22718 29582
rect 22782 29518 22788 29582
rect 22168 29512 22788 29518
rect 22984 29718 23196 29724
rect 22984 29654 23126 29718
rect 23190 29654 23196 29718
rect 22984 29582 23196 29654
rect 22984 29518 22990 29582
rect 23054 29518 23196 29582
rect 22984 29512 23196 29518
rect 23392 29718 23604 29724
rect 23392 29654 23398 29718
rect 23462 29654 23604 29718
rect 23392 29582 23604 29654
rect 23392 29518 23398 29582
rect 23462 29518 23604 29582
rect 23392 29512 23604 29518
rect 28288 29512 28636 29996
rect 190128 29512 190340 29996
rect 195024 29990 195236 30132
rect 195024 29926 195166 29990
rect 195230 29926 195236 29990
rect 195024 29920 195236 29926
rect 195432 29990 195644 30132
rect 195432 29926 195438 29990
rect 195502 29926 195644 29990
rect 195432 29920 195644 29926
rect 195840 30192 196052 30404
rect 196248 30398 196460 30404
rect 196248 30334 196254 30398
rect 196318 30334 196460 30398
rect 196248 30192 196460 30334
rect 196656 30398 196868 30540
rect 196656 30334 196662 30398
rect 196726 30334 196868 30398
rect 196656 30328 196868 30334
rect 198968 30192 199588 30268
rect 195840 30132 195916 30192
rect 196248 30132 196324 30192
rect 198968 30132 199044 30192
rect 199512 30132 199588 30192
rect 195840 29990 196052 30132
rect 195840 29926 195846 29990
rect 195910 29926 196052 29990
rect 195840 29920 196052 29926
rect 196248 29920 196460 30132
rect 196656 30126 196868 30132
rect 196656 30062 196662 30126
rect 196726 30062 196868 30126
rect 196656 29990 196868 30062
rect 196656 29926 196798 29990
rect 196862 29926 196868 29990
rect 196656 29920 196868 29926
rect 198832 29920 199044 30132
rect 199104 30126 199452 30132
rect 199104 30062 199110 30126
rect 199174 30062 199452 30126
rect 199104 29990 199452 30062
rect 199104 29926 199110 29990
rect 199174 29926 199382 29990
rect 199446 29926 199452 29990
rect 199104 29920 199452 29926
rect 199512 30126 199860 30132
rect 199512 30062 199790 30126
rect 199854 30062 199860 30126
rect 199512 30056 199860 30062
rect 199512 29996 199724 30056
rect 199920 29996 200268 30132
rect 199512 29990 200268 29996
rect 199512 29926 199926 29990
rect 199990 29926 200268 29990
rect 199512 29920 200268 29926
rect 200464 29990 200676 30132
rect 200464 29926 200606 29990
rect 200670 29926 200676 29990
rect 200464 29920 200676 29926
rect 196248 29860 196324 29920
rect 195976 29784 196324 29860
rect 195976 29724 196052 29784
rect 195024 29718 195236 29724
rect 195024 29654 195166 29718
rect 195230 29654 195236 29718
rect 195024 29582 195236 29654
rect 195024 29518 195166 29582
rect 195230 29518 195236 29582
rect 195024 29512 195236 29518
rect 195432 29718 195644 29724
rect 195432 29654 195438 29718
rect 195502 29654 195644 29718
rect 195432 29582 195644 29654
rect 195432 29518 195438 29582
rect 195502 29518 195644 29582
rect 195432 29512 195644 29518
rect 195840 29718 196460 29724
rect 195840 29654 195846 29718
rect 195910 29654 196460 29718
rect 195840 29648 196460 29654
rect 195840 29582 196052 29648
rect 195840 29518 195846 29582
rect 195910 29518 196052 29582
rect 195840 29512 196052 29518
rect 196248 29512 196460 29648
rect 196656 29718 199180 29724
rect 196656 29654 196798 29718
rect 196862 29654 199110 29718
rect 199174 29654 199180 29718
rect 196656 29648 199180 29654
rect 196656 29582 196868 29648
rect 196656 29518 196662 29582
rect 196726 29518 196868 29582
rect 196656 29512 196868 29518
rect 28424 29452 28500 29512
rect 190264 29452 190340 29512
rect 18088 29310 18300 29316
rect 18088 29246 18230 29310
rect 18294 29246 18300 29310
rect 1224 29174 1844 29180
rect 1224 29110 1230 29174
rect 1294 29110 1844 29174
rect 1224 29104 1844 29110
rect 18088 29174 18300 29246
rect 18088 29110 18230 29174
rect 18294 29110 18300 29174
rect 18088 29104 18300 29110
rect 18496 29310 19116 29316
rect 18496 29246 18910 29310
rect 18974 29246 19116 29310
rect 18496 29240 19116 29246
rect 18496 29104 18708 29240
rect 18904 29180 19116 29240
rect 19312 29310 19524 29316
rect 19312 29246 19318 29310
rect 19382 29246 19524 29310
rect 18904 29174 19252 29180
rect 18904 29110 18910 29174
rect 18974 29110 19252 29174
rect 18904 29104 19252 29110
rect 19312 29174 19524 29246
rect 19312 29110 19454 29174
rect 19518 29110 19524 29174
rect 19312 29104 19524 29110
rect 19720 29310 19932 29316
rect 19720 29246 19862 29310
rect 19926 29246 19932 29310
rect 19720 29104 19932 29246
rect 21760 29310 21972 29316
rect 21760 29246 21902 29310
rect 21966 29246 21972 29310
rect 21760 29174 21972 29246
rect 21760 29110 21766 29174
rect 21830 29110 21972 29174
rect 21760 29104 21972 29110
rect 22168 29310 22380 29316
rect 22168 29246 22310 29310
rect 22374 29246 22380 29310
rect 22168 29104 22380 29246
rect 22576 29310 22788 29316
rect 22576 29246 22718 29310
rect 22782 29246 22788 29310
rect 22576 29174 22788 29246
rect 22576 29110 22582 29174
rect 22646 29110 22788 29174
rect 22576 29104 22788 29110
rect 22984 29310 23196 29316
rect 22984 29246 22990 29310
rect 23054 29246 23196 29310
rect 22984 29174 23196 29246
rect 22984 29110 23126 29174
rect 23190 29110 23196 29174
rect 22984 29104 23196 29110
rect 23392 29310 23604 29316
rect 23392 29246 23398 29310
rect 23462 29246 23604 29310
rect 23392 29174 23604 29246
rect 23392 29110 23534 29174
rect 23598 29110 23604 29174
rect 23392 29104 23604 29110
rect 28288 29240 28636 29452
rect 190128 29240 190340 29452
rect 198968 29376 199588 29452
rect 198968 29316 199044 29376
rect 199512 29316 199588 29376
rect 195024 29310 195236 29316
rect 195024 29246 195166 29310
rect 195230 29246 195236 29310
rect 28288 29180 28364 29240
rect 190128 29180 190204 29240
rect 1632 29092 1844 29104
rect 1632 29036 1702 29092
rect 1758 29036 1844 29092
rect 1632 28968 1844 29036
rect 19176 29044 19252 29104
rect 19720 29044 19796 29104
rect 19176 28968 19796 29044
rect 28288 28968 28636 29180
rect 190128 28968 190340 29180
rect 195024 29174 195236 29246
rect 195024 29110 195166 29174
rect 195230 29110 195236 29174
rect 195024 29104 195236 29110
rect 195432 29310 195644 29316
rect 195432 29246 195438 29310
rect 195502 29246 195644 29310
rect 195432 29174 195644 29246
rect 195432 29110 195438 29174
rect 195502 29110 195644 29174
rect 195432 29104 195644 29110
rect 195840 29310 196052 29316
rect 195840 29246 195846 29310
rect 195910 29246 196052 29310
rect 195840 29174 196052 29246
rect 195840 29110 195846 29174
rect 195910 29110 196052 29174
rect 195840 29104 196052 29110
rect 196248 29174 196460 29316
rect 196248 29110 196254 29174
rect 196318 29110 196460 29174
rect 196248 29104 196460 29110
rect 196656 29310 196868 29316
rect 196656 29246 196662 29310
rect 196726 29246 196868 29310
rect 196656 29174 196868 29246
rect 196656 29110 196662 29174
rect 196726 29110 196868 29174
rect 196656 29104 196868 29110
rect 198832 29174 199044 29316
rect 198832 29110 198838 29174
rect 198902 29110 199044 29174
rect 198832 29104 199044 29110
rect 199104 29310 199452 29316
rect 199104 29246 199382 29310
rect 199446 29246 199452 29310
rect 199104 29174 199452 29246
rect 199104 29110 199246 29174
rect 199310 29110 199452 29174
rect 199104 29104 199452 29110
rect 199512 29310 199860 29316
rect 199512 29246 199790 29310
rect 199854 29246 199860 29310
rect 199512 29240 199860 29246
rect 199512 29180 199724 29240
rect 199920 29180 200268 29316
rect 199512 29104 200268 29180
rect 200464 29310 200676 29316
rect 200464 29246 200606 29310
rect 200670 29246 200676 29310
rect 200464 29174 200676 29246
rect 200464 29110 200470 29174
rect 200534 29110 200676 29174
rect 200464 29104 200676 29110
rect 216784 29092 216996 29180
rect 216784 29036 216908 29092
rect 216964 29044 216996 29092
rect 216964 29038 217540 29044
rect 216964 29036 217470 29038
rect 216784 28974 217470 29036
rect 217534 28974 217540 29038
rect 216784 28968 217540 28974
rect 28288 28908 28364 28968
rect 190128 28908 190204 28968
rect 21760 28902 21972 28908
rect 21760 28838 21766 28902
rect 21830 28838 21972 28902
rect 21760 28766 21972 28838
rect 21760 28702 21902 28766
rect 21966 28702 21972 28766
rect 21760 28696 21972 28702
rect 22168 28766 22380 28908
rect 22168 28702 22310 28766
rect 22374 28702 22380 28766
rect 22168 28696 22380 28702
rect 22576 28902 22788 28908
rect 22576 28838 22582 28902
rect 22646 28838 22788 28902
rect 22576 28766 22788 28838
rect 22576 28702 22718 28766
rect 22782 28702 22788 28766
rect 22576 28696 22788 28702
rect 22984 28902 23196 28908
rect 22984 28838 23126 28902
rect 23190 28838 23196 28902
rect 22984 28766 23196 28838
rect 22984 28702 22990 28766
rect 23054 28702 23196 28766
rect 22984 28696 23196 28702
rect 23392 28902 23604 28908
rect 23392 28838 23534 28902
rect 23598 28838 23604 28902
rect 23392 28766 23604 28838
rect 23392 28702 23398 28766
rect 23462 28702 23604 28766
rect 23392 28696 23604 28702
rect 28288 28696 28636 28908
rect 190128 28696 190340 28908
rect 195024 28902 195236 28908
rect 195024 28838 195166 28902
rect 195230 28838 195236 28902
rect 195024 28766 195236 28838
rect 195024 28702 195030 28766
rect 195094 28702 195236 28766
rect 195024 28696 195236 28702
rect 195432 28902 195644 28908
rect 195432 28838 195438 28902
rect 195502 28838 195644 28902
rect 195432 28766 195644 28838
rect 195432 28702 195438 28766
rect 195502 28702 195644 28766
rect 195432 28696 195644 28702
rect 195840 28902 196052 28908
rect 195840 28838 195846 28902
rect 195910 28838 196052 28902
rect 195840 28772 196052 28838
rect 196248 28902 196460 28908
rect 196248 28838 196254 28902
rect 196318 28838 196460 28902
rect 196248 28772 196460 28838
rect 195840 28696 196460 28772
rect 196656 28902 196868 28908
rect 196656 28838 196662 28902
rect 196726 28838 196868 28902
rect 196656 28766 196868 28838
rect 196656 28702 196798 28766
rect 196862 28702 196868 28766
rect 196656 28696 196868 28702
rect 28424 28636 28500 28696
rect 190264 28636 190340 28696
rect 196248 28636 196324 28696
rect 18632 28630 18980 28636
rect 18632 28566 18910 28630
rect 18974 28566 18980 28630
rect 18632 28560 18980 28566
rect 18632 28500 18708 28560
rect 18088 28494 18300 28500
rect 18088 28430 18230 28494
rect 18294 28430 18300 28494
rect 18088 28364 18300 28430
rect 18496 28424 19116 28500
rect 18088 28358 18436 28364
rect 18088 28294 18094 28358
rect 18158 28294 18366 28358
rect 18430 28294 18436 28358
rect 18088 28288 18436 28294
rect 18496 28288 18708 28424
rect 18904 28364 19116 28424
rect 19312 28494 19524 28500
rect 19312 28430 19454 28494
rect 19518 28430 19524 28494
rect 18904 28358 19252 28364
rect 18904 28294 19046 28358
rect 19110 28294 19252 28358
rect 18904 28288 19252 28294
rect 19312 28358 19524 28430
rect 19312 28294 19318 28358
rect 19382 28294 19454 28358
rect 19518 28294 19524 28358
rect 19312 28288 19524 28294
rect 19720 28358 19932 28500
rect 19720 28294 19862 28358
rect 19926 28294 19932 28358
rect 19720 28288 19932 28294
rect 21760 28494 21972 28500
rect 21760 28430 21902 28494
rect 21966 28430 21972 28494
rect 21760 28358 21972 28430
rect 21760 28294 21902 28358
rect 21966 28294 21972 28358
rect 21760 28288 21972 28294
rect 22168 28494 22788 28500
rect 22168 28430 22310 28494
rect 22374 28430 22718 28494
rect 22782 28430 22788 28494
rect 22168 28424 22788 28430
rect 22168 28364 22380 28424
rect 22168 28358 22516 28364
rect 22168 28294 22446 28358
rect 22510 28294 22516 28358
rect 22168 28288 22516 28294
rect 22576 28288 22788 28424
rect 22984 28494 23196 28500
rect 22984 28430 22990 28494
rect 23054 28430 23196 28494
rect 22984 28358 23196 28430
rect 22984 28294 22990 28358
rect 23054 28294 23196 28358
rect 22984 28288 23196 28294
rect 23392 28494 23604 28500
rect 23392 28430 23398 28494
rect 23462 28430 23604 28494
rect 23392 28358 23604 28430
rect 28288 28424 28636 28636
rect 190128 28424 190340 28636
rect 195976 28560 196324 28636
rect 198968 28560 199588 28636
rect 195976 28500 196052 28560
rect 198968 28500 199044 28560
rect 199512 28500 199588 28560
rect 28560 28364 28636 28424
rect 190264 28364 190340 28424
rect 23392 28294 23398 28358
rect 23462 28294 23604 28358
rect 23392 28288 23604 28294
rect 19176 28228 19252 28288
rect 19720 28228 19796 28288
rect 2720 28152 3748 28228
rect 19176 28152 19796 28228
rect 28288 28152 28636 28364
rect 190128 28152 190340 28364
rect 195024 28494 195236 28500
rect 195024 28430 195030 28494
rect 195094 28430 195236 28494
rect 195024 28358 195236 28430
rect 195024 28294 195166 28358
rect 195230 28294 195236 28358
rect 195024 28288 195236 28294
rect 195432 28494 195644 28500
rect 195432 28430 195438 28494
rect 195502 28430 195644 28494
rect 195432 28358 195644 28430
rect 195432 28294 195438 28358
rect 195502 28294 195644 28358
rect 195432 28288 195644 28294
rect 195840 28424 196460 28500
rect 195840 28288 196052 28424
rect 196248 28358 196460 28424
rect 196248 28294 196390 28358
rect 196454 28294 196460 28358
rect 196248 28288 196460 28294
rect 196656 28494 196868 28500
rect 196656 28430 196798 28494
rect 196862 28430 196868 28494
rect 196656 28358 196868 28430
rect 196656 28294 196798 28358
rect 196862 28294 196868 28358
rect 196656 28288 196868 28294
rect 198832 28494 199044 28500
rect 198832 28430 198838 28494
rect 198902 28430 199044 28494
rect 198832 28358 199044 28430
rect 198832 28294 198974 28358
rect 199038 28294 199044 28358
rect 198832 28288 199044 28294
rect 199104 28494 199452 28500
rect 199104 28430 199246 28494
rect 199310 28430 199452 28494
rect 199104 28358 199452 28430
rect 199104 28294 199382 28358
rect 199446 28294 199452 28358
rect 199104 28288 199452 28294
rect 199512 28364 199724 28500
rect 199920 28364 200268 28500
rect 199512 28288 200268 28364
rect 200464 28494 200676 28500
rect 200464 28430 200470 28494
rect 200534 28430 200676 28494
rect 200464 28358 200676 28430
rect 200464 28294 200470 28358
rect 200534 28294 200676 28358
rect 200464 28288 200676 28294
rect 199376 28228 199452 28288
rect 200464 28228 200540 28288
rect 199376 28152 200540 28228
rect 2720 28092 2932 28152
rect 1942 28086 2932 28092
rect 1904 28022 1910 28086
rect 1974 28022 2932 28086
rect 1942 28016 2932 28022
rect 3400 28016 3748 28152
rect 28288 28092 28364 28152
rect 190128 28092 190204 28152
rect 18398 28086 19388 28092
rect 18360 28022 18366 28086
rect 18430 28022 19318 28086
rect 19382 28022 19388 28086
rect 18398 28016 19388 28022
rect 21760 28086 21972 28092
rect 21760 28022 21902 28086
rect 21966 28022 21972 28086
rect 21760 27950 21972 28022
rect 21760 27886 21766 27950
rect 21830 27886 21972 27950
rect 21760 27880 21972 27886
rect 22168 27950 22380 28092
rect 22478 28086 22788 28092
rect 22440 28022 22446 28086
rect 22510 28022 22788 28086
rect 22478 28016 22788 28022
rect 22168 27886 22174 27950
rect 22238 27886 22380 27950
rect 22168 27880 22380 27886
rect 22576 27950 22788 28016
rect 22576 27886 22582 27950
rect 22646 27886 22788 27950
rect 22576 27880 22788 27886
rect 22984 28086 23196 28092
rect 22984 28022 22990 28086
rect 23054 28022 23196 28086
rect 22984 27950 23196 28022
rect 22984 27886 23126 27950
rect 23190 27886 23196 27950
rect 22984 27880 23196 27886
rect 23392 28086 23604 28092
rect 23392 28022 23398 28086
rect 23462 28022 23604 28086
rect 23392 27950 23604 28022
rect 23392 27886 23398 27950
rect 23462 27886 23604 27950
rect 23392 27880 23604 27886
rect 28288 27880 28636 28092
rect 190128 27880 190340 28092
rect 195024 28086 195236 28092
rect 195024 28022 195166 28086
rect 195230 28022 195236 28086
rect 195024 27950 195236 28022
rect 195024 27886 195166 27950
rect 195230 27886 195236 27950
rect 195024 27880 195236 27886
rect 195432 28086 195644 28092
rect 195432 28022 195438 28086
rect 195502 28022 195644 28086
rect 195432 27950 195644 28022
rect 195432 27886 195438 27950
rect 195502 27886 195644 27950
rect 195432 27880 195644 27886
rect 195840 27950 196052 28092
rect 195840 27886 195982 27950
rect 196046 27886 196052 27950
rect 195840 27880 196052 27886
rect 196248 28086 196460 28092
rect 196248 28022 196390 28086
rect 196454 28022 196460 28086
rect 196248 27880 196460 28022
rect 196656 28086 196868 28092
rect 196656 28022 196798 28086
rect 196862 28022 196868 28086
rect 196656 27950 196868 28022
rect 196656 27886 196798 27950
rect 196862 27886 196868 27950
rect 196656 27880 196868 27886
rect 28424 27820 28500 27880
rect 190128 27820 190204 27880
rect 196248 27820 196324 27880
rect 16864 27744 18164 27820
rect 16864 27684 16940 27744
rect 18088 27684 18164 27744
rect 19584 27744 21836 27820
rect 19584 27684 19660 27744
rect 21760 27684 21836 27744
rect 16592 27608 16940 27684
rect 1224 27542 1980 27548
rect 1224 27478 1230 27542
rect 1294 27478 1910 27542
rect 1974 27478 1980 27542
rect 1224 27472 1980 27478
rect 16592 27472 16804 27608
rect 17000 27548 17212 27684
rect 18088 27678 18300 27684
rect 18088 27614 18094 27678
rect 18158 27614 18300 27678
rect 17000 27472 18028 27548
rect 18088 27472 18300 27614
rect 18496 27678 19116 27684
rect 18496 27614 19046 27678
rect 19110 27614 19116 27678
rect 18496 27608 19116 27614
rect 18496 27472 18708 27608
rect 18904 27472 19116 27608
rect 19312 27678 19660 27684
rect 19312 27614 19454 27678
rect 19518 27614 19660 27678
rect 19312 27608 19660 27614
rect 19720 27678 19932 27684
rect 19720 27614 19862 27678
rect 19926 27614 19932 27678
rect 19312 27542 19524 27608
rect 19312 27478 19454 27542
rect 19518 27478 19524 27542
rect 19312 27472 19524 27478
rect 19720 27542 19932 27614
rect 19720 27478 19726 27542
rect 19790 27478 19932 27542
rect 19720 27472 19932 27478
rect 21760 27678 21972 27684
rect 21760 27614 21766 27678
rect 21830 27614 21972 27678
rect 21760 27472 21972 27614
rect 22168 27678 22380 27684
rect 22168 27614 22174 27678
rect 22238 27614 22380 27678
rect 22168 27548 22380 27614
rect 22576 27678 22788 27684
rect 22576 27614 22582 27678
rect 22646 27614 22788 27678
rect 22576 27548 22788 27614
rect 22168 27542 22788 27548
rect 22168 27478 22310 27542
rect 22374 27478 22788 27542
rect 22168 27472 22788 27478
rect 22984 27678 23196 27684
rect 22984 27614 23126 27678
rect 23190 27614 23196 27678
rect 22984 27542 23196 27614
rect 22984 27478 23126 27542
rect 23190 27478 23196 27542
rect 22984 27472 23196 27478
rect 23392 27678 23604 27684
rect 23392 27614 23398 27678
rect 23462 27614 23604 27678
rect 23392 27542 23604 27614
rect 28288 27608 28636 27820
rect 190128 27608 190340 27820
rect 195976 27744 196324 27820
rect 198968 27744 199588 27820
rect 195976 27684 196052 27744
rect 198968 27684 199044 27744
rect 199512 27684 199588 27744
rect 200328 27744 201492 27820
rect 200328 27684 200404 27744
rect 201416 27684 201492 27744
rect 28424 27548 28500 27608
rect 190264 27548 190340 27608
rect 23392 27478 23398 27542
rect 23462 27478 23604 27542
rect 23392 27472 23604 27478
rect 1632 27412 1844 27472
rect 1632 27356 1702 27412
rect 1758 27356 1844 27412
rect 1632 27200 1844 27356
rect 17952 27412 18028 27472
rect 18496 27412 18572 27472
rect 21896 27412 21972 27472
rect 17952 27336 18572 27412
rect 21760 27270 21972 27412
rect 22304 27412 22380 27472
rect 22304 27336 22652 27412
rect 28288 27336 28636 27548
rect 190128 27336 190340 27548
rect 195024 27678 195236 27684
rect 195024 27614 195166 27678
rect 195230 27614 195236 27678
rect 195024 27542 195236 27614
rect 195024 27478 195030 27542
rect 195094 27478 195236 27542
rect 195024 27472 195236 27478
rect 195432 27678 195644 27684
rect 195432 27614 195438 27678
rect 195502 27614 195644 27678
rect 195432 27542 195644 27614
rect 195432 27478 195438 27542
rect 195502 27478 195644 27542
rect 195432 27472 195644 27478
rect 195840 27678 196460 27684
rect 195840 27614 195982 27678
rect 196046 27614 196460 27678
rect 195840 27608 196460 27614
rect 195840 27472 196052 27608
rect 196248 27542 196460 27608
rect 196248 27478 196390 27542
rect 196454 27478 196460 27542
rect 196248 27472 196460 27478
rect 196656 27678 196868 27684
rect 196656 27614 196798 27678
rect 196862 27614 196868 27678
rect 196656 27472 196868 27614
rect 198832 27678 199044 27684
rect 198832 27614 198974 27678
rect 199038 27614 199044 27678
rect 198832 27472 199044 27614
rect 199104 27678 199452 27684
rect 199104 27614 199382 27678
rect 199446 27614 199452 27678
rect 199104 27472 199452 27614
rect 199512 27548 199724 27684
rect 199920 27608 200404 27684
rect 200464 27678 200676 27684
rect 200464 27614 200470 27678
rect 200534 27614 200676 27678
rect 199920 27548 200268 27608
rect 199512 27472 200268 27548
rect 200464 27548 200676 27614
rect 200464 27542 201356 27548
rect 200464 27478 200470 27542
rect 200534 27478 201356 27542
rect 200464 27472 201356 27478
rect 201416 27472 201764 27684
rect 201824 27472 202036 27684
rect 196792 27412 196868 27472
rect 199512 27412 199588 27472
rect 22576 27276 22652 27336
rect 28560 27276 28636 27336
rect 190264 27276 190340 27336
rect 21760 27206 21902 27270
rect 21966 27206 21972 27270
rect 21760 27200 21972 27206
rect 22168 27270 22380 27276
rect 22168 27206 22310 27270
rect 22374 27206 22380 27270
rect 22168 27064 22380 27206
rect 22576 27064 22788 27276
rect 22984 27270 23196 27276
rect 22984 27206 23126 27270
rect 23190 27206 23196 27270
rect 22984 27134 23196 27206
rect 22984 27070 23126 27134
rect 23190 27070 23196 27134
rect 22984 27064 23196 27070
rect 23392 27270 23604 27276
rect 23392 27206 23398 27270
rect 23462 27206 23604 27270
rect 23392 27134 23604 27206
rect 23392 27070 23534 27134
rect 23598 27070 23604 27134
rect 23392 27064 23604 27070
rect 22576 27004 22652 27064
rect 21760 26998 21972 27004
rect 21760 26934 21902 26998
rect 21966 26934 21972 26998
rect 2720 26792 3748 26868
rect 2720 26732 2932 26792
rect 544 26726 2932 26732
rect 544 26662 550 26726
rect 614 26662 2932 26726
rect 544 26656 2932 26662
rect 3400 26656 3748 26792
rect 21760 26656 21972 26934
rect 22168 26726 22380 27004
rect 22576 26732 22788 27004
rect 22478 26726 22788 26732
rect 22168 26662 22174 26726
rect 22238 26662 22380 26726
rect 22440 26662 22446 26726
rect 22510 26662 22788 26726
rect 22168 26656 22380 26662
rect 22478 26656 22788 26662
rect 22984 26862 23196 26868
rect 22984 26798 23126 26862
rect 23190 26798 23196 26862
rect 22984 26656 23196 26798
rect 23392 26862 23604 26868
rect 23392 26798 23534 26862
rect 23598 26798 23604 26862
rect 23392 26656 23604 26798
rect 28288 26792 28636 27276
rect 190128 26792 190340 27276
rect 195024 27270 195236 27276
rect 195024 27206 195030 27270
rect 195094 27206 195236 27270
rect 195024 27134 195236 27206
rect 195024 27070 195166 27134
rect 195230 27070 195236 27134
rect 195024 27064 195236 27070
rect 195432 27270 195644 27276
rect 195432 27206 195438 27270
rect 195502 27206 195644 27270
rect 195432 27134 195644 27206
rect 195432 27070 195574 27134
rect 195638 27070 195644 27134
rect 195432 27064 195644 27070
rect 195840 27064 196052 27276
rect 196248 27270 196460 27276
rect 196248 27206 196390 27270
rect 196454 27206 196460 27270
rect 196248 27064 196460 27206
rect 196656 27270 196868 27412
rect 199006 27406 199588 27412
rect 198968 27342 198974 27406
rect 199038 27342 199588 27406
rect 199006 27336 199588 27342
rect 201280 27412 201356 27472
rect 201824 27412 201900 27472
rect 201280 27336 201900 27412
rect 216784 27412 216996 27548
rect 216784 27356 216908 27412
rect 216964 27406 217540 27412
rect 216964 27356 217470 27406
rect 216784 27342 217470 27356
rect 217534 27342 217540 27406
rect 216784 27336 217540 27342
rect 196656 27206 196798 27270
rect 196862 27206 196868 27270
rect 196656 27200 196868 27206
rect 216784 27200 216996 27336
rect 195840 27004 195916 27064
rect 196248 27004 196324 27064
rect 28288 26732 28364 26792
rect 190264 26732 190340 26792
rect 21896 26596 21972 26656
rect 21760 26454 21972 26596
rect 22984 26596 23060 26656
rect 23392 26596 23468 26656
rect 21760 26390 21902 26454
rect 21966 26390 21972 26454
rect 21760 26384 21972 26390
rect 22168 26454 22516 26460
rect 22168 26390 22174 26454
rect 22238 26390 22446 26454
rect 22510 26390 22516 26454
rect 22168 26384 22516 26390
rect 22168 26324 22380 26384
rect 19176 26248 19796 26324
rect 22168 26248 22516 26324
rect 22576 26248 22788 26460
rect 19176 26188 19252 26248
rect 19720 26188 19796 26248
rect 22304 26188 22380 26248
rect 18496 26046 18708 26188
rect 18496 25982 18638 26046
rect 18702 25982 18708 26046
rect 18496 25976 18708 25982
rect 18904 26112 19252 26188
rect 19312 26182 19524 26188
rect 19312 26118 19454 26182
rect 19518 26118 19524 26182
rect 18904 25976 19116 26112
rect 19312 25910 19524 26118
rect 19312 25846 19454 25910
rect 19518 25846 19524 25910
rect 19312 25840 19524 25846
rect 19720 26182 19932 26188
rect 19720 26118 19726 26182
rect 19790 26118 19932 26182
rect 19720 25910 19932 26118
rect 21760 26182 21972 26188
rect 21760 26118 21902 26182
rect 21966 26118 21972 26182
rect 21760 26046 21972 26118
rect 21760 25982 21766 26046
rect 21830 25982 21972 26046
rect 21760 25976 21972 25982
rect 22168 26046 22380 26188
rect 22440 26188 22516 26248
rect 22712 26188 22788 26248
rect 22440 26112 22788 26188
rect 22168 25982 22174 26046
rect 22238 25982 22380 26046
rect 22168 25976 22380 25982
rect 22576 26046 22788 26112
rect 22576 25982 22582 26046
rect 22646 25982 22788 26046
rect 22576 25976 22788 25982
rect 22984 26248 23196 26596
rect 23392 26248 23604 26596
rect 28288 26590 28636 26732
rect 28288 26526 28566 26590
rect 28630 26526 28636 26590
rect 28288 26318 28636 26526
rect 28288 26254 28566 26318
rect 28630 26254 28636 26318
rect 22984 26188 23060 26248
rect 23392 26188 23468 26248
rect 19720 25846 19726 25910
rect 19790 25846 19932 25910
rect 19720 25840 19932 25846
rect 22984 25840 23196 26188
rect 23392 25840 23604 26188
rect 28288 26182 28636 26254
rect 28288 26118 28430 26182
rect 28494 26118 28636 26182
rect 28288 26112 28636 26118
rect 190128 26590 190340 26732
rect 195024 26862 195236 26868
rect 195024 26798 195166 26862
rect 195230 26798 195236 26862
rect 195024 26656 195236 26798
rect 195160 26596 195236 26656
rect 190128 26526 190270 26590
rect 190334 26526 190340 26590
rect 190128 26318 190340 26526
rect 190128 26254 190270 26318
rect 190334 26254 190340 26318
rect 190128 26182 190340 26254
rect 195024 26248 195236 26596
rect 195160 26188 195236 26248
rect 190128 26118 190270 26182
rect 190334 26118 190340 26182
rect 190128 26112 190340 26118
rect 23120 25780 23196 25840
rect 23528 25780 23604 25840
rect 1632 25732 1844 25780
rect 1632 25676 1702 25732
rect 1758 25676 1844 25732
rect 1632 25644 1844 25676
rect 21760 25774 21972 25780
rect 21760 25710 21766 25774
rect 21830 25710 21972 25774
rect 1224 25638 2796 25644
rect 18806 25638 19388 25644
rect 1224 25574 1230 25638
rect 1294 25574 2796 25638
rect 18768 25574 18774 25638
rect 18838 25574 19318 25638
rect 19382 25574 19388 25638
rect 1224 25568 2796 25574
rect 18806 25568 19388 25574
rect 21760 25638 21972 25710
rect 21760 25574 21902 25638
rect 21966 25574 21972 25638
rect 21760 25568 21972 25574
rect 22168 25774 22380 25780
rect 22168 25710 22174 25774
rect 22238 25710 22380 25774
rect 2720 25508 2796 25568
rect 2720 25236 2932 25508
rect 3400 25236 3748 25508
rect 17408 25432 18572 25508
rect 17408 25372 17484 25432
rect 18496 25372 18572 25432
rect 19176 25502 19796 25508
rect 19176 25438 19726 25502
rect 19790 25438 19796 25502
rect 19176 25432 19796 25438
rect 22168 25432 22380 25710
rect 22576 25774 22788 25780
rect 22576 25710 22582 25774
rect 22646 25710 22788 25774
rect 22576 25508 22788 25710
rect 22984 25638 23196 25780
rect 22984 25574 23126 25638
rect 23190 25574 23196 25638
rect 22984 25568 23196 25574
rect 23392 25638 23604 25780
rect 23392 25574 23398 25638
rect 23462 25574 23604 25638
rect 23392 25568 23604 25574
rect 28288 25910 28636 25916
rect 28288 25846 28430 25910
rect 28494 25846 28636 25910
rect 28288 25774 28636 25846
rect 28288 25710 28294 25774
rect 28358 25710 28636 25774
rect 28288 25568 28636 25710
rect 190128 25910 190340 25916
rect 190128 25846 190270 25910
rect 190334 25846 190340 25910
rect 190128 25568 190340 25846
rect 195024 25840 195236 26188
rect 195432 26862 195644 26868
rect 195432 26798 195574 26862
rect 195638 26798 195644 26862
rect 195432 26656 195644 26798
rect 195840 26732 196052 27004
rect 196248 26732 196460 27004
rect 195840 26726 196460 26732
rect 195840 26662 196390 26726
rect 196454 26662 196460 26726
rect 195840 26656 196460 26662
rect 196656 26998 196868 27004
rect 196656 26934 196798 26998
rect 196862 26934 196868 26998
rect 196656 26656 196868 26934
rect 195432 26596 195508 26656
rect 196656 26596 196732 26656
rect 195432 26248 195644 26596
rect 195840 26324 196052 26460
rect 196248 26454 196460 26460
rect 196248 26390 196390 26454
rect 196454 26390 196460 26454
rect 195840 26248 196188 26324
rect 195432 26188 195508 26248
rect 195976 26188 196052 26248
rect 195432 25840 195644 26188
rect 195840 25976 196052 26188
rect 196112 26188 196188 26248
rect 196248 26248 196460 26390
rect 196656 26454 196868 26596
rect 196656 26390 196798 26454
rect 196862 26390 196868 26454
rect 196656 26384 196868 26390
rect 198968 26248 199588 26324
rect 196248 26188 196324 26248
rect 198968 26188 199044 26248
rect 199512 26188 199588 26248
rect 196112 26112 196460 26188
rect 196248 26046 196460 26112
rect 196248 25982 196254 26046
rect 196318 25982 196460 26046
rect 196248 25976 196460 25982
rect 196656 26182 196868 26188
rect 196656 26118 196798 26182
rect 196862 26118 196868 26182
rect 196656 26046 196868 26118
rect 196656 25982 196662 26046
rect 196726 25982 196868 26046
rect 196656 25976 196868 25982
rect 198832 26182 199044 26188
rect 198832 26118 198974 26182
rect 199038 26118 199044 26182
rect 198832 25840 199044 26118
rect 199104 25910 199452 26188
rect 199512 26046 199724 26188
rect 199512 25982 199654 26046
rect 199718 25982 199724 26046
rect 199512 25976 199724 25982
rect 199920 26182 200540 26188
rect 199920 26118 200470 26182
rect 200534 26118 200540 26182
rect 199920 26112 200540 26118
rect 199920 26052 200268 26112
rect 199920 26046 201356 26052
rect 199920 25982 200198 26046
rect 200262 25982 201286 26046
rect 201350 25982 201356 26046
rect 199920 25976 201356 25982
rect 199104 25846 199382 25910
rect 199446 25846 199452 25910
rect 199104 25840 199452 25846
rect 195160 25780 195236 25840
rect 195568 25780 195644 25840
rect 195024 25638 195236 25780
rect 195024 25574 195030 25638
rect 195094 25574 195236 25638
rect 195024 25568 195236 25574
rect 195432 25638 195644 25780
rect 195432 25574 195438 25638
rect 195502 25574 195644 25638
rect 195432 25568 195644 25574
rect 22440 25432 22788 25508
rect 28288 25508 28364 25568
rect 190128 25508 190204 25568
rect 28288 25502 28636 25508
rect 28288 25438 28294 25502
rect 28358 25438 28636 25502
rect 19176 25372 19252 25432
rect 22440 25372 22516 25432
rect 2720 25160 3748 25236
rect 17136 25296 17484 25372
rect 17136 25230 17348 25296
rect 17136 25166 17142 25230
rect 17206 25166 17348 25230
rect 17136 25160 17348 25166
rect 17544 25236 17756 25372
rect 18496 25366 18844 25372
rect 18496 25302 18638 25366
rect 18702 25302 18774 25366
rect 18838 25302 18844 25366
rect 18496 25296 18844 25302
rect 18904 25296 19252 25372
rect 19312 25366 19524 25372
rect 19312 25302 19318 25366
rect 19382 25302 19454 25366
rect 19518 25302 19524 25366
rect 17544 25230 18436 25236
rect 17544 25166 17550 25230
rect 17614 25166 18436 25230
rect 17544 25160 18436 25166
rect 18496 25160 18708 25296
rect 18904 25236 19116 25296
rect 18904 25160 19252 25236
rect 19312 25160 19524 25302
rect 19720 25160 19932 25372
rect 21760 25366 21972 25372
rect 21760 25302 21902 25366
rect 21966 25302 21972 25366
rect 21760 25230 21972 25302
rect 21760 25166 21902 25230
rect 21966 25166 21972 25230
rect 21760 25160 21972 25166
rect 22168 25296 22516 25372
rect 22168 25236 22380 25296
rect 22576 25236 22788 25372
rect 22168 25160 22788 25236
rect 22984 25366 23196 25372
rect 22984 25302 23126 25366
rect 23190 25302 23196 25366
rect 22984 25160 23196 25302
rect 23392 25366 23604 25372
rect 23392 25302 23398 25366
rect 23462 25302 23604 25366
rect 23392 25230 23604 25302
rect 28288 25296 28636 25438
rect 190128 25296 190340 25508
rect 195840 25432 196052 25780
rect 196248 25774 196460 25780
rect 196248 25710 196254 25774
rect 196318 25710 196460 25774
rect 196248 25508 196460 25710
rect 196656 25774 196868 25780
rect 196656 25710 196662 25774
rect 196726 25710 196868 25774
rect 196656 25638 196868 25710
rect 196656 25574 196662 25638
rect 196726 25574 196868 25638
rect 196656 25568 196868 25574
rect 216784 25774 217540 25780
rect 216784 25732 217470 25774
rect 216784 25676 216908 25732
rect 216964 25710 217470 25732
rect 217534 25710 217540 25774
rect 216964 25704 217540 25710
rect 216964 25676 216996 25704
rect 216784 25568 216996 25676
rect 195976 25372 196052 25432
rect 196112 25432 196460 25508
rect 196112 25372 196188 25432
rect 196384 25372 196460 25432
rect 199784 25432 200948 25508
rect 199784 25372 199860 25432
rect 200872 25372 200948 25432
rect 28424 25236 28500 25296
rect 190264 25236 190340 25296
rect 23392 25166 23398 25230
rect 23462 25166 23604 25230
rect 23392 25160 23604 25166
rect 18360 25100 18436 25160
rect 18904 25100 18980 25160
rect 18360 25024 18980 25100
rect 19176 25100 19252 25160
rect 19720 25100 19796 25160
rect 19176 25024 19796 25100
rect 28288 25024 28636 25236
rect 190128 25024 190340 25236
rect 195024 25366 195236 25372
rect 195024 25302 195030 25366
rect 195094 25302 195236 25366
rect 195024 25230 195236 25302
rect 195024 25166 195030 25230
rect 195094 25166 195236 25230
rect 195024 25160 195236 25166
rect 195432 25366 195644 25372
rect 195432 25302 195438 25366
rect 195502 25302 195644 25366
rect 195432 25160 195644 25302
rect 195840 25296 196188 25372
rect 195840 25160 196052 25296
rect 196248 25160 196460 25372
rect 196656 25366 196868 25372
rect 196656 25302 196662 25366
rect 196726 25302 196868 25366
rect 196656 25160 196868 25302
rect 198832 25160 199044 25372
rect 199104 25366 199452 25372
rect 199104 25302 199382 25366
rect 199446 25302 199452 25366
rect 199104 25230 199452 25302
rect 199104 25166 199382 25230
rect 199446 25166 199452 25230
rect 199104 25160 199452 25166
rect 199512 25366 199860 25372
rect 199512 25302 199654 25366
rect 199718 25302 199860 25366
rect 199512 25296 199860 25302
rect 199920 25366 200268 25372
rect 199920 25302 200198 25366
rect 200262 25302 200268 25366
rect 199512 25160 199724 25296
rect 199920 25230 200268 25302
rect 199920 25166 199926 25230
rect 199990 25166 200268 25230
rect 199920 25160 200268 25166
rect 200872 25236 201084 25372
rect 201280 25366 201492 25372
rect 201280 25302 201286 25366
rect 201350 25302 201492 25366
rect 201280 25236 201492 25302
rect 200872 25230 201220 25236
rect 200872 25166 201150 25230
rect 201214 25166 201220 25230
rect 200872 25160 201220 25166
rect 201280 25230 204076 25236
rect 201280 25166 204006 25230
rect 204070 25166 204076 25230
rect 201280 25160 204076 25166
rect 198968 25100 199044 25160
rect 199512 25100 199588 25160
rect 198968 25024 199588 25100
rect 28288 24964 28364 25024
rect 190264 24964 190340 25024
rect 28288 24828 28636 24964
rect 23392 24822 24556 24828
rect 23392 24758 23398 24822
rect 23462 24758 24556 24822
rect 23392 24752 24556 24758
rect 23392 24556 23604 24752
rect 23158 24550 23604 24556
rect 23120 24486 23126 24550
rect 23190 24486 23604 24550
rect 23158 24480 23604 24486
rect 24208 24692 24556 24752
rect 28016 24752 28636 24828
rect 190128 24828 190340 24964
rect 199414 24958 199996 24964
rect 199376 24894 199382 24958
rect 199446 24894 199926 24958
rect 199990 24894 199996 24958
rect 199414 24888 199996 24894
rect 204000 24958 204212 24964
rect 204000 24894 204006 24958
rect 204070 24894 204212 24958
rect 190128 24752 190748 24828
rect 204000 24822 204212 24894
rect 204000 24758 204142 24822
rect 204206 24758 204212 24822
rect 204000 24752 204212 24758
rect 28016 24692 28228 24752
rect 24208 24616 27140 24692
rect 28016 24686 29996 24692
rect 28016 24622 29926 24686
rect 29990 24622 29996 24686
rect 28016 24616 29996 24622
rect 190400 24616 190748 24752
rect 24208 24480 24556 24616
rect 26928 24556 27140 24616
rect 203428 24562 203512 24566
rect 203395 24557 203512 24562
rect 26928 24480 29044 24556
rect 203395 24501 203400 24557
rect 203456 24501 203512 24557
rect 203395 24496 203512 24501
rect 203428 24492 203512 24496
rect 28968 24420 29044 24480
rect 28968 24284 29316 24420
rect 29414 24414 30540 24420
rect 30638 24414 31084 24420
rect 29376 24350 29382 24414
rect 29446 24350 30540 24414
rect 30600 24350 30606 24414
rect 30670 24350 31084 24414
rect 29414 24344 30540 24350
rect 30638 24344 31084 24350
rect 29648 24284 29860 24344
rect 28968 24208 29860 24284
rect 30328 24284 30540 24344
rect 30872 24284 31084 24344
rect 31552 24344 32988 24420
rect 31552 24284 31764 24344
rect 30328 24208 31764 24284
rect 32096 24278 32444 24344
rect 32096 24214 32238 24278
rect 32302 24214 32444 24278
rect 32096 24208 32444 24214
rect 32776 24278 32988 24344
rect 32776 24214 32918 24278
rect 32982 24214 32988 24278
rect 32776 24208 32988 24214
rect 33456 24344 34892 24420
rect 33456 24278 33668 24344
rect 33456 24214 33462 24278
rect 33526 24214 33668 24278
rect 33456 24208 33668 24214
rect 34000 24278 34212 24344
rect 34000 24214 34142 24278
rect 34206 24214 34212 24278
rect 34000 24208 34212 24214
rect 34680 24284 34892 24344
rect 35224 24284 35572 24420
rect 35904 24344 36796 24420
rect 35904 24284 36116 24344
rect 34680 24278 36116 24284
rect 34680 24214 35502 24278
rect 35566 24214 36116 24278
rect 34680 24208 36116 24214
rect 36584 24284 36796 24344
rect 37128 24284 37340 24420
rect 37808 24344 39244 24420
rect 39342 24414 39924 24420
rect 39304 24350 39310 24414
rect 39374 24350 39924 24414
rect 39342 24344 39924 24350
rect 37808 24284 38020 24344
rect 36584 24278 38020 24284
rect 36584 24214 37134 24278
rect 37198 24214 38020 24278
rect 36584 24208 38020 24214
rect 38352 24278 38564 24344
rect 38352 24214 38494 24278
rect 38558 24214 38564 24278
rect 38352 24208 38564 24214
rect 39032 24284 39244 24344
rect 39576 24284 39924 24344
rect 40256 24344 41148 24420
rect 40256 24284 40468 24344
rect 39032 24208 40468 24284
rect 40936 24284 41148 24344
rect 41480 24284 41692 24420
rect 42160 24344 43596 24420
rect 42160 24284 42372 24344
rect 40936 24278 42372 24284
rect 40936 24214 40942 24278
rect 41006 24214 41622 24278
rect 41686 24214 42372 24278
rect 40936 24208 42372 24214
rect 42704 24278 43052 24344
rect 42704 24214 42846 24278
rect 42910 24214 43052 24278
rect 42704 24208 43052 24214
rect 43384 24284 43596 24344
rect 44064 24344 45500 24420
rect 44064 24284 44276 24344
rect 43384 24208 44276 24284
rect 44608 24278 44820 24344
rect 44608 24214 44614 24278
rect 44678 24214 44820 24278
rect 44608 24208 44820 24214
rect 45288 24284 45500 24344
rect 45832 24284 46180 24420
rect 46512 24344 47404 24420
rect 46512 24284 46724 24344
rect 45288 24278 46724 24284
rect 45288 24214 45430 24278
rect 45494 24214 46724 24278
rect 45288 24208 46724 24214
rect 47192 24284 47404 24344
rect 47736 24284 47948 24420
rect 48416 24344 49852 24420
rect 48416 24284 48628 24344
rect 47192 24278 47948 24284
rect 48046 24278 48628 24284
rect 47192 24214 47198 24278
rect 47262 24214 47948 24278
rect 48008 24214 48014 24278
rect 48078 24214 48628 24278
rect 47192 24208 47948 24214
rect 48046 24208 48628 24214
rect 48960 24208 49172 24344
rect 49640 24284 49852 24344
rect 50184 24284 50532 24420
rect 49640 24278 50532 24284
rect 49640 24214 49646 24278
rect 49710 24214 50462 24278
rect 50526 24214 50532 24278
rect 49640 24208 50532 24214
rect 50864 24344 51756 24420
rect 50864 24278 51076 24344
rect 50864 24214 50870 24278
rect 50934 24214 51076 24278
rect 50864 24208 51076 24214
rect 51544 24284 51756 24344
rect 52088 24284 52300 24420
rect 52768 24344 53660 24420
rect 52768 24284 52980 24344
rect 51544 24278 52980 24284
rect 51544 24214 51686 24278
rect 51750 24214 52910 24278
rect 52974 24214 52980 24278
rect 51544 24208 52980 24214
rect 53312 24284 53660 24344
rect 53992 24284 54204 24420
rect 54672 24344 56108 24420
rect 54672 24284 54884 24344
rect 53312 24278 54884 24284
rect 53312 24214 54678 24278
rect 54742 24214 54884 24278
rect 53312 24208 54884 24214
rect 55216 24278 55428 24344
rect 55216 24214 55358 24278
rect 55422 24214 55428 24278
rect 55216 24208 55428 24214
rect 55896 24284 56108 24344
rect 56440 24284 56788 24420
rect 57120 24344 58012 24420
rect 58110 24414 58556 24420
rect 58072 24350 58078 24414
rect 58142 24350 58556 24414
rect 58110 24344 58556 24350
rect 57120 24284 57332 24344
rect 55896 24278 57332 24284
rect 55896 24214 56582 24278
rect 56646 24214 57332 24278
rect 55896 24208 57332 24214
rect 57800 24284 58012 24344
rect 58344 24284 58556 24344
rect 59024 24344 60460 24420
rect 59024 24284 59236 24344
rect 57800 24208 59236 24284
rect 59568 24278 59780 24344
rect 59568 24214 59710 24278
rect 59774 24214 59780 24278
rect 59568 24208 59780 24214
rect 60248 24284 60460 24344
rect 60792 24284 61140 24420
rect 61472 24284 61684 24420
rect 60248 24278 61684 24284
rect 60248 24214 60390 24278
rect 60454 24214 61614 24278
rect 61678 24214 61684 24278
rect 60248 24208 61684 24214
rect 62152 24284 62364 24420
rect 62696 24284 62908 24420
rect 63376 24344 64812 24420
rect 63376 24284 63588 24344
rect 62152 24278 63588 24284
rect 62152 24214 62158 24278
rect 62222 24214 62838 24278
rect 62902 24214 63588 24278
rect 62152 24208 63588 24214
rect 63920 24278 64268 24344
rect 63920 24214 64062 24278
rect 64126 24214 64268 24278
rect 63920 24208 64268 24214
rect 64600 24284 64812 24344
rect 65280 24344 66716 24420
rect 65280 24284 65492 24344
rect 64600 24208 65492 24284
rect 65824 24208 66036 24344
rect 66504 24284 66716 24344
rect 67048 24284 67396 24420
rect 67728 24284 67940 24420
rect 66504 24278 67940 24284
rect 66504 24214 66646 24278
rect 66710 24214 67870 24278
rect 67934 24214 67940 24278
rect 66504 24208 67940 24214
rect 68408 24284 68620 24420
rect 68952 24284 69164 24420
rect 68408 24278 69164 24284
rect 68408 24214 68414 24278
rect 68478 24214 69094 24278
rect 69158 24214 69164 24278
rect 68408 24208 69164 24214
rect 69632 24344 70388 24420
rect 69632 24278 69844 24344
rect 69632 24214 69638 24278
rect 69702 24214 69844 24278
rect 69632 24208 69844 24214
rect 70176 24278 70388 24344
rect 70176 24214 70318 24278
rect 70382 24214 70388 24278
rect 70176 24208 70388 24214
rect 70856 24284 71068 24420
rect 71400 24284 71748 24420
rect 72080 24344 72972 24420
rect 72080 24284 72292 24344
rect 70856 24278 72292 24284
rect 70856 24214 70862 24278
rect 70926 24214 71678 24278
rect 71742 24214 72292 24278
rect 70856 24208 72292 24214
rect 72760 24284 72972 24344
rect 73304 24284 73516 24420
rect 73984 24344 74876 24420
rect 73984 24284 74196 24344
rect 72760 24278 74196 24284
rect 72760 24214 73446 24278
rect 73510 24214 74196 24278
rect 72760 24208 74196 24214
rect 74528 24278 74876 24344
rect 74528 24214 74670 24278
rect 74734 24214 74876 24278
rect 74528 24208 74876 24214
rect 75208 24278 75420 24420
rect 75208 24214 75214 24278
rect 75278 24214 75420 24278
rect 75208 24208 75420 24214
rect 75888 24344 77324 24420
rect 75888 24278 76100 24344
rect 75888 24214 75894 24278
rect 75958 24214 76100 24278
rect 75888 24208 76100 24214
rect 76432 24278 76644 24344
rect 76432 24214 76574 24278
rect 76638 24214 76644 24278
rect 76432 24208 76644 24214
rect 77112 24284 77324 24344
rect 77656 24284 78004 24420
rect 78336 24344 79228 24420
rect 78336 24284 78548 24344
rect 77112 24278 78548 24284
rect 77112 24214 78342 24278
rect 78406 24214 78548 24278
rect 77112 24208 78548 24214
rect 79016 24284 79228 24344
rect 79560 24284 79772 24420
rect 80240 24344 80996 24420
rect 80240 24284 80452 24344
rect 80784 24284 80996 24344
rect 79016 24278 80452 24284
rect 80550 24278 80996 24284
rect 79016 24214 79566 24278
rect 79630 24214 80452 24278
rect 80512 24214 80518 24278
rect 80582 24214 80996 24278
rect 79016 24208 80452 24214
rect 80550 24208 80996 24214
rect 81464 24284 81676 24420
rect 82008 24284 82356 24420
rect 82688 24344 83580 24420
rect 82688 24284 82900 24344
rect 81464 24278 82900 24284
rect 81464 24214 82014 24278
rect 82078 24214 82900 24278
rect 81464 24208 82900 24214
rect 83368 24284 83580 24344
rect 83912 24284 84124 24420
rect 84592 24344 86028 24420
rect 84592 24284 84804 24344
rect 83368 24278 84804 24284
rect 83368 24214 83374 24278
rect 83438 24214 84598 24278
rect 84662 24214 84804 24278
rect 83368 24208 84804 24214
rect 85136 24284 85484 24344
rect 85816 24284 86028 24344
rect 86496 24344 87932 24420
rect 86496 24284 86708 24344
rect 85136 24278 85756 24284
rect 85136 24214 85686 24278
rect 85750 24214 85756 24278
rect 85136 24208 85756 24214
rect 85816 24278 86708 24284
rect 85816 24214 86502 24278
rect 86566 24214 86708 24278
rect 85816 24208 86708 24214
rect 87040 24208 87252 24344
rect 87720 24284 87932 24344
rect 88264 24284 88612 24420
rect 88944 24344 89836 24420
rect 88944 24284 89156 24344
rect 87720 24278 89156 24284
rect 87720 24214 88406 24278
rect 88470 24214 89086 24278
rect 89150 24214 89156 24278
rect 87720 24208 89156 24214
rect 89624 24284 89836 24344
rect 90168 24284 90380 24420
rect 90848 24344 92284 24420
rect 90848 24284 91060 24344
rect 89624 24278 91060 24284
rect 89624 24214 89766 24278
rect 89830 24214 91060 24278
rect 89624 24208 91060 24214
rect 91392 24208 91604 24344
rect 92072 24284 92284 24344
rect 92616 24284 92964 24420
rect 93296 24344 94188 24420
rect 93296 24284 93508 24344
rect 92072 24278 93508 24284
rect 92072 24214 92078 24278
rect 92142 24214 93508 24278
rect 92072 24208 93508 24214
rect 93976 24284 94188 24344
rect 94520 24284 94732 24420
rect 95200 24284 95412 24420
rect 93976 24278 95412 24284
rect 93976 24214 94662 24278
rect 94726 24214 95342 24278
rect 95406 24214 95412 24278
rect 93976 24208 95412 24214
rect 95744 24344 96636 24420
rect 95744 24278 96092 24344
rect 95744 24214 95750 24278
rect 95814 24214 96092 24278
rect 95744 24208 96092 24214
rect 96424 24284 96636 24344
rect 97104 24344 98540 24420
rect 97104 24284 97316 24344
rect 96424 24278 97316 24284
rect 96424 24214 97110 24278
rect 97174 24214 97316 24278
rect 96424 24208 97316 24214
rect 97648 24278 97860 24344
rect 97648 24214 97790 24278
rect 97854 24214 97860 24278
rect 97648 24208 97860 24214
rect 98328 24284 98540 24344
rect 98872 24344 100444 24420
rect 98872 24284 99220 24344
rect 98328 24208 99220 24284
rect 99552 24208 99764 24344
rect 100232 24284 100444 24344
rect 100776 24284 100988 24420
rect 101456 24284 101668 24420
rect 100232 24278 101668 24284
rect 100232 24214 100782 24278
rect 100846 24214 101598 24278
rect 101662 24214 101668 24278
rect 100232 24208 101668 24214
rect 102000 24344 102892 24420
rect 102000 24278 102212 24344
rect 102000 24214 102142 24278
rect 102206 24214 102212 24278
rect 102000 24208 102212 24214
rect 102680 24284 102892 24344
rect 103224 24344 104116 24420
rect 103224 24284 103572 24344
rect 102680 24278 103572 24284
rect 102680 24214 103366 24278
rect 103430 24214 103572 24278
rect 102680 24208 103572 24214
rect 103904 24278 104116 24344
rect 103904 24214 104046 24278
rect 104110 24214 104116 24278
rect 103904 24208 104116 24214
rect 104584 24284 104796 24420
rect 105128 24284 105340 24420
rect 105808 24344 107244 24420
rect 105808 24284 106020 24344
rect 104584 24278 106020 24284
rect 104584 24214 104590 24278
rect 104654 24214 105270 24278
rect 105334 24214 106020 24278
rect 104584 24208 106020 24214
rect 106352 24208 106700 24344
rect 107032 24284 107244 24344
rect 107712 24344 109148 24420
rect 107712 24284 107924 24344
rect 107032 24208 107924 24284
rect 108256 24208 108468 24344
rect 108936 24284 109148 24344
rect 109480 24284 109828 24420
rect 110160 24284 110372 24420
rect 108936 24278 110372 24284
rect 108936 24214 109622 24278
rect 109686 24214 110302 24278
rect 110366 24214 110372 24278
rect 108936 24208 110372 24214
rect 110840 24284 111052 24420
rect 111384 24284 111596 24420
rect 112064 24344 112820 24420
rect 112064 24284 112276 24344
rect 110840 24278 112276 24284
rect 110840 24214 110846 24278
rect 110910 24214 111526 24278
rect 111590 24214 112276 24278
rect 110840 24208 112276 24214
rect 112608 24278 112820 24344
rect 112608 24214 112750 24278
rect 112814 24214 112820 24278
rect 112608 24208 112820 24214
rect 113288 24284 113500 24420
rect 113832 24284 114180 24420
rect 114278 24414 115404 24420
rect 114240 24350 114246 24414
rect 114310 24350 115404 24414
rect 114278 24344 115404 24350
rect 114512 24284 114724 24344
rect 113288 24278 114724 24284
rect 113288 24214 113294 24278
rect 113358 24214 114724 24278
rect 113288 24208 114724 24214
rect 115192 24284 115404 24344
rect 115736 24284 115948 24420
rect 116416 24344 117308 24420
rect 116416 24284 116628 24344
rect 115192 24278 116628 24284
rect 115192 24214 115334 24278
rect 115398 24214 116628 24278
rect 115192 24208 116628 24214
rect 116960 24278 117308 24344
rect 116960 24214 117102 24278
rect 117166 24214 117308 24278
rect 116960 24208 117308 24214
rect 117640 24284 117852 24420
rect 118320 24344 119756 24420
rect 118320 24284 118532 24344
rect 117640 24278 118532 24284
rect 117640 24214 117646 24278
rect 117710 24214 118532 24278
rect 117640 24208 118532 24214
rect 118864 24278 119076 24344
rect 118864 24214 119006 24278
rect 119070 24214 119076 24278
rect 118864 24208 119076 24214
rect 119544 24284 119756 24344
rect 120088 24284 120436 24420
rect 120768 24344 121660 24420
rect 120768 24284 120980 24344
rect 119544 24278 120980 24284
rect 119544 24214 120230 24278
rect 120294 24214 120980 24278
rect 119544 24208 120980 24214
rect 121448 24284 121660 24344
rect 121992 24284 122204 24420
rect 122672 24344 123428 24420
rect 122672 24284 122884 24344
rect 123216 24284 123428 24344
rect 121448 24278 122884 24284
rect 122982 24278 123428 24284
rect 121448 24214 121998 24278
rect 122062 24214 122884 24278
rect 122944 24214 122950 24278
rect 123014 24214 123428 24278
rect 121448 24208 122884 24214
rect 122982 24208 123428 24214
rect 123896 24284 124108 24420
rect 124440 24284 124788 24420
rect 125120 24344 126012 24420
rect 125120 24284 125332 24344
rect 123896 24278 125332 24284
rect 123896 24214 123902 24278
rect 123966 24214 124446 24278
rect 124510 24214 125332 24278
rect 123896 24208 125332 24214
rect 125800 24284 126012 24344
rect 126344 24284 126556 24420
rect 125800 24278 126556 24284
rect 125800 24214 125806 24278
rect 125870 24214 126556 24278
rect 125800 24208 126556 24214
rect 127024 24344 128460 24420
rect 127024 24278 127236 24344
rect 127024 24214 127030 24278
rect 127094 24214 127236 24278
rect 127024 24208 127236 24214
rect 127568 24208 127916 24344
rect 128248 24284 128460 24344
rect 128928 24344 130364 24420
rect 128928 24284 129140 24344
rect 128248 24278 129140 24284
rect 128248 24214 128934 24278
rect 128998 24214 129140 24278
rect 128248 24208 129140 24214
rect 129472 24208 129684 24344
rect 130152 24284 130364 24344
rect 130696 24344 132268 24420
rect 130696 24284 131044 24344
rect 130152 24278 131044 24284
rect 130152 24214 130294 24278
rect 130358 24214 131044 24278
rect 130152 24208 131044 24214
rect 131376 24208 131588 24344
rect 132056 24284 132268 24344
rect 132600 24284 132812 24420
rect 131686 24278 132812 24284
rect 131648 24214 131654 24278
rect 131718 24214 132812 24278
rect 131686 24208 132812 24214
rect 133280 24344 134716 24420
rect 133280 24278 133492 24344
rect 133280 24214 133286 24278
rect 133350 24214 133492 24278
rect 133280 24208 133492 24214
rect 133824 24208 134036 24344
rect 134504 24284 134716 24344
rect 135048 24284 135396 24420
rect 134504 24278 135396 24284
rect 134504 24214 134510 24278
rect 134574 24214 135190 24278
rect 135254 24214 135396 24278
rect 134504 24208 135396 24214
rect 135728 24344 136620 24420
rect 136718 24414 137164 24420
rect 136680 24350 136686 24414
rect 136750 24350 137164 24414
rect 136718 24344 137164 24350
rect 135728 24278 135940 24344
rect 135728 24214 135734 24278
rect 135798 24214 135940 24278
rect 135728 24208 135940 24214
rect 136408 24284 136620 24344
rect 136952 24284 137164 24344
rect 137632 24344 139068 24420
rect 137632 24284 137844 24344
rect 136408 24208 137844 24284
rect 138176 24278 138524 24344
rect 138176 24214 138182 24278
rect 138246 24214 138524 24278
rect 138176 24208 138524 24214
rect 138856 24284 139068 24344
rect 139536 24344 140972 24420
rect 139536 24284 139748 24344
rect 138856 24278 139748 24284
rect 138856 24214 139542 24278
rect 139606 24214 139748 24278
rect 138856 24208 139748 24214
rect 140080 24278 140292 24344
rect 140080 24214 140222 24278
rect 140286 24214 140292 24278
rect 140080 24208 140292 24214
rect 140760 24284 140972 24344
rect 141304 24344 142876 24420
rect 141304 24284 141652 24344
rect 140760 24278 141924 24284
rect 140760 24214 141854 24278
rect 141918 24214 141924 24278
rect 140760 24208 141924 24214
rect 141984 24208 142196 24344
rect 142664 24284 142876 24344
rect 143208 24284 143420 24420
rect 143888 24344 145324 24420
rect 145422 24414 146004 24420
rect 145384 24350 145390 24414
rect 145454 24350 146004 24414
rect 145422 24344 146004 24350
rect 143888 24284 144100 24344
rect 142664 24278 144100 24284
rect 142664 24214 143214 24278
rect 143278 24214 144030 24278
rect 144094 24214 144100 24278
rect 142664 24208 144100 24214
rect 144432 24208 144644 24344
rect 145112 24284 145324 24344
rect 145656 24284 146004 24344
rect 146336 24284 146548 24420
rect 145112 24278 146548 24284
rect 145112 24214 146478 24278
rect 146542 24214 146548 24278
rect 145112 24208 146548 24214
rect 147016 24284 147228 24420
rect 147560 24284 147772 24420
rect 148240 24344 149132 24420
rect 148240 24284 148452 24344
rect 147016 24278 148452 24284
rect 147016 24214 147022 24278
rect 147086 24214 147702 24278
rect 147766 24214 148452 24278
rect 147016 24208 148452 24214
rect 148784 24284 149132 24344
rect 149464 24284 149676 24420
rect 150144 24344 151580 24420
rect 150144 24284 150356 24344
rect 150688 24284 150900 24344
rect 148784 24278 150356 24284
rect 150454 24278 150900 24284
rect 148784 24214 149062 24278
rect 149126 24214 150356 24278
rect 150416 24214 150422 24278
rect 150486 24214 150900 24278
rect 148784 24208 150356 24214
rect 150454 24208 150900 24214
rect 151368 24284 151580 24344
rect 151912 24344 152804 24420
rect 151912 24284 152260 24344
rect 151368 24278 152260 24284
rect 151368 24214 152054 24278
rect 152118 24214 152260 24278
rect 151368 24208 152260 24214
rect 152592 24278 152804 24344
rect 152592 24214 152734 24278
rect 152798 24214 152804 24278
rect 152592 24208 152804 24214
rect 153272 24284 153484 24420
rect 153816 24284 154028 24420
rect 154496 24344 155252 24420
rect 154496 24284 154708 24344
rect 153272 24278 154708 24284
rect 153272 24214 153278 24278
rect 153342 24214 154502 24278
rect 154566 24214 154708 24278
rect 153272 24208 154708 24214
rect 155040 24278 155252 24344
rect 155040 24214 155182 24278
rect 155246 24214 155252 24278
rect 155040 24208 155252 24214
rect 155720 24284 155932 24420
rect 156264 24344 157836 24420
rect 156264 24284 156612 24344
rect 155720 24278 156612 24284
rect 155720 24214 155726 24278
rect 155790 24214 156612 24278
rect 155720 24208 156612 24214
rect 156944 24278 157156 24344
rect 156944 24214 156950 24278
rect 157014 24214 157156 24278
rect 156944 24208 157156 24214
rect 157624 24284 157836 24344
rect 158168 24284 158380 24420
rect 158848 24344 160284 24420
rect 158848 24284 159060 24344
rect 157624 24278 159060 24284
rect 157624 24214 158174 24278
rect 158238 24214 159060 24278
rect 157624 24208 159060 24214
rect 159392 24278 159740 24344
rect 159392 24214 159534 24278
rect 159598 24214 159740 24278
rect 159392 24208 159740 24214
rect 160072 24278 160284 24344
rect 160072 24214 160214 24278
rect 160278 24214 160284 24278
rect 160072 24208 160284 24214
rect 160752 24344 162188 24420
rect 160752 24278 160964 24344
rect 160752 24214 160758 24278
rect 160822 24214 160964 24278
rect 160752 24208 160964 24214
rect 161296 24278 161508 24344
rect 161296 24214 161438 24278
rect 161502 24214 161508 24278
rect 161296 24208 161508 24214
rect 161976 24284 162188 24344
rect 162520 24344 164092 24420
rect 162520 24284 162868 24344
rect 161976 24208 162868 24284
rect 163200 24278 163412 24344
rect 163200 24214 163206 24278
rect 163270 24214 163412 24278
rect 163200 24208 163412 24214
rect 163880 24284 164092 24344
rect 164424 24284 164636 24420
rect 165104 24344 165860 24420
rect 165104 24284 165316 24344
rect 165648 24284 165860 24344
rect 163880 24278 165316 24284
rect 165414 24278 165860 24284
rect 163880 24214 164430 24278
rect 164494 24214 165316 24278
rect 165376 24214 165382 24278
rect 165446 24214 165860 24278
rect 163880 24208 165316 24214
rect 165414 24208 165860 24214
rect 166328 24284 166540 24420
rect 166872 24344 168444 24420
rect 166872 24284 167220 24344
rect 166328 24278 167220 24284
rect 166328 24214 166878 24278
rect 166942 24214 167220 24278
rect 166328 24208 167220 24214
rect 167552 24208 167764 24344
rect 168232 24284 168444 24344
rect 168776 24284 168988 24420
rect 169456 24344 170892 24420
rect 169456 24284 169668 24344
rect 168232 24278 169668 24284
rect 168232 24214 168238 24278
rect 168302 24214 169462 24278
rect 169526 24214 169668 24278
rect 168232 24208 169668 24214
rect 170000 24284 170348 24344
rect 170680 24284 170892 24344
rect 171360 24284 171572 24420
rect 170000 24278 170620 24284
rect 170000 24214 170550 24278
rect 170614 24214 170620 24278
rect 170000 24208 170620 24214
rect 170680 24278 171572 24284
rect 170680 24214 171366 24278
rect 171430 24214 171572 24278
rect 170680 24208 171572 24214
rect 171904 24344 172796 24420
rect 171904 24278 172116 24344
rect 171904 24214 171910 24278
rect 171974 24214 172116 24278
rect 171904 24208 172116 24214
rect 172584 24284 172796 24344
rect 173128 24284 173476 24420
rect 173808 24344 174700 24420
rect 173808 24284 174020 24344
rect 172584 24278 174020 24284
rect 172584 24214 173270 24278
rect 173334 24214 174020 24278
rect 172584 24208 174020 24214
rect 174488 24284 174700 24344
rect 175032 24284 175244 24420
rect 175712 24344 177148 24420
rect 175712 24284 175924 24344
rect 174488 24278 175924 24284
rect 174488 24214 175174 24278
rect 175238 24214 175924 24278
rect 174488 24208 175924 24214
rect 176256 24208 176468 24344
rect 176936 24284 177148 24344
rect 177480 24284 177828 24420
rect 178160 24344 179052 24420
rect 179150 24414 179596 24420
rect 179112 24350 179118 24414
rect 179182 24350 179596 24414
rect 179150 24344 179596 24350
rect 178160 24284 178372 24344
rect 176936 24278 178372 24284
rect 176936 24214 176942 24278
rect 177006 24214 178166 24278
rect 178230 24214 178372 24278
rect 176936 24208 178372 24214
rect 178840 24284 179052 24344
rect 179384 24284 179596 24344
rect 180064 24344 181500 24420
rect 180064 24284 180276 24344
rect 178840 24278 180276 24284
rect 178840 24214 180206 24278
rect 180270 24214 180276 24278
rect 178840 24208 180276 24214
rect 180608 24208 180956 24344
rect 181288 24284 181500 24344
rect 181968 24344 183404 24420
rect 181968 24284 182180 24344
rect 181288 24278 182180 24284
rect 181288 24214 181430 24278
rect 181494 24214 182180 24278
rect 181288 24208 182180 24214
rect 182512 24208 182724 24344
rect 183192 24284 183404 24344
rect 183736 24284 184084 24420
rect 184416 24344 185308 24420
rect 184416 24284 184628 24344
rect 183192 24278 184628 24284
rect 183192 24214 183198 24278
rect 183262 24214 184628 24278
rect 183192 24208 184628 24214
rect 185096 24284 185308 24344
rect 185640 24284 185852 24420
rect 186320 24344 187756 24420
rect 186320 24284 186532 24344
rect 185096 24278 186532 24284
rect 185096 24214 185646 24278
rect 185710 24214 186462 24278
rect 186526 24214 186532 24278
rect 185096 24208 186532 24214
rect 186864 24208 187076 24344
rect 187544 24284 187756 24344
rect 188088 24284 188436 24420
rect 188768 24414 195100 24420
rect 188768 24350 195030 24414
rect 195094 24350 195100 24414
rect 188768 24344 195100 24350
rect 188768 24284 188980 24344
rect 187544 24278 188980 24284
rect 187544 24214 187686 24278
rect 187750 24214 188910 24278
rect 188974 24214 188980 24278
rect 187544 24208 188980 24214
rect 189448 24208 189660 24344
rect 204408 24301 204620 24420
rect 204408 24245 204482 24301
rect 204538 24284 204620 24301
rect 204538 24245 218764 24284
rect 203194 24232 203260 24235
rect 203532 24232 203598 24235
rect 203194 24230 203598 24232
rect 203194 24174 203199 24230
rect 203255 24174 203537 24230
rect 203593 24174 203598 24230
rect 204408 24208 218764 24245
rect 203194 24172 203598 24174
rect 203194 24169 203260 24172
rect 203532 24169 203598 24172
rect 1632 24052 1844 24148
rect 1632 24012 1702 24052
rect 1224 24006 1702 24012
rect 1224 23942 1230 24006
rect 1294 23996 1702 24006
rect 1758 23996 1844 24052
rect 216784 24142 217540 24148
rect 216784 24078 217470 24142
rect 217534 24078 217540 24142
rect 216784 24072 217540 24078
rect 216784 24052 216996 24072
rect 1294 23942 1844 23996
rect 1224 23936 1844 23942
rect 2720 23876 2932 24012
rect 3400 23876 3748 24012
rect 544 23870 3748 23876
rect 544 23806 550 23870
rect 614 23806 3748 23870
rect 544 23800 3748 23806
rect 15096 24006 17212 24012
rect 15096 23942 17142 24006
rect 17206 23942 17212 24006
rect 15096 23936 17212 23942
rect 216784 23996 216908 24052
rect 216964 23996 216996 24052
rect 216784 23936 216996 23996
rect 15096 23870 15308 23936
rect 15096 23806 15238 23870
rect 15302 23806 15308 23870
rect 15096 23800 15308 23806
rect 29104 23734 29724 23740
rect 29104 23670 29382 23734
rect 29446 23670 29724 23734
rect 29104 23664 29724 23670
rect 29104 23528 29452 23664
rect 29512 23598 29724 23664
rect 29512 23534 29654 23598
rect 29718 23534 29724 23598
rect 29512 23528 29724 23534
rect 30464 23734 31084 23740
rect 30464 23670 30606 23734
rect 30670 23670 31084 23734
rect 30464 23664 31084 23670
rect 30464 23528 30676 23664
rect 30736 23528 31084 23664
rect 31688 23604 31900 23740
rect 32096 23734 32308 23740
rect 32096 23670 32238 23734
rect 32302 23670 32308 23734
rect 32096 23604 32308 23670
rect 31688 23528 32308 23604
rect 32912 23734 33124 23740
rect 32912 23670 32918 23734
rect 32982 23670 33124 23734
rect 32912 23604 33124 23670
rect 33320 23734 33532 23740
rect 33320 23670 33462 23734
rect 33526 23670 33532 23734
rect 33320 23604 33532 23670
rect 32912 23528 33532 23604
rect 34136 23734 34756 23740
rect 34136 23670 34142 23734
rect 34206 23670 34756 23734
rect 34136 23664 34756 23670
rect 34136 23528 34348 23664
rect 34544 23598 34756 23664
rect 34544 23534 34686 23598
rect 34750 23534 34756 23598
rect 34544 23528 34756 23534
rect 35360 23734 35980 23740
rect 35360 23670 35502 23734
rect 35566 23670 35980 23734
rect 35360 23664 35980 23670
rect 35360 23528 35572 23664
rect 35768 23528 35980 23664
rect 36584 23604 36932 23740
rect 36992 23734 37204 23740
rect 36992 23670 37134 23734
rect 37198 23670 37204 23734
rect 36992 23604 37204 23670
rect 36584 23528 37204 23604
rect 37944 23734 38564 23740
rect 37944 23670 38494 23734
rect 38558 23670 38564 23734
rect 37944 23664 38564 23670
rect 37944 23528 38156 23664
rect 38216 23528 38564 23664
rect 39168 23734 39788 23740
rect 39168 23670 39310 23734
rect 39374 23670 39788 23734
rect 39168 23664 39788 23670
rect 39168 23528 39380 23664
rect 39576 23598 39788 23664
rect 39576 23534 39718 23598
rect 39782 23534 39788 23598
rect 39576 23528 39788 23534
rect 40392 23734 41012 23740
rect 40392 23670 40942 23734
rect 41006 23670 41012 23734
rect 40392 23664 41012 23670
rect 40392 23528 40604 23664
rect 40800 23528 41012 23664
rect 41616 23734 41828 23740
rect 41616 23670 41622 23734
rect 41686 23670 41828 23734
rect 41616 23604 41828 23670
rect 42024 23604 42236 23740
rect 41616 23528 42236 23604
rect 42840 23734 43460 23740
rect 42840 23670 42846 23734
rect 42910 23670 43460 23734
rect 42840 23664 43460 23670
rect 42840 23528 43052 23664
rect 43248 23528 43460 23664
rect 44064 23734 44684 23740
rect 44064 23670 44614 23734
rect 44678 23670 44684 23734
rect 44064 23664 44684 23670
rect 44064 23528 44412 23664
rect 44472 23528 44684 23664
rect 45424 23734 45636 23740
rect 45424 23670 45430 23734
rect 45494 23670 45636 23734
rect 45424 23604 45636 23670
rect 45696 23604 46044 23740
rect 45424 23598 46044 23604
rect 45424 23534 45430 23598
rect 45494 23534 46044 23598
rect 45424 23528 46044 23534
rect 46648 23734 47268 23740
rect 46648 23670 47198 23734
rect 47262 23670 47268 23734
rect 46648 23664 47268 23670
rect 46648 23528 46860 23664
rect 47056 23604 47268 23664
rect 47872 23734 48492 23740
rect 47872 23670 48014 23734
rect 48078 23670 48492 23734
rect 47872 23664 48492 23670
rect 47872 23604 48084 23664
rect 47056 23528 48084 23604
rect 48280 23528 48492 23664
rect 49096 23734 49716 23740
rect 49096 23670 49646 23734
rect 49710 23670 49716 23734
rect 49096 23664 49716 23670
rect 49096 23604 49308 23664
rect 49096 23598 49444 23604
rect 49096 23534 49374 23598
rect 49438 23534 49444 23598
rect 49096 23528 49444 23534
rect 49504 23528 49716 23664
rect 50320 23734 50940 23740
rect 50320 23670 50462 23734
rect 50526 23670 50870 23734
rect 50934 23670 50940 23734
rect 50320 23664 50940 23670
rect 50320 23528 50668 23664
rect 50728 23528 50940 23664
rect 51680 23734 52300 23740
rect 51680 23670 51686 23734
rect 51750 23670 52300 23734
rect 51680 23664 52300 23670
rect 51680 23528 51892 23664
rect 51952 23528 52300 23664
rect 52904 23734 53524 23740
rect 52904 23670 52910 23734
rect 52974 23670 53524 23734
rect 52904 23664 53524 23670
rect 52904 23528 53116 23664
rect 53312 23528 53524 23664
rect 54128 23604 54340 23740
rect 54536 23734 54748 23740
rect 54536 23670 54678 23734
rect 54742 23670 54748 23734
rect 54536 23604 54748 23670
rect 54128 23598 54748 23604
rect 54128 23534 54270 23598
rect 54334 23534 54748 23598
rect 54128 23528 54748 23534
rect 55352 23734 55972 23740
rect 55352 23670 55358 23734
rect 55422 23670 55972 23734
rect 55352 23664 55972 23670
rect 55352 23528 55564 23664
rect 55760 23528 55972 23664
rect 56576 23734 57196 23740
rect 56576 23670 56582 23734
rect 56646 23670 57196 23734
rect 56576 23664 57196 23670
rect 56576 23528 56788 23664
rect 56984 23528 57196 23664
rect 57800 23734 58420 23740
rect 57800 23670 58078 23734
rect 58142 23670 58420 23734
rect 57800 23664 58420 23670
rect 57800 23528 58148 23664
rect 58208 23528 58420 23664
rect 59160 23734 59780 23740
rect 59160 23670 59710 23734
rect 59774 23670 59780 23734
rect 59160 23664 59780 23670
rect 59160 23528 59372 23664
rect 59432 23528 59780 23664
rect 60384 23734 61004 23740
rect 60384 23670 60390 23734
rect 60454 23670 61004 23734
rect 60384 23664 61004 23670
rect 60384 23528 60596 23664
rect 60792 23598 61004 23664
rect 60792 23534 60798 23598
rect 60862 23534 61004 23598
rect 60792 23528 61004 23534
rect 61608 23734 62228 23740
rect 61608 23670 61614 23734
rect 61678 23670 62158 23734
rect 62222 23670 62228 23734
rect 61608 23664 62228 23670
rect 61608 23528 61820 23664
rect 62016 23528 62228 23664
rect 62832 23734 63044 23740
rect 62832 23670 62838 23734
rect 62902 23670 63044 23734
rect 62832 23604 63044 23670
rect 63240 23604 63452 23740
rect 62832 23528 63452 23604
rect 64056 23734 64676 23740
rect 64056 23670 64062 23734
rect 64126 23670 64676 23734
rect 64056 23664 64676 23670
rect 64056 23528 64268 23664
rect 64464 23604 64676 23664
rect 65280 23604 65628 23740
rect 65688 23604 65900 23740
rect 64464 23598 65900 23604
rect 64464 23534 64606 23598
rect 64670 23534 65900 23598
rect 64464 23528 65900 23534
rect 66640 23734 66852 23740
rect 66640 23670 66646 23734
rect 66710 23670 66852 23734
rect 66640 23604 66852 23670
rect 66912 23604 67260 23740
rect 66640 23528 67260 23604
rect 67864 23734 68484 23740
rect 67864 23670 67870 23734
rect 67934 23670 68414 23734
rect 68478 23670 68484 23734
rect 67864 23664 68484 23670
rect 67864 23528 68076 23664
rect 68272 23528 68484 23664
rect 69088 23734 69708 23740
rect 69088 23670 69094 23734
rect 69158 23670 69638 23734
rect 69702 23670 69708 23734
rect 69088 23664 69708 23670
rect 69088 23528 69300 23664
rect 69496 23528 69708 23664
rect 70312 23734 70932 23740
rect 70312 23670 70318 23734
rect 70382 23670 70862 23734
rect 70926 23670 70932 23734
rect 70312 23664 70932 23670
rect 70312 23598 70524 23664
rect 70312 23534 70318 23598
rect 70382 23534 70524 23598
rect 70312 23528 70524 23534
rect 70720 23528 70932 23664
rect 71536 23734 72156 23740
rect 71536 23670 71678 23734
rect 71742 23670 72156 23734
rect 71536 23664 72156 23670
rect 71536 23528 71884 23664
rect 71944 23528 72156 23664
rect 72896 23734 73516 23740
rect 72896 23670 73446 23734
rect 73510 23670 73516 23734
rect 72896 23664 73516 23670
rect 72896 23528 73108 23664
rect 73168 23528 73516 23664
rect 74120 23734 75284 23740
rect 74120 23670 74670 23734
rect 74734 23670 75214 23734
rect 75278 23670 75284 23734
rect 74120 23664 75284 23670
rect 74120 23528 74332 23664
rect 74528 23604 74740 23664
rect 75344 23604 75556 23740
rect 75752 23734 75964 23740
rect 75752 23670 75894 23734
rect 75958 23670 75964 23734
rect 75752 23604 75964 23670
rect 74528 23598 75964 23604
rect 74528 23534 75350 23598
rect 75414 23534 75964 23598
rect 74528 23528 75964 23534
rect 76568 23734 77188 23740
rect 76568 23670 76574 23734
rect 76638 23670 77188 23734
rect 76568 23664 77188 23670
rect 76568 23528 76780 23664
rect 76976 23528 77188 23664
rect 77792 23734 78412 23740
rect 77792 23670 78342 23734
rect 78406 23670 78412 23734
rect 77792 23664 78412 23670
rect 77792 23528 78004 23664
rect 78200 23528 78412 23664
rect 79016 23734 79636 23740
rect 79016 23670 79566 23734
rect 79630 23670 79636 23734
rect 79016 23664 79636 23670
rect 79016 23528 79364 23664
rect 79424 23528 79636 23664
rect 80376 23734 80996 23740
rect 80376 23670 80518 23734
rect 80582 23670 80996 23734
rect 80376 23664 80996 23670
rect 80376 23528 80588 23664
rect 80648 23604 80996 23664
rect 81600 23734 82220 23740
rect 81600 23670 82014 23734
rect 82078 23670 82220 23734
rect 81600 23664 82220 23670
rect 81600 23604 81812 23664
rect 80648 23528 81812 23604
rect 82008 23528 82220 23664
rect 82824 23734 83444 23740
rect 82824 23670 83374 23734
rect 83438 23670 83444 23734
rect 82824 23664 83444 23670
rect 82824 23528 83036 23664
rect 83232 23528 83444 23664
rect 84048 23604 84260 23740
rect 84456 23734 84668 23740
rect 84456 23670 84598 23734
rect 84662 23670 84668 23734
rect 84456 23604 84668 23670
rect 84048 23598 84668 23604
rect 84048 23534 84190 23598
rect 84254 23534 84668 23598
rect 84048 23528 84668 23534
rect 85272 23734 85892 23740
rect 85272 23670 85686 23734
rect 85750 23670 85892 23734
rect 85272 23664 85892 23670
rect 85272 23528 85484 23664
rect 85680 23528 85892 23664
rect 86496 23734 87116 23740
rect 86496 23670 86502 23734
rect 86566 23670 87116 23734
rect 86496 23664 87116 23670
rect 86496 23528 86844 23664
rect 86904 23528 87116 23664
rect 87856 23604 88068 23740
rect 88128 23734 88476 23740
rect 88128 23670 88406 23734
rect 88470 23670 88476 23734
rect 88128 23604 88476 23670
rect 87856 23528 88476 23604
rect 89080 23734 89700 23740
rect 89798 23734 90924 23740
rect 89080 23670 89086 23734
rect 89150 23670 89700 23734
rect 89760 23670 89766 23734
rect 89830 23670 90924 23734
rect 89080 23664 89700 23670
rect 89798 23664 90924 23670
rect 89080 23528 89292 23664
rect 89488 23598 89700 23664
rect 89488 23534 89630 23598
rect 89694 23534 89700 23598
rect 89488 23528 89700 23534
rect 90304 23528 90516 23664
rect 90712 23528 90924 23664
rect 91528 23734 93100 23740
rect 91528 23670 92078 23734
rect 92142 23670 93100 23734
rect 91528 23664 93100 23670
rect 91528 23528 91740 23664
rect 91936 23528 92148 23664
rect 92752 23604 93100 23664
rect 93160 23604 93372 23740
rect 92752 23528 93372 23604
rect 94112 23734 94732 23740
rect 94112 23670 94662 23734
rect 94726 23670 94732 23734
rect 94112 23664 94732 23670
rect 94112 23528 94324 23664
rect 94384 23528 94732 23664
rect 95336 23734 95956 23740
rect 95336 23670 95342 23734
rect 95406 23670 95750 23734
rect 95814 23670 95956 23734
rect 95336 23664 95956 23670
rect 95336 23598 95548 23664
rect 95336 23534 95342 23598
rect 95406 23534 95548 23598
rect 95336 23528 95548 23534
rect 95744 23528 95956 23664
rect 96560 23604 96772 23740
rect 96968 23734 97180 23740
rect 96968 23670 97110 23734
rect 97174 23670 97180 23734
rect 96968 23604 97180 23670
rect 96560 23528 97180 23604
rect 97784 23734 98404 23740
rect 97784 23670 97790 23734
rect 97854 23670 98404 23734
rect 97784 23664 98404 23670
rect 97784 23528 97996 23664
rect 98192 23604 98404 23664
rect 99008 23664 99628 23740
rect 99008 23604 99220 23664
rect 98192 23528 99220 23604
rect 99416 23598 99628 23664
rect 99416 23534 99558 23598
rect 99622 23534 99628 23598
rect 99416 23528 99628 23534
rect 100232 23604 100580 23740
rect 100640 23734 100852 23740
rect 100640 23670 100782 23734
rect 100846 23670 100852 23734
rect 100640 23604 100852 23670
rect 100232 23528 100852 23604
rect 101592 23734 102212 23740
rect 101592 23670 101598 23734
rect 101662 23670 102142 23734
rect 102206 23670 102212 23734
rect 101592 23664 102212 23670
rect 101592 23528 101804 23664
rect 101864 23528 102212 23664
rect 102816 23734 103436 23740
rect 102816 23670 103366 23734
rect 103430 23670 103436 23734
rect 102816 23664 103436 23670
rect 102816 23528 103028 23664
rect 103224 23528 103436 23664
rect 104040 23734 104660 23740
rect 104040 23670 104046 23734
rect 104110 23670 104590 23734
rect 104654 23670 104660 23734
rect 104040 23664 104660 23670
rect 104040 23528 104252 23664
rect 104448 23528 104660 23664
rect 105264 23734 105476 23740
rect 105264 23670 105270 23734
rect 105334 23670 105476 23734
rect 105264 23604 105476 23670
rect 105672 23604 105884 23740
rect 106488 23664 107108 23740
rect 106488 23604 106700 23664
rect 105264 23598 106700 23604
rect 105264 23534 105270 23598
rect 105334 23534 106700 23598
rect 105264 23528 106700 23534
rect 106896 23604 107108 23664
rect 107712 23664 108332 23740
rect 107712 23604 108060 23664
rect 106896 23528 108060 23604
rect 108120 23528 108332 23664
rect 109072 23604 109284 23740
rect 109344 23734 109692 23740
rect 109344 23670 109622 23734
rect 109686 23670 109692 23734
rect 109344 23604 109692 23670
rect 109072 23528 109692 23604
rect 110296 23734 110916 23740
rect 110296 23670 110302 23734
rect 110366 23670 110846 23734
rect 110910 23670 110916 23734
rect 110296 23664 110916 23670
rect 110296 23598 110508 23664
rect 110296 23534 110302 23598
rect 110366 23534 110508 23598
rect 110296 23528 110508 23534
rect 110704 23528 110916 23664
rect 111520 23734 112140 23740
rect 111520 23670 111526 23734
rect 111590 23670 112140 23734
rect 111520 23664 112140 23670
rect 111520 23528 111732 23664
rect 111928 23528 112140 23664
rect 112744 23734 112956 23740
rect 112744 23670 112750 23734
rect 112814 23670 112956 23734
rect 112744 23604 112956 23670
rect 113152 23734 113364 23740
rect 113152 23670 113294 23734
rect 113358 23670 113364 23734
rect 113152 23604 113364 23670
rect 112744 23528 113364 23604
rect 113968 23734 114588 23740
rect 113968 23670 114246 23734
rect 114310 23670 114588 23734
rect 113968 23664 114588 23670
rect 113968 23528 114316 23664
rect 114376 23598 114588 23664
rect 114376 23534 114518 23598
rect 114582 23534 114588 23598
rect 114376 23528 114588 23534
rect 115328 23734 115948 23740
rect 115328 23670 115334 23734
rect 115398 23670 115948 23734
rect 115328 23664 115948 23670
rect 115328 23528 115540 23664
rect 115600 23528 115948 23664
rect 116552 23734 117716 23740
rect 116552 23670 117102 23734
rect 117166 23670 117646 23734
rect 117710 23670 117716 23734
rect 116552 23664 117716 23670
rect 116552 23528 116764 23664
rect 116960 23604 117172 23664
rect 117776 23604 117988 23740
rect 118184 23604 118396 23740
rect 116960 23528 118396 23604
rect 119000 23734 119620 23740
rect 119000 23670 119006 23734
rect 119070 23670 119620 23734
rect 119000 23664 119620 23670
rect 119000 23604 119212 23664
rect 119000 23598 119348 23604
rect 119000 23534 119278 23598
rect 119342 23534 119348 23598
rect 119000 23528 119348 23534
rect 119408 23528 119620 23664
rect 120224 23734 120844 23740
rect 120224 23670 120230 23734
rect 120294 23670 120844 23734
rect 120224 23664 120844 23670
rect 120224 23528 120436 23664
rect 120632 23528 120844 23664
rect 121448 23604 121796 23740
rect 121856 23734 122068 23740
rect 121856 23670 121998 23734
rect 122062 23670 122068 23734
rect 121856 23604 122068 23670
rect 121448 23528 122068 23604
rect 122808 23734 123972 23740
rect 122808 23670 122950 23734
rect 123014 23670 123902 23734
rect 123966 23670 123972 23734
rect 122808 23664 123972 23670
rect 124032 23734 124652 23740
rect 124032 23670 124446 23734
rect 124510 23670 124652 23734
rect 124032 23664 124652 23670
rect 122808 23528 123020 23664
rect 123080 23528 123428 23664
rect 124032 23528 124244 23664
rect 124440 23598 124652 23664
rect 124440 23534 124582 23598
rect 124646 23534 124652 23598
rect 124440 23528 124652 23534
rect 125256 23604 125468 23740
rect 125664 23734 126692 23740
rect 125664 23670 125806 23734
rect 125870 23670 126692 23734
rect 125664 23664 126692 23670
rect 125664 23604 125876 23664
rect 125256 23528 125876 23604
rect 126480 23604 126692 23664
rect 126888 23734 127100 23740
rect 126888 23670 127030 23734
rect 127094 23670 127100 23734
rect 126888 23604 127100 23670
rect 127704 23664 128324 23740
rect 127704 23604 127916 23664
rect 126480 23528 127916 23604
rect 128112 23528 128324 23664
rect 128928 23734 129276 23740
rect 128928 23670 128934 23734
rect 128998 23670 129276 23734
rect 128928 23604 129276 23670
rect 129336 23604 129548 23740
rect 128928 23528 129548 23604
rect 130288 23734 130500 23740
rect 130288 23670 130294 23734
rect 130358 23670 130500 23734
rect 130288 23604 130500 23670
rect 130560 23604 130908 23740
rect 130288 23598 130908 23604
rect 130288 23534 130294 23598
rect 130358 23534 130908 23598
rect 130288 23528 130908 23534
rect 131512 23734 132132 23740
rect 131512 23670 131654 23734
rect 131718 23670 132132 23734
rect 131512 23664 132132 23670
rect 131512 23528 131724 23664
rect 131920 23604 132132 23664
rect 132736 23734 133356 23740
rect 132736 23670 133286 23734
rect 133350 23670 133356 23734
rect 132736 23664 133356 23670
rect 132736 23604 132948 23664
rect 131920 23528 132948 23604
rect 133144 23528 133356 23664
rect 133960 23604 134172 23740
rect 134368 23734 134580 23740
rect 134368 23670 134510 23734
rect 134574 23670 134580 23734
rect 134368 23604 134580 23670
rect 133960 23598 134580 23604
rect 133960 23534 134102 23598
rect 134166 23534 134580 23598
rect 133960 23528 134580 23534
rect 135184 23734 135804 23740
rect 135184 23670 135190 23734
rect 135254 23670 135734 23734
rect 135798 23670 135804 23734
rect 135184 23664 135804 23670
rect 135184 23528 135532 23664
rect 135592 23528 135804 23664
rect 136544 23734 137164 23740
rect 136544 23670 136686 23734
rect 136750 23670 137164 23734
rect 136544 23664 137164 23670
rect 136544 23528 136756 23664
rect 136816 23528 137164 23664
rect 137768 23734 138388 23740
rect 137768 23670 138182 23734
rect 138246 23670 138388 23734
rect 137768 23664 138388 23670
rect 137768 23528 137980 23664
rect 138176 23528 138388 23664
rect 138992 23604 139204 23740
rect 139400 23734 139612 23740
rect 139400 23670 139542 23734
rect 139606 23670 139612 23734
rect 139400 23604 139612 23670
rect 138992 23598 139612 23604
rect 138992 23534 139134 23598
rect 139198 23534 139612 23598
rect 138992 23528 139612 23534
rect 140216 23734 140836 23740
rect 140216 23670 140222 23734
rect 140286 23670 140836 23734
rect 140216 23664 140836 23670
rect 140216 23528 140428 23664
rect 140624 23528 140836 23664
rect 141440 23734 142060 23740
rect 141440 23670 141854 23734
rect 141918 23670 142060 23734
rect 141440 23664 142060 23670
rect 141440 23528 141652 23664
rect 141848 23528 142060 23664
rect 142664 23604 143012 23740
rect 143072 23734 143284 23740
rect 143072 23670 143214 23734
rect 143278 23670 143284 23734
rect 143072 23604 143284 23670
rect 142664 23528 143284 23604
rect 144024 23734 144644 23740
rect 144024 23670 144030 23734
rect 144094 23670 144644 23734
rect 144024 23664 144644 23670
rect 144024 23528 144236 23664
rect 144296 23528 144644 23664
rect 145248 23734 145868 23740
rect 145248 23670 145390 23734
rect 145454 23670 145868 23734
rect 145248 23664 145868 23670
rect 145248 23528 145460 23664
rect 145656 23598 145868 23664
rect 145656 23534 145662 23598
rect 145726 23534 145868 23598
rect 145656 23528 145868 23534
rect 146472 23734 147092 23740
rect 146472 23670 146478 23734
rect 146542 23670 147022 23734
rect 147086 23670 147092 23734
rect 146472 23664 147092 23670
rect 146472 23528 146684 23664
rect 146880 23528 147092 23664
rect 147696 23734 147908 23740
rect 147696 23670 147702 23734
rect 147766 23670 147908 23734
rect 147696 23604 147908 23670
rect 148104 23604 148316 23740
rect 147696 23528 148316 23604
rect 148920 23734 149540 23740
rect 148920 23670 149062 23734
rect 149126 23670 149540 23734
rect 148920 23664 149540 23670
rect 148920 23528 149132 23664
rect 149328 23598 149540 23664
rect 149328 23534 149470 23598
rect 149534 23534 149540 23598
rect 149328 23528 149540 23534
rect 150144 23734 150764 23740
rect 150144 23670 150422 23734
rect 150486 23670 150764 23734
rect 150144 23664 150764 23670
rect 150144 23528 150492 23664
rect 150552 23528 150764 23664
rect 151504 23604 151716 23740
rect 151776 23734 152124 23740
rect 151776 23670 152054 23734
rect 152118 23670 152124 23734
rect 151776 23604 152124 23670
rect 151504 23528 152124 23604
rect 152728 23734 153348 23740
rect 152728 23670 152734 23734
rect 152798 23670 153278 23734
rect 153342 23670 153348 23734
rect 152728 23664 153348 23670
rect 152728 23528 152940 23664
rect 153136 23528 153348 23664
rect 153952 23734 154572 23740
rect 153952 23670 154502 23734
rect 154566 23670 154572 23734
rect 153952 23664 154572 23670
rect 153952 23528 154164 23664
rect 154360 23528 154572 23664
rect 155176 23734 155388 23740
rect 155176 23670 155182 23734
rect 155246 23670 155388 23734
rect 155176 23604 155388 23670
rect 155584 23734 155796 23740
rect 155584 23670 155726 23734
rect 155790 23670 155796 23734
rect 155584 23604 155796 23670
rect 155176 23598 155796 23604
rect 155176 23534 155182 23598
rect 155246 23534 155796 23598
rect 155176 23528 155796 23534
rect 156400 23604 156748 23740
rect 156808 23734 157020 23740
rect 156808 23670 156950 23734
rect 157014 23670 157020 23734
rect 156808 23604 157020 23670
rect 156400 23528 157020 23604
rect 157760 23734 158380 23740
rect 157760 23670 158174 23734
rect 158238 23670 158380 23734
rect 157760 23664 158380 23670
rect 157760 23528 157972 23664
rect 158032 23528 158380 23664
rect 158984 23734 159604 23740
rect 158984 23670 159534 23734
rect 159598 23670 159604 23734
rect 158984 23664 159604 23670
rect 158984 23528 159196 23664
rect 159392 23528 159604 23664
rect 160208 23734 160420 23740
rect 160208 23670 160214 23734
rect 160278 23670 160420 23734
rect 160208 23604 160420 23670
rect 160616 23734 160828 23740
rect 160616 23670 160758 23734
rect 160822 23670 160828 23734
rect 160616 23604 160828 23670
rect 160208 23598 160828 23604
rect 160208 23534 160214 23598
rect 160278 23534 160828 23598
rect 160208 23528 160828 23534
rect 161432 23734 162052 23740
rect 161432 23670 161438 23734
rect 161502 23670 162052 23734
rect 161432 23664 162052 23670
rect 161432 23528 161644 23664
rect 161840 23528 162052 23664
rect 162656 23734 163276 23740
rect 162656 23670 163206 23734
rect 163270 23670 163276 23734
rect 162656 23664 163276 23670
rect 162656 23528 162868 23664
rect 163064 23528 163276 23664
rect 163880 23604 164228 23740
rect 164288 23734 164500 23740
rect 164288 23670 164430 23734
rect 164494 23670 164500 23734
rect 164288 23604 164500 23670
rect 163880 23598 164500 23604
rect 163880 23534 164158 23598
rect 164222 23534 164500 23598
rect 163880 23528 164500 23534
rect 165240 23734 165860 23740
rect 165240 23670 165382 23734
rect 165446 23670 165860 23734
rect 165240 23664 165860 23670
rect 165240 23528 165452 23664
rect 165512 23604 165860 23664
rect 166464 23734 167084 23740
rect 166464 23670 166878 23734
rect 166942 23670 167084 23734
rect 166464 23664 167084 23670
rect 166464 23604 166676 23664
rect 165512 23528 166676 23604
rect 166872 23528 167084 23664
rect 167688 23604 167900 23740
rect 168096 23734 168308 23740
rect 168096 23670 168238 23734
rect 168302 23670 168308 23734
rect 168096 23604 168308 23670
rect 167688 23528 168308 23604
rect 168912 23604 169124 23740
rect 169320 23734 169532 23740
rect 169320 23670 169462 23734
rect 169526 23670 169532 23734
rect 169320 23604 169532 23670
rect 168912 23528 169532 23604
rect 170136 23734 170756 23740
rect 170136 23670 170550 23734
rect 170614 23670 170756 23734
rect 170136 23664 170756 23670
rect 170136 23598 170348 23664
rect 170136 23534 170142 23598
rect 170206 23534 170348 23598
rect 170136 23528 170348 23534
rect 170544 23528 170756 23664
rect 171360 23734 171980 23740
rect 171360 23670 171366 23734
rect 171430 23670 171910 23734
rect 171974 23670 171980 23734
rect 171360 23664 171980 23670
rect 171360 23528 171708 23664
rect 171768 23528 171980 23664
rect 172720 23604 172932 23740
rect 172992 23734 173340 23740
rect 172992 23670 173270 23734
rect 173334 23670 173340 23734
rect 172992 23604 173340 23670
rect 172720 23528 173340 23604
rect 173944 23664 174564 23740
rect 173944 23528 174156 23664
rect 174352 23604 174564 23664
rect 175168 23734 175788 23740
rect 175168 23670 175174 23734
rect 175238 23670 175788 23734
rect 175168 23664 175788 23670
rect 175168 23604 175380 23664
rect 174352 23598 175380 23604
rect 174352 23534 174494 23598
rect 174558 23534 175380 23598
rect 174352 23528 175380 23534
rect 175576 23528 175788 23664
rect 176392 23734 177012 23740
rect 176392 23670 176942 23734
rect 177006 23670 177012 23734
rect 176392 23664 177012 23670
rect 176392 23528 176604 23664
rect 176800 23528 177012 23664
rect 177616 23734 178236 23740
rect 177616 23670 178166 23734
rect 178230 23670 178236 23734
rect 177616 23664 178236 23670
rect 177616 23528 177964 23664
rect 178024 23528 178236 23664
rect 178976 23734 179596 23740
rect 178976 23670 179118 23734
rect 179182 23670 179596 23734
rect 178976 23664 179596 23670
rect 178976 23528 179188 23664
rect 179248 23528 179596 23664
rect 180200 23734 180820 23740
rect 180200 23670 180206 23734
rect 180270 23670 180820 23734
rect 180200 23664 180820 23670
rect 180200 23598 180412 23664
rect 180200 23534 180206 23598
rect 180270 23534 180412 23598
rect 180200 23528 180412 23534
rect 180608 23528 180820 23664
rect 181424 23734 181636 23740
rect 181424 23670 181430 23734
rect 181494 23670 181636 23734
rect 181424 23604 181636 23670
rect 181832 23604 182044 23740
rect 181424 23528 182044 23604
rect 182648 23734 183268 23740
rect 182648 23670 183198 23734
rect 183262 23670 183268 23734
rect 182648 23664 183268 23670
rect 182648 23528 182860 23664
rect 183056 23604 183268 23664
rect 183872 23664 184492 23740
rect 183872 23604 184084 23664
rect 183056 23528 184084 23604
rect 184280 23598 184492 23664
rect 184280 23534 184422 23598
rect 184486 23534 184492 23598
rect 184280 23528 184492 23534
rect 185096 23604 185444 23740
rect 185504 23734 185716 23740
rect 185504 23670 185646 23734
rect 185710 23670 185716 23734
rect 185504 23604 185716 23670
rect 185096 23528 185716 23604
rect 186456 23734 187076 23740
rect 186456 23670 186462 23734
rect 186526 23670 187076 23734
rect 186456 23664 187076 23670
rect 186456 23528 186668 23664
rect 186728 23528 187076 23664
rect 187680 23734 188300 23740
rect 187680 23670 187686 23734
rect 187750 23670 188300 23734
rect 187680 23664 188300 23670
rect 187680 23528 187892 23664
rect 188088 23528 188300 23664
rect 188904 23734 189116 23740
rect 188904 23670 188910 23734
rect 188974 23670 189116 23734
rect 188904 23528 189116 23670
rect 201182 23598 204212 23604
rect 201144 23534 201150 23598
rect 201214 23534 204212 23598
rect 201182 23528 204212 23534
rect 204000 23326 204212 23528
rect 204000 23262 204006 23326
rect 204070 23262 204212 23326
rect 204000 23256 204212 23262
rect 15205 23246 15271 23249
rect 23747 23246 23813 23249
rect 15205 23244 23813 23246
rect 15205 23188 15210 23244
rect 15266 23188 23752 23244
rect 23808 23188 23813 23244
rect 15205 23186 23813 23188
rect 15205 23183 15271 23186
rect 23747 23183 23813 23186
rect 2103 22885 2109 22949
rect 2173 22947 2179 22949
rect 2173 22887 29381 22947
rect 2173 22885 2179 22887
rect 203114 22674 203180 22677
rect 203532 22674 203598 22677
rect 203114 22672 203598 22674
rect 2720 22576 3748 22652
rect 2720 22516 2932 22576
rect 1632 22440 2932 22516
rect 3400 22440 3748 22576
rect 15096 22646 17620 22652
rect 15096 22582 17550 22646
rect 17614 22582 17620 22646
rect 203114 22616 203119 22672
rect 203175 22616 203537 22672
rect 203593 22616 203598 22672
rect 203114 22614 203598 22616
rect 203114 22611 203180 22614
rect 203532 22611 203598 22614
rect 15096 22576 17620 22582
rect 204408 22601 218764 22652
rect 15096 22510 15308 22576
rect 15096 22446 15102 22510
rect 15166 22446 15308 22510
rect 15096 22440 15308 22446
rect 204408 22545 204482 22601
rect 204538 22576 218764 22601
rect 204538 22545 204620 22576
rect 204408 22440 204620 22545
rect 1632 22380 1844 22440
rect 216784 22380 216996 22516
rect 1224 22374 1844 22380
rect 1224 22310 1230 22374
rect 1294 22372 1844 22374
rect 1294 22316 1702 22372
rect 1758 22316 1844 22372
rect 1294 22310 1844 22316
rect 1224 22304 1844 22310
rect 1632 22168 1844 22304
rect 20400 22244 20612 22380
rect 21760 22374 21972 22380
rect 21760 22310 21902 22374
rect 21966 22310 21972 22374
rect 21760 22244 21972 22310
rect 216784 22374 217540 22380
rect 216784 22372 217470 22374
rect 216784 22316 216908 22372
rect 216964 22316 217470 22372
rect 216784 22310 217470 22316
rect 217534 22310 217540 22374
rect 216784 22304 217540 22310
rect 20400 22238 21972 22244
rect 20400 22174 21766 22238
rect 21830 22174 21972 22238
rect 20400 22168 21972 22174
rect 29920 22238 32716 22244
rect 29920 22174 29926 22238
rect 29990 22174 32716 22238
rect 29920 22168 32716 22174
rect 29920 22102 30268 22168
rect 29920 22038 29926 22102
rect 29990 22038 30268 22102
rect 29920 22032 30268 22038
rect 31280 22032 31492 22168
rect 32504 22108 32716 22168
rect 33728 22168 35164 22244
rect 33728 22108 33940 22168
rect 32504 22032 33940 22108
rect 34952 22108 35164 22168
rect 36176 22168 37748 22244
rect 36176 22108 36388 22168
rect 34952 22102 36388 22108
rect 34952 22038 35094 22102
rect 35158 22038 36388 22102
rect 34952 22032 36388 22038
rect 37400 22108 37748 22168
rect 38760 22108 38972 22244
rect 39984 22168 41420 22244
rect 39984 22108 40196 22168
rect 37400 22102 40196 22108
rect 37400 22038 39990 22102
rect 40054 22038 40196 22102
rect 37400 22032 40196 22038
rect 41208 22108 41420 22168
rect 42432 22168 43868 22244
rect 42432 22108 42644 22168
rect 41208 22032 42644 22108
rect 43656 22108 43868 22168
rect 44880 22168 47676 22244
rect 44880 22108 45228 22168
rect 43656 22102 45228 22108
rect 43656 22038 44886 22102
rect 44950 22038 45228 22102
rect 43656 22032 45228 22038
rect 46240 22032 46452 22168
rect 47464 22108 47676 22168
rect 48688 22168 50124 22244
rect 48688 22108 48900 22168
rect 47464 22032 48900 22108
rect 49912 22108 50124 22168
rect 51136 22108 51484 22244
rect 52496 22168 53932 22244
rect 52496 22108 52708 22168
rect 49912 22102 52708 22108
rect 49912 22038 50054 22102
rect 50118 22038 52708 22102
rect 49912 22032 52708 22038
rect 53720 22108 53932 22168
rect 54944 22168 56380 22244
rect 54944 22108 55156 22168
rect 53720 22102 55156 22108
rect 53720 22038 55086 22102
rect 55150 22038 55156 22102
rect 53720 22032 55156 22038
rect 56168 22108 56380 22168
rect 57392 22168 60188 22244
rect 57392 22108 57604 22168
rect 56168 22032 57604 22108
rect 58616 22108 58964 22168
rect 59976 22108 60188 22168
rect 61200 22168 62636 22244
rect 61200 22108 61412 22168
rect 58616 22102 59780 22108
rect 58616 22038 59710 22102
rect 59774 22038 59780 22102
rect 58616 22032 59780 22038
rect 59976 22032 61412 22108
rect 62424 22108 62636 22168
rect 63648 22168 65084 22244
rect 63648 22108 63860 22168
rect 62424 22032 63860 22108
rect 64872 22108 65084 22168
rect 66096 22168 68892 22244
rect 66096 22108 66444 22168
rect 64872 22102 66444 22108
rect 64872 22038 64878 22102
rect 64942 22038 66444 22102
rect 64872 22032 66444 22038
rect 67456 22032 67668 22168
rect 68680 22108 68892 22168
rect 69904 22168 71340 22244
rect 69904 22108 70116 22168
rect 68680 22102 70116 22108
rect 68680 22038 70046 22102
rect 70110 22038 70116 22102
rect 68680 22032 70116 22038
rect 71128 22108 71340 22168
rect 72352 22168 75148 22244
rect 72352 22108 72700 22168
rect 71128 22032 72700 22108
rect 73712 22032 73924 22168
rect 74936 22108 75148 22168
rect 76160 22168 77596 22244
rect 76160 22108 76372 22168
rect 74936 22102 76372 22108
rect 74936 22038 75078 22102
rect 75142 22038 76372 22102
rect 74936 22032 76372 22038
rect 77384 22108 77596 22168
rect 78608 22168 80180 22244
rect 78608 22108 78820 22168
rect 77384 22032 78820 22108
rect 79832 22108 80180 22168
rect 81192 22108 81404 22244
rect 82416 22168 83852 22244
rect 82416 22108 82628 22168
rect 79832 22102 82628 22108
rect 79832 22038 79838 22102
rect 79902 22038 82628 22102
rect 79832 22032 82628 22038
rect 83640 22108 83852 22168
rect 84864 22168 86300 22244
rect 84864 22108 85076 22168
rect 83640 22102 85076 22108
rect 83640 22038 85006 22102
rect 85070 22038 85076 22102
rect 83640 22032 85076 22038
rect 86088 22108 86300 22168
rect 87312 22108 87660 22244
rect 88672 22168 90108 22244
rect 88672 22108 88884 22168
rect 86088 22032 88884 22108
rect 89896 22108 90108 22168
rect 91120 22168 92556 22244
rect 91120 22108 91332 22168
rect 89896 22102 91332 22108
rect 89896 22038 90038 22102
rect 90102 22038 91332 22102
rect 89896 22032 91332 22038
rect 92344 22108 92556 22168
rect 93568 22168 96364 22244
rect 93568 22108 93916 22168
rect 94928 22108 95140 22168
rect 92344 22032 93916 22108
rect 94830 22102 95140 22108
rect 94792 22038 94798 22102
rect 94862 22038 95140 22102
rect 94830 22032 95140 22038
rect 96152 22108 96364 22168
rect 97376 22168 98812 22244
rect 97376 22108 97588 22168
rect 96152 22032 97588 22108
rect 98600 22108 98812 22168
rect 99824 22168 102620 22244
rect 99824 22108 100036 22168
rect 98600 22102 100036 22108
rect 98600 22038 99966 22102
rect 100030 22038 100036 22102
rect 98600 22032 100036 22038
rect 101048 22032 101396 22168
rect 102408 22108 102620 22168
rect 103632 22168 105068 22244
rect 103632 22108 103844 22168
rect 102408 22032 103844 22108
rect 104856 22108 105068 22168
rect 106080 22168 107516 22244
rect 106080 22108 106292 22168
rect 104856 22102 106292 22108
rect 104856 22038 104998 22102
rect 105062 22038 106292 22102
rect 104856 22032 106292 22038
rect 107304 22108 107516 22168
rect 108528 22168 111324 22244
rect 108528 22108 108876 22168
rect 107304 22032 108876 22108
rect 109888 22102 110100 22168
rect 109888 22038 110030 22102
rect 110094 22038 110100 22102
rect 109888 22032 110100 22038
rect 111112 22108 111324 22168
rect 112336 22168 113772 22244
rect 112336 22108 112548 22168
rect 111112 22032 112548 22108
rect 113560 22108 113772 22168
rect 114784 22108 115132 22244
rect 116144 22168 117580 22244
rect 116144 22108 116356 22168
rect 113560 22102 116356 22108
rect 113560 22038 114790 22102
rect 114854 22038 116356 22102
rect 113560 22032 116356 22038
rect 117368 22108 117580 22168
rect 118592 22168 120028 22244
rect 118592 22108 118804 22168
rect 117368 22032 118804 22108
rect 119816 22108 120028 22168
rect 121040 22168 122612 22244
rect 121040 22108 121252 22168
rect 119816 22102 121252 22108
rect 119816 22038 119958 22102
rect 120022 22038 121252 22102
rect 119816 22032 121252 22038
rect 122264 22108 122612 22168
rect 123624 22108 123836 22244
rect 124848 22168 126284 22244
rect 124848 22108 125060 22168
rect 122264 22102 125060 22108
rect 122264 22038 124990 22102
rect 125054 22038 125060 22102
rect 122264 22032 125060 22038
rect 126072 22108 126284 22168
rect 127296 22168 128732 22244
rect 127296 22108 127508 22168
rect 126072 22032 127508 22108
rect 128520 22108 128732 22168
rect 129744 22168 132540 22244
rect 129744 22108 130092 22168
rect 128520 22102 130092 22108
rect 128520 22038 129750 22102
rect 129814 22038 130092 22102
rect 128520 22032 130092 22038
rect 131104 22032 131316 22168
rect 132328 22108 132540 22168
rect 133552 22168 134988 22244
rect 133552 22108 133764 22168
rect 132328 22032 133764 22108
rect 134776 22108 134988 22168
rect 136000 22168 138796 22244
rect 136000 22108 136348 22168
rect 134776 22102 136348 22108
rect 134776 22038 134918 22102
rect 134982 22038 136348 22102
rect 134776 22032 136348 22038
rect 137360 22032 137572 22168
rect 138584 22108 138796 22168
rect 139808 22168 141244 22244
rect 139808 22108 140020 22168
rect 138584 22102 140020 22108
rect 138584 22038 139950 22102
rect 140014 22038 140020 22102
rect 138584 22032 140020 22038
rect 141032 22108 141244 22168
rect 142256 22168 143828 22244
rect 142256 22108 142468 22168
rect 141032 22032 142468 22108
rect 143480 22108 143828 22168
rect 144840 22108 145052 22244
rect 146064 22168 147500 22244
rect 146064 22108 146276 22168
rect 143480 22102 146276 22108
rect 143480 22038 144846 22102
rect 144910 22038 146276 22102
rect 143480 22032 146276 22038
rect 147288 22108 147500 22168
rect 148512 22168 149948 22244
rect 148512 22108 148724 22168
rect 147288 22032 148724 22108
rect 149736 22108 149948 22168
rect 150960 22108 151308 22244
rect 152320 22168 153756 22244
rect 152320 22108 152532 22168
rect 149736 22102 152532 22108
rect 149736 22038 149742 22102
rect 149806 22038 152532 22102
rect 149736 22032 152532 22038
rect 153544 22108 153756 22168
rect 154768 22168 156204 22244
rect 154768 22108 154980 22168
rect 153544 22102 154980 22108
rect 153544 22038 154910 22102
rect 154974 22038 154980 22102
rect 153544 22032 154980 22038
rect 155992 22108 156204 22168
rect 157216 22168 160012 22244
rect 157216 22108 157564 22168
rect 155992 22032 157564 22108
rect 158576 22032 158788 22168
rect 159800 22108 160012 22168
rect 161024 22168 162460 22244
rect 161024 22108 161236 22168
rect 159800 22102 161236 22108
rect 159800 22038 159942 22102
rect 160006 22038 161236 22102
rect 159800 22032 161236 22038
rect 162248 22108 162460 22168
rect 163472 22168 166268 22244
rect 163472 22108 163684 22168
rect 162248 22032 163684 22108
rect 164696 22102 165044 22168
rect 164696 22038 164838 22102
rect 164902 22038 165044 22102
rect 164696 22032 165044 22038
rect 166056 22108 166268 22168
rect 167280 22168 168716 22244
rect 167280 22108 167492 22168
rect 166056 22032 167492 22108
rect 168504 22108 168716 22168
rect 169728 22168 171164 22244
rect 169728 22108 169940 22168
rect 168504 22102 169940 22108
rect 168504 22038 169870 22102
rect 169934 22038 169940 22102
rect 168504 22032 169940 22038
rect 170952 22108 171164 22168
rect 172176 22168 174972 22244
rect 172176 22108 172524 22168
rect 170952 22032 172524 22108
rect 173536 22032 173748 22168
rect 174760 22108 174972 22168
rect 175984 22168 177420 22244
rect 175984 22108 176196 22168
rect 174760 22102 176196 22108
rect 174760 22038 174902 22102
rect 174966 22038 176196 22102
rect 174760 22032 176196 22038
rect 177208 22108 177420 22168
rect 178432 22168 181228 22244
rect 178432 22108 178780 22168
rect 179792 22108 180004 22168
rect 177208 22032 178780 22108
rect 179694 22102 180004 22108
rect 179656 22038 179662 22102
rect 179726 22038 180004 22102
rect 179694 22032 180004 22038
rect 181016 22108 181228 22168
rect 182240 22168 183676 22244
rect 182240 22108 182452 22168
rect 181016 22032 182452 22108
rect 183464 22108 183676 22168
rect 184688 22168 186260 22244
rect 184688 22108 184900 22168
rect 183464 22102 184900 22108
rect 183464 22038 184694 22102
rect 184758 22038 184900 22102
rect 183464 22032 184900 22038
rect 185912 22108 186260 22168
rect 187272 22108 187484 22244
rect 188496 22108 188708 22244
rect 216784 22168 216996 22304
rect 185912 22032 188708 22108
rect 204000 22102 204212 22108
rect 204000 22038 204142 22102
rect 204206 22038 204212 22102
rect 204000 21966 204212 22038
rect 204000 21902 204142 21966
rect 204206 21902 204212 21966
rect 204000 21896 204212 21902
rect 204408 21488 218764 21564
rect 204408 21473 204620 21488
rect 204408 21417 204482 21473
rect 204538 21417 204620 21473
rect 203034 21404 203100 21407
rect 203532 21404 203598 21407
rect 203034 21402 203598 21404
rect 203034 21346 203039 21402
rect 203095 21346 203537 21402
rect 203593 21346 203598 21402
rect 204408 21352 204620 21417
rect 203034 21344 203598 21346
rect 203034 21341 203100 21344
rect 203532 21341 203598 21344
rect 2720 21080 3748 21156
rect 2720 21020 2932 21080
rect 544 21014 2932 21020
rect 544 20950 550 21014
rect 614 20950 2932 21014
rect 544 20944 2932 20950
rect 3400 20944 3748 21080
rect 15096 21150 15308 21156
rect 15096 21086 15238 21150
rect 15302 21086 15308 21150
rect 15096 21014 15308 21086
rect 15096 20950 15238 21014
rect 15302 20950 15308 21014
rect 15096 20944 15308 20950
rect 20400 20884 20612 21020
rect 21760 21014 23196 21020
rect 21760 20950 23126 21014
rect 23190 20950 23196 21014
rect 21760 20944 23196 20950
rect 21760 20884 21972 20944
rect 20400 20878 21972 20884
rect 20400 20814 20542 20878
rect 20606 20814 21972 20878
rect 20400 20808 21972 20814
rect 1224 20742 1844 20748
rect 1224 20678 1230 20742
rect 1294 20692 1844 20742
rect 1294 20678 1702 20692
rect 1224 20672 1702 20678
rect 1632 20636 1702 20672
rect 1758 20636 1844 20692
rect 1632 20612 1844 20636
rect 204000 20742 204212 20748
rect 204000 20678 204006 20742
rect 204070 20678 204212 20742
rect 1632 20606 2796 20612
rect 1632 20542 2726 20606
rect 2790 20542 2796 20606
rect 1632 20536 2796 20542
rect 204000 20606 204212 20678
rect 204000 20542 204006 20606
rect 204070 20542 204212 20606
rect 204000 20536 204212 20542
rect 216784 20692 216996 20748
rect 216784 20636 216908 20692
rect 216964 20636 216996 20692
rect 216784 20612 216996 20636
rect 216784 20606 217540 20612
rect 216784 20542 217470 20606
rect 217534 20542 217540 20606
rect 216784 20536 217540 20542
rect 15205 20418 15271 20421
rect 27448 20418 27514 20421
rect 15205 20416 27514 20418
rect 15205 20360 15210 20416
rect 15266 20360 27453 20416
rect 27509 20360 27514 20416
rect 15205 20358 27514 20360
rect 15205 20355 15271 20358
rect 27448 20355 27514 20358
rect 202954 19846 203020 19849
rect 203532 19846 203598 19849
rect 202954 19844 203598 19846
rect 2720 19790 3748 19796
rect 2720 19726 2726 19790
rect 2790 19726 3748 19790
rect 2720 19720 3748 19726
rect 2720 19584 2932 19720
rect 3400 19584 3748 19720
rect 15096 19790 15308 19796
rect 15096 19726 15102 19790
rect 15166 19726 15308 19790
rect 202954 19788 202959 19844
rect 203015 19788 203537 19844
rect 203593 19788 203598 19844
rect 202954 19786 203598 19788
rect 202954 19783 203020 19786
rect 203532 19783 203598 19786
rect 15096 19654 15308 19726
rect 204408 19773 204620 19796
rect 204408 19717 204482 19773
rect 204538 19717 204620 19773
rect 29863 19660 29961 19692
rect 34855 19660 34953 19692
rect 39847 19660 39945 19692
rect 44839 19660 44937 19692
rect 49831 19660 49929 19692
rect 54823 19660 54921 19692
rect 59815 19660 59913 19692
rect 64807 19660 64905 19692
rect 69799 19660 69897 19692
rect 74791 19660 74889 19692
rect 79783 19660 79881 19692
rect 84775 19660 84873 19692
rect 89767 19660 89865 19692
rect 94759 19660 94857 19692
rect 99751 19660 99849 19692
rect 104743 19660 104841 19692
rect 109735 19660 109833 19692
rect 114727 19660 114825 19692
rect 119719 19660 119817 19692
rect 124711 19660 124809 19692
rect 129703 19660 129801 19692
rect 134695 19660 134793 19692
rect 139687 19660 139785 19692
rect 144679 19660 144777 19692
rect 149671 19660 149769 19692
rect 154663 19660 154761 19692
rect 159655 19660 159753 19692
rect 164647 19660 164745 19692
rect 169639 19660 169737 19692
rect 174631 19660 174729 19692
rect 179623 19660 179721 19692
rect 184615 19660 184713 19692
rect 204408 19660 204620 19717
rect 15096 19590 15102 19654
rect 15166 19590 15308 19654
rect 15096 19584 15308 19590
rect 29784 19654 30094 19660
rect 34816 19654 35164 19660
rect 29784 19590 29926 19654
rect 29990 19590 30062 19654
rect 30126 19590 30132 19654
rect 34816 19590 34958 19654
rect 35022 19590 35094 19654
rect 35158 19590 35164 19654
rect 29784 19584 30094 19590
rect 34816 19584 35164 19590
rect 39712 19654 40060 19660
rect 39712 19590 39854 19654
rect 39918 19590 39990 19654
rect 40054 19590 40060 19654
rect 39712 19584 40060 19590
rect 44744 19654 45054 19660
rect 49776 19654 50124 19660
rect 44744 19590 44886 19654
rect 44950 19590 45022 19654
rect 45086 19590 45092 19654
rect 49776 19590 49918 19654
rect 49982 19590 50054 19654
rect 50118 19590 50124 19654
rect 44744 19584 45054 19590
rect 49776 19584 50124 19590
rect 54808 19654 55156 19660
rect 54808 19590 54950 19654
rect 55014 19590 55086 19654
rect 55150 19590 55156 19654
rect 54808 19584 55156 19590
rect 59704 19654 60014 19660
rect 64736 19654 65046 19660
rect 69768 19654 70116 19660
rect 59704 19590 59710 19654
rect 59774 19590 59982 19654
rect 60046 19590 60052 19654
rect 64736 19590 64878 19654
rect 64942 19590 65014 19654
rect 65078 19590 65084 19654
rect 69768 19590 69910 19654
rect 69974 19590 70046 19654
rect 70110 19590 70116 19654
rect 59704 19584 60014 19590
rect 64736 19584 65046 19590
rect 69768 19584 70116 19590
rect 74664 19654 75148 19660
rect 74664 19590 74942 19654
rect 75006 19590 75078 19654
rect 75142 19590 75148 19654
rect 74664 19584 75148 19590
rect 79696 19654 80006 19660
rect 84728 19654 85076 19660
rect 79696 19590 79838 19654
rect 79902 19590 79974 19654
rect 80038 19590 80044 19654
rect 84728 19590 84870 19654
rect 84934 19590 85006 19654
rect 85070 19590 85076 19654
rect 79696 19584 80006 19590
rect 84728 19584 85076 19590
rect 89760 19654 90108 19660
rect 89760 19590 89902 19654
rect 89966 19590 90038 19654
rect 90102 19590 90108 19654
rect 89760 19584 90108 19590
rect 94656 19654 94966 19660
rect 99688 19654 100036 19660
rect 94656 19590 94798 19654
rect 94862 19590 94934 19654
rect 94998 19590 95004 19654
rect 99688 19590 99830 19654
rect 99894 19590 99966 19654
rect 100030 19590 100036 19654
rect 94656 19584 94966 19590
rect 99688 19584 100036 19590
rect 104720 19654 105068 19660
rect 104720 19590 104862 19654
rect 104926 19590 104998 19654
rect 105062 19590 105068 19654
rect 104720 19584 105068 19590
rect 109616 19654 110100 19660
rect 109616 19590 109894 19654
rect 109958 19590 110030 19654
rect 110094 19590 110100 19654
rect 109616 19584 110100 19590
rect 114648 19654 114958 19660
rect 119680 19654 120028 19660
rect 114648 19590 114790 19654
rect 114854 19590 114926 19654
rect 114990 19590 114996 19654
rect 119680 19590 119822 19654
rect 119886 19590 119958 19654
rect 120022 19590 120028 19654
rect 114648 19584 114958 19590
rect 119680 19584 120028 19590
rect 124576 19654 125060 19660
rect 124576 19590 124854 19654
rect 124918 19590 124990 19654
rect 125054 19590 125060 19654
rect 124576 19584 125060 19590
rect 129608 19654 129918 19660
rect 134640 19654 134988 19660
rect 129608 19590 129750 19654
rect 129814 19590 129886 19654
rect 129950 19590 129956 19654
rect 134640 19590 134782 19654
rect 134846 19590 134918 19654
rect 134982 19590 134988 19654
rect 129608 19584 129918 19590
rect 134640 19584 134988 19590
rect 139672 19654 140020 19660
rect 139672 19590 139814 19654
rect 139878 19590 139950 19654
rect 140014 19590 140020 19654
rect 139672 19584 140020 19590
rect 144568 19654 144878 19660
rect 149600 19654 149910 19660
rect 154632 19654 154980 19660
rect 144568 19590 144710 19654
rect 144774 19590 144846 19654
rect 144910 19590 144916 19654
rect 149600 19590 149742 19654
rect 149806 19590 149878 19654
rect 149942 19590 149948 19654
rect 154632 19590 154774 19654
rect 154838 19590 154910 19654
rect 154974 19590 154980 19654
rect 144568 19584 144878 19590
rect 149600 19584 149910 19590
rect 154632 19584 154980 19590
rect 159528 19654 160012 19660
rect 159528 19590 159806 19654
rect 159870 19590 159942 19654
rect 160006 19590 160012 19654
rect 159528 19584 160012 19590
rect 164560 19654 164908 19660
rect 164560 19590 164702 19654
rect 164766 19590 164838 19654
rect 164902 19590 164908 19654
rect 164560 19584 164908 19590
rect 169592 19654 169940 19660
rect 169592 19590 169734 19654
rect 169798 19590 169870 19654
rect 169934 19590 169940 19654
rect 169592 19584 169940 19590
rect 174624 19654 174972 19660
rect 174624 19590 174766 19654
rect 174830 19590 174902 19654
rect 174966 19590 174972 19654
rect 174624 19584 174972 19590
rect 179520 19654 179830 19660
rect 184552 19654 184764 19660
rect 179520 19590 179662 19654
rect 179726 19590 179798 19654
rect 179862 19590 179868 19654
rect 184552 19590 184558 19654
rect 184622 19590 184694 19654
rect 184758 19590 184764 19654
rect 179520 19584 179830 19590
rect 184552 19584 184764 19590
rect 204408 19584 218764 19660
rect 20400 19518 21972 19524
rect 20400 19454 21766 19518
rect 21830 19454 21972 19518
rect 20400 19448 21972 19454
rect 20400 19312 20612 19448
rect 21760 19382 21972 19448
rect 21760 19318 21766 19382
rect 21830 19318 21972 19382
rect 21760 19312 21972 19318
rect 204000 19246 204212 19252
rect 204000 19182 204142 19246
rect 204206 19182 204212 19246
rect 204000 19116 204212 19182
rect 1632 19012 1844 19116
rect 204000 19110 204348 19116
rect 204000 19046 204278 19110
rect 204342 19046 204348 19110
rect 204000 19040 204348 19046
rect 216784 19110 217540 19116
rect 216784 19046 217470 19110
rect 217534 19046 217540 19110
rect 216784 19040 217540 19046
rect 1632 18980 1702 19012
rect 1224 18974 1702 18980
rect 1224 18910 1230 18974
rect 1294 18956 1702 18974
rect 1758 18956 1844 19012
rect 216784 19012 216996 19040
rect 1294 18910 1844 18956
rect 15205 19004 15271 19007
rect 27696 19004 27762 19007
rect 15205 19002 27762 19004
rect 15205 18946 15210 19002
rect 15266 18946 27701 19002
rect 27757 18946 27762 19002
rect 15205 18944 27762 18946
rect 15205 18941 15271 18944
rect 27696 18941 27762 18944
rect 29648 18974 29996 18980
rect 1224 18904 1844 18910
rect 29648 18910 29654 18974
rect 29718 18910 29996 18974
rect 29648 18838 29996 18910
rect 29648 18774 29790 18838
rect 29854 18774 29996 18838
rect 29648 18768 29996 18774
rect 34680 18974 34892 18980
rect 34680 18910 34686 18974
rect 34750 18910 34892 18974
rect 34680 18838 34892 18910
rect 34680 18774 34686 18838
rect 34750 18774 34892 18838
rect 34680 18768 34892 18774
rect 39712 18974 39924 18980
rect 39712 18910 39718 18974
rect 39782 18910 39924 18974
rect 39712 18838 39924 18910
rect 39712 18774 39718 18838
rect 39782 18774 39924 18838
rect 39712 18768 39924 18774
rect 44744 18974 45500 18980
rect 49406 18974 49852 18980
rect 54302 18974 54884 18980
rect 44744 18910 45430 18974
rect 45494 18910 45500 18974
rect 49368 18910 49374 18974
rect 49438 18910 49852 18974
rect 54264 18910 54270 18974
rect 54334 18910 54884 18974
rect 44744 18904 45500 18910
rect 49406 18904 49852 18910
rect 54302 18904 54884 18910
rect 44744 18838 44956 18904
rect 44744 18774 44750 18838
rect 44814 18774 44956 18838
rect 44744 18768 44956 18774
rect 49640 18838 49852 18904
rect 49640 18774 49646 18838
rect 49710 18774 49852 18838
rect 49640 18768 49852 18774
rect 54672 18838 54884 18904
rect 54672 18774 54678 18838
rect 54742 18774 54884 18838
rect 54672 18768 54884 18774
rect 59704 18974 60868 18980
rect 59704 18910 60798 18974
rect 60862 18910 60868 18974
rect 59704 18904 60868 18910
rect 64600 18974 64948 18980
rect 64600 18910 64606 18974
rect 64670 18910 64948 18974
rect 59704 18838 59916 18904
rect 59704 18774 59710 18838
rect 59774 18774 59916 18838
rect 59704 18768 59916 18774
rect 64600 18838 64948 18910
rect 64600 18774 64878 18838
rect 64942 18774 64948 18838
rect 64600 18768 64948 18774
rect 69632 18974 70388 18980
rect 69632 18910 70318 18974
rect 70382 18910 70388 18974
rect 69632 18904 70388 18910
rect 74664 18974 75420 18980
rect 74664 18910 75350 18974
rect 75414 18910 75420 18974
rect 74664 18904 75420 18910
rect 69632 18838 69844 18904
rect 69632 18774 69774 18838
rect 69838 18774 69844 18838
rect 69632 18768 69844 18774
rect 74664 18838 74876 18904
rect 74664 18774 74670 18838
rect 74734 18774 74876 18838
rect 74664 18768 74876 18774
rect 79696 18838 79908 18980
rect 84222 18974 84804 18980
rect 84184 18910 84190 18974
rect 84254 18910 84804 18974
rect 84222 18904 84804 18910
rect 79696 18774 79702 18838
rect 79766 18774 79908 18838
rect 79696 18768 79908 18774
rect 84592 18838 84804 18904
rect 84592 18774 84734 18838
rect 84798 18774 84804 18838
rect 84592 18768 84804 18774
rect 89624 18974 89836 18980
rect 89624 18910 89630 18974
rect 89694 18910 89836 18974
rect 89624 18838 89836 18910
rect 89624 18774 89766 18838
rect 89830 18774 89836 18838
rect 89624 18768 89836 18774
rect 94656 18974 95412 18980
rect 94656 18910 95342 18974
rect 95406 18910 95412 18974
rect 94656 18904 95412 18910
rect 99552 18974 99900 18980
rect 99552 18910 99558 18974
rect 99622 18910 99900 18974
rect 94656 18838 94868 18904
rect 94656 18774 94798 18838
rect 94862 18774 94868 18838
rect 94656 18768 94868 18774
rect 99552 18838 99900 18910
rect 99552 18774 99694 18838
rect 99758 18774 99900 18838
rect 99552 18768 99900 18774
rect 104584 18974 105340 18980
rect 104584 18910 105270 18974
rect 105334 18910 105340 18974
rect 104584 18904 105340 18910
rect 109616 18974 110372 18980
rect 109616 18910 110302 18974
rect 110366 18910 110372 18974
rect 109616 18904 110372 18910
rect 114512 18974 114860 18980
rect 119310 18974 119756 18980
rect 114512 18910 114518 18974
rect 114582 18910 114860 18974
rect 119272 18910 119278 18974
rect 119342 18910 119756 18974
rect 104584 18838 104796 18904
rect 104584 18774 104590 18838
rect 104654 18774 104796 18838
rect 104584 18768 104796 18774
rect 109616 18838 109828 18904
rect 109616 18774 109758 18838
rect 109822 18774 109828 18838
rect 109616 18768 109828 18774
rect 114512 18838 114860 18910
rect 119310 18904 119756 18910
rect 114512 18774 114790 18838
rect 114854 18774 114860 18838
rect 114512 18768 114860 18774
rect 119544 18838 119756 18904
rect 119544 18774 119550 18838
rect 119614 18774 119756 18838
rect 119544 18768 119756 18774
rect 124576 18974 124788 18980
rect 124576 18910 124582 18974
rect 124646 18910 124788 18974
rect 124576 18838 124788 18910
rect 124576 18774 124582 18838
rect 124646 18774 124788 18838
rect 124576 18768 124788 18774
rect 129608 18974 130364 18980
rect 134134 18974 134716 18980
rect 139166 18974 139748 18980
rect 129608 18910 130294 18974
rect 130358 18910 130364 18974
rect 134096 18910 134102 18974
rect 134166 18910 134716 18974
rect 139128 18910 139134 18974
rect 139198 18910 139748 18974
rect 129608 18904 130364 18910
rect 134134 18904 134716 18910
rect 139166 18904 139748 18910
rect 129608 18838 129820 18904
rect 129608 18774 129614 18838
rect 129678 18774 129820 18838
rect 129608 18768 129820 18774
rect 134504 18838 134716 18904
rect 134504 18774 134510 18838
rect 134574 18774 134716 18838
rect 134504 18768 134716 18774
rect 139536 18838 139748 18904
rect 139536 18774 139542 18838
rect 139606 18774 139748 18838
rect 139536 18768 139748 18774
rect 144568 18974 145732 18980
rect 144568 18910 145662 18974
rect 145726 18910 145732 18974
rect 144568 18904 145732 18910
rect 149464 18974 149812 18980
rect 149464 18910 149470 18974
rect 149534 18910 149812 18974
rect 144568 18838 144780 18904
rect 144568 18774 144574 18838
rect 144638 18774 144780 18838
rect 144568 18768 144780 18774
rect 149464 18838 149812 18910
rect 149464 18774 149606 18838
rect 149670 18774 149812 18838
rect 149464 18768 149812 18774
rect 154496 18974 155252 18980
rect 154496 18910 155182 18974
rect 155246 18910 155252 18974
rect 154496 18904 155252 18910
rect 159528 18974 160284 18980
rect 164190 18974 164772 18980
rect 159528 18910 160214 18974
rect 160278 18910 160284 18974
rect 164152 18910 164158 18974
rect 164222 18910 164772 18974
rect 159528 18904 160284 18910
rect 164190 18904 164772 18910
rect 154496 18838 154708 18904
rect 154496 18774 154638 18838
rect 154702 18774 154708 18838
rect 154496 18768 154708 18774
rect 159528 18838 159740 18904
rect 159528 18774 159534 18838
rect 159598 18774 159740 18838
rect 159528 18768 159740 18774
rect 164560 18838 164772 18904
rect 164560 18774 164566 18838
rect 164630 18774 164772 18838
rect 164560 18768 164772 18774
rect 169456 18974 170212 18980
rect 169456 18910 170142 18974
rect 170206 18910 170212 18974
rect 169456 18904 170212 18910
rect 174488 18974 174700 18980
rect 174488 18910 174494 18974
rect 174558 18910 174700 18974
rect 169456 18838 169668 18904
rect 169456 18774 169598 18838
rect 169662 18774 169668 18838
rect 169456 18768 169668 18774
rect 174488 18838 174700 18910
rect 174488 18774 174630 18838
rect 174694 18774 174700 18838
rect 174488 18768 174700 18774
rect 179520 18974 180276 18980
rect 179520 18910 180206 18974
rect 180270 18910 180276 18974
rect 179520 18904 180276 18910
rect 184416 18974 184764 18980
rect 184416 18910 184422 18974
rect 184486 18910 184764 18974
rect 179520 18838 179732 18904
rect 179520 18774 179662 18838
rect 179726 18774 179732 18838
rect 179520 18768 179732 18774
rect 184416 18838 184764 18910
rect 216784 18956 216908 19012
rect 216964 18956 216996 19012
rect 216784 18904 216996 18956
rect 184416 18774 184422 18838
rect 184486 18774 184764 18838
rect 184416 18768 184764 18774
rect 204408 18645 204620 18708
rect 204408 18589 204482 18645
rect 204538 18589 204620 18645
rect 202874 18576 202940 18579
rect 203532 18576 203598 18579
rect 202874 18574 203598 18576
rect 202874 18518 202879 18574
rect 202935 18518 203537 18574
rect 203593 18518 203598 18574
rect 202874 18516 203598 18518
rect 202874 18513 202940 18516
rect 203532 18513 203598 18516
rect 204408 18572 204620 18589
rect 204408 18496 218764 18572
rect 544 18430 2932 18436
rect 544 18366 550 18430
rect 614 18366 2932 18430
rect 544 18360 2932 18366
rect 2720 18164 2932 18360
rect 3400 18164 3748 18436
rect 2720 18088 3748 18164
rect 15096 18430 15308 18436
rect 15096 18366 15238 18430
rect 15302 18366 15308 18430
rect 15096 18158 15308 18366
rect 15096 18094 15238 18158
rect 15302 18094 15308 18158
rect 15096 18088 15308 18094
rect 20400 18158 21972 18164
rect 20400 18094 20542 18158
rect 20606 18094 21972 18158
rect 20400 18088 21972 18094
rect 29784 18158 29996 18164
rect 29784 18094 29790 18158
rect 29854 18094 29996 18158
rect 29784 18088 29996 18094
rect 34680 18158 34892 18164
rect 34680 18094 34686 18158
rect 34750 18094 34892 18158
rect 34680 18088 34892 18094
rect 20400 18022 20612 18088
rect 20400 17958 20406 18022
rect 20470 17958 20612 18022
rect 20400 17952 20612 17958
rect 21760 17952 21972 18088
rect 29793 18022 29996 18088
rect 29793 17982 29926 18022
rect 29920 17958 29926 17982
rect 29990 17958 29996 18022
rect 34785 18022 34892 18088
rect 34785 17982 34822 18022
rect 29920 17952 29996 17958
rect 34816 17958 34822 17982
rect 34886 17958 34892 18022
rect 34816 17952 34892 17958
rect 39712 18158 39924 18164
rect 39712 18094 39718 18158
rect 39782 18094 39924 18158
rect 39712 18022 39924 18094
rect 44744 18158 44956 18164
rect 44744 18094 44750 18158
rect 44814 18094 44956 18158
rect 44744 18088 44956 18094
rect 49640 18158 49988 18164
rect 49640 18094 49646 18158
rect 49710 18094 49988 18158
rect 49640 18088 49988 18094
rect 54672 18158 54884 18164
rect 54672 18094 54678 18158
rect 54742 18094 54884 18158
rect 54672 18088 54884 18094
rect 59704 18158 59916 18164
rect 59704 18094 59710 18158
rect 59774 18094 59916 18158
rect 59704 18088 59916 18094
rect 39712 17958 39718 18022
rect 39782 17958 39924 18022
rect 44769 18022 44956 18088
rect 44769 17982 44886 18022
rect 39712 17952 39924 17958
rect 44880 17958 44886 17982
rect 44950 17958 44956 18022
rect 49761 18022 49988 18088
rect 49761 17982 49782 18022
rect 44880 17952 44956 17958
rect 49776 17958 49782 17982
rect 49846 17958 49988 18022
rect 54753 18022 54884 18088
rect 54753 17982 54814 18022
rect 49776 17952 49988 17958
rect 54808 17958 54814 17982
rect 54878 17958 54884 18022
rect 59745 18022 59916 18088
rect 59745 17982 59846 18022
rect 54808 17952 54884 17958
rect 59840 17958 59846 17982
rect 59910 17958 59916 18022
rect 59840 17952 59916 17958
rect 64736 18158 64948 18164
rect 64736 18094 64878 18158
rect 64942 18094 64948 18158
rect 64736 18022 64948 18094
rect 69632 18158 69844 18164
rect 69632 18094 69774 18158
rect 69838 18094 69844 18158
rect 69632 18088 69844 18094
rect 74664 18158 74876 18164
rect 74664 18094 74670 18158
rect 74734 18094 74876 18158
rect 74664 18088 74876 18094
rect 79696 18158 84804 18164
rect 79696 18094 79702 18158
rect 79766 18094 84734 18158
rect 84798 18094 84804 18158
rect 79696 18088 84804 18094
rect 89624 18158 89836 18164
rect 89624 18094 89766 18158
rect 89830 18094 89836 18158
rect 89624 18088 89836 18094
rect 94656 18158 94868 18164
rect 94656 18094 94798 18158
rect 94862 18094 94868 18158
rect 94656 18088 94868 18094
rect 64736 17958 64742 18022
rect 64806 17958 64948 18022
rect 69729 18022 69844 18088
rect 69729 17982 69774 18022
rect 64736 17952 64948 17958
rect 69768 17958 69774 17982
rect 69838 17958 69844 18022
rect 74721 18022 74876 18088
rect 74721 17982 74806 18022
rect 69768 17952 69844 17958
rect 74800 17958 74806 17982
rect 74870 17958 74876 18022
rect 79713 18022 79908 18088
rect 79713 17982 79838 18022
rect 74800 17952 74876 17958
rect 79832 17958 79838 17982
rect 79902 17958 79908 18022
rect 84705 18022 84804 18088
rect 84705 17982 84734 18022
rect 79832 17952 79908 17958
rect 84728 17958 84734 17982
rect 84798 17958 84804 18022
rect 89697 18022 89836 18088
rect 89697 17982 89766 18022
rect 84728 17952 84804 17958
rect 89760 17958 89766 17982
rect 89830 17958 89836 18022
rect 94689 18022 94868 18088
rect 94689 17982 94798 18022
rect 89760 17952 89836 17958
rect 94792 17958 94798 17982
rect 94862 17958 94868 18022
rect 94792 17952 94868 17958
rect 99552 18158 99900 18164
rect 99552 18094 99694 18158
rect 99758 18094 99900 18158
rect 99552 18022 99900 18094
rect 104584 18158 104796 18164
rect 104584 18094 104590 18158
rect 104654 18094 104796 18158
rect 104584 18088 104796 18094
rect 109616 18158 109828 18164
rect 109616 18094 109758 18158
rect 109822 18094 109828 18158
rect 109616 18088 109828 18094
rect 114648 18158 114860 18164
rect 114648 18094 114790 18158
rect 114854 18094 114860 18158
rect 114648 18088 114860 18094
rect 119544 18158 119756 18164
rect 119544 18094 119550 18158
rect 119614 18094 119756 18158
rect 119544 18088 119756 18094
rect 124576 18158 124788 18164
rect 124576 18094 124582 18158
rect 124646 18094 124788 18158
rect 124576 18088 124788 18094
rect 129608 18158 129820 18164
rect 129608 18094 129614 18158
rect 129678 18094 129820 18158
rect 129608 18088 129820 18094
rect 134504 18158 134852 18164
rect 134504 18094 134510 18158
rect 134574 18094 134852 18158
rect 134504 18088 134852 18094
rect 139536 18158 139748 18164
rect 139536 18094 139542 18158
rect 139606 18094 139748 18158
rect 139536 18088 139748 18094
rect 144568 18158 144780 18164
rect 144568 18094 144574 18158
rect 144638 18094 144780 18158
rect 144568 18088 144780 18094
rect 149600 18158 149812 18164
rect 149600 18094 149606 18158
rect 149670 18094 149812 18158
rect 149600 18088 149812 18094
rect 154496 18158 154708 18164
rect 154496 18094 154638 18158
rect 154702 18094 154708 18158
rect 154496 18088 154708 18094
rect 159528 18158 159740 18164
rect 159528 18094 159534 18158
rect 159598 18094 159740 18158
rect 159528 18088 159740 18094
rect 99552 17958 99558 18022
rect 99622 17958 99900 18022
rect 104673 18022 104796 18088
rect 104673 17982 104726 18022
rect 99552 17952 99900 17958
rect 104720 17958 104726 17982
rect 104790 17958 104796 18022
rect 109665 18022 109828 18088
rect 109665 17982 109758 18022
rect 104720 17952 104796 17958
rect 109752 17958 109758 17982
rect 109822 17958 109828 18022
rect 114657 18022 114860 18088
rect 114657 17982 114790 18022
rect 109752 17952 109828 17958
rect 114784 17958 114790 17982
rect 114854 17958 114860 18022
rect 119649 18022 119756 18088
rect 119649 17982 119686 18022
rect 114784 17952 114860 17958
rect 119680 17958 119686 17982
rect 119750 17958 119756 18022
rect 124641 18022 124788 18088
rect 124641 17982 124718 18022
rect 119680 17952 119756 17958
rect 124712 17958 124718 17982
rect 124782 17958 124788 18022
rect 129633 18022 129820 18088
rect 129633 17982 129750 18022
rect 124712 17952 124788 17958
rect 129744 17958 129750 17982
rect 129814 17958 129820 18022
rect 134625 18022 134852 18088
rect 134625 17982 134646 18022
rect 129744 17952 129820 17958
rect 134640 17958 134646 17982
rect 134710 17958 134852 18022
rect 139617 18022 139748 18088
rect 139617 17982 139678 18022
rect 134640 17952 134852 17958
rect 139672 17958 139678 17982
rect 139742 17958 139748 18022
rect 144609 18022 144780 18088
rect 144609 17982 144710 18022
rect 139672 17952 139748 17958
rect 144704 17958 144710 17982
rect 144774 17958 144780 18022
rect 149601 18022 149812 18088
rect 149601 17982 149742 18022
rect 144704 17952 144780 17958
rect 149736 17958 149742 17982
rect 149806 17958 149812 18022
rect 154593 18022 154708 18088
rect 154593 17982 154638 18022
rect 149736 17952 149812 17958
rect 154632 17958 154638 17982
rect 154702 17958 154708 18022
rect 159585 18022 159740 18088
rect 159585 17982 159670 18022
rect 154632 17952 154708 17958
rect 159664 17958 159670 17982
rect 159734 17958 159740 18022
rect 159664 17952 159740 17958
rect 164560 18158 164772 18164
rect 164560 18094 164566 18158
rect 164630 18094 164772 18158
rect 164560 18022 164772 18094
rect 169456 18158 169668 18164
rect 169456 18094 169598 18158
rect 169662 18094 169668 18158
rect 169456 18088 169668 18094
rect 174488 18158 174700 18164
rect 174488 18094 174630 18158
rect 174694 18094 174700 18158
rect 174488 18088 174700 18094
rect 179520 18158 179732 18164
rect 179520 18094 179662 18158
rect 179726 18094 179732 18158
rect 179520 18088 179732 18094
rect 164560 17958 164566 18022
rect 164630 17958 164772 18022
rect 169569 18022 169668 18088
rect 169569 17982 169598 18022
rect 164560 17952 164772 17958
rect 169592 17958 169598 17982
rect 169662 17958 169668 18022
rect 174561 18022 174700 18088
rect 174561 17982 174630 18022
rect 169592 17952 169668 17958
rect 174624 17958 174630 17982
rect 174694 17958 174700 18022
rect 179553 18022 179732 18088
rect 179553 17982 179662 18022
rect 174624 17952 174700 17958
rect 179656 17958 179662 17982
rect 179726 17958 179732 18022
rect 179656 17952 179732 17958
rect 184416 18158 184764 18164
rect 184416 18094 184422 18158
rect 184486 18094 184764 18158
rect 184416 18022 184764 18094
rect 184416 17958 184422 18022
rect 184486 17958 184764 18022
rect 184416 17952 184764 17958
rect 29512 17756 29724 17892
rect 29920 17886 30132 17892
rect 29920 17822 30062 17886
rect 30126 17822 30132 17886
rect 29920 17816 30132 17822
rect 29920 17758 29996 17816
rect 29512 17700 29560 17756
rect 29616 17700 29724 17756
rect 29512 17620 29724 17700
rect 29793 17660 29996 17758
rect 28968 17614 29724 17620
rect 15205 17590 15271 17593
rect 27572 17590 27638 17593
rect 15205 17588 27638 17590
rect 15205 17532 15210 17588
rect 15266 17532 27577 17588
rect 27633 17532 27638 17588
rect 28968 17550 28974 17614
rect 29038 17550 29724 17614
rect 28968 17544 29724 17550
rect 15205 17530 27638 17532
rect 15205 17527 15271 17530
rect 27572 17527 27638 17530
rect 29920 17484 29996 17660
rect 34408 17777 34620 17892
rect 34816 17886 35028 17892
rect 34816 17822 34958 17886
rect 35022 17822 35028 17886
rect 34816 17816 35028 17822
rect 34408 17756 34629 17777
rect 34816 17758 34892 17816
rect 34408 17700 34552 17756
rect 34608 17700 34629 17756
rect 34408 17679 34629 17700
rect 34408 17614 34620 17679
rect 34785 17660 34892 17758
rect 34408 17550 34550 17614
rect 34614 17550 34620 17614
rect 34408 17544 34620 17550
rect 34816 17620 34892 17660
rect 39440 17756 39652 17892
rect 39440 17700 39544 17756
rect 39600 17700 39652 17756
rect 34816 17614 34990 17620
rect 39440 17614 39652 17700
rect 34816 17550 34958 17614
rect 35022 17550 35028 17614
rect 39440 17550 39446 17614
rect 39510 17550 39652 17614
rect 34816 17544 34990 17550
rect 39440 17544 39652 17550
rect 39712 17886 39924 17892
rect 39712 17822 39854 17886
rect 39918 17822 39924 17886
rect 39712 17614 39924 17822
rect 44472 17756 44684 17892
rect 44880 17886 45092 17892
rect 44880 17822 45022 17886
rect 45086 17822 45092 17886
rect 44880 17816 45092 17822
rect 44880 17758 44956 17816
rect 44472 17700 44536 17756
rect 44592 17700 44684 17756
rect 44472 17620 44684 17700
rect 44769 17660 44956 17758
rect 39712 17550 39854 17614
rect 39918 17550 39924 17614
rect 39712 17544 39924 17550
rect 44200 17614 44684 17620
rect 44200 17550 44206 17614
rect 44270 17550 44684 17614
rect 44200 17544 44684 17550
rect 44880 17484 44956 17660
rect 49504 17777 49580 17892
rect 49776 17886 49988 17892
rect 49776 17822 49918 17886
rect 49982 17822 49988 17886
rect 49504 17756 49605 17777
rect 49776 17758 49988 17822
rect 49504 17700 49528 17756
rect 49584 17700 49605 17756
rect 49504 17679 49605 17700
rect 49504 17614 49580 17679
rect 49761 17660 49988 17758
rect 49504 17550 49510 17614
rect 49574 17550 49580 17614
rect 49504 17544 49580 17550
rect 49776 17614 49988 17660
rect 49776 17550 49918 17614
rect 49982 17550 49988 17614
rect 49776 17544 49988 17550
rect 54400 17756 54612 17892
rect 54808 17886 55020 17892
rect 54808 17822 54950 17886
rect 55014 17822 55020 17886
rect 54808 17816 55020 17822
rect 54808 17758 54884 17816
rect 54400 17700 54520 17756
rect 54576 17700 54612 17756
rect 54400 17614 54612 17700
rect 54753 17660 54884 17758
rect 54400 17550 54542 17614
rect 54606 17550 54612 17614
rect 54400 17544 54612 17550
rect 54808 17620 54884 17660
rect 59432 17756 59644 17892
rect 59840 17886 60052 17892
rect 59840 17822 59982 17886
rect 60046 17822 60052 17886
rect 59840 17816 60052 17822
rect 59840 17758 59916 17816
rect 59432 17700 59512 17756
rect 59568 17700 59644 17756
rect 59432 17620 59644 17700
rect 59745 17660 59916 17758
rect 54808 17614 54982 17620
rect 59296 17614 59644 17620
rect 54808 17550 54950 17614
rect 55014 17550 55020 17614
rect 59296 17550 59302 17614
rect 59366 17550 59644 17614
rect 54808 17544 54982 17550
rect 59296 17544 59644 17550
rect 59840 17484 59916 17660
rect 64464 17756 64676 17892
rect 64464 17700 64504 17756
rect 64560 17700 64676 17756
rect 64464 17614 64676 17700
rect 64464 17550 64470 17614
rect 64534 17550 64676 17614
rect 64464 17544 64676 17550
rect 64736 17886 65084 17892
rect 64736 17822 65014 17886
rect 65078 17822 65084 17886
rect 64736 17816 65084 17822
rect 64736 17614 64948 17816
rect 64736 17550 64878 17614
rect 64942 17550 64948 17614
rect 64736 17544 64948 17550
rect 69360 17777 69572 17892
rect 69768 17886 69980 17892
rect 69768 17822 69910 17886
rect 69974 17822 69980 17886
rect 69768 17816 69980 17822
rect 69360 17756 69573 17777
rect 69768 17758 69844 17816
rect 69360 17700 69496 17756
rect 69552 17700 69573 17756
rect 69360 17679 69573 17700
rect 69360 17614 69572 17679
rect 69729 17660 69844 17758
rect 69360 17550 69502 17614
rect 69566 17550 69572 17614
rect 69360 17544 69572 17550
rect 69768 17620 69844 17660
rect 74392 17756 74604 17892
rect 74800 17886 75012 17892
rect 74800 17822 74942 17886
rect 75006 17822 75012 17886
rect 74800 17816 75012 17822
rect 74800 17758 74876 17816
rect 74392 17700 74488 17756
rect 74544 17700 74604 17756
rect 69768 17614 69942 17620
rect 74392 17614 74604 17700
rect 74721 17660 74876 17758
rect 69768 17550 69910 17614
rect 69974 17550 69980 17614
rect 74392 17550 74398 17614
rect 74462 17550 74604 17614
rect 69768 17544 69942 17550
rect 74392 17544 74604 17550
rect 74800 17484 74876 17660
rect 79424 17756 79636 17892
rect 79832 17886 80044 17892
rect 79832 17822 79974 17886
rect 80038 17822 80044 17886
rect 79832 17816 80044 17822
rect 79832 17758 79908 17816
rect 79424 17700 79480 17756
rect 79536 17700 79636 17756
rect 79424 17614 79636 17700
rect 79713 17660 79908 17758
rect 79424 17550 79430 17614
rect 79494 17550 79636 17614
rect 79424 17544 79636 17550
rect 79832 17484 79908 17660
rect 84320 17777 84532 17892
rect 84728 17886 84940 17892
rect 84728 17822 84870 17886
rect 84934 17822 84940 17886
rect 84728 17816 84940 17822
rect 84320 17756 84549 17777
rect 84728 17758 84804 17816
rect 84320 17700 84472 17756
rect 84528 17700 84549 17756
rect 84320 17679 84549 17700
rect 84320 17614 84532 17679
rect 84705 17660 84804 17758
rect 84320 17550 84326 17614
rect 84390 17550 84532 17614
rect 84320 17544 84532 17550
rect 84728 17620 84804 17660
rect 89352 17756 89564 17892
rect 89760 17886 89972 17892
rect 89760 17822 89902 17886
rect 89966 17822 89972 17886
rect 89760 17816 89972 17822
rect 89760 17758 89836 17816
rect 89352 17700 89464 17756
rect 89520 17700 89564 17756
rect 84728 17614 84902 17620
rect 89352 17614 89564 17700
rect 89697 17660 89836 17758
rect 84728 17550 84870 17614
rect 84934 17550 84940 17614
rect 89352 17550 89358 17614
rect 89422 17550 89564 17614
rect 84728 17544 84902 17550
rect 89352 17544 89564 17550
rect 89760 17484 89836 17660
rect 94384 17756 94596 17892
rect 94792 17886 95004 17892
rect 94792 17822 94934 17886
rect 94998 17822 95004 17886
rect 94792 17816 95004 17822
rect 94792 17758 94868 17816
rect 94384 17700 94456 17756
rect 94512 17700 94596 17756
rect 94384 17614 94596 17700
rect 94689 17660 94868 17758
rect 94384 17550 94390 17614
rect 94454 17550 94596 17614
rect 94384 17544 94596 17550
rect 94792 17484 94868 17660
rect 99416 17777 99492 17892
rect 99688 17886 99900 17892
rect 99688 17822 99830 17886
rect 99894 17822 99900 17886
rect 99416 17756 99525 17777
rect 99688 17758 99900 17822
rect 99416 17700 99448 17756
rect 99504 17700 99525 17756
rect 99416 17679 99525 17700
rect 99416 17614 99492 17679
rect 99681 17660 99900 17758
rect 99416 17550 99422 17614
rect 99486 17550 99492 17614
rect 99416 17544 99492 17550
rect 99688 17614 99900 17660
rect 99688 17550 99694 17614
rect 99758 17550 99900 17614
rect 99688 17544 99900 17550
rect 104312 17756 104524 17892
rect 104720 17886 104932 17892
rect 104720 17822 104862 17886
rect 104926 17822 104932 17886
rect 104720 17816 104932 17822
rect 104720 17758 104796 17816
rect 104312 17700 104440 17756
rect 104496 17700 104524 17756
rect 104312 17614 104524 17700
rect 104673 17660 104796 17758
rect 104312 17550 104318 17614
rect 104382 17550 104524 17614
rect 104312 17544 104524 17550
rect 104720 17484 104796 17660
rect 109344 17756 109556 17892
rect 109752 17886 109964 17892
rect 109752 17822 109894 17886
rect 109958 17822 109964 17886
rect 109752 17816 109964 17822
rect 109752 17758 109828 17816
rect 109344 17700 109432 17756
rect 109488 17700 109556 17756
rect 109344 17620 109556 17700
rect 109665 17660 109828 17758
rect 109072 17614 109556 17620
rect 109072 17550 109078 17614
rect 109142 17550 109556 17614
rect 109072 17544 109556 17550
rect 109752 17484 109828 17660
rect 114376 17756 114588 17892
rect 114784 17886 114996 17892
rect 114784 17822 114926 17886
rect 114990 17822 114996 17886
rect 114784 17816 114996 17822
rect 114784 17758 114860 17816
rect 114376 17700 114424 17756
rect 114480 17700 114588 17756
rect 114376 17614 114588 17700
rect 114657 17660 114860 17758
rect 114376 17550 114382 17614
rect 114446 17550 114588 17614
rect 114376 17544 114588 17550
rect 114784 17484 114860 17660
rect 119272 17777 119484 17892
rect 119680 17886 119892 17892
rect 119680 17822 119822 17886
rect 119886 17822 119892 17886
rect 119680 17816 119892 17822
rect 119272 17756 119493 17777
rect 119680 17758 119756 17816
rect 119272 17700 119416 17756
rect 119472 17700 119493 17756
rect 119272 17679 119493 17700
rect 119272 17614 119484 17679
rect 119649 17660 119756 17758
rect 119272 17550 119278 17614
rect 119342 17550 119484 17614
rect 119272 17544 119484 17550
rect 119680 17620 119756 17660
rect 124304 17756 124516 17892
rect 124712 17886 124924 17892
rect 124712 17822 124854 17886
rect 124918 17822 124924 17886
rect 124712 17816 124924 17822
rect 124712 17758 124788 17816
rect 124304 17700 124408 17756
rect 124464 17700 124516 17756
rect 119680 17614 119854 17620
rect 124304 17614 124516 17700
rect 124641 17660 124788 17758
rect 119680 17550 119822 17614
rect 119886 17550 119892 17614
rect 124304 17550 124310 17614
rect 124374 17550 124516 17614
rect 119680 17544 119854 17550
rect 124304 17544 124516 17550
rect 124712 17484 124788 17660
rect 129336 17756 129548 17892
rect 129744 17886 129956 17892
rect 129744 17822 129886 17886
rect 129950 17822 129956 17886
rect 129744 17816 129956 17822
rect 129744 17758 129820 17816
rect 129336 17700 129400 17756
rect 129456 17700 129548 17756
rect 129336 17614 129548 17700
rect 129633 17660 129820 17758
rect 129336 17550 129342 17614
rect 129406 17550 129548 17614
rect 129336 17544 129548 17550
rect 129744 17484 129820 17660
rect 134368 17777 134444 17892
rect 134640 17886 134852 17892
rect 134640 17822 134782 17886
rect 134846 17822 134852 17886
rect 134368 17756 134469 17777
rect 134640 17758 134852 17822
rect 134368 17700 134392 17756
rect 134448 17700 134469 17756
rect 134368 17679 134469 17700
rect 134368 17614 134444 17679
rect 134625 17660 134852 17758
rect 134368 17550 134374 17614
rect 134438 17550 134444 17614
rect 134368 17544 134444 17550
rect 134640 17614 134852 17660
rect 134640 17550 134782 17614
rect 134846 17550 134852 17614
rect 134640 17544 134852 17550
rect 139264 17756 139476 17892
rect 139672 17886 139884 17892
rect 139672 17822 139814 17886
rect 139878 17822 139884 17886
rect 139672 17816 139884 17822
rect 139672 17758 139748 17816
rect 139264 17700 139384 17756
rect 139440 17700 139476 17756
rect 139264 17614 139476 17700
rect 139617 17660 139748 17758
rect 139264 17550 139270 17614
rect 139334 17550 139476 17614
rect 139264 17544 139476 17550
rect 139672 17484 139748 17660
rect 144296 17756 144508 17892
rect 144704 17886 144916 17892
rect 144704 17822 144846 17886
rect 144910 17822 144916 17886
rect 144704 17816 144916 17822
rect 144704 17758 144780 17816
rect 144296 17700 144376 17756
rect 144432 17700 144508 17756
rect 144296 17614 144508 17700
rect 144609 17660 144780 17758
rect 144296 17550 144302 17614
rect 144366 17550 144508 17614
rect 144296 17544 144508 17550
rect 144704 17484 144780 17660
rect 149328 17756 149540 17892
rect 149736 17886 149948 17892
rect 149736 17822 149878 17886
rect 149942 17822 149948 17886
rect 149736 17816 149948 17822
rect 149736 17758 149812 17816
rect 149328 17700 149368 17756
rect 149424 17700 149540 17756
rect 149328 17620 149540 17700
rect 149601 17660 149812 17758
rect 149056 17614 149540 17620
rect 149056 17550 149062 17614
rect 149126 17550 149540 17614
rect 149056 17544 149540 17550
rect 149736 17484 149812 17660
rect 154224 17777 154436 17892
rect 154632 17886 154844 17892
rect 154632 17822 154774 17886
rect 154838 17822 154844 17886
rect 154632 17816 154844 17822
rect 154224 17756 154437 17777
rect 154632 17758 154708 17816
rect 154224 17700 154360 17756
rect 154416 17700 154437 17756
rect 154224 17679 154437 17700
rect 154224 17614 154436 17679
rect 154593 17660 154708 17758
rect 154224 17550 154230 17614
rect 154294 17550 154436 17614
rect 154224 17544 154436 17550
rect 154632 17620 154708 17660
rect 159256 17756 159468 17892
rect 159664 17886 159876 17892
rect 159664 17822 159806 17886
rect 159870 17822 159876 17886
rect 159664 17816 159876 17822
rect 159664 17758 159740 17816
rect 159256 17700 159352 17756
rect 159408 17700 159468 17756
rect 154632 17614 154806 17620
rect 159256 17614 159468 17700
rect 159585 17660 159740 17758
rect 154632 17550 154774 17614
rect 154838 17550 154844 17614
rect 159256 17550 159262 17614
rect 159326 17550 159468 17614
rect 154632 17544 154806 17550
rect 159256 17544 159468 17550
rect 159664 17484 159740 17660
rect 164288 17756 164500 17892
rect 164288 17700 164344 17756
rect 164400 17700 164500 17756
rect 164288 17614 164500 17700
rect 164288 17550 164294 17614
rect 164358 17550 164500 17614
rect 164288 17544 164500 17550
rect 164560 17886 164772 17892
rect 164560 17822 164702 17886
rect 164766 17822 164772 17886
rect 164560 17614 164772 17822
rect 164560 17550 164702 17614
rect 164766 17550 164772 17614
rect 164560 17544 164772 17550
rect 169184 17777 169396 17892
rect 169592 17886 169804 17892
rect 169592 17822 169734 17886
rect 169798 17822 169804 17886
rect 169592 17816 169804 17822
rect 169184 17756 169413 17777
rect 169592 17758 169668 17816
rect 169184 17700 169336 17756
rect 169392 17700 169413 17756
rect 169184 17679 169413 17700
rect 169184 17614 169396 17679
rect 169569 17660 169668 17758
rect 169184 17550 169190 17614
rect 169254 17550 169396 17614
rect 169184 17544 169396 17550
rect 169592 17620 169668 17660
rect 174216 17756 174428 17892
rect 174624 17886 174836 17892
rect 174624 17822 174766 17886
rect 174830 17822 174836 17886
rect 174624 17816 174836 17822
rect 174624 17758 174700 17816
rect 174216 17700 174328 17756
rect 174384 17700 174428 17756
rect 169592 17614 169766 17620
rect 174216 17614 174428 17700
rect 174561 17660 174700 17758
rect 169592 17550 169734 17614
rect 169798 17550 169804 17614
rect 174216 17550 174222 17614
rect 174286 17550 174428 17614
rect 169592 17544 169766 17550
rect 174216 17544 174428 17550
rect 174624 17484 174700 17660
rect 179248 17756 179460 17892
rect 179656 17886 179868 17892
rect 179656 17822 179798 17886
rect 179862 17822 179868 17886
rect 179656 17816 179868 17822
rect 179656 17758 179732 17816
rect 179248 17700 179320 17756
rect 179376 17700 179460 17756
rect 179248 17614 179460 17700
rect 179553 17660 179732 17758
rect 179248 17550 179254 17614
rect 179318 17550 179460 17614
rect 179248 17544 179460 17550
rect 179656 17484 179732 17660
rect 184280 17777 184356 17892
rect 184552 17886 184764 17892
rect 184552 17822 184558 17886
rect 184622 17822 184764 17886
rect 184280 17756 184389 17777
rect 184552 17758 184764 17822
rect 184280 17700 184312 17756
rect 184368 17700 184389 17756
rect 184280 17679 184389 17700
rect 184280 17614 184356 17679
rect 184545 17660 184764 17758
rect 204000 17886 204212 17892
rect 204000 17822 204006 17886
rect 204070 17822 204212 17886
rect 204000 17750 204212 17822
rect 204000 17686 204142 17750
rect 204206 17686 204212 17750
rect 204000 17680 204212 17686
rect 184280 17550 184286 17614
rect 184350 17550 184356 17614
rect 184280 17544 184356 17550
rect 184552 17614 184764 17660
rect 184552 17550 184558 17614
rect 184622 17550 184764 17614
rect 184552 17544 184764 17550
rect 1632 17348 1844 17484
rect 29822 17478 29996 17484
rect 44782 17478 44956 17484
rect 59742 17478 59916 17484
rect 74702 17478 74876 17484
rect 79734 17478 79908 17484
rect 89662 17478 89836 17484
rect 94694 17478 94868 17484
rect 104622 17478 104796 17484
rect 109654 17478 109828 17484
rect 114686 17478 114860 17484
rect 124614 17478 124788 17484
rect 129646 17478 129820 17484
rect 139574 17478 139748 17484
rect 144606 17478 144780 17484
rect 149638 17478 149812 17484
rect 159566 17478 159740 17484
rect 174526 17478 174700 17484
rect 179558 17478 179732 17484
rect 29784 17414 29790 17478
rect 29854 17414 29996 17478
rect 44744 17414 44750 17478
rect 44814 17414 44956 17478
rect 59704 17414 59710 17478
rect 59774 17414 59916 17478
rect 74664 17414 74670 17478
rect 74734 17414 74876 17478
rect 79696 17414 79702 17478
rect 79766 17414 79908 17478
rect 89624 17414 89630 17478
rect 89694 17414 89836 17478
rect 94656 17414 94662 17478
rect 94726 17414 94868 17478
rect 104584 17414 104590 17478
rect 104654 17414 104796 17478
rect 109616 17414 109622 17478
rect 109686 17414 109828 17478
rect 114648 17414 114654 17478
rect 114718 17414 114860 17478
rect 124576 17414 124582 17478
rect 124646 17414 124788 17478
rect 129608 17414 129614 17478
rect 129678 17414 129820 17478
rect 139536 17414 139542 17478
rect 139606 17414 139748 17478
rect 144568 17414 144574 17478
rect 144638 17414 144780 17478
rect 149600 17414 149606 17478
rect 149670 17414 149812 17478
rect 159528 17414 159534 17478
rect 159598 17414 159740 17478
rect 174488 17414 174494 17478
rect 174558 17414 174700 17478
rect 179520 17414 179526 17478
rect 179590 17414 179732 17478
rect 29822 17408 29996 17414
rect 44782 17408 44956 17414
rect 59742 17408 59916 17414
rect 74702 17408 74876 17414
rect 79734 17408 79908 17414
rect 89662 17408 89836 17414
rect 94694 17408 94868 17414
rect 104622 17408 104796 17414
rect 109654 17408 109828 17414
rect 114686 17408 114860 17414
rect 124614 17408 124788 17414
rect 129646 17408 129820 17414
rect 139574 17408 139748 17414
rect 144606 17408 144780 17414
rect 149638 17408 149812 17414
rect 159566 17408 159740 17414
rect 174526 17408 174700 17414
rect 179558 17408 179732 17414
rect 1224 17342 1844 17348
rect 1224 17278 1230 17342
rect 1294 17332 1844 17342
rect 1294 17278 1702 17332
rect 1224 17276 1702 17278
rect 1758 17276 1844 17332
rect 1224 17272 1844 17276
rect 1632 17136 1844 17272
rect 216784 17332 216996 17484
rect 216784 17276 216908 17332
rect 216964 17276 216996 17332
rect 216784 17212 216996 17276
rect 49776 17206 49988 17212
rect 49776 17142 49918 17206
rect 49982 17142 49988 17206
rect 49776 17136 49988 17142
rect 134640 17206 134852 17212
rect 134640 17142 134782 17206
rect 134846 17142 134852 17206
rect 134640 17136 134852 17142
rect 216784 17206 217540 17212
rect 216784 17142 217470 17206
rect 217534 17142 217540 17206
rect 216784 17136 217540 17142
rect 49776 17076 49852 17136
rect 134640 17076 134716 17136
rect 29648 17070 29860 17076
rect 29648 17006 29790 17070
rect 29854 17006 29860 17070
rect 15096 16934 15308 16940
rect 15096 16870 15102 16934
rect 15166 16870 15308 16934
rect 15096 16798 15308 16870
rect 29648 16934 29860 17006
rect 29648 16870 29790 16934
rect 29854 16870 29860 16934
rect 29648 16864 29860 16870
rect 34544 17070 35028 17076
rect 34544 17006 34958 17070
rect 35022 17006 35028 17070
rect 34544 17000 35028 17006
rect 39576 17070 39924 17076
rect 39576 17006 39854 17070
rect 39918 17006 39924 17070
rect 39576 17000 39924 17006
rect 44608 17070 44820 17076
rect 44608 17006 44750 17070
rect 44814 17006 44820 17070
rect 34544 16940 34892 17000
rect 39576 16940 39788 17000
rect 34544 16934 35028 16940
rect 34544 16870 34958 16934
rect 35022 16870 35028 16934
rect 34544 16864 35028 16870
rect 39576 16934 39924 16940
rect 39576 16870 39854 16934
rect 39918 16870 39924 16934
rect 39576 16864 39924 16870
rect 44608 16934 44820 17006
rect 44608 16870 44614 16934
rect 44678 16870 44820 16934
rect 44608 16864 44820 16870
rect 49640 17070 50124 17076
rect 49640 17006 50054 17070
rect 50118 17006 50124 17070
rect 49640 17000 50124 17006
rect 54536 17070 55020 17076
rect 54536 17006 54950 17070
rect 55014 17006 55020 17070
rect 54536 17000 55020 17006
rect 59568 17070 59780 17076
rect 59568 17006 59710 17070
rect 59774 17006 59780 17070
rect 49640 16940 49852 17000
rect 54536 16940 54748 17000
rect 49640 16934 49950 16940
rect 54536 16934 55020 16940
rect 49640 16870 49918 16934
rect 49982 16870 49988 16934
rect 54536 16870 54950 16934
rect 55014 16870 55020 16934
rect 49640 16864 49950 16870
rect 54536 16864 55020 16870
rect 59568 16934 59780 17006
rect 59568 16870 59574 16934
rect 59638 16870 59780 16934
rect 59568 16864 59780 16870
rect 64600 17070 64948 17076
rect 64600 17006 64878 17070
rect 64942 17006 64948 17070
rect 64600 17000 64948 17006
rect 69496 17070 69980 17076
rect 69496 17006 69910 17070
rect 69974 17006 69980 17070
rect 69496 17000 69980 17006
rect 74528 17070 74740 17076
rect 74528 17006 74670 17070
rect 74734 17006 74740 17070
rect 64600 16940 64812 17000
rect 69496 16940 69844 17000
rect 64600 16934 64948 16940
rect 64600 16870 64878 16934
rect 64942 16870 64948 16934
rect 64600 16864 64948 16870
rect 69496 16934 69980 16940
rect 69496 16870 69910 16934
rect 69974 16870 69980 16934
rect 69496 16864 69980 16870
rect 74528 16934 74740 17006
rect 79560 17070 79772 17076
rect 79560 17006 79702 17070
rect 79766 17006 79772 17070
rect 79560 16940 79772 17006
rect 84456 17070 84940 17076
rect 84456 17006 84870 17070
rect 84934 17006 84940 17070
rect 84456 17000 84940 17006
rect 89488 17070 89700 17076
rect 89488 17006 89630 17070
rect 89694 17006 89700 17070
rect 84456 16940 84804 17000
rect 79326 16934 80044 16940
rect 74528 16870 74670 16934
rect 74734 16870 74740 16934
rect 79288 16870 79294 16934
rect 79358 16870 79974 16934
rect 80038 16870 80044 16934
rect 74528 16864 74740 16870
rect 79326 16864 80044 16870
rect 84456 16934 84940 16940
rect 84456 16870 84870 16934
rect 84934 16870 84940 16934
rect 84456 16864 84940 16870
rect 89488 16934 89700 17006
rect 89488 16870 89630 16934
rect 89694 16870 89700 16934
rect 89488 16864 89700 16870
rect 94520 17070 94732 17076
rect 94520 17006 94662 17070
rect 94726 17006 94732 17070
rect 94520 16940 94732 17006
rect 99552 17070 99764 17076
rect 99552 17006 99694 17070
rect 99758 17006 99764 17070
rect 99552 16940 99764 17006
rect 104448 17070 104660 17076
rect 104448 17006 104590 17070
rect 104654 17006 104660 17070
rect 94520 16934 95004 16940
rect 94520 16870 94934 16934
rect 94998 16870 95004 16934
rect 94520 16864 95004 16870
rect 99552 16934 99900 16940
rect 99552 16870 99694 16934
rect 99758 16870 99830 16934
rect 99894 16870 99900 16934
rect 99552 16864 99900 16870
rect 104448 16934 104660 17006
rect 104448 16870 104454 16934
rect 104518 16870 104660 16934
rect 104448 16864 104660 16870
rect 109480 17070 109692 17076
rect 109480 17006 109622 17070
rect 109686 17006 109692 17070
rect 109480 16934 109692 17006
rect 109480 16870 109486 16934
rect 109550 16870 109692 16934
rect 109480 16864 109692 16870
rect 114512 17070 114724 17076
rect 114512 17006 114654 17070
rect 114718 17006 114724 17070
rect 114512 16934 114724 17006
rect 114512 16870 114654 16934
rect 114718 16870 114724 16934
rect 114512 16864 114724 16870
rect 119408 17070 119892 17076
rect 119408 17006 119822 17070
rect 119886 17006 119892 17070
rect 119408 17000 119892 17006
rect 124440 17070 124652 17076
rect 124440 17006 124582 17070
rect 124646 17006 124652 17070
rect 119408 16940 119756 17000
rect 124440 16940 124652 17006
rect 129472 17070 129684 17076
rect 129472 17006 129614 17070
rect 129678 17006 129684 17070
rect 129472 16940 129684 17006
rect 134504 17070 134988 17076
rect 134504 17006 134918 17070
rect 134982 17006 134988 17070
rect 134504 17000 134988 17006
rect 139400 17070 139612 17076
rect 139400 17006 139542 17070
rect 139606 17006 139612 17070
rect 134504 16940 134716 17000
rect 139400 16940 139612 17006
rect 144432 17070 144644 17076
rect 144432 17006 144574 17070
rect 144638 17006 144644 17070
rect 144432 16940 144644 17006
rect 149464 17070 149676 17076
rect 149464 17006 149606 17070
rect 149670 17006 149676 17070
rect 119408 16934 119892 16940
rect 119408 16870 119550 16934
rect 119614 16870 119822 16934
rect 119886 16870 119892 16934
rect 119408 16864 119892 16870
rect 124440 16934 124924 16940
rect 124440 16870 124854 16934
rect 124918 16870 124924 16934
rect 124440 16864 124924 16870
rect 129472 16934 129956 16940
rect 129472 16870 129886 16934
rect 129950 16870 129956 16934
rect 129472 16864 129956 16870
rect 134504 16934 134814 16940
rect 139400 16934 139884 16940
rect 134504 16870 134782 16934
rect 134846 16870 134852 16934
rect 139400 16870 139814 16934
rect 139878 16870 139884 16934
rect 134504 16864 134814 16870
rect 139400 16864 139884 16870
rect 144432 16934 144916 16940
rect 144432 16870 144846 16934
rect 144910 16870 144916 16934
rect 144432 16864 144916 16870
rect 149464 16934 149676 17006
rect 149464 16870 149470 16934
rect 149534 16870 149676 16934
rect 149464 16864 149676 16870
rect 154360 17070 154844 17076
rect 154360 17006 154774 17070
rect 154838 17006 154844 17070
rect 154360 17000 154844 17006
rect 159392 17070 159604 17076
rect 159392 17006 159534 17070
rect 159598 17006 159604 17070
rect 154360 16940 154708 17000
rect 154360 16934 154844 16940
rect 154360 16870 154774 16934
rect 154838 16870 154844 16934
rect 154360 16864 154844 16870
rect 159392 16934 159604 17006
rect 159392 16870 159534 16934
rect 159598 16870 159604 16934
rect 159392 16864 159604 16870
rect 164424 17070 164772 17076
rect 164424 17006 164702 17070
rect 164766 17006 164772 17070
rect 164424 17000 164772 17006
rect 169320 17070 169804 17076
rect 169320 17006 169734 17070
rect 169798 17006 169804 17070
rect 169320 17000 169804 17006
rect 174352 17070 174564 17076
rect 174352 17006 174494 17070
rect 174558 17006 174564 17070
rect 164424 16940 164636 17000
rect 164424 16934 164772 16940
rect 164424 16870 164702 16934
rect 164766 16870 164772 16934
rect 164424 16864 164772 16870
rect 169320 16934 169668 17000
rect 169320 16870 169462 16934
rect 169526 16870 169668 16934
rect 169320 16864 169668 16870
rect 174352 16940 174564 17006
rect 179384 17070 179596 17076
rect 179384 17006 179526 17070
rect 179590 17006 179596 17070
rect 179384 16940 179596 17006
rect 184416 17070 184628 17076
rect 184416 17006 184558 17070
rect 184622 17006 184628 17070
rect 184416 16940 184628 17006
rect 202794 17018 202860 17021
rect 203532 17018 203598 17021
rect 202794 17016 203598 17018
rect 202794 16960 202799 17016
rect 202855 16960 203537 17016
rect 203593 16960 203598 17016
rect 202794 16958 203598 16960
rect 202794 16955 202860 16958
rect 203532 16955 203598 16958
rect 204408 16945 204620 17076
rect 174352 16934 174836 16940
rect 174352 16870 174766 16934
rect 174830 16870 174836 16934
rect 174352 16864 174836 16870
rect 179384 16934 179868 16940
rect 179384 16870 179798 16934
rect 179862 16870 179868 16934
rect 179384 16864 179868 16870
rect 184416 16934 184764 16940
rect 184416 16870 184558 16934
rect 184622 16870 184694 16934
rect 184758 16870 184764 16934
rect 184416 16864 184764 16870
rect 204408 16889 204482 16945
rect 204538 16940 204620 16945
rect 204538 16889 218764 16940
rect 204408 16864 218764 16889
rect 15096 16734 15102 16798
rect 15166 16734 15308 16798
rect 15096 16728 15308 16734
rect 20400 16532 20612 16804
rect 21760 16798 21972 16804
rect 21760 16734 21766 16798
rect 21830 16734 21972 16798
rect 21760 16532 21972 16734
rect 20400 16526 21972 16532
rect 20400 16462 21766 16526
rect 21830 16462 21972 16526
rect 20400 16456 21972 16462
rect 29648 16526 29996 16532
rect 29648 16462 29926 16526
rect 29990 16462 29996 16526
rect 29648 16456 29996 16462
rect 34544 16526 34892 16532
rect 34544 16462 34822 16526
rect 34886 16462 34892 16526
rect 29648 16390 29860 16456
rect 29648 16326 29654 16390
rect 29718 16326 29860 16390
rect 29648 16320 29860 16326
rect 34544 16390 34892 16462
rect 34544 16326 34822 16390
rect 34886 16326 34892 16390
rect 34544 16320 34892 16326
rect 39576 16526 39788 16532
rect 39576 16462 39718 16526
rect 39782 16462 39788 16526
rect 39576 16390 39788 16462
rect 39576 16326 39718 16390
rect 39782 16326 39788 16390
rect 39576 16320 39788 16326
rect 44608 16526 44956 16532
rect 44608 16462 44886 16526
rect 44950 16462 44956 16526
rect 44608 16456 44956 16462
rect 49504 16526 49852 16532
rect 49504 16462 49782 16526
rect 49846 16462 49852 16526
rect 44608 16390 44820 16456
rect 44608 16326 44750 16390
rect 44814 16326 44820 16390
rect 44608 16320 44820 16326
rect 49504 16390 49852 16462
rect 49504 16326 49782 16390
rect 49846 16326 49852 16390
rect 49504 16320 49852 16326
rect 54536 16526 54884 16532
rect 54536 16462 54814 16526
rect 54878 16462 54884 16526
rect 54536 16456 54884 16462
rect 59568 16526 59916 16532
rect 59568 16462 59846 16526
rect 59910 16462 59916 16526
rect 59568 16456 59916 16462
rect 64600 16526 64812 16532
rect 64600 16462 64742 16526
rect 64806 16462 64812 16526
rect 54536 16396 54748 16456
rect 54536 16390 54884 16396
rect 54536 16326 54814 16390
rect 54878 16326 54884 16390
rect 54536 16320 54884 16326
rect 59568 16390 59780 16456
rect 59568 16326 59710 16390
rect 59774 16326 59780 16390
rect 59568 16320 59780 16326
rect 64600 16390 64812 16462
rect 64600 16326 64742 16390
rect 64806 16326 64812 16390
rect 64600 16320 64812 16326
rect 69496 16526 69844 16532
rect 69496 16462 69774 16526
rect 69838 16462 69844 16526
rect 69496 16456 69844 16462
rect 74528 16526 74876 16532
rect 74528 16462 74806 16526
rect 74870 16462 74876 16526
rect 74528 16456 74876 16462
rect 79560 16526 79908 16532
rect 79560 16462 79838 16526
rect 79902 16462 79908 16526
rect 79560 16456 79908 16462
rect 84456 16526 84804 16532
rect 84456 16462 84734 16526
rect 84798 16462 84804 16526
rect 69496 16396 69708 16456
rect 69496 16390 69844 16396
rect 69496 16326 69774 16390
rect 69838 16326 69844 16390
rect 69496 16320 69844 16326
rect 74528 16390 74740 16456
rect 74528 16326 74534 16390
rect 74598 16326 74740 16390
rect 74528 16320 74740 16326
rect 79560 16390 79772 16456
rect 79560 16326 79702 16390
rect 79766 16326 79772 16390
rect 79560 16320 79772 16326
rect 84456 16390 84804 16462
rect 84456 16326 84598 16390
rect 84662 16326 84804 16390
rect 84456 16320 84804 16326
rect 89488 16526 89836 16532
rect 89488 16462 89766 16526
rect 89830 16462 89836 16526
rect 89488 16456 89836 16462
rect 94520 16526 94868 16532
rect 94520 16462 94798 16526
rect 94862 16462 94868 16526
rect 94520 16456 94868 16462
rect 99552 16526 99764 16532
rect 99552 16462 99558 16526
rect 99622 16462 99764 16526
rect 89488 16390 89700 16456
rect 89488 16326 89494 16390
rect 89558 16326 89700 16390
rect 89488 16320 89700 16326
rect 94520 16390 94732 16456
rect 94520 16326 94662 16390
rect 94726 16326 94732 16390
rect 94520 16320 94732 16326
rect 99552 16390 99764 16462
rect 99552 16326 99558 16390
rect 99622 16326 99764 16390
rect 99552 16320 99764 16326
rect 104448 16526 104796 16532
rect 104448 16462 104726 16526
rect 104790 16462 104796 16526
rect 104448 16456 104796 16462
rect 109480 16526 109828 16532
rect 109480 16462 109758 16526
rect 109822 16462 109828 16526
rect 109480 16456 109828 16462
rect 114512 16526 114860 16532
rect 114512 16462 114790 16526
rect 114854 16462 114860 16526
rect 114512 16456 114860 16462
rect 119408 16526 119756 16532
rect 119408 16462 119686 16526
rect 119750 16462 119756 16526
rect 104448 16390 104660 16456
rect 104448 16326 104590 16390
rect 104654 16326 104660 16390
rect 104448 16320 104660 16326
rect 109480 16390 109692 16456
rect 109480 16326 109622 16390
rect 109686 16326 109692 16390
rect 109480 16320 109692 16326
rect 114512 16390 114724 16456
rect 114512 16326 114518 16390
rect 114582 16326 114724 16390
rect 114512 16320 114724 16326
rect 119408 16390 119756 16462
rect 119408 16326 119686 16390
rect 119750 16326 119756 16390
rect 119408 16320 119756 16326
rect 124440 16526 124788 16532
rect 124440 16462 124718 16526
rect 124782 16462 124788 16526
rect 124440 16456 124788 16462
rect 129472 16526 129820 16532
rect 129472 16462 129750 16526
rect 129814 16462 129820 16526
rect 129472 16456 129820 16462
rect 134368 16526 134716 16532
rect 134368 16462 134646 16526
rect 134710 16462 134716 16526
rect 124440 16390 124652 16456
rect 124440 16326 124582 16390
rect 124646 16326 124652 16390
rect 124440 16320 124652 16326
rect 129472 16390 129684 16456
rect 129472 16326 129614 16390
rect 129678 16326 129684 16390
rect 129472 16320 129684 16326
rect 134368 16390 134716 16462
rect 134368 16326 134646 16390
rect 134710 16326 134716 16390
rect 134368 16320 134716 16326
rect 139400 16526 139748 16532
rect 139400 16462 139678 16526
rect 139742 16462 139748 16526
rect 139400 16456 139748 16462
rect 144432 16526 144780 16532
rect 144432 16462 144710 16526
rect 144774 16462 144780 16526
rect 144432 16456 144780 16462
rect 149464 16526 149812 16532
rect 149464 16462 149742 16526
rect 149806 16462 149812 16526
rect 149464 16456 149812 16462
rect 154360 16526 154708 16532
rect 154360 16462 154638 16526
rect 154702 16462 154708 16526
rect 154360 16456 154708 16462
rect 159392 16526 159740 16532
rect 159392 16462 159670 16526
rect 159734 16462 159740 16526
rect 159392 16456 159740 16462
rect 164424 16526 164636 16532
rect 164424 16462 164566 16526
rect 164630 16462 164636 16526
rect 139400 16390 139612 16456
rect 139400 16326 139542 16390
rect 139606 16326 139612 16390
rect 139400 16320 139612 16326
rect 144432 16390 144644 16456
rect 144432 16326 144574 16390
rect 144638 16326 144644 16390
rect 144432 16320 144644 16326
rect 149464 16390 149676 16456
rect 149464 16326 149606 16390
rect 149670 16326 149676 16390
rect 149464 16320 149676 16326
rect 154360 16390 154572 16456
rect 154360 16326 154502 16390
rect 154566 16326 154572 16390
rect 154360 16320 154572 16326
rect 159392 16390 159604 16456
rect 159392 16326 159398 16390
rect 159462 16326 159604 16390
rect 159392 16320 159604 16326
rect 164424 16390 164636 16462
rect 164424 16326 164566 16390
rect 164630 16326 164636 16390
rect 164424 16320 164636 16326
rect 169320 16526 169668 16532
rect 169320 16462 169598 16526
rect 169662 16462 169668 16526
rect 169320 16390 169668 16462
rect 169320 16326 169598 16390
rect 169662 16326 169668 16390
rect 169320 16320 169668 16326
rect 174352 16526 174700 16532
rect 174352 16462 174630 16526
rect 174694 16462 174700 16526
rect 174352 16456 174700 16462
rect 179384 16526 179732 16532
rect 179384 16462 179662 16526
rect 179726 16462 179732 16526
rect 179384 16456 179732 16462
rect 184416 16526 184628 16532
rect 184416 16462 184422 16526
rect 184486 16462 184628 16526
rect 174352 16390 174564 16456
rect 174352 16326 174494 16390
rect 174558 16326 174564 16390
rect 174352 16320 174564 16326
rect 179384 16390 179596 16456
rect 179384 16326 179526 16390
rect 179590 16326 179596 16390
rect 179384 16320 179596 16326
rect 184416 16390 184628 16462
rect 184416 16326 184422 16390
rect 184486 16326 184628 16390
rect 184416 16320 184628 16326
rect 204000 16526 204310 16532
rect 204000 16462 204278 16526
rect 204342 16462 204348 16526
rect 204000 16456 204310 16462
rect 29784 16254 29996 16260
rect 29784 16190 29790 16254
rect 29854 16190 29996 16254
rect 29784 16124 29996 16190
rect 34680 16254 34990 16260
rect 39712 16254 39924 16260
rect 44646 16254 44956 16260
rect 34680 16190 34958 16254
rect 35022 16190 35028 16254
rect 39712 16190 39854 16254
rect 39918 16190 39924 16254
rect 44608 16190 44614 16254
rect 44678 16190 44956 16254
rect 34680 16184 34990 16190
rect 34680 16124 34892 16184
rect 39712 16124 39924 16190
rect 44646 16184 44956 16190
rect 44744 16124 44956 16184
rect 29648 16048 29996 16124
rect 29648 15852 29860 16048
rect 29278 15846 29860 15852
rect 29240 15782 29246 15846
rect 29310 15782 29860 15846
rect 29278 15776 29860 15782
rect 34544 15776 34892 16124
rect 39576 16048 39924 16124
rect 44608 16048 44956 16124
rect 49640 16254 50086 16260
rect 54672 16254 54982 16260
rect 59606 16254 59916 16260
rect 49640 16190 50054 16254
rect 50118 16190 50124 16254
rect 54672 16190 54950 16254
rect 55014 16190 55020 16254
rect 59568 16190 59574 16254
rect 59638 16190 59916 16254
rect 49640 16184 50086 16190
rect 54672 16184 54982 16190
rect 59606 16184 59916 16190
rect 49640 16048 49988 16184
rect 54672 16124 54884 16184
rect 59704 16124 59916 16184
rect 54536 16048 54884 16124
rect 59568 16048 59916 16124
rect 64600 16254 64948 16260
rect 64600 16190 64878 16254
rect 64942 16190 64948 16254
rect 64600 16048 64948 16190
rect 69632 16254 69942 16260
rect 74664 16254 74876 16260
rect 69632 16190 69910 16254
rect 69974 16190 69980 16254
rect 74664 16190 74670 16254
rect 74734 16190 74876 16254
rect 69632 16184 69942 16190
rect 39576 15776 39788 16048
rect 44608 15776 44820 16048
rect 49640 15988 49852 16048
rect 49640 15982 49988 15988
rect 49640 15918 49918 15982
rect 49982 15918 49988 15982
rect 49640 15912 49988 15918
rect 49640 15776 49852 15912
rect 54536 15776 54748 16048
rect 59568 15776 59780 16048
rect 64600 15776 64812 16048
rect 69496 15994 69572 16124
rect 69632 16048 69844 16184
rect 74664 16124 74876 16190
rect 79696 16254 80006 16260
rect 84592 16254 84902 16260
rect 89624 16254 89836 16260
rect 79696 16190 79974 16254
rect 80038 16190 80044 16254
rect 84592 16190 84870 16254
rect 84934 16190 84940 16254
rect 89624 16190 89630 16254
rect 89694 16190 89836 16254
rect 79696 16184 80006 16190
rect 84592 16184 84902 16190
rect 79696 16124 79908 16184
rect 84592 16124 84804 16184
rect 89624 16124 89836 16190
rect 94656 16254 94966 16260
rect 99552 16254 99900 16260
rect 104486 16254 104796 16260
rect 109518 16254 109828 16260
rect 94656 16190 94934 16254
rect 94998 16190 95004 16254
rect 99552 16190 99830 16254
rect 99894 16190 99900 16254
rect 104448 16190 104454 16254
rect 104518 16190 104796 16254
rect 109480 16190 109486 16254
rect 109550 16190 109828 16254
rect 94656 16184 94966 16190
rect 94656 16124 94868 16184
rect 69768 15994 69844 16048
rect 69496 15896 69844 15994
rect 69496 15776 69572 15896
rect 69768 15776 69844 15896
rect 74528 16048 74876 16124
rect 79288 16118 79908 16124
rect 79288 16054 79294 16118
rect 79358 16054 79908 16118
rect 79288 16048 79908 16054
rect 74528 15776 74740 16048
rect 79560 15776 79772 16048
rect 84456 15776 84804 16124
rect 89488 16048 89836 16124
rect 94520 16048 94868 16124
rect 99552 16118 99900 16190
rect 104486 16184 104796 16190
rect 109518 16184 109828 16190
rect 104584 16124 104796 16184
rect 109616 16124 109828 16184
rect 114648 16254 114860 16260
rect 114648 16190 114654 16254
rect 114718 16190 114860 16254
rect 114648 16124 114860 16190
rect 119544 16254 119854 16260
rect 124576 16254 124886 16260
rect 129608 16254 129918 16260
rect 134504 16254 134950 16260
rect 139536 16254 139846 16260
rect 144568 16254 144878 16260
rect 149464 16254 149812 16260
rect 119544 16190 119822 16254
rect 119886 16190 119892 16254
rect 124576 16190 124854 16254
rect 124918 16190 124924 16254
rect 129608 16190 129886 16254
rect 129950 16190 129956 16254
rect 134504 16190 134918 16254
rect 134982 16190 134988 16254
rect 139536 16190 139814 16254
rect 139878 16190 139884 16254
rect 144568 16190 144846 16254
rect 144910 16190 144916 16254
rect 149464 16190 149470 16254
rect 149534 16190 149812 16254
rect 119544 16184 119854 16190
rect 124576 16184 124886 16190
rect 129608 16184 129918 16190
rect 134504 16184 134950 16190
rect 139536 16184 139846 16190
rect 144568 16184 144878 16190
rect 119544 16124 119756 16184
rect 124576 16124 124788 16184
rect 129608 16124 129820 16184
rect 99552 16054 99694 16118
rect 99758 16054 99900 16118
rect 99552 16048 99900 16054
rect 104448 16048 104796 16124
rect 109480 16048 109828 16124
rect 114512 16048 114860 16124
rect 119408 16118 119756 16124
rect 119408 16054 119550 16118
rect 119614 16054 119756 16118
rect 89488 15776 89700 16048
rect 94520 15776 94732 16048
rect 99552 15776 99764 16048
rect 104448 15776 104660 16048
rect 109480 15776 109692 16048
rect 114512 15776 114724 16048
rect 119408 15776 119756 16054
rect 124440 16048 124788 16124
rect 129472 16048 129820 16124
rect 134504 16048 134852 16184
rect 139536 16124 139748 16184
rect 144568 16124 144780 16184
rect 139400 16048 139748 16124
rect 144432 16048 144780 16124
rect 149464 16048 149812 16190
rect 154496 16254 154806 16260
rect 159528 16254 159740 16260
rect 154496 16190 154774 16254
rect 154838 16190 154844 16254
rect 159528 16190 159534 16254
rect 159598 16190 159740 16254
rect 154496 16184 154806 16190
rect 124440 15776 124652 16048
rect 129472 15776 129684 16048
rect 134504 15988 134716 16048
rect 134504 15982 134852 15988
rect 134504 15918 134782 15982
rect 134846 15918 134852 15982
rect 134504 15912 134852 15918
rect 134504 15776 134716 15912
rect 139400 15776 139612 16048
rect 144432 15776 144644 16048
rect 149464 15776 149676 16048
rect 154360 15994 154436 16124
rect 154496 16048 154708 16184
rect 159528 16124 159740 16190
rect 164560 16254 164772 16260
rect 164560 16190 164702 16254
rect 164766 16190 164772 16254
rect 164560 16124 164772 16190
rect 169456 16254 169668 16260
rect 169456 16190 169462 16254
rect 169526 16190 169668 16254
rect 169456 16124 169668 16190
rect 174488 16254 174798 16260
rect 179520 16254 179830 16260
rect 184416 16254 184764 16260
rect 174488 16190 174766 16254
rect 174830 16190 174836 16254
rect 179520 16190 179798 16254
rect 179862 16190 179868 16254
rect 184416 16190 184694 16254
rect 184758 16190 184764 16254
rect 174488 16184 174798 16190
rect 179520 16184 179830 16190
rect 174488 16124 174700 16184
rect 179520 16124 179732 16184
rect 154632 15994 154708 16048
rect 154360 15896 154708 15994
rect 154360 15776 154436 15896
rect 154632 15776 154708 15896
rect 159392 16048 159740 16124
rect 164424 16048 164772 16124
rect 159392 15776 159604 16048
rect 164424 15776 164636 16048
rect 169320 15776 169668 16124
rect 174352 16048 174700 16124
rect 179384 16048 179732 16124
rect 184416 16118 184764 16190
rect 204000 16254 204212 16456
rect 204000 16190 204006 16254
rect 204070 16190 204212 16254
rect 204000 16184 204212 16190
rect 184416 16054 184558 16118
rect 184622 16054 184764 16118
rect 184416 16048 184764 16054
rect 174352 15776 174564 16048
rect 179384 15776 179596 16048
rect 184416 15852 184628 16048
rect 184416 15846 189252 15852
rect 184416 15782 189182 15846
rect 189246 15782 189252 15846
rect 184416 15776 189252 15782
rect 204408 15817 218764 15852
rect 204408 15761 204482 15817
rect 204538 15776 218764 15817
rect 204538 15761 204620 15776
rect 202714 15748 202780 15751
rect 203532 15748 203598 15751
rect 202714 15746 203598 15748
rect 1632 15652 1844 15716
rect 202714 15690 202719 15746
rect 202775 15690 203537 15746
rect 203593 15690 203598 15746
rect 202714 15688 203598 15690
rect 202714 15685 202780 15688
rect 203532 15685 203598 15688
rect 1632 15596 1702 15652
rect 1758 15596 1844 15652
rect 204408 15640 204620 15761
rect 216784 15710 217540 15716
rect 216784 15652 217470 15710
rect 1632 15580 1844 15596
rect 216784 15596 216908 15652
rect 216964 15646 217470 15652
rect 217534 15646 217540 15710
rect 216964 15640 217540 15646
rect 216964 15596 216996 15640
rect 1224 15574 2252 15580
rect 1224 15510 1230 15574
rect 1294 15510 2252 15574
rect 1224 15504 2252 15510
rect 2040 15368 2252 15504
rect 15096 15574 15308 15580
rect 29550 15574 29860 15580
rect 15096 15510 15238 15574
rect 15302 15510 15308 15574
rect 29512 15510 29518 15574
rect 29582 15510 29654 15574
rect 29718 15510 29860 15574
rect 15096 15438 15308 15510
rect 29550 15504 29860 15510
rect 34544 15574 34892 15580
rect 34544 15510 34822 15574
rect 34886 15510 34892 15574
rect 34544 15504 34892 15510
rect 39576 15574 39788 15580
rect 39576 15510 39718 15574
rect 39782 15510 39788 15574
rect 39576 15504 39788 15510
rect 44608 15574 44820 15580
rect 44608 15510 44750 15574
rect 44814 15510 44820 15574
rect 44608 15504 44820 15510
rect 49640 15574 49852 15580
rect 49640 15510 49782 15574
rect 49846 15510 49852 15574
rect 49640 15504 49852 15510
rect 54536 15574 54846 15580
rect 59568 15574 59780 15580
rect 54536 15510 54814 15574
rect 54878 15510 54884 15574
rect 59568 15510 59710 15574
rect 59774 15510 59780 15574
rect 54536 15504 54846 15510
rect 59568 15504 59780 15510
rect 64600 15574 64812 15580
rect 64600 15510 64742 15574
rect 64806 15510 64812 15574
rect 64600 15504 64812 15510
rect 69496 15574 69844 15580
rect 69496 15510 69774 15574
rect 69838 15510 69844 15574
rect 69496 15504 69844 15510
rect 74528 15574 74740 15580
rect 74528 15510 74534 15574
rect 74598 15510 74740 15574
rect 74528 15504 74740 15510
rect 79560 15574 79772 15580
rect 79560 15510 79702 15574
rect 79766 15510 79772 15574
rect 79560 15504 79772 15510
rect 84592 15574 84804 15580
rect 84592 15510 84598 15574
rect 84662 15510 84804 15574
rect 84592 15504 84804 15510
rect 89488 15574 89700 15580
rect 89488 15510 89494 15574
rect 89558 15510 89700 15574
rect 89488 15504 89700 15510
rect 94520 15574 94732 15580
rect 94520 15510 94662 15574
rect 94726 15510 94732 15574
rect 94520 15504 94732 15510
rect 99552 15574 99764 15580
rect 99552 15510 99558 15574
rect 99622 15510 99764 15574
rect 99552 15504 99764 15510
rect 104448 15574 104796 15580
rect 104448 15510 104590 15574
rect 104654 15510 104796 15574
rect 104448 15504 104796 15510
rect 109480 15574 109692 15580
rect 109480 15510 109622 15574
rect 109686 15510 109692 15574
rect 109480 15504 109692 15510
rect 114512 15574 114724 15580
rect 114512 15510 114518 15574
rect 114582 15510 114724 15574
rect 114512 15504 114724 15510
rect 119408 15574 119756 15580
rect 119408 15510 119686 15574
rect 119750 15510 119756 15574
rect 119408 15504 119756 15510
rect 124440 15574 124652 15580
rect 124440 15510 124582 15574
rect 124646 15510 124652 15574
rect 124440 15504 124652 15510
rect 129472 15574 129684 15580
rect 129472 15510 129614 15574
rect 129678 15510 129684 15574
rect 129472 15504 129684 15510
rect 134504 15574 134716 15580
rect 134504 15510 134646 15574
rect 134710 15510 134716 15574
rect 134504 15504 134716 15510
rect 139400 15574 139612 15580
rect 139400 15510 139542 15574
rect 139606 15510 139612 15574
rect 139400 15504 139612 15510
rect 144432 15574 144644 15580
rect 144432 15510 144574 15574
rect 144638 15510 144644 15574
rect 144432 15504 144644 15510
rect 149464 15574 149676 15580
rect 149464 15510 149606 15574
rect 149670 15510 149676 15574
rect 149464 15504 149676 15510
rect 154360 15574 154708 15580
rect 154360 15510 154502 15574
rect 154566 15510 154708 15574
rect 154360 15504 154708 15510
rect 159392 15574 159604 15580
rect 159392 15510 159398 15574
rect 159462 15510 159604 15574
rect 159392 15504 159604 15510
rect 164424 15574 164636 15580
rect 164424 15510 164566 15574
rect 164630 15510 164636 15574
rect 164424 15504 164636 15510
rect 169456 15574 169668 15580
rect 169456 15510 169598 15574
rect 169662 15510 169668 15574
rect 169456 15504 169668 15510
rect 174352 15574 174564 15580
rect 174352 15510 174494 15574
rect 174558 15510 174564 15574
rect 174352 15504 174564 15510
rect 179384 15574 179596 15580
rect 179384 15510 179526 15574
rect 179590 15510 179596 15574
rect 179384 15504 179596 15510
rect 184416 15574 189116 15580
rect 184416 15510 184422 15574
rect 184486 15510 189046 15574
rect 189110 15510 189116 15574
rect 184416 15504 189116 15510
rect 216784 15504 216996 15596
rect 29688 15480 29786 15504
rect 34680 15480 34778 15504
rect 39672 15480 39770 15504
rect 44664 15480 44762 15504
rect 49656 15480 49754 15504
rect 54648 15480 54746 15504
rect 59640 15480 59738 15504
rect 64632 15480 64730 15504
rect 69624 15480 69722 15504
rect 74616 15480 74714 15504
rect 79608 15480 79706 15504
rect 84600 15480 84698 15504
rect 89592 15480 89690 15504
rect 94584 15480 94682 15504
rect 99576 15480 99674 15504
rect 104568 15480 104666 15504
rect 109560 15480 109658 15504
rect 114552 15480 114650 15504
rect 119544 15480 119642 15504
rect 124536 15480 124634 15504
rect 129528 15480 129626 15504
rect 134520 15480 134618 15504
rect 139512 15480 139610 15504
rect 144504 15480 144602 15504
rect 149496 15480 149594 15504
rect 154488 15480 154586 15504
rect 159480 15480 159578 15504
rect 164472 15480 164570 15504
rect 169464 15480 169562 15504
rect 174456 15480 174554 15504
rect 179448 15480 179546 15504
rect 184440 15480 184538 15504
rect 15096 15374 15238 15438
rect 15302 15374 15308 15438
rect 15096 15368 15308 15374
rect 20400 15302 21972 15308
rect 20400 15238 20406 15302
rect 20470 15238 21972 15302
rect 20400 15232 21972 15238
rect 20400 15096 20612 15232
rect 21760 15166 21972 15232
rect 21760 15102 21902 15166
rect 21966 15102 21972 15166
rect 21760 15096 21972 15102
rect 28016 15166 29588 15172
rect 28016 15102 29518 15166
rect 29582 15102 29588 15166
rect 28016 15096 29588 15102
rect 189040 15166 189388 15172
rect 189040 15102 189046 15166
rect 189110 15102 189388 15166
rect 0 14960 2524 15036
rect 28016 14960 28228 15096
rect 189040 14960 189388 15102
rect 204000 15030 204212 15036
rect 204000 14966 204142 15030
rect 204206 14966 204212 15030
rect 2176 14903 2524 14960
rect 2176 14847 2326 14903
rect 2382 14847 2524 14903
rect 2176 14824 2524 14847
rect 204000 14824 204212 14966
rect 544 14214 1980 14220
rect 544 14150 550 14214
rect 614 14150 1980 14214
rect 544 14144 1980 14150
rect 1904 14084 1980 14144
rect 202634 14190 202700 14193
rect 203532 14190 203598 14193
rect 202634 14188 203598 14190
rect 202634 14132 202639 14188
rect 202695 14132 203537 14188
rect 203593 14132 203598 14188
rect 202634 14130 203598 14132
rect 202634 14127 202700 14130
rect 203532 14127 203598 14130
rect 204408 14144 218764 14220
rect 204408 14117 204620 14144
rect 1632 13972 1844 14084
rect 1904 14008 2252 14084
rect 1632 13948 1702 13972
rect 1224 13942 1702 13948
rect 1224 13878 1230 13942
rect 1294 13916 1702 13942
rect 1758 13916 1844 13972
rect 1294 13878 1844 13916
rect 1224 13872 1844 13878
rect 2040 13872 2252 14008
rect 15096 14078 15308 14084
rect 15096 14014 15102 14078
rect 15166 14014 15308 14078
rect 15096 13872 15308 14014
rect 28016 14078 29316 14084
rect 28016 14014 29246 14078
rect 29310 14014 29316 14078
rect 28016 14008 29316 14014
rect 189040 14078 189388 14084
rect 189040 14014 189182 14078
rect 189246 14014 189388 14078
rect 20400 13812 20612 13948
rect 21760 13942 21972 13948
rect 21760 13878 21766 13942
rect 21830 13878 21972 13942
rect 21760 13812 21972 13878
rect 28016 13872 28228 14008
rect 189040 13872 189388 14014
rect 204408 14061 204482 14117
rect 204538 14061 204620 14117
rect 204408 14008 204620 14061
rect 216784 14078 217540 14084
rect 216784 14014 217470 14078
rect 217534 14014 217540 14078
rect 216784 14008 217540 14014
rect 216784 13972 216996 14008
rect 216784 13916 216908 13972
rect 216964 13916 216996 13972
rect 216784 13872 216996 13916
rect 20400 13806 21972 13812
rect 20400 13742 20406 13806
rect 20470 13742 21972 13806
rect 20400 13736 21972 13742
rect 204000 13670 204212 13676
rect 204000 13606 204006 13670
rect 204070 13606 204212 13670
rect 204000 13464 204212 13606
rect 0 13328 2660 13404
rect 2584 13268 2660 13328
rect 5440 13308 5652 13404
rect 5440 13268 5511 13308
rect 0 13203 2524 13268
rect 0 13192 2326 13203
rect 2176 13147 2326 13192
rect 2382 13147 2524 13203
rect 2584 13252 5511 13268
rect 5567 13252 5652 13308
rect 2584 13192 5652 13252
rect 2176 13056 2524 13147
rect 2040 12582 2252 12724
rect 2040 12518 2046 12582
rect 2110 12518 2252 12582
rect 2040 12512 2252 12518
rect 15096 12718 15308 12724
rect 15096 12654 15238 12718
rect 15302 12654 15308 12718
rect 15096 12512 15308 12654
rect 20400 12446 21972 12452
rect 20400 12382 21902 12446
rect 21966 12382 21972 12446
rect 20400 12376 21972 12382
rect 1224 12310 2116 12316
rect 1224 12246 1230 12310
rect 1294 12292 2046 12310
rect 1294 12246 1702 12292
rect 1224 12240 1702 12246
rect 1632 12236 1702 12240
rect 1758 12246 2046 12292
rect 2110 12246 2116 12310
rect 1758 12240 2116 12246
rect 20400 12240 20612 12376
rect 21760 12240 21972 12376
rect 216784 12292 216996 12316
rect 1758 12236 1844 12240
rect 1632 12104 1844 12236
rect 216784 12236 216908 12292
rect 216964 12236 216996 12292
rect 216784 12180 216996 12236
rect 216784 12174 217540 12180
rect 216784 12110 217470 12174
rect 217534 12110 217540 12174
rect 216784 12104 217540 12110
rect 20400 11086 21972 11092
rect 20400 11022 20406 11086
rect 20470 11022 21972 11086
rect 20400 11016 21972 11022
rect 20400 10880 20612 11016
rect 21760 10880 21972 11016
rect 1224 10678 1844 10684
rect 1224 10614 1230 10678
rect 1294 10614 1844 10678
rect 1224 10612 1844 10614
rect 1224 10608 1702 10612
rect 1632 10556 1702 10608
rect 1758 10556 1844 10612
rect 1632 10472 1844 10556
rect 216784 10612 216996 10684
rect 216784 10556 216908 10612
rect 216964 10556 216996 10612
rect 216784 10548 216996 10556
rect 216784 10542 217540 10548
rect 216784 10478 217470 10542
rect 217534 10478 217540 10542
rect 216784 10472 217540 10478
rect 1224 9046 1844 9052
rect 1224 8982 1230 9046
rect 1294 8982 1844 9046
rect 1224 8976 1844 8982
rect 1632 8932 1844 8976
rect 1632 8876 1702 8932
rect 1758 8876 1844 8932
rect 1632 8840 1844 8876
rect 216784 8932 216996 9052
rect 216784 8876 216908 8932
rect 216964 8916 216996 8932
rect 216964 8910 217540 8916
rect 216964 8876 217470 8910
rect 216784 8846 217470 8876
rect 217534 8846 217540 8910
rect 216784 8840 217540 8846
rect 1632 7252 1844 7284
rect 1632 7196 1702 7252
rect 1758 7196 1844 7252
rect 1632 7148 1844 7196
rect 1224 7142 1844 7148
rect 1224 7078 1230 7142
rect 1294 7078 1844 7142
rect 1224 7072 1844 7078
rect 216784 7278 217540 7284
rect 216784 7252 217470 7278
rect 216784 7196 216908 7252
rect 216964 7214 217470 7252
rect 217534 7214 217540 7278
rect 216964 7208 217540 7214
rect 216964 7196 216996 7208
rect 216784 7072 216996 7196
rect 1632 5572 1844 5652
rect 1632 5516 1702 5572
rect 1758 5516 1844 5572
rect 1224 5510 1844 5516
rect 1224 5446 1230 5510
rect 1294 5446 1844 5510
rect 1224 5440 1844 5446
rect 216784 5646 217540 5652
rect 216784 5582 217470 5646
rect 217534 5582 217540 5646
rect 216784 5576 217540 5582
rect 216784 5572 216996 5576
rect 216784 5516 216908 5572
rect 216964 5516 216996 5572
rect 216784 5440 216996 5516
rect 1632 3892 1844 4020
rect 1632 3884 1702 3892
rect 1224 3878 1702 3884
rect 1224 3814 1230 3878
rect 1294 3836 1702 3878
rect 1758 3836 1844 3892
rect 1294 3814 1844 3836
rect 1224 3808 1844 3814
rect 216784 4014 217540 4020
rect 216784 3950 217470 4014
rect 217534 3950 217540 4014
rect 216784 3944 217540 3950
rect 216784 3892 216996 3944
rect 216784 3836 216908 3892
rect 216964 3836 216996 3892
rect 216784 3808 216996 3836
rect 16864 3672 18300 3748
rect 16864 3606 17076 3672
rect 16864 3542 16870 3606
rect 16934 3542 17076 3606
rect 16864 3536 17076 3542
rect 18088 3612 18300 3672
rect 19176 3612 19388 3748
rect 20400 3672 21836 3748
rect 20400 3612 20612 3672
rect 18088 3536 20612 3612
rect 21488 3612 21836 3672
rect 22712 3612 22924 3748
rect 23936 3672 26460 3748
rect 23936 3612 24148 3672
rect 21488 3536 24148 3612
rect 25024 3536 25236 3672
rect 26248 3612 26460 3672
rect 27336 3612 27684 3748
rect 28560 3672 29996 3748
rect 28560 3612 28772 3672
rect 26248 3536 28772 3612
rect 29784 3612 29996 3672
rect 30872 3612 31084 3748
rect 32096 3672 34620 3748
rect 32096 3612 32308 3672
rect 29784 3536 32308 3612
rect 33184 3536 33396 3672
rect 34408 3612 34620 3672
rect 35496 3672 38156 3748
rect 35496 3612 35844 3672
rect 34408 3536 35844 3612
rect 36720 3536 36932 3672
rect 37944 3612 38156 3672
rect 39032 3612 39244 3748
rect 40256 3672 41692 3748
rect 40256 3612 40468 3672
rect 37944 3536 40468 3612
rect 41344 3612 41692 3672
rect 42568 3612 42780 3748
rect 43792 3672 46316 3748
rect 43792 3612 44004 3672
rect 41344 3536 44004 3612
rect 44880 3536 45092 3672
rect 46104 3612 46316 3672
rect 47192 3612 47540 3748
rect 48416 3672 49852 3748
rect 48416 3612 48628 3672
rect 46104 3536 48628 3612
rect 49640 3612 49852 3672
rect 50728 3612 50940 3748
rect 51952 3672 54476 3748
rect 51952 3612 52164 3672
rect 49640 3536 52164 3612
rect 53040 3536 53252 3672
rect 54264 3612 54476 3672
rect 55352 3612 55700 3748
rect 56576 3672 58012 3748
rect 56576 3612 56788 3672
rect 54264 3536 56788 3612
rect 57800 3612 58012 3672
rect 58888 3612 59100 3748
rect 60112 3672 61548 3748
rect 60112 3612 60324 3672
rect 57800 3536 60324 3612
rect 61200 3536 61548 3672
rect 16456 2776 16668 2932
rect 16456 2720 16548 2776
rect 16604 2720 16668 2776
rect 16456 2654 16668 2720
rect 16456 2590 16462 2654
rect 16526 2590 16668 2654
rect 16456 2584 16668 2590
rect 17680 2776 17892 2932
rect 17680 2720 17716 2776
rect 17772 2720 17892 2776
rect 18768 2776 18980 2932
rect 18768 2720 18884 2776
rect 18940 2720 18980 2776
rect 17680 2699 17793 2720
rect 17680 2654 17756 2699
rect 17680 2590 17686 2654
rect 17750 2590 17756 2654
rect 17680 2584 17756 2590
rect 18768 2654 18980 2720
rect 18768 2590 18774 2654
rect 18838 2590 18980 2654
rect 18768 2584 18980 2590
rect 19992 2776 20204 2932
rect 21216 2797 21428 2932
rect 22440 2797 22516 2932
rect 19992 2720 20052 2776
rect 20108 2720 20204 2776
rect 19992 2654 20204 2720
rect 21199 2776 21428 2797
rect 21199 2720 21220 2776
rect 21276 2720 21428 2776
rect 22367 2776 22516 2797
rect 22367 2720 22388 2776
rect 22444 2720 22516 2776
rect 21199 2699 21297 2720
rect 21216 2660 21292 2699
rect 22367 2660 22516 2720
rect 19992 2590 19998 2654
rect 20062 2590 20204 2654
rect 19992 2584 20204 2590
rect 21080 2654 21292 2660
rect 21080 2590 21086 2654
rect 21150 2590 21292 2654
rect 21080 2584 21292 2590
rect 22304 2654 22516 2660
rect 22304 2590 22310 2654
rect 22374 2590 22516 2654
rect 22304 2584 22516 2590
rect 23528 2776 23740 2932
rect 24752 2797 24828 2932
rect 23528 2720 23556 2776
rect 23612 2720 23740 2776
rect 24703 2776 24828 2797
rect 24703 2720 24724 2776
rect 24780 2720 24828 2776
rect 23528 2699 23633 2720
rect 23528 2654 23604 2699
rect 24703 2660 24828 2720
rect 23528 2590 23534 2654
rect 23598 2590 23604 2654
rect 23528 2584 23604 2590
rect 24616 2654 24828 2660
rect 24616 2590 24622 2654
rect 24686 2590 24828 2654
rect 24616 2584 24828 2590
rect 25840 2776 26052 2932
rect 27064 2797 27140 2932
rect 28288 2797 28364 2932
rect 29376 2797 29588 2932
rect 30600 2797 30676 2932
rect 25840 2720 25892 2776
rect 25948 2720 26052 2776
rect 25840 2654 26052 2720
rect 27039 2776 27140 2797
rect 27039 2720 27060 2776
rect 27116 2720 27140 2776
rect 27039 2660 27140 2720
rect 28207 2776 28364 2797
rect 28207 2720 28228 2776
rect 28284 2720 28364 2776
rect 28207 2660 28364 2720
rect 29375 2776 29588 2797
rect 29375 2720 29396 2776
rect 29452 2720 29588 2776
rect 30543 2776 30676 2797
rect 30543 2720 30564 2776
rect 30620 2720 30676 2776
rect 29375 2699 29473 2720
rect 29376 2660 29452 2699
rect 30543 2660 30676 2720
rect 25840 2590 25982 2654
rect 26046 2590 26052 2654
rect 25840 2584 26052 2590
rect 26928 2654 27140 2660
rect 26928 2590 27070 2654
rect 27134 2590 27140 2654
rect 26928 2584 27140 2590
rect 28152 2654 28364 2660
rect 28152 2590 28294 2654
rect 28358 2590 28364 2654
rect 28152 2584 28364 2590
rect 29240 2654 29452 2660
rect 29240 2590 29246 2654
rect 29310 2590 29452 2654
rect 29240 2584 29452 2590
rect 30464 2654 30676 2660
rect 30464 2590 30606 2654
rect 30670 2590 30676 2654
rect 30464 2584 30676 2590
rect 31688 2776 31900 2932
rect 32912 2797 32988 2932
rect 34136 2797 34212 2932
rect 35224 2797 35436 2932
rect 36448 2797 36524 2932
rect 31688 2720 31732 2776
rect 31788 2720 31900 2776
rect 32879 2776 32988 2797
rect 32879 2720 32900 2776
rect 32956 2720 32988 2776
rect 31688 2699 31809 2720
rect 31688 2654 31764 2699
rect 32879 2660 32988 2720
rect 34047 2776 34212 2797
rect 34047 2720 34068 2776
rect 34124 2720 34212 2776
rect 34047 2660 34212 2720
rect 35215 2776 35436 2797
rect 35215 2720 35236 2776
rect 35292 2720 35436 2776
rect 36383 2776 36524 2797
rect 36383 2720 36404 2776
rect 36460 2720 36524 2776
rect 35215 2699 35313 2720
rect 35224 2660 35300 2699
rect 36383 2660 36524 2720
rect 31688 2590 31694 2654
rect 31758 2590 31764 2654
rect 31688 2584 31764 2590
rect 32776 2654 32988 2660
rect 32776 2590 32782 2654
rect 32846 2590 32988 2654
rect 32776 2584 32988 2590
rect 34000 2654 34212 2660
rect 34000 2590 34006 2654
rect 34070 2590 34212 2654
rect 34000 2584 34212 2590
rect 35088 2654 35300 2660
rect 35088 2590 35094 2654
rect 35158 2590 35300 2654
rect 35088 2584 35300 2590
rect 36312 2654 36524 2660
rect 36312 2590 36454 2654
rect 36518 2590 36524 2654
rect 36312 2584 36524 2590
rect 37536 2776 37748 2932
rect 38760 2797 38836 2932
rect 39984 2797 40060 2932
rect 41072 2797 41284 2932
rect 42296 2797 42372 2932
rect 37536 2720 37572 2776
rect 37628 2720 37748 2776
rect 38719 2776 38836 2797
rect 38719 2720 38740 2776
rect 38796 2720 38836 2776
rect 37536 2699 37649 2720
rect 37536 2654 37612 2699
rect 38719 2660 38836 2720
rect 39887 2776 40060 2797
rect 39887 2720 39908 2776
rect 39964 2720 40060 2776
rect 39887 2660 40060 2720
rect 41055 2776 41284 2797
rect 41055 2720 41076 2776
rect 41132 2720 41284 2776
rect 42223 2776 42372 2797
rect 42223 2720 42244 2776
rect 42300 2720 42372 2776
rect 41055 2699 41153 2720
rect 41072 2660 41148 2699
rect 42223 2660 42372 2720
rect 37536 2590 37542 2654
rect 37606 2590 37612 2654
rect 37536 2584 37612 2590
rect 38624 2654 38836 2660
rect 38624 2590 38630 2654
rect 38694 2590 38836 2654
rect 38624 2584 38836 2590
rect 39848 2654 40060 2660
rect 39848 2590 39854 2654
rect 39918 2590 40060 2654
rect 39848 2584 40060 2590
rect 40936 2654 41148 2660
rect 40936 2590 40942 2654
rect 41006 2590 41148 2654
rect 40936 2584 41148 2590
rect 42160 2654 42372 2660
rect 42160 2590 42302 2654
rect 42366 2590 42372 2654
rect 42160 2584 42372 2590
rect 43384 2776 43596 2932
rect 44608 2797 44684 2932
rect 43384 2720 43412 2776
rect 43468 2720 43596 2776
rect 44559 2776 44684 2797
rect 44559 2720 44580 2776
rect 44636 2720 44684 2776
rect 43384 2699 43489 2720
rect 43384 2654 43460 2699
rect 44559 2660 44684 2720
rect 43384 2590 43390 2654
rect 43454 2590 43460 2654
rect 43384 2584 43460 2590
rect 44472 2654 44684 2660
rect 44472 2590 44614 2654
rect 44678 2590 44684 2654
rect 44472 2584 44684 2590
rect 45696 2776 45908 2932
rect 46920 2797 46996 2932
rect 48144 2797 48220 2932
rect 49232 2797 49444 2932
rect 50456 2797 50532 2932
rect 45696 2720 45748 2776
rect 45804 2720 45908 2776
rect 45696 2654 45908 2720
rect 46895 2776 46996 2797
rect 46895 2720 46916 2776
rect 46972 2720 46996 2776
rect 46895 2660 46996 2720
rect 48063 2776 48220 2797
rect 48063 2720 48084 2776
rect 48140 2720 48220 2776
rect 48063 2660 48220 2720
rect 49231 2776 49444 2797
rect 49231 2720 49252 2776
rect 49308 2720 49444 2776
rect 50399 2776 50532 2797
rect 50399 2720 50420 2776
rect 50476 2720 50532 2776
rect 49231 2699 49329 2720
rect 49232 2660 49308 2699
rect 50399 2660 50532 2720
rect 45696 2590 45838 2654
rect 45902 2590 45908 2654
rect 45696 2584 45908 2590
rect 46784 2654 46996 2660
rect 46784 2590 46926 2654
rect 46990 2590 46996 2654
rect 46784 2584 46996 2590
rect 48008 2654 48220 2660
rect 48008 2590 48014 2654
rect 48078 2590 48220 2654
rect 48008 2584 48220 2590
rect 49096 2654 49308 2660
rect 49096 2590 49102 2654
rect 49166 2590 49308 2654
rect 49096 2584 49308 2590
rect 50320 2654 50532 2660
rect 50320 2590 50326 2654
rect 50390 2590 50532 2654
rect 50320 2584 50532 2590
rect 51544 2776 51756 2932
rect 52768 2797 52844 2932
rect 53992 2797 54068 2932
rect 55080 2797 55292 2932
rect 56304 2797 56380 2932
rect 51544 2720 51588 2776
rect 51644 2720 51756 2776
rect 52735 2776 52844 2797
rect 52735 2720 52756 2776
rect 52812 2720 52844 2776
rect 51544 2699 51665 2720
rect 51544 2654 51620 2699
rect 52735 2660 52844 2720
rect 53903 2776 54068 2797
rect 53903 2720 53924 2776
rect 53980 2720 54068 2776
rect 53903 2660 54068 2720
rect 55071 2776 55292 2797
rect 55071 2720 55092 2776
rect 55148 2720 55292 2776
rect 56239 2776 56380 2797
rect 56239 2720 56260 2776
rect 56316 2720 56380 2776
rect 55071 2699 55169 2720
rect 55080 2660 55156 2699
rect 56239 2660 56380 2720
rect 51544 2590 51550 2654
rect 51614 2590 51620 2654
rect 51544 2584 51620 2590
rect 52632 2654 52844 2660
rect 52632 2590 52774 2654
rect 52838 2590 52844 2654
rect 52632 2584 52844 2590
rect 53856 2654 54068 2660
rect 53856 2590 53862 2654
rect 53926 2590 54068 2654
rect 53856 2584 54068 2590
rect 54944 2654 55156 2660
rect 54944 2590 54950 2654
rect 55014 2590 55156 2654
rect 54944 2584 55156 2590
rect 56168 2654 56380 2660
rect 56168 2590 56174 2654
rect 56238 2590 56380 2654
rect 56168 2584 56380 2590
rect 57392 2776 57604 2932
rect 58616 2797 58692 2932
rect 59840 2797 59916 2932
rect 60928 2797 61140 2932
rect 57392 2720 57428 2776
rect 57484 2720 57604 2776
rect 58575 2776 58692 2797
rect 58575 2720 58596 2776
rect 58652 2720 58692 2776
rect 57392 2699 57505 2720
rect 57392 2654 57468 2699
rect 58575 2660 58692 2720
rect 59743 2776 59916 2797
rect 59743 2720 59764 2776
rect 59820 2720 59916 2776
rect 59743 2660 59916 2720
rect 60911 2776 61140 2797
rect 60911 2720 60932 2776
rect 60988 2720 61140 2776
rect 60911 2699 61009 2720
rect 60928 2660 61004 2699
rect 57392 2590 57398 2654
rect 57462 2590 57468 2654
rect 57392 2584 57468 2590
rect 58480 2654 58692 2660
rect 58480 2590 58622 2654
rect 58686 2590 58692 2654
rect 58480 2584 58692 2590
rect 59704 2654 59916 2660
rect 59704 2590 59846 2654
rect 59910 2590 59916 2654
rect 59704 2584 59916 2590
rect 60792 2654 61004 2660
rect 60792 2590 60798 2654
rect 60862 2590 61004 2654
rect 60792 2584 61004 2590
rect 15289 2522 15355 2525
rect 15289 2520 18158 2522
rect 15289 2464 15294 2520
rect 15350 2464 18158 2520
rect 15289 2462 18158 2464
rect 15289 2459 15355 2462
rect 1224 2246 1844 2252
rect 1224 2182 1230 2246
rect 1294 2212 1844 2246
rect 1294 2182 1702 2212
rect 1224 2176 1702 2182
rect 1632 2156 1702 2176
rect 1758 2156 1844 2212
rect 1632 2116 1844 2156
rect 16864 2116 17076 2252
rect 18088 2116 18300 2252
rect 1632 2040 1980 2116
rect 16864 2040 17212 2116
rect 18088 2040 18844 2116
rect 1904 1980 1980 2040
rect 17136 1980 17212 2040
rect 18768 1980 18844 2040
rect 19176 2040 19388 2252
rect 20400 2040 20612 2252
rect 21488 2116 21836 2252
rect 21488 2040 22244 2116
rect 19176 1980 19252 2040
rect 1904 1876 2116 1980
rect 1904 1820 2038 1876
rect 2094 1820 2116 1876
rect 1904 1768 2116 1820
rect 3672 1876 3884 1980
rect 3672 1838 3718 1876
rect 3672 1774 3678 1838
rect 3774 1820 3884 1876
rect 3742 1774 3884 1820
rect 3672 1768 3884 1774
rect 5304 1876 5516 1980
rect 5304 1820 5398 1876
rect 5454 1838 5516 1876
rect 5304 1774 5446 1820
rect 5510 1774 5516 1838
rect 5304 1768 5516 1774
rect 6936 1876 7284 1980
rect 6936 1838 7078 1876
rect 6936 1774 6942 1838
rect 7006 1820 7078 1838
rect 7134 1820 7284 1876
rect 7006 1774 7284 1820
rect 6936 1768 7284 1774
rect 8704 1876 8916 1980
rect 8704 1838 8758 1876
rect 8704 1774 8710 1838
rect 8814 1820 8916 1876
rect 8774 1774 8916 1820
rect 8704 1768 8916 1774
rect 10336 1876 10548 1980
rect 10336 1820 10438 1876
rect 10494 1838 10548 1876
rect 10336 1774 10478 1820
rect 10542 1774 10548 1838
rect 10336 1768 10548 1774
rect 11968 1876 12316 1980
rect 11968 1838 12118 1876
rect 11968 1774 12110 1838
rect 12174 1774 12316 1876
rect 11968 1768 12316 1774
rect 13736 1876 13948 1980
rect 13736 1838 13798 1876
rect 13736 1774 13742 1838
rect 13854 1820 13948 1876
rect 13806 1774 13948 1820
rect 13736 1768 13948 1774
rect 15368 1876 15580 1980
rect 15368 1820 15478 1876
rect 15534 1838 15580 1876
rect 15368 1774 15510 1820
rect 15574 1774 15580 1838
rect 15368 1768 15580 1774
rect 17136 1876 17348 1980
rect 17136 1838 17158 1876
rect 17136 1774 17142 1838
rect 17214 1820 17348 1876
rect 17206 1774 17348 1820
rect 17136 1768 17348 1774
rect 18768 1904 19252 1980
rect 20400 1980 20476 2040
rect 22168 1980 22244 2040
rect 22712 2040 22924 2252
rect 23936 2040 24148 2252
rect 25024 2116 25236 2252
rect 26248 2116 26460 2252
rect 25024 2040 25508 2116
rect 26248 2040 27276 2116
rect 22712 1980 22788 2040
rect 23936 1980 24012 2040
rect 18768 1876 18980 1904
rect 18768 1820 18838 1876
rect 18894 1844 18980 1876
rect 20400 1876 20612 1980
rect 18894 1838 19116 1844
rect 18894 1820 19046 1838
rect 18768 1774 19046 1820
rect 19110 1774 19116 1838
rect 18768 1768 19116 1774
rect 20400 1838 20518 1876
rect 20400 1774 20406 1838
rect 20470 1820 20518 1838
rect 20574 1820 20612 1876
rect 20470 1774 20612 1820
rect 20400 1768 20612 1774
rect 22168 1904 22788 1980
rect 22168 1876 22380 1904
rect 22168 1838 22198 1876
rect 22168 1774 22174 1838
rect 22254 1820 22380 1876
rect 22238 1774 22380 1820
rect 22168 1768 22380 1774
rect 23800 1876 24012 1980
rect 23800 1820 23878 1876
rect 23934 1838 24012 1876
rect 23934 1820 23942 1838
rect 23800 1774 23942 1820
rect 24006 1774 24012 1838
rect 23800 1768 24012 1774
rect 25432 1980 25508 2040
rect 27200 1980 27276 2040
rect 27336 2040 27684 2252
rect 28560 2116 28772 2252
rect 29784 2116 29996 2252
rect 28560 2040 28908 2116
rect 29784 2040 30540 2116
rect 27336 1980 27412 2040
rect 25432 1876 25644 1980
rect 25432 1838 25558 1876
rect 25432 1774 25438 1838
rect 25502 1820 25558 1838
rect 25614 1820 25644 1876
rect 25502 1774 25644 1820
rect 25432 1768 25644 1774
rect 27200 1876 27412 1980
rect 27200 1838 27238 1876
rect 27200 1774 27206 1838
rect 27294 1820 27412 1876
rect 27270 1774 27412 1820
rect 27200 1768 27412 1774
rect 28832 1980 28908 2040
rect 30464 1980 30540 2040
rect 30872 2040 31084 2252
rect 32096 2040 32308 2252
rect 33184 2116 33396 2252
rect 33184 2040 33940 2116
rect 30872 1980 30948 2040
rect 28832 1876 29044 1980
rect 28832 1838 28918 1876
rect 28832 1774 28838 1838
rect 28902 1820 28918 1838
rect 28974 1820 29044 1876
rect 28902 1774 29044 1820
rect 28832 1768 29044 1774
rect 30464 1904 30948 1980
rect 32232 1980 32308 2040
rect 33864 1980 33940 2040
rect 34408 2040 34620 2252
rect 35496 2040 35844 2252
rect 36720 2116 36932 2252
rect 36720 2040 37340 2116
rect 34408 1980 34484 2040
rect 35768 1980 35844 2040
rect 30464 1876 30676 1904
rect 30464 1838 30598 1876
rect 30464 1774 30470 1838
rect 30534 1820 30598 1838
rect 30654 1820 30676 1876
rect 30534 1774 30676 1820
rect 30464 1768 30676 1774
rect 32232 1876 32444 1980
rect 32232 1820 32278 1876
rect 32334 1838 32444 1876
rect 32334 1820 32374 1838
rect 32232 1774 32374 1820
rect 32438 1774 32444 1838
rect 32232 1768 32444 1774
rect 33864 1904 34484 1980
rect 33864 1876 34076 1904
rect 33864 1838 33958 1876
rect 33864 1774 33870 1838
rect 33934 1820 33958 1838
rect 34014 1820 34076 1876
rect 33934 1774 34076 1820
rect 33864 1768 34076 1774
rect 35496 1876 35844 1980
rect 35496 1838 35638 1876
rect 35496 1774 35502 1838
rect 35566 1820 35638 1838
rect 35694 1820 35844 1876
rect 35566 1774 35844 1820
rect 35496 1768 35844 1774
rect 37264 1980 37340 2040
rect 37944 2040 38156 2252
rect 39032 2040 39244 2252
rect 40256 2116 40468 2252
rect 40256 2040 40604 2116
rect 37944 1980 38020 2040
rect 39032 1980 39108 2040
rect 37264 1904 38020 1980
rect 37264 1876 37476 1904
rect 37264 1838 37318 1876
rect 37264 1774 37270 1838
rect 37374 1820 37476 1876
rect 37334 1774 37476 1820
rect 37264 1768 37476 1774
rect 38896 1876 39108 1980
rect 38896 1838 38998 1876
rect 38896 1774 38902 1838
rect 38966 1820 38998 1838
rect 39054 1820 39108 1876
rect 38966 1774 39108 1820
rect 38896 1768 39108 1774
rect 40528 1980 40604 2040
rect 41344 2040 41692 2252
rect 42568 2040 42780 2252
rect 43792 2040 44004 2252
rect 44880 2116 45092 2252
rect 44880 2040 45772 2116
rect 41344 1980 41420 2040
rect 42568 1980 42644 2040
rect 40528 1904 41420 1980
rect 42296 1904 42644 1980
rect 43928 1980 44004 2040
rect 45696 1980 45772 2040
rect 46104 2040 46316 2252
rect 47192 2040 47540 2252
rect 48416 2116 48628 2252
rect 48416 2040 49036 2116
rect 46104 1980 46180 2040
rect 40528 1876 40876 1904
rect 40528 1820 40678 1876
rect 40734 1838 40876 1876
rect 40734 1820 40806 1838
rect 40528 1774 40806 1820
rect 40870 1774 40876 1838
rect 40528 1768 40876 1774
rect 42296 1876 42508 1904
rect 42296 1820 42358 1876
rect 42414 1838 42508 1876
rect 42414 1820 42438 1838
rect 42296 1774 42438 1820
rect 42502 1774 42508 1838
rect 42296 1768 42508 1774
rect 43928 1876 44140 1980
rect 43928 1838 44038 1876
rect 43928 1774 43934 1838
rect 43998 1820 44038 1838
rect 44094 1820 44140 1876
rect 43998 1774 44140 1820
rect 43928 1768 44140 1774
rect 45696 1904 46180 1980
rect 47328 1980 47404 2040
rect 48960 1980 49036 2040
rect 49640 2040 49852 2252
rect 50728 2040 50940 2252
rect 51952 2116 52164 2252
rect 51952 2040 52436 2116
rect 49640 1980 49716 2040
rect 45696 1876 45908 1904
rect 45696 1838 45718 1876
rect 45696 1774 45702 1838
rect 45774 1820 45908 1876
rect 45766 1774 45908 1820
rect 45696 1768 45908 1774
rect 47328 1876 47540 1980
rect 47328 1820 47398 1876
rect 47454 1838 47540 1876
rect 47454 1820 47470 1838
rect 47328 1774 47470 1820
rect 47534 1774 47540 1838
rect 47328 1768 47540 1774
rect 48960 1904 49716 1980
rect 50728 1980 50804 2040
rect 52360 1980 52436 2040
rect 53040 2040 53252 2252
rect 54264 2040 54476 2252
rect 55352 2116 55700 2252
rect 55352 2040 55836 2116
rect 53040 1980 53116 2040
rect 54264 1980 54340 2040
rect 48960 1876 49172 1904
rect 48960 1838 49078 1876
rect 48960 1774 48966 1838
rect 49030 1820 49078 1838
rect 49134 1820 49172 1876
rect 49030 1774 49172 1820
rect 48960 1768 49172 1774
rect 50728 1876 50940 1980
rect 50728 1838 50758 1876
rect 50728 1774 50734 1838
rect 50814 1820 50940 1876
rect 50798 1774 50940 1820
rect 50728 1768 50940 1774
rect 52360 1904 53116 1980
rect 53992 1904 54340 1980
rect 55760 1980 55836 2040
rect 56576 2040 56788 2252
rect 57800 2040 58012 2252
rect 58888 2040 59100 2252
rect 60112 2116 60324 2252
rect 60112 2040 60868 2116
rect 56576 1980 56652 2040
rect 57800 1980 57876 2040
rect 55760 1904 56652 1980
rect 57392 1904 57876 1980
rect 59024 1980 59100 2040
rect 60792 1980 60868 2040
rect 61200 2040 61548 2252
rect 216784 2212 216996 2252
rect 216784 2156 216908 2212
rect 216964 2156 216996 2212
rect 216784 2116 216996 2156
rect 216784 2110 217540 2116
rect 216784 2046 217470 2110
rect 217534 2046 217540 2110
rect 216784 2040 217540 2046
rect 61200 1980 61276 2040
rect 52360 1876 52572 1904
rect 52360 1838 52438 1876
rect 52360 1774 52366 1838
rect 52430 1820 52438 1838
rect 52494 1820 52572 1876
rect 52430 1774 52572 1820
rect 52360 1768 52572 1774
rect 53992 1876 54204 1904
rect 53992 1820 54118 1876
rect 54174 1838 54204 1876
rect 53992 1774 54134 1820
rect 54198 1774 54204 1838
rect 53992 1768 54204 1774
rect 55760 1876 55972 1904
rect 55760 1820 55798 1876
rect 55854 1838 55972 1876
rect 55854 1820 55902 1838
rect 55760 1774 55902 1820
rect 55966 1774 55972 1838
rect 55760 1768 55972 1774
rect 57392 1876 57604 1904
rect 57392 1820 57478 1876
rect 57534 1844 57604 1876
rect 59024 1876 59236 1980
rect 57534 1838 57740 1844
rect 57534 1820 57670 1838
rect 57392 1774 57670 1820
rect 57734 1774 57740 1838
rect 57392 1768 57740 1774
rect 59024 1820 59158 1876
rect 59214 1838 59236 1876
rect 59024 1774 59166 1820
rect 59230 1774 59236 1838
rect 59024 1768 59236 1774
rect 60792 1904 61276 1980
rect 60792 1876 61004 1904
rect 60792 1820 60838 1876
rect 60894 1844 61004 1876
rect 62424 1876 62636 1980
rect 60894 1838 61140 1844
rect 60894 1820 61070 1838
rect 60792 1774 61070 1820
rect 61134 1774 61140 1838
rect 60792 1768 61140 1774
rect 62424 1838 62518 1876
rect 62424 1774 62430 1838
rect 62494 1820 62518 1838
rect 62574 1820 62636 1876
rect 62494 1774 62636 1820
rect 62424 1768 62636 1774
rect 64056 1876 64404 1980
rect 64056 1838 64198 1876
rect 64056 1774 64062 1838
rect 64126 1820 64198 1838
rect 64254 1820 64404 1876
rect 64126 1774 64404 1820
rect 64056 1768 64404 1774
rect 65824 1876 66036 1980
rect 65824 1820 65878 1876
rect 65934 1838 66036 1876
rect 65934 1820 65966 1838
rect 65824 1774 65966 1820
rect 66030 1774 66036 1838
rect 65824 1768 66036 1774
rect 67456 1876 67668 1980
rect 67456 1838 67558 1876
rect 67456 1774 67462 1838
rect 67526 1820 67558 1838
rect 67614 1820 67668 1876
rect 67526 1774 67668 1820
rect 67456 1768 67668 1774
rect 69088 1876 69436 1980
rect 69088 1838 69238 1876
rect 69088 1774 69230 1838
rect 69294 1774 69436 1876
rect 69088 1768 69436 1774
rect 70856 1876 71068 1980
rect 70856 1838 70918 1876
rect 70856 1774 70862 1838
rect 70974 1820 71068 1876
rect 70926 1774 71068 1820
rect 70856 1768 71068 1774
rect 72488 1876 72700 1980
rect 72488 1838 72598 1876
rect 72488 1774 72494 1838
rect 72558 1820 72598 1838
rect 72654 1820 72700 1876
rect 72558 1774 72700 1820
rect 72488 1768 72700 1774
rect 74256 1876 74468 1980
rect 74256 1838 74278 1876
rect 74256 1774 74262 1838
rect 74334 1820 74468 1876
rect 74326 1774 74468 1820
rect 74256 1768 74468 1774
rect 75888 1876 76100 1980
rect 75888 1838 75958 1876
rect 75888 1774 75894 1838
rect 76014 1820 76100 1876
rect 75958 1774 76100 1820
rect 75888 1768 76100 1774
rect 77520 1876 77732 1980
rect 77520 1820 77638 1876
rect 77694 1838 77732 1876
rect 77520 1774 77662 1820
rect 77726 1774 77732 1838
rect 77520 1768 77732 1774
rect 79288 1876 79500 1980
rect 79288 1838 79318 1876
rect 79288 1774 79294 1838
rect 79374 1820 79500 1876
rect 79358 1774 79500 1820
rect 79288 1768 79500 1774
rect 80920 1876 81132 1980
rect 80920 1838 80998 1876
rect 80920 1774 80926 1838
rect 80990 1820 80998 1838
rect 81054 1820 81132 1876
rect 80990 1774 81132 1820
rect 80920 1768 81132 1774
rect 82552 1876 82764 1980
rect 82552 1820 82678 1876
rect 82734 1838 82764 1876
rect 82552 1774 82694 1820
rect 82758 1774 82764 1838
rect 82552 1768 82764 1774
rect 84320 1876 84532 1980
rect 84320 1820 84358 1876
rect 84414 1844 84532 1876
rect 85952 1876 86164 1980
rect 84414 1838 84668 1844
rect 84414 1820 84598 1838
rect 84320 1774 84598 1820
rect 84662 1774 84668 1838
rect 84320 1768 84668 1774
rect 85952 1838 86038 1876
rect 85952 1774 85958 1838
rect 86022 1820 86038 1838
rect 86094 1820 86164 1876
rect 86022 1774 86164 1820
rect 85952 1768 86164 1774
rect 87584 1876 87796 1980
rect 87584 1820 87718 1876
rect 87774 1838 87796 1876
rect 87584 1774 87726 1820
rect 87790 1774 87796 1838
rect 87584 1768 87796 1774
rect 89352 1876 89564 1980
rect 89352 1820 89398 1876
rect 89454 1838 89564 1876
rect 89454 1820 89494 1838
rect 89352 1774 89494 1820
rect 89558 1774 89564 1838
rect 89352 1768 89564 1774
rect 90984 1876 91196 1980
rect 90984 1820 91078 1876
rect 91134 1838 91196 1876
rect 90984 1774 91126 1820
rect 91190 1774 91196 1838
rect 90984 1768 91196 1774
rect 92616 1876 92964 1980
rect 92616 1838 92758 1876
rect 92616 1774 92622 1838
rect 92686 1820 92758 1838
rect 92814 1820 92964 1876
rect 92686 1774 92964 1820
rect 92616 1768 92964 1774
rect 94384 1876 94596 1980
rect 94384 1820 94438 1876
rect 94494 1844 94596 1876
rect 96016 1876 96228 1980
rect 94494 1838 94732 1844
rect 94494 1820 94662 1838
rect 94384 1774 94662 1820
rect 94726 1774 94732 1838
rect 94384 1768 94732 1774
rect 96016 1820 96118 1876
rect 96174 1838 96228 1876
rect 96016 1774 96158 1820
rect 96222 1774 96228 1838
rect 96016 1768 96228 1774
rect 97648 1876 97996 1980
rect 97648 1838 97798 1876
rect 97648 1774 97790 1838
rect 97854 1774 97996 1876
rect 97648 1768 97996 1774
rect 99416 1876 99628 1980
rect 99416 1820 99478 1876
rect 99534 1838 99628 1876
rect 99534 1820 99558 1838
rect 99416 1774 99558 1820
rect 99622 1774 99628 1838
rect 99416 1768 99628 1774
rect 101048 1876 101260 1980
rect 101048 1820 101158 1876
rect 101214 1838 101260 1876
rect 101048 1774 101190 1820
rect 101254 1774 101260 1838
rect 101048 1768 101260 1774
rect 102816 1876 103028 1980
rect 102816 1820 102838 1876
rect 102894 1838 103028 1876
rect 102894 1820 102958 1838
rect 102816 1774 102958 1820
rect 103022 1774 103028 1838
rect 102816 1768 103028 1774
rect 104448 1876 104660 1980
rect 104448 1838 104518 1876
rect 104448 1774 104454 1838
rect 104574 1820 104660 1876
rect 104518 1774 104660 1820
rect 104448 1768 104660 1774
rect 106080 1876 106292 1980
rect 106080 1820 106198 1876
rect 106254 1838 106292 1876
rect 106080 1774 106222 1820
rect 106286 1774 106292 1838
rect 106080 1768 106292 1774
rect 107848 1876 108060 1980
rect 107848 1838 107878 1876
rect 107848 1774 107854 1838
rect 107934 1820 108060 1876
rect 107918 1774 108060 1820
rect 107848 1768 108060 1774
rect 109480 1876 109692 1980
rect 109480 1838 109558 1876
rect 109480 1774 109486 1838
rect 109550 1820 109558 1838
rect 109614 1820 109692 1876
rect 109550 1774 109692 1820
rect 109480 1768 109692 1774
rect 111112 1876 111324 1980
rect 111112 1838 111238 1876
rect 111112 1774 111118 1838
rect 111182 1820 111238 1838
rect 111294 1820 111324 1876
rect 111182 1774 111324 1820
rect 111112 1768 111324 1774
rect 112880 1876 113092 1980
rect 112880 1838 112918 1876
rect 112880 1774 112886 1838
rect 112974 1820 113092 1876
rect 112950 1774 113092 1820
rect 112880 1768 113092 1774
rect 114512 1876 114724 1980
rect 114512 1820 114598 1876
rect 114654 1838 114724 1876
rect 114512 1774 114654 1820
rect 114718 1774 114724 1838
rect 114512 1768 114724 1774
rect 116144 1876 116356 1980
rect 116144 1838 116278 1876
rect 116144 1774 116150 1838
rect 116214 1820 116278 1838
rect 116334 1820 116356 1876
rect 116214 1774 116356 1820
rect 116144 1768 116356 1774
rect 117912 1876 118124 1980
rect 117912 1838 117958 1876
rect 117912 1774 117918 1838
rect 118014 1820 118124 1876
rect 117982 1774 118124 1820
rect 117912 1768 118124 1774
rect 119544 1876 119756 1980
rect 119544 1820 119638 1876
rect 119694 1838 119756 1876
rect 119544 1774 119686 1820
rect 119750 1774 119756 1838
rect 119544 1768 119756 1774
rect 121176 1876 121524 1980
rect 121176 1820 121318 1876
rect 121374 1838 121524 1876
rect 121374 1820 121454 1838
rect 121176 1774 121454 1820
rect 121518 1774 121524 1838
rect 121176 1768 121524 1774
rect 122944 1876 123156 1980
rect 122944 1838 122998 1876
rect 122944 1774 122950 1838
rect 123054 1820 123156 1876
rect 123014 1774 123156 1820
rect 122944 1768 123156 1774
rect 124576 1876 124788 1980
rect 124576 1820 124678 1876
rect 124734 1838 124788 1876
rect 124576 1774 124718 1820
rect 124782 1774 124788 1838
rect 124576 1768 124788 1774
rect 126208 1876 126556 1980
rect 126208 1838 126358 1876
rect 126208 1774 126214 1838
rect 126278 1820 126358 1838
rect 126414 1820 126556 1876
rect 126278 1774 126556 1820
rect 126208 1768 126556 1774
rect 127976 1876 128188 1980
rect 127976 1838 128038 1876
rect 127976 1774 127982 1838
rect 128094 1820 128188 1876
rect 128046 1774 128188 1820
rect 127976 1768 128188 1774
rect 129608 1876 129820 1980
rect 129608 1838 129718 1876
rect 129608 1774 129614 1838
rect 129678 1820 129718 1838
rect 129774 1820 129820 1876
rect 129678 1774 129820 1820
rect 129608 1768 129820 1774
rect 131376 1876 131588 1980
rect 131376 1838 131398 1876
rect 131376 1774 131382 1838
rect 131454 1820 131588 1876
rect 131446 1774 131588 1820
rect 131376 1768 131588 1774
rect 133008 1876 133220 1980
rect 133008 1820 133078 1876
rect 133134 1838 133220 1876
rect 133134 1820 133150 1838
rect 133008 1774 133150 1820
rect 133214 1774 133220 1838
rect 133008 1768 133220 1774
rect 134640 1876 134852 1980
rect 134640 1838 134758 1876
rect 134640 1774 134646 1838
rect 134710 1820 134758 1838
rect 134814 1820 134852 1876
rect 134710 1774 134852 1820
rect 134640 1768 134852 1774
rect 136408 1876 136620 1980
rect 136408 1838 136438 1876
rect 136408 1774 136414 1838
rect 136494 1820 136620 1876
rect 136478 1774 136620 1820
rect 136408 1768 136620 1774
rect 138040 1876 138252 1980
rect 138040 1820 138118 1876
rect 138174 1838 138252 1876
rect 138174 1820 138182 1838
rect 138040 1774 138182 1820
rect 138246 1774 138252 1838
rect 138040 1768 138252 1774
rect 139672 1876 139884 1980
rect 139672 1838 139798 1876
rect 139672 1774 139678 1838
rect 139742 1820 139798 1838
rect 139854 1820 139884 1876
rect 139742 1774 139884 1820
rect 139672 1768 139884 1774
rect 141440 1876 141652 1980
rect 141440 1838 141478 1876
rect 141440 1774 141446 1838
rect 141534 1820 141652 1876
rect 141510 1774 141652 1820
rect 141440 1768 141652 1774
rect 143072 1876 143284 1980
rect 143072 1820 143158 1876
rect 143214 1838 143284 1876
rect 143072 1774 143214 1820
rect 143278 1774 143284 1838
rect 143072 1768 143284 1774
rect 144704 1876 144916 1980
rect 144704 1838 144838 1876
rect 144704 1774 144710 1838
rect 144774 1820 144838 1838
rect 144894 1820 144916 1876
rect 144774 1774 144916 1820
rect 144704 1768 144916 1774
rect 146472 1876 146684 1980
rect 146472 1838 146518 1876
rect 146472 1774 146478 1838
rect 146574 1820 146684 1876
rect 146542 1774 146684 1820
rect 146472 1768 146684 1774
rect 148104 1876 148316 1980
rect 148104 1838 148198 1876
rect 148104 1774 148110 1838
rect 148174 1820 148198 1838
rect 148254 1820 148316 1876
rect 148174 1774 148316 1820
rect 148104 1768 148316 1774
rect 149736 1876 150084 1980
rect 149736 1820 149878 1876
rect 149934 1838 150084 1876
rect 149934 1820 150014 1838
rect 149736 1774 150014 1820
rect 150078 1774 150084 1838
rect 149736 1768 150084 1774
rect 151504 1876 151716 1980
rect 151504 1820 151558 1876
rect 151614 1838 151716 1876
rect 151614 1820 151646 1838
rect 151504 1774 151646 1820
rect 151710 1774 151716 1838
rect 151504 1768 151716 1774
rect 153136 1876 153348 1980
rect 153136 1838 153238 1876
rect 153136 1774 153142 1838
rect 153206 1820 153238 1838
rect 153294 1820 153348 1876
rect 153206 1774 153348 1820
rect 153136 1768 153348 1774
rect 154768 1876 155116 1980
rect 154768 1838 154918 1876
rect 154768 1774 154910 1838
rect 154974 1774 155116 1876
rect 154768 1768 155116 1774
rect 156536 1876 156748 1980
rect 156536 1820 156598 1876
rect 156654 1838 156748 1876
rect 156654 1820 156678 1838
rect 156536 1774 156678 1820
rect 156742 1774 156748 1838
rect 156536 1768 156748 1774
rect 158168 1876 158380 1980
rect 158168 1838 158278 1876
rect 158168 1774 158174 1838
rect 158238 1820 158278 1838
rect 158334 1820 158380 1876
rect 158238 1774 158380 1820
rect 158168 1768 158380 1774
rect 159936 1876 160148 1980
rect 159936 1838 159958 1876
rect 159936 1774 159942 1838
rect 160014 1820 160148 1876
rect 160006 1774 160148 1820
rect 159936 1768 160148 1774
rect 161568 1876 161780 1980
rect 161568 1820 161638 1876
rect 161694 1838 161780 1876
rect 161694 1820 161710 1838
rect 161568 1774 161710 1820
rect 161774 1774 161780 1838
rect 161568 1768 161780 1774
rect 163200 1876 163412 1980
rect 163200 1838 163318 1876
rect 163200 1774 163206 1838
rect 163270 1820 163318 1838
rect 163374 1820 163412 1876
rect 163270 1774 163412 1820
rect 163200 1768 163412 1774
rect 164968 1876 165180 1980
rect 164968 1838 164998 1876
rect 164968 1774 164974 1838
rect 165054 1820 165180 1876
rect 165038 1774 165180 1820
rect 164968 1768 165180 1774
rect 166600 1876 166812 1980
rect 166600 1838 166678 1876
rect 166600 1774 166606 1838
rect 166670 1820 166678 1838
rect 166734 1820 166812 1876
rect 166670 1774 166812 1820
rect 166600 1768 166812 1774
rect 168232 1876 168444 1980
rect 168232 1820 168358 1876
rect 168414 1838 168444 1876
rect 168232 1774 168374 1820
rect 168438 1774 168444 1838
rect 168232 1768 168444 1774
rect 170000 1876 170212 1980
rect 170000 1820 170038 1876
rect 170094 1838 170212 1876
rect 170094 1820 170142 1838
rect 170000 1774 170142 1820
rect 170206 1774 170212 1838
rect 170000 1768 170212 1774
rect 171632 1876 171844 1980
rect 171632 1838 171718 1876
rect 171632 1774 171638 1838
rect 171702 1820 171718 1838
rect 171774 1820 171844 1876
rect 171702 1774 171844 1820
rect 171632 1768 171844 1774
rect 173264 1876 173476 1980
rect 173264 1820 173398 1876
rect 173454 1838 173476 1876
rect 173264 1774 173406 1820
rect 173470 1774 173476 1838
rect 173264 1768 173476 1774
rect 175032 1876 175244 1980
rect 175032 1820 175078 1876
rect 175134 1838 175244 1876
rect 175134 1820 175174 1838
rect 175032 1774 175174 1820
rect 175238 1774 175244 1838
rect 175032 1768 175244 1774
rect 176664 1876 176876 1980
rect 176664 1838 176758 1876
rect 176664 1774 176670 1838
rect 176734 1820 176758 1838
rect 176814 1820 176876 1876
rect 176734 1774 176876 1820
rect 176664 1768 176876 1774
rect 178296 1876 178644 1980
rect 178296 1774 178438 1876
rect 178494 1838 178644 1876
rect 178502 1774 178644 1838
rect 178296 1768 178644 1774
rect 180064 1876 180276 1980
rect 180064 1820 180118 1876
rect 180174 1838 180276 1876
rect 180174 1820 180206 1838
rect 180064 1774 180206 1820
rect 180270 1774 180276 1838
rect 180064 1768 180276 1774
rect 181696 1876 181908 1980
rect 181696 1838 181798 1876
rect 181696 1774 181702 1838
rect 181766 1820 181798 1838
rect 181854 1820 181908 1876
rect 181766 1774 181908 1820
rect 181696 1768 181908 1774
rect 183328 1876 183676 1980
rect 183328 1838 183478 1876
rect 183328 1774 183470 1838
rect 183534 1774 183676 1876
rect 183328 1768 183676 1774
rect 185096 1876 185308 1980
rect 185096 1838 185158 1876
rect 185096 1774 185102 1838
rect 185214 1820 185308 1876
rect 185166 1774 185308 1820
rect 185096 1768 185308 1774
rect 186728 1876 186940 1980
rect 186728 1820 186838 1876
rect 186894 1838 186940 1876
rect 186728 1774 186870 1820
rect 186934 1774 186940 1838
rect 186728 1768 186940 1774
rect 188496 1876 188708 1980
rect 188496 1820 188518 1876
rect 188574 1838 188708 1876
rect 188574 1820 188638 1838
rect 188496 1774 188638 1820
rect 188702 1774 188708 1838
rect 188496 1768 188708 1774
rect 190128 1876 190340 1980
rect 190128 1838 190198 1876
rect 190128 1774 190134 1838
rect 190254 1820 190340 1876
rect 190198 1774 190340 1820
rect 190128 1768 190340 1774
rect 191760 1876 191972 1980
rect 191760 1820 191878 1876
rect 191934 1838 191972 1876
rect 191760 1774 191902 1820
rect 191966 1774 191972 1838
rect 191760 1768 191972 1774
rect 193528 1876 193740 1980
rect 193528 1820 193558 1876
rect 193614 1838 193740 1876
rect 193614 1820 193670 1838
rect 193528 1774 193670 1820
rect 193734 1774 193740 1838
rect 193528 1768 193740 1774
rect 195160 1876 195372 1980
rect 195160 1838 195238 1876
rect 195160 1774 195166 1838
rect 195230 1820 195238 1838
rect 195294 1820 195372 1876
rect 195230 1774 195372 1820
rect 195160 1768 195372 1774
rect 196792 1876 197004 1980
rect 196792 1820 196918 1876
rect 196974 1838 197004 1876
rect 196792 1774 196934 1820
rect 196998 1774 197004 1838
rect 196792 1768 197004 1774
rect 198560 1876 198772 1980
rect 198560 1820 198598 1876
rect 198654 1838 198772 1876
rect 198654 1820 198702 1838
rect 198560 1774 198702 1820
rect 198766 1774 198772 1838
rect 198560 1768 198772 1774
rect 200192 1876 200404 1980
rect 200192 1838 200278 1876
rect 200192 1774 200198 1838
rect 200262 1820 200278 1838
rect 200334 1820 200404 1876
rect 200262 1774 200404 1820
rect 200192 1768 200404 1774
rect 201824 1876 202036 1980
rect 201824 1820 201958 1876
rect 202014 1838 202036 1876
rect 201824 1774 201966 1820
rect 202030 1774 202036 1838
rect 201824 1768 202036 1774
rect 203592 1876 203804 1980
rect 203592 1838 203638 1876
rect 203592 1774 203598 1838
rect 203694 1820 203804 1876
rect 203662 1774 203804 1820
rect 203592 1768 203804 1774
rect 205224 1876 205436 1980
rect 205224 1838 205318 1876
rect 205224 1774 205230 1838
rect 205294 1820 205318 1838
rect 205374 1820 205436 1876
rect 205294 1774 205436 1820
rect 205224 1768 205436 1774
rect 206856 1876 207204 1980
rect 206856 1820 206998 1876
rect 207054 1838 207204 1876
rect 207054 1820 207134 1838
rect 206856 1774 207134 1820
rect 207198 1774 207204 1838
rect 206856 1768 207204 1774
rect 208624 1876 208836 1980
rect 208624 1838 208678 1876
rect 208624 1774 208630 1838
rect 208734 1820 208836 1876
rect 208694 1774 208836 1820
rect 208624 1768 208836 1774
rect 210256 1876 210468 1980
rect 210256 1820 210358 1876
rect 210414 1838 210468 1876
rect 210256 1774 210398 1820
rect 210462 1774 210468 1838
rect 210256 1768 210468 1774
rect 211888 1876 212236 1980
rect 211888 1838 212038 1876
rect 211888 1774 211894 1838
rect 211958 1820 212038 1838
rect 212094 1820 212236 1876
rect 211958 1774 212236 1820
rect 211888 1768 212236 1774
rect 213656 1876 213868 1980
rect 213656 1838 213718 1876
rect 213656 1774 213662 1838
rect 213774 1820 213868 1876
rect 213726 1774 213868 1820
rect 213656 1768 213868 1774
rect 215288 1876 215500 1980
rect 215288 1820 215398 1876
rect 215454 1838 215500 1876
rect 215288 1774 215430 1820
rect 215494 1774 215500 1838
rect 215288 1768 215500 1774
rect 952 1294 217812 1300
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 3678 1294
rect 3742 1230 5446 1294
rect 5510 1230 6942 1294
rect 7006 1230 8710 1294
rect 8774 1230 10478 1294
rect 10542 1230 12110 1294
rect 12174 1230 13742 1294
rect 13806 1230 15510 1294
rect 15574 1230 17142 1294
rect 17206 1230 19046 1294
rect 19110 1230 20406 1294
rect 20470 1230 22174 1294
rect 22238 1230 23942 1294
rect 24006 1230 25438 1294
rect 25502 1230 27206 1294
rect 27270 1230 28838 1294
rect 28902 1230 30470 1294
rect 30534 1230 32374 1294
rect 32438 1230 33870 1294
rect 33934 1230 35502 1294
rect 35566 1230 37270 1294
rect 37334 1230 38902 1294
rect 38966 1230 40806 1294
rect 40870 1230 42438 1294
rect 42502 1230 43934 1294
rect 43998 1230 45702 1294
rect 45766 1230 47470 1294
rect 47534 1230 48966 1294
rect 49030 1230 50734 1294
rect 50798 1230 52366 1294
rect 52430 1230 54134 1294
rect 54198 1230 55902 1294
rect 55966 1230 57670 1294
rect 57734 1230 59166 1294
rect 59230 1230 61070 1294
rect 61134 1230 62430 1294
rect 62494 1230 64062 1294
rect 64126 1230 65966 1294
rect 66030 1230 67462 1294
rect 67526 1230 69230 1294
rect 69294 1230 70862 1294
rect 70926 1230 72494 1294
rect 72558 1230 74262 1294
rect 74326 1230 75894 1294
rect 75958 1230 77662 1294
rect 77726 1230 79294 1294
rect 79358 1230 80926 1294
rect 80990 1230 82694 1294
rect 82758 1230 84598 1294
rect 84662 1230 85958 1294
rect 86022 1230 87726 1294
rect 87790 1230 89494 1294
rect 89558 1230 91126 1294
rect 91190 1230 92622 1294
rect 92686 1230 94662 1294
rect 94726 1230 96158 1294
rect 96222 1230 97790 1294
rect 97854 1230 99558 1294
rect 99622 1230 101190 1294
rect 101254 1230 102958 1294
rect 103022 1230 104454 1294
rect 104518 1230 106222 1294
rect 106286 1230 107854 1294
rect 107918 1230 109486 1294
rect 109550 1230 111118 1294
rect 111182 1230 112886 1294
rect 112950 1230 114654 1294
rect 114718 1230 116150 1294
rect 116214 1230 117918 1294
rect 117982 1230 119686 1294
rect 119750 1230 121454 1294
rect 121518 1230 122950 1294
rect 123014 1230 124718 1294
rect 124782 1230 126214 1294
rect 126278 1230 127982 1294
rect 128046 1230 129614 1294
rect 129678 1230 131382 1294
rect 131446 1230 133150 1294
rect 133214 1230 134646 1294
rect 134710 1230 136414 1294
rect 136478 1230 138182 1294
rect 138246 1230 139678 1294
rect 139742 1230 141446 1294
rect 141510 1230 143214 1294
rect 143278 1230 144710 1294
rect 144774 1230 146478 1294
rect 146542 1230 148110 1294
rect 148174 1230 150014 1294
rect 150078 1230 151646 1294
rect 151710 1230 153142 1294
rect 153206 1230 154910 1294
rect 154974 1230 156678 1294
rect 156742 1230 158174 1294
rect 158238 1230 159942 1294
rect 160006 1230 161710 1294
rect 161774 1230 163206 1294
rect 163270 1230 164974 1294
rect 165038 1230 166606 1294
rect 166670 1230 168374 1294
rect 168438 1230 170142 1294
rect 170206 1230 171638 1294
rect 171702 1230 173406 1294
rect 173470 1230 175174 1294
rect 175238 1230 176670 1294
rect 176734 1230 178438 1294
rect 178502 1230 180206 1294
rect 180270 1230 181702 1294
rect 181766 1230 183470 1294
rect 183534 1230 185102 1294
rect 185166 1230 186870 1294
rect 186934 1230 188638 1294
rect 188702 1230 190134 1294
rect 190198 1230 191902 1294
rect 191966 1230 193670 1294
rect 193734 1230 195166 1294
rect 195230 1230 196934 1294
rect 196998 1230 198702 1294
rect 198766 1230 200198 1294
rect 200262 1230 201966 1294
rect 202030 1230 203598 1294
rect 203662 1230 205230 1294
rect 205294 1230 207134 1294
rect 207198 1230 208630 1294
rect 208694 1230 210398 1294
rect 210462 1230 211894 1294
rect 211958 1230 213662 1294
rect 213726 1230 215430 1294
rect 215494 1230 217470 1294
rect 217534 1230 217606 1294
rect 217670 1230 217742 1294
rect 217806 1230 217812 1294
rect 952 1158 217812 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 217470 1158
rect 217534 1094 217606 1158
rect 217670 1094 217742 1158
rect 217806 1094 217812 1158
rect 952 1022 217812 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 217470 1022
rect 217534 958 217606 1022
rect 217670 958 217742 1022
rect 217806 958 217812 1022
rect 952 952 217812 958
rect 272 614 218492 620
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 16870 614
rect 16934 550 218150 614
rect 218214 550 218286 614
rect 218350 550 218422 614
rect 218486 550 218492 614
rect 272 478 218492 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 218150 478
rect 218214 414 218286 478
rect 218350 414 218422 478
rect 218486 414 218492 478
rect 272 342 218492 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 218150 342
rect 218214 278 218286 342
rect 218350 278 218422 342
rect 218486 278 218492 342
rect 272 272 218492 278
<< via3 >>
rect 278 143758 342 143822
rect 414 143758 478 143822
rect 550 143758 614 143822
rect 218150 143758 218214 143822
rect 218286 143758 218350 143822
rect 218422 143758 218486 143822
rect 278 143622 342 143686
rect 414 143622 478 143686
rect 550 143622 614 143686
rect 218150 143622 218214 143686
rect 218286 143622 218350 143686
rect 218422 143622 218486 143686
rect 278 143486 342 143550
rect 414 143486 478 143550
rect 550 143486 614 143550
rect 198158 143486 198222 143550
rect 218150 143486 218214 143550
rect 218286 143486 218350 143550
rect 218422 143486 218486 143550
rect 958 143078 1022 143142
rect 1094 143078 1158 143142
rect 1230 143078 1294 143142
rect 217470 143078 217534 143142
rect 217606 143078 217670 143142
rect 217742 143078 217806 143142
rect 958 142942 1022 143006
rect 1094 142942 1158 143006
rect 1230 142942 1294 143006
rect 217470 142942 217534 143006
rect 217606 142942 217670 143006
rect 217742 142942 217806 143006
rect 958 142806 1022 142870
rect 1094 142806 1158 142870
rect 1230 142806 1294 142870
rect 1910 142806 1974 142870
rect 3678 142806 3742 142870
rect 5446 142806 5510 142870
rect 7214 142806 7278 142870
rect 8710 142806 8774 142870
rect 10478 142806 10542 142870
rect 12246 142806 12310 142870
rect 13742 142806 13806 142870
rect 15374 142806 15438 142870
rect 17142 142806 17206 142870
rect 18910 142806 18974 142870
rect 20406 142806 20470 142870
rect 22174 142806 22238 142870
rect 23942 142806 24006 142870
rect 25438 142806 25502 142870
rect 27206 142806 27270 142870
rect 28974 142806 29038 142870
rect 30470 142806 30534 142870
rect 32238 142806 32302 142870
rect 33870 142806 33934 142870
rect 35502 142806 35566 142870
rect 37406 142806 37470 142870
rect 38902 142806 38966 142870
rect 40670 142806 40734 142870
rect 42438 142806 42502 142870
rect 43934 142806 43998 142870
rect 45702 142806 45766 142870
rect 47470 142806 47534 142870
rect 48966 142806 49030 142870
rect 50734 142806 50798 142870
rect 52366 142806 52430 142870
rect 53998 142806 54062 142870
rect 55902 142806 55966 142870
rect 57398 142806 57462 142870
rect 59166 142806 59230 142870
rect 60934 142806 60998 142870
rect 62430 142806 62494 142870
rect 64062 142806 64126 142870
rect 65966 142806 66030 142870
rect 67462 142806 67526 142870
rect 69366 142806 69430 142870
rect 70862 142806 70926 142870
rect 72494 142806 72558 142870
rect 74262 142806 74326 142870
rect 75894 142806 75958 142870
rect 77662 142806 77726 142870
rect 79430 142806 79494 142870
rect 80926 142806 80990 142870
rect 82694 142806 82758 142870
rect 84598 142806 84662 142870
rect 85958 142806 86022 142870
rect 87726 142806 87790 142870
rect 89494 142806 89558 142870
rect 90990 142806 91054 142870
rect 92894 142806 92958 142870
rect 94390 142806 94454 142870
rect 96158 142806 96222 142870
rect 97790 142806 97854 142870
rect 99558 142806 99622 142870
rect 101190 142806 101254 142870
rect 102958 142806 103022 142870
rect 104454 142806 104518 142870
rect 106222 142806 106286 142870
rect 107854 142806 107918 142870
rect 109622 142806 109686 142870
rect 111118 142806 111182 142870
rect 112886 142806 112950 142870
rect 114654 142806 114718 142870
rect 116150 142806 116214 142870
rect 117918 142806 117982 142870
rect 119686 142806 119750 142870
rect 121318 142806 121382 142870
rect 122950 142806 123014 142870
rect 124718 142806 124782 142870
rect 126214 142806 126278 142870
rect 127982 142806 128046 142870
rect 129614 142806 129678 142870
rect 131382 142806 131446 142870
rect 133150 142806 133214 142870
rect 134646 142806 134710 142870
rect 136414 142806 136478 142870
rect 138182 142806 138246 142870
rect 139678 142806 139742 142870
rect 141446 142806 141510 142870
rect 143214 142806 143278 142870
rect 144710 142806 144774 142870
rect 146478 142806 146542 142870
rect 148110 142806 148174 142870
rect 149742 142806 149806 142870
rect 151646 142806 151710 142870
rect 153142 142806 153206 142870
rect 154774 142806 154838 142870
rect 156678 142806 156742 142870
rect 158174 142806 158238 142870
rect 159942 142806 160006 142870
rect 161710 142806 161774 142870
rect 163206 142806 163270 142870
rect 164974 142806 165038 142870
rect 166606 142806 166670 142870
rect 168238 142806 168302 142870
rect 170142 142806 170206 142870
rect 171638 142806 171702 142870
rect 173406 142806 173470 142870
rect 175174 142806 175238 142870
rect 176670 142806 176734 142870
rect 178438 142806 178502 142870
rect 180206 142806 180270 142870
rect 181702 142806 181766 142870
rect 183334 142806 183398 142870
rect 185102 142806 185166 142870
rect 186734 142806 186798 142870
rect 188638 142806 188702 142870
rect 190134 142806 190198 142870
rect 191902 142806 191966 142870
rect 193670 142806 193734 142870
rect 195166 142806 195230 142870
rect 196934 142806 196998 142870
rect 198838 142806 198902 142870
rect 200198 142806 200262 142870
rect 201966 142806 202030 142870
rect 203598 142806 203662 142870
rect 205230 142806 205294 142870
rect 206862 142806 206926 142870
rect 208630 142806 208694 142870
rect 210398 142806 210462 142870
rect 212030 142806 212094 142870
rect 213662 142806 213726 142870
rect 215430 142806 215494 142870
rect 217470 142806 217534 142870
rect 217606 142806 217670 142870
rect 217742 142806 217806 142870
rect 1910 142398 1974 142462
rect 3678 142398 3742 142462
rect 5446 142398 5510 142462
rect 7214 142398 7278 142462
rect 8710 142398 8774 142462
rect 10478 142398 10542 142462
rect 12246 142398 12310 142462
rect 13742 142398 13806 142462
rect 15374 142398 15438 142462
rect 17142 142398 17206 142462
rect 18910 142398 18974 142462
rect 20406 142398 20470 142462
rect 22174 142398 22238 142462
rect 23942 142398 24006 142462
rect 25438 142398 25502 142462
rect 27206 142398 27270 142462
rect 28974 142398 29038 142462
rect 30470 142398 30534 142462
rect 32238 142398 32302 142462
rect 33870 142398 33934 142462
rect 35502 142398 35566 142462
rect 37406 142398 37470 142462
rect 38902 142398 38966 142462
rect 40670 142398 40734 142462
rect 42438 142398 42502 142462
rect 43934 142398 43998 142462
rect 45702 142398 45766 142462
rect 47470 142398 47534 142462
rect 48966 142398 49030 142462
rect 50734 142398 50798 142462
rect 52366 142398 52430 142462
rect 53998 142398 54062 142462
rect 55902 142398 55966 142462
rect 57398 142398 57462 142462
rect 59166 142398 59230 142462
rect 60934 142398 60998 142462
rect 62430 142398 62494 142462
rect 64062 142398 64126 142462
rect 65966 142398 66030 142462
rect 67462 142398 67526 142462
rect 69366 142398 69430 142462
rect 70862 142398 70926 142462
rect 72494 142398 72558 142462
rect 74262 142398 74326 142462
rect 75894 142398 75958 142462
rect 77662 142398 77726 142462
rect 79430 142398 79494 142462
rect 80926 142398 80990 142462
rect 82694 142398 82758 142462
rect 84598 142398 84662 142462
rect 85958 142398 86022 142462
rect 87726 142398 87790 142462
rect 89494 142398 89558 142462
rect 90990 142398 91054 142462
rect 92894 142398 92958 142462
rect 94390 142398 94454 142462
rect 96158 142398 96222 142462
rect 97790 142398 97854 142462
rect 99558 142398 99622 142462
rect 101190 142398 101254 142462
rect 102958 142398 103022 142462
rect 104454 142398 104518 142462
rect 106222 142398 106286 142462
rect 107854 142398 107918 142462
rect 109622 142398 109686 142462
rect 111118 142398 111182 142462
rect 112886 142398 112950 142462
rect 114654 142398 114718 142462
rect 116150 142398 116214 142462
rect 117918 142398 117982 142462
rect 119686 142398 119750 142462
rect 121318 142398 121382 142462
rect 122950 142398 123014 142462
rect 124718 142398 124782 142462
rect 126214 142398 126278 142462
rect 127982 142398 128046 142462
rect 129614 142398 129678 142462
rect 131382 142398 131446 142462
rect 133150 142398 133214 142462
rect 134646 142398 134710 142462
rect 136414 142398 136478 142462
rect 138182 142398 138246 142462
rect 139678 142398 139742 142462
rect 141446 142398 141510 142462
rect 143214 142398 143278 142462
rect 144710 142398 144774 142462
rect 146478 142398 146542 142462
rect 148110 142398 148174 142462
rect 149742 142398 149806 142462
rect 151646 142398 151710 142462
rect 153142 142398 153206 142462
rect 154774 142398 154838 142462
rect 156678 142398 156742 142462
rect 158174 142398 158238 142462
rect 159942 142398 160006 142462
rect 161710 142398 161774 142462
rect 163206 142398 163270 142462
rect 164974 142398 165038 142462
rect 166606 142398 166670 142462
rect 168238 142398 168302 142462
rect 170142 142398 170206 142462
rect 171638 142398 171702 142462
rect 173406 142398 173470 142462
rect 175174 142398 175238 142462
rect 176670 142398 176734 142462
rect 178438 142398 178502 142462
rect 180206 142398 180270 142462
rect 181702 142398 181766 142462
rect 183334 142398 183398 142462
rect 185102 142398 185166 142462
rect 186734 142398 186798 142462
rect 188638 142398 188702 142462
rect 190134 142398 190198 142462
rect 191902 142398 191966 142462
rect 193670 142398 193734 142462
rect 195166 142398 195230 142462
rect 196934 142398 196998 142462
rect 198838 142398 198902 142462
rect 200198 142398 200262 142462
rect 199246 142262 199310 142326
rect 201966 142398 202030 142462
rect 200470 142262 200534 142326
rect 203598 142398 203662 142462
rect 205230 142398 205294 142462
rect 206862 142398 206926 142462
rect 208630 142398 208694 142462
rect 210398 142398 210462 142462
rect 212030 142398 212094 142462
rect 213662 142398 213726 142462
rect 215430 142398 215494 142462
rect 199246 141990 199310 142054
rect 198294 141854 198358 141918
rect 200470 141990 200534 142054
rect 1230 141718 1294 141782
rect 217470 141718 217534 141782
rect 198566 141446 198630 141510
rect 199926 141446 199990 141510
rect 201014 141472 201078 141510
rect 201014 141446 201034 141472
rect 201034 141446 201078 141472
rect 198158 140630 198222 140694
rect 198158 140494 198222 140558
rect 217470 139950 217534 140014
rect 1230 139814 1294 139878
rect 198294 139814 198358 139878
rect 197886 139678 197950 139742
rect 198158 138454 198222 138518
rect 196662 138318 196726 138382
rect 217470 138318 217534 138382
rect 1230 138182 1294 138246
rect 197886 137094 197950 137158
rect 197886 136822 197950 136886
rect 1230 136686 1294 136750
rect 217470 136550 217534 136614
rect 196662 135598 196726 135662
rect 198022 135462 198086 135526
rect 203326 135190 203390 135254
rect 216790 135190 216854 135254
rect 1230 134918 1294 134982
rect 216790 134918 216854 134982
rect 217470 134782 217534 134846
rect 197886 134238 197950 134302
rect 196662 134102 196726 134166
rect 203462 133830 203526 133894
rect 203598 133830 203662 133894
rect 218150 133830 218214 133894
rect 1230 133150 1294 133214
rect 217470 133286 217534 133350
rect 29518 133150 29582 133214
rect 29926 133014 29990 133078
rect 34414 133150 34478 133214
rect 34822 133014 34886 133078
rect 39446 133150 39510 133214
rect 39854 133014 39918 133078
rect 44478 133150 44542 133214
rect 44886 133014 44950 133078
rect 49510 133150 49574 133214
rect 49918 133014 49982 133078
rect 54542 133150 54606 133214
rect 54814 133014 54878 133078
rect 59438 133150 59502 133214
rect 59846 133014 59910 133078
rect 64470 133150 64534 133214
rect 64742 133014 64806 133078
rect 69502 133150 69566 133214
rect 74534 133150 74598 133214
rect 69910 133014 69974 133078
rect 74806 133014 74870 133078
rect 79566 133150 79630 133214
rect 79838 133014 79902 133078
rect 84326 133150 84390 133214
rect 89358 133150 89422 133214
rect 84870 133014 84934 133078
rect 94526 133150 94590 133214
rect 89902 133014 89966 133078
rect 99422 133150 99486 133214
rect 94934 133014 94998 133078
rect 99830 133014 99894 133078
rect 104318 133150 104382 133214
rect 104726 133014 104790 133078
rect 109350 133150 109414 133214
rect 114382 133150 114446 133214
rect 109894 133014 109958 133078
rect 114790 133014 114854 133078
rect 119278 133150 119342 133214
rect 119686 133014 119750 133078
rect 124310 133150 124374 133214
rect 124718 133014 124782 133078
rect 129342 133150 129406 133214
rect 129750 133014 129814 133078
rect 134374 133150 134438 133214
rect 134782 133014 134846 133078
rect 139406 133150 139470 133214
rect 139678 133014 139742 133078
rect 144302 133150 144366 133214
rect 144710 133014 144774 133078
rect 149334 133150 149398 133214
rect 149742 133014 149806 133078
rect 154366 133150 154430 133214
rect 159398 133150 159462 133214
rect 154774 133014 154838 133078
rect 164430 133150 164494 133214
rect 159806 133014 159870 133078
rect 164702 133014 164766 133078
rect 169190 133150 169254 133214
rect 174222 133150 174286 133214
rect 169734 133014 169798 133078
rect 179390 133150 179454 133214
rect 174766 133014 174830 133078
rect 184286 133150 184350 133214
rect 179798 133014 179862 133078
rect 184558 133014 184622 133078
rect 29790 132606 29854 132670
rect 34686 132606 34750 132670
rect 39718 132606 39782 132670
rect 44750 132606 44814 132670
rect 49646 132606 49710 132670
rect 54678 132606 54742 132670
rect 59710 132606 59774 132670
rect 64878 132606 64942 132670
rect 69774 132606 69838 132670
rect 74670 132606 74734 132670
rect 79702 132606 79766 132670
rect 84734 132606 84798 132670
rect 89766 132606 89830 132670
rect 94798 132606 94862 132670
rect 99694 132606 99758 132670
rect 104590 132606 104654 132670
rect 109758 132606 109822 132670
rect 114790 132606 114854 132670
rect 119550 132606 119614 132670
rect 124582 132606 124646 132670
rect 129614 132606 129678 132670
rect 134646 132606 134710 132670
rect 139542 132606 139606 132670
rect 144574 132606 144638 132670
rect 149606 132606 149670 132670
rect 154638 132606 154702 132670
rect 159670 132606 159734 132670
rect 164566 132606 164630 132670
rect 169598 132606 169662 132670
rect 174630 132606 174694 132670
rect 198022 132742 198086 132806
rect 203462 132742 203526 132806
rect 179662 132606 179726 132670
rect 184422 132606 184486 132670
rect 196526 132606 196590 132670
rect 203326 132606 203390 132670
rect 203326 132470 203390 132534
rect 203462 132470 203526 132534
rect 29790 131926 29854 131990
rect 29654 131790 29718 131854
rect 34686 131926 34750 131990
rect 39718 131926 39782 131990
rect 35774 131790 35838 131854
rect 44750 131926 44814 131990
rect 39718 131790 39782 131854
rect 44342 131790 44406 131854
rect 49646 131926 49710 131990
rect 54678 131926 54742 131990
rect 50734 131790 50798 131854
rect 54678 131790 54742 131854
rect 59710 131926 59774 131990
rect 64878 131926 64942 131990
rect 60798 131790 60862 131854
rect 69774 131926 69838 131990
rect 64606 131790 64670 131854
rect 69230 131790 69294 131854
rect 74670 131926 74734 131990
rect 79702 131926 79766 131990
rect 84734 131926 84798 131990
rect 74670 131790 74734 131854
rect 79294 131790 79358 131854
rect 84190 131790 84254 131854
rect 89766 131926 89830 131990
rect 89630 131790 89694 131854
rect 94798 131926 94862 131990
rect 94662 131790 94726 131854
rect 99694 131926 99758 131990
rect 104590 131926 104654 131990
rect 99558 131790 99622 131854
rect 104318 131790 104382 131854
rect 109758 131926 109822 131990
rect 114790 131926 114854 131990
rect 109622 131790 109686 131854
rect 114246 131790 114310 131854
rect 119550 131926 119614 131990
rect 124582 131926 124646 131990
rect 120230 131790 120294 131854
rect 129614 131926 129678 131990
rect 124582 131790 124646 131854
rect 129206 131790 129270 131854
rect 134646 131926 134710 131990
rect 139542 131926 139606 131990
rect 135598 131790 135662 131854
rect 139542 131790 139606 131854
rect 144574 131926 144638 131990
rect 149606 131926 149670 131990
rect 145254 131790 145318 131854
rect 154638 131926 154702 131990
rect 149470 131790 149534 131854
rect 154094 131790 154158 131854
rect 159670 131926 159734 131990
rect 164566 131926 164630 131990
rect 169598 131926 169662 131990
rect 174630 131926 174694 131990
rect 160214 131790 160278 131854
rect 165518 131790 165582 131854
rect 170142 131790 170206 131854
rect 174494 131790 174558 131854
rect 179662 131926 179726 131990
rect 179526 131790 179590 131854
rect 184422 131926 184486 131990
rect 184422 131790 184486 131854
rect 1230 131518 1294 131582
rect 217470 131518 217534 131582
rect 196662 131382 196726 131446
rect 203462 131382 203526 131446
rect 29926 131246 29990 131310
rect 29926 131110 29990 131174
rect 34822 131246 34886 131310
rect 34958 131110 35022 131174
rect 39854 131246 39918 131310
rect 39990 131110 40054 131174
rect 44886 131246 44950 131310
rect 44886 131110 44950 131174
rect 49918 131246 49982 131310
rect 49918 131110 49982 131174
rect 54814 131246 54878 131310
rect 54814 131110 54878 131174
rect 59846 131246 59910 131310
rect 64742 131246 64806 131310
rect 59982 131110 60046 131174
rect 64878 131110 64942 131174
rect 69910 131246 69974 131310
rect 69910 131110 69974 131174
rect 74806 131246 74870 131310
rect 74942 131110 75006 131174
rect 79838 131246 79902 131310
rect 79838 131110 79902 131174
rect 84870 131246 84934 131310
rect 84870 131110 84934 131174
rect 89902 131246 89966 131310
rect 89902 131110 89966 131174
rect 94934 131246 94998 131310
rect 99830 131246 99894 131310
rect 94934 131110 94998 131174
rect 99830 131110 99894 131174
rect 104726 131246 104790 131310
rect 104862 131110 104926 131174
rect 109894 131246 109958 131310
rect 109894 131110 109958 131174
rect 114654 131246 114718 131310
rect 114654 131110 114718 131174
rect 119686 131246 119750 131310
rect 119822 131110 119886 131174
rect 124718 131246 124782 131310
rect 124854 131110 124918 131174
rect 129750 131246 129814 131310
rect 129750 131110 129814 131174
rect 134782 131246 134846 131310
rect 134782 131110 134846 131174
rect 139678 131246 139742 131310
rect 139814 131110 139878 131174
rect 144710 131246 144774 131310
rect 149742 131246 149806 131310
rect 144846 131110 144910 131174
rect 149606 131110 149670 131174
rect 154774 131246 154838 131310
rect 154774 131110 154838 131174
rect 159806 131246 159870 131310
rect 159806 131110 159870 131174
rect 164702 131246 164766 131310
rect 164702 131110 164766 131174
rect 169734 131246 169798 131310
rect 169734 131110 169798 131174
rect 174766 131246 174830 131310
rect 174630 131110 174694 131174
rect 179798 131246 179862 131310
rect 184558 131246 184622 131310
rect 179798 131110 179862 131174
rect 197886 131246 197950 131310
rect 184694 131110 184758 131174
rect 203598 131110 203662 131174
rect 203598 130974 203662 131038
rect 196526 130022 196590 130086
rect 1230 129750 1294 129814
rect 196526 129750 196590 129814
rect 217470 129886 217534 129950
rect 203326 129750 203390 129814
rect 203462 129614 203526 129678
rect 218150 129614 218214 129678
rect 29926 128662 29990 128726
rect 28838 128526 28902 128590
rect 34958 128662 35022 128726
rect 39990 128662 40054 128726
rect 44886 128662 44950 128726
rect 49918 128662 49982 128726
rect 54814 128662 54878 128726
rect 59982 128662 60046 128726
rect 64878 128662 64942 128726
rect 69910 128662 69974 128726
rect 74942 128662 75006 128726
rect 79838 128662 79902 128726
rect 84870 128662 84934 128726
rect 89902 128662 89966 128726
rect 94934 128662 94998 128726
rect 99830 128662 99894 128726
rect 104862 128662 104926 128726
rect 109894 128662 109958 128726
rect 114654 128662 114718 128726
rect 119822 128662 119886 128726
rect 124854 128662 124918 128726
rect 129750 128662 129814 128726
rect 134782 128662 134846 128726
rect 139814 128662 139878 128726
rect 144846 128662 144910 128726
rect 149606 128662 149670 128726
rect 154774 128662 154838 128726
rect 159806 128662 159870 128726
rect 164702 128662 164766 128726
rect 169734 128662 169798 128726
rect 174630 128662 174694 128726
rect 179798 128662 179862 128726
rect 184694 128662 184758 128726
rect 190406 128526 190470 128590
rect 197886 128526 197950 128590
rect 196662 128390 196726 128454
rect 203598 128390 203662 128454
rect 1230 128118 1294 128182
rect 217470 128254 217534 128318
rect 216493 127845 216557 127909
rect 29654 127166 29718 127230
rect 29654 127030 29718 127094
rect 30878 127030 30942 127094
rect 31694 127030 31758 127094
rect 32918 127030 32982 127094
rect 33462 127030 33526 127094
rect 34142 127030 34206 127094
rect 34686 127030 34750 127094
rect 35774 127166 35838 127230
rect 35910 127030 35974 127094
rect 36590 127030 36654 127094
rect 37134 127030 37198 127094
rect 38086 127030 38150 127094
rect 39718 127166 39782 127230
rect 39446 127030 39510 127094
rect 40398 127030 40462 127094
rect 41622 127030 41686 127094
rect 42166 127030 42230 127094
rect 42982 127030 43046 127094
rect 43254 127030 43318 127094
rect 44342 127166 44406 127230
rect 44614 127030 44678 127094
rect 45430 127030 45494 127094
rect 45974 127030 46038 127094
rect 46654 127030 46718 127094
rect 46790 127030 46854 127094
rect 48422 127030 48486 127094
rect 49102 127030 49166 127094
rect 50734 127166 50798 127230
rect 50326 127030 50390 127094
rect 50870 127030 50934 127094
rect 52230 127030 52294 127094
rect 52774 127030 52838 127094
rect 53318 127030 53382 127094
rect 54678 127166 54742 127230
rect 54134 127030 54198 127094
rect 54678 127030 54742 127094
rect 55358 127030 55422 127094
rect 55902 127030 55966 127094
rect 57126 127030 57190 127094
rect 57806 127030 57870 127094
rect 59574 127030 59638 127094
rect 60798 127166 60862 127230
rect 60934 127030 60998 127094
rect 61478 127030 61542 127094
rect 61614 127030 61678 127094
rect 62158 127030 62222 127094
rect 62838 127030 62902 127094
rect 63382 127030 63446 127094
rect 64606 127166 64670 127230
rect 64062 127030 64126 127094
rect 65694 127030 65758 127094
rect 66646 127030 66710 127094
rect 67190 127030 67254 127094
rect 67326 127030 67390 127094
rect 68414 127030 68478 127094
rect 69230 127166 69294 127230
rect 69094 127030 69158 127094
rect 69638 127030 69702 127094
rect 70318 127030 70382 127094
rect 70862 127030 70926 127094
rect 71950 127030 72014 127094
rect 72902 127030 72966 127094
rect 74670 127166 74734 127230
rect 74126 127030 74190 127094
rect 75214 127030 75278 127094
rect 75350 127030 75414 127094
rect 75894 127030 75958 127094
rect 76574 127030 76638 127094
rect 77118 127030 77182 127094
rect 77798 127030 77862 127094
rect 78342 127030 78406 127094
rect 79294 127166 79358 127230
rect 79566 127030 79630 127094
rect 80926 127030 80990 127094
rect 81470 127030 81534 127094
rect 81606 127030 81670 127094
rect 82014 127030 82078 127094
rect 82830 127030 82894 127094
rect 84190 127166 84254 127230
rect 84054 127030 84118 127094
rect 84598 127030 84662 127094
rect 85278 127030 85342 127094
rect 85822 127030 85886 127094
rect 86502 127030 86566 127094
rect 87046 127030 87110 127094
rect 88406 127030 88470 127094
rect 89630 127166 89694 127230
rect 89222 127030 89286 127094
rect 90310 127030 90374 127094
rect 90854 127030 90918 127094
rect 91534 127030 91598 127094
rect 92758 127030 92822 127094
rect 93302 127030 93366 127094
rect 94662 127166 94726 127230
rect 94662 127030 94726 127094
rect 95342 127030 95406 127094
rect 95750 127030 95814 127094
rect 96566 127030 96630 127094
rect 97110 127030 97174 127094
rect 97926 127030 97990 127094
rect 99558 127166 99622 127230
rect 99558 127030 99622 127094
rect 100238 127030 100302 127094
rect 100510 127030 100574 127094
rect 102006 127030 102070 127094
rect 103366 127030 103430 127094
rect 104318 127166 104382 127230
rect 104046 127030 104110 127094
rect 104590 127030 104654 127094
rect 105270 127030 105334 127094
rect 105814 127030 105878 127094
rect 106494 127030 106558 127094
rect 108126 127030 108190 127094
rect 109622 127166 109686 127230
rect 109214 127030 109278 127094
rect 110302 127030 110366 127094
rect 110846 127030 110910 127094
rect 111526 127030 111590 127094
rect 112070 127030 112134 127094
rect 112750 127030 112814 127094
rect 113294 127030 113358 127094
rect 114246 127166 114310 127230
rect 114518 127030 114582 127094
rect 115742 127030 115806 127094
rect 116558 127030 116622 127094
rect 117646 127030 117710 127094
rect 117782 127030 117846 127094
rect 118326 127030 118390 127094
rect 119006 127030 119070 127094
rect 119550 127030 119614 127094
rect 120230 127166 120294 127230
rect 120774 127030 120838 127094
rect 121454 127030 121518 127094
rect 121998 127030 122062 127094
rect 124582 127166 124646 127230
rect 122950 127030 123014 127094
rect 123902 127030 123966 127094
rect 124310 127030 124374 127094
rect 125262 127030 125326 127094
rect 125806 127030 125870 127094
rect 126486 127030 126550 127094
rect 127030 127030 127094 127094
rect 128254 127030 128318 127094
rect 129206 127166 129270 127230
rect 128934 127030 128998 127094
rect 129478 127030 129542 127094
rect 130294 127030 130358 127094
rect 130838 127030 130902 127094
rect 132062 127030 132126 127094
rect 133286 127030 133350 127094
rect 133966 127030 134030 127094
rect 134510 127030 134574 127094
rect 135598 127166 135662 127230
rect 135190 127030 135254 127094
rect 135462 127030 135526 127094
rect 137094 127030 137158 127094
rect 138182 127030 138246 127094
rect 139542 127166 139606 127230
rect 139542 127030 139606 127094
rect 140358 127030 140422 127094
rect 141446 127030 141510 127094
rect 141990 127030 142054 127094
rect 142670 127030 142734 127094
rect 144438 127030 144502 127094
rect 145254 127166 145318 127230
rect 145254 127030 145318 127094
rect 146478 127030 146542 127094
rect 147022 127030 147086 127094
rect 147702 127030 147766 127094
rect 148246 127030 148310 127094
rect 149470 127166 149534 127230
rect 150150 127030 150214 127094
rect 151510 127030 151574 127094
rect 151918 127030 151982 127094
rect 153278 127030 153342 127094
rect 154094 127166 154158 127230
rect 153958 127030 154022 127094
rect 154502 127030 154566 127094
rect 155182 127030 155246 127094
rect 155726 127030 155790 127094
rect 156678 127030 156742 127094
rect 157902 127030 157966 127094
rect 158990 127030 159054 127094
rect 160214 127166 160278 127230
rect 160214 127030 160278 127094
rect 160758 127030 160822 127094
rect 161982 127030 162046 127094
rect 163206 127030 163270 127094
rect 163886 127030 163950 127094
rect 164430 127030 164494 127094
rect 165518 127166 165582 127230
rect 165382 127030 165446 127094
rect 166334 127030 166398 127094
rect 166470 127030 166534 127094
rect 168238 127030 168302 127094
rect 168918 127030 168982 127094
rect 169462 127030 169526 127094
rect 170142 127166 170206 127230
rect 170686 127030 170750 127094
rect 171366 127030 171430 127094
rect 171910 127030 171974 127094
rect 173134 127030 173198 127094
rect 174494 127166 174558 127230
rect 174494 127030 174558 127094
rect 175174 127030 175238 127094
rect 175718 127030 175782 127094
rect 176942 127030 177006 127094
rect 178166 127030 178230 127094
rect 179526 127166 179590 127230
rect 178982 127030 179046 127094
rect 180206 127030 180270 127094
rect 180614 127030 180678 127094
rect 181430 127030 181494 127094
rect 181974 127030 182038 127094
rect 183198 127030 183262 127094
rect 184014 127030 184078 127094
rect 184422 127166 184486 127230
rect 184286 127030 184350 127094
rect 184966 127030 185030 127094
rect 185238 127030 185302 127094
rect 185374 127030 185438 127094
rect 187006 127030 187070 127094
rect 188230 127030 188294 127094
rect 188910 127030 188974 127094
rect 189454 127030 189518 127094
rect 149470 126894 149534 126958
rect 203462 126894 203526 126958
rect 218150 126894 218214 126958
rect 1230 126486 1294 126550
rect 29654 126622 29718 126686
rect 30878 126622 30942 126686
rect 31694 126622 31758 126686
rect 28838 126350 28902 126414
rect 32918 126622 32982 126686
rect 33462 126622 33526 126686
rect 34142 126622 34206 126686
rect 34686 126622 34750 126686
rect 35910 126622 35974 126686
rect 36590 126622 36654 126686
rect 37134 126622 37198 126686
rect 38086 126622 38150 126686
rect 39446 126622 39510 126686
rect 40398 126622 40462 126686
rect 41622 126622 41686 126686
rect 42166 126622 42230 126686
rect 42982 126622 43046 126686
rect 43254 126622 43318 126686
rect 44614 126622 44678 126686
rect 45430 126622 45494 126686
rect 45974 126622 46038 126686
rect 46654 126622 46718 126686
rect 46790 126622 46854 126686
rect 48422 126622 48486 126686
rect 49102 126622 49166 126686
rect 50326 126622 50390 126686
rect 50870 126622 50934 126686
rect 52230 126622 52294 126686
rect 52774 126622 52838 126686
rect 53318 126622 53382 126686
rect 54134 126622 54198 126686
rect 54678 126622 54742 126686
rect 55358 126622 55422 126686
rect 55902 126622 55966 126686
rect 57126 126622 57190 126686
rect 57806 126622 57870 126686
rect 59574 126622 59638 126686
rect 60934 126622 60998 126686
rect 61478 126622 61542 126686
rect 61614 126622 61678 126686
rect 62158 126622 62222 126686
rect 62838 126622 62902 126686
rect 63382 126622 63446 126686
rect 64062 126622 64126 126686
rect 65694 126622 65758 126686
rect 66646 126622 66710 126686
rect 67190 126622 67254 126686
rect 67326 126622 67390 126686
rect 68414 126622 68478 126686
rect 69094 126622 69158 126686
rect 69638 126622 69702 126686
rect 70318 126622 70382 126686
rect 70862 126622 70926 126686
rect 71950 126622 72014 126686
rect 72902 126622 72966 126686
rect 74126 126622 74190 126686
rect 75214 126622 75278 126686
rect 75350 126622 75414 126686
rect 75894 126622 75958 126686
rect 76574 126622 76638 126686
rect 77118 126622 77182 126686
rect 77798 126622 77862 126686
rect 78342 126622 78406 126686
rect 79566 126622 79630 126686
rect 80926 126622 80990 126686
rect 81470 126622 81534 126686
rect 81606 126622 81670 126686
rect 82014 126622 82078 126686
rect 82830 126622 82894 126686
rect 84054 126622 84118 126686
rect 84598 126622 84662 126686
rect 85278 126622 85342 126686
rect 85822 126622 85886 126686
rect 86502 126622 86566 126686
rect 87046 126622 87110 126686
rect 88406 126622 88470 126686
rect 90310 126622 90374 126686
rect 89222 126486 89286 126550
rect 90854 126622 90918 126686
rect 91534 126622 91598 126686
rect 92758 126622 92822 126686
rect 93302 126622 93366 126686
rect 94662 126622 94726 126686
rect 95342 126622 95406 126686
rect 95750 126622 95814 126686
rect 96566 126622 96630 126686
rect 97110 126622 97174 126686
rect 97926 126486 97990 126550
rect 99558 126622 99622 126686
rect 100238 126622 100302 126686
rect 100510 126622 100574 126686
rect 102006 126622 102070 126686
rect 103366 126622 103430 126686
rect 104046 126622 104110 126686
rect 104590 126622 104654 126686
rect 105270 126622 105334 126686
rect 105814 126622 105878 126686
rect 106494 126622 106558 126686
rect 108126 126622 108190 126686
rect 109214 126622 109278 126686
rect 110302 126622 110366 126686
rect 110846 126622 110910 126686
rect 111526 126622 111590 126686
rect 112070 126622 112134 126686
rect 112750 126622 112814 126686
rect 113294 126622 113358 126686
rect 114518 126622 114582 126686
rect 115742 126622 115806 126686
rect 116558 126622 116622 126686
rect 117646 126622 117710 126686
rect 117782 126622 117846 126686
rect 118326 126622 118390 126686
rect 119006 126622 119070 126686
rect 119550 126622 119614 126686
rect 120774 126622 120838 126686
rect 121454 126622 121518 126686
rect 121998 126622 122062 126686
rect 122950 126622 123014 126686
rect 123902 126622 123966 126686
rect 124446 126622 124510 126686
rect 125262 126622 125326 126686
rect 125806 126622 125870 126686
rect 126486 126622 126550 126686
rect 127030 126622 127094 126686
rect 128254 126622 128318 126686
rect 128934 126622 128998 126686
rect 129478 126622 129542 126686
rect 130294 126622 130358 126686
rect 130838 126622 130902 126686
rect 132062 126622 132126 126686
rect 133286 126622 133350 126686
rect 133966 126622 134030 126686
rect 134510 126622 134574 126686
rect 135190 126622 135254 126686
rect 135462 126622 135526 126686
rect 137094 126622 137158 126686
rect 138182 126622 138246 126686
rect 139542 126622 139606 126686
rect 140358 126622 140422 126686
rect 141446 126622 141510 126686
rect 141990 126622 142054 126686
rect 142670 126622 142734 126686
rect 144438 126622 144502 126686
rect 145254 126622 145318 126686
rect 146478 126622 146542 126686
rect 147022 126622 147086 126686
rect 147702 126622 147766 126686
rect 148246 126622 148310 126686
rect 149470 126622 149534 126686
rect 150150 126622 150214 126686
rect 151510 126622 151574 126686
rect 151918 126622 151982 126686
rect 153278 126622 153342 126686
rect 153958 126622 154022 126686
rect 154502 126622 154566 126686
rect 155182 126622 155246 126686
rect 155726 126622 155790 126686
rect 156678 126622 156742 126686
rect 157902 126486 157966 126550
rect 158990 126622 159054 126686
rect 160214 126622 160278 126686
rect 160758 126622 160822 126686
rect 161982 126622 162046 126686
rect 163206 126622 163270 126686
rect 163886 126622 163950 126686
rect 164430 126622 164494 126686
rect 165382 126622 165446 126686
rect 166334 126622 166398 126686
rect 166470 126622 166534 126686
rect 168238 126622 168302 126686
rect 168918 126622 168982 126686
rect 169462 126622 169526 126686
rect 170686 126622 170750 126686
rect 171366 126622 171430 126686
rect 171910 126622 171974 126686
rect 173134 126622 173198 126686
rect 174494 126622 174558 126686
rect 175174 126622 175238 126686
rect 175718 126622 175782 126686
rect 176942 126622 177006 126686
rect 178166 126622 178230 126686
rect 178982 126622 179046 126686
rect 180206 126622 180270 126686
rect 180614 126622 180678 126686
rect 181430 126622 181494 126686
rect 181974 126622 182038 126686
rect 183198 126622 183262 126686
rect 184014 126622 184078 126686
rect 184286 126622 184350 126686
rect 184966 126622 185030 126686
rect 185238 126622 185302 126686
rect 185374 126622 185438 126686
rect 187006 126622 187070 126686
rect 188230 126622 188294 126686
rect 188910 126622 188974 126686
rect 189454 126622 189518 126686
rect 191494 126486 191558 126550
rect 190406 126350 190470 126414
rect 28294 126214 28358 126278
rect 217470 126350 217534 126414
rect 190406 126214 190470 126278
rect 191494 126214 191558 126278
rect 196526 126214 196590 126278
rect 194894 126078 194958 126142
rect 195166 126078 195230 126142
rect 28294 125942 28358 126006
rect 28294 125806 28358 125870
rect 21902 125534 21966 125598
rect 22310 125534 22374 125598
rect 22446 125534 22510 125598
rect 28566 125670 28630 125734
rect 190406 125942 190470 126006
rect 190134 125670 190198 125734
rect 194894 125670 194958 125734
rect 195166 125670 195230 125734
rect 28294 125398 28358 125462
rect 28566 125398 28630 125462
rect 21902 125262 21966 125326
rect 21766 125126 21830 125190
rect 22310 125262 22374 125326
rect 22446 125262 22510 125326
rect 1230 124854 1294 124918
rect 21766 124854 21830 124918
rect 21766 124718 21830 124782
rect 22718 124718 22782 124782
rect 22990 124718 23054 124782
rect 23398 124718 23462 124782
rect 28430 125262 28494 125326
rect 28430 124990 28494 125054
rect 190134 125262 190198 125326
rect 190270 125262 190334 125326
rect 190270 124990 190334 125054
rect 21766 124446 21830 124510
rect 21902 124310 21966 124374
rect 22718 124446 22782 124510
rect 22446 124310 22510 124374
rect 22990 124446 23054 124510
rect 23126 124310 23190 124374
rect 23398 124446 23462 124510
rect 23398 124310 23462 124374
rect 196662 125670 196726 125734
rect 196798 125534 196862 125598
rect 216790 125398 216854 125462
rect 196798 125262 196862 125326
rect 196662 125126 196726 125190
rect 195166 124718 195230 124782
rect 195438 124718 195502 124782
rect 195982 124718 196046 124782
rect 196118 124718 196182 124782
rect 196662 124854 196726 124918
rect 196662 124718 196726 124782
rect 216790 124854 216854 124918
rect 217470 124718 217534 124782
rect 195166 124446 195230 124510
rect 195030 124310 195094 124374
rect 195438 124446 195502 124510
rect 195574 124310 195638 124374
rect 195982 124446 196046 124510
rect 196118 124446 196182 124510
rect 195982 124310 196046 124374
rect 196118 124310 196182 124374
rect 196662 124446 196726 124510
rect 196798 124310 196862 124374
rect 21902 124038 21966 124102
rect 21766 123902 21830 123966
rect 22446 124038 22510 124102
rect 22174 123902 22238 123966
rect 22582 123902 22646 123966
rect 23126 124038 23190 124102
rect 22990 123902 23054 123966
rect 23398 124038 23462 124102
rect 23534 123902 23598 123966
rect 195030 124038 195094 124102
rect 195166 123902 195230 123966
rect 195574 124038 195638 124102
rect 195438 123902 195502 123966
rect 195982 124038 196046 124102
rect 196118 124038 196182 124102
rect 196254 123902 196318 123966
rect 196798 124038 196862 124102
rect 196662 123902 196726 123966
rect 218150 123902 218214 123966
rect 21766 123630 21830 123694
rect 21766 123494 21830 123558
rect 22174 123630 22238 123694
rect 22582 123630 22646 123694
rect 22446 123494 22510 123558
rect 22582 123494 22646 123558
rect 22990 123630 23054 123694
rect 23126 123494 23190 123558
rect 23534 123630 23598 123694
rect 23534 123494 23598 123558
rect 195166 123630 195230 123694
rect 195166 123494 195230 123558
rect 195438 123630 195502 123694
rect 195574 123494 195638 123558
rect 196254 123630 196318 123694
rect 195982 123494 196046 123558
rect 196118 123494 196182 123558
rect 196662 123630 196726 123694
rect 196798 123494 196862 123558
rect 1230 123222 1294 123286
rect 21766 123222 21830 123286
rect 22446 123222 22510 123286
rect 22582 123222 22646 123286
rect 22310 123086 22374 123150
rect 22446 123086 22510 123150
rect 23126 123222 23190 123286
rect 22990 123086 23054 123150
rect 23534 123222 23598 123286
rect 23398 123086 23462 123150
rect 195166 123222 195230 123286
rect 195166 123086 195230 123150
rect 195574 123222 195638 123286
rect 195438 123086 195502 123150
rect 195982 123222 196046 123286
rect 196118 123222 196182 123286
rect 196254 123086 196318 123150
rect 196798 123222 196862 123286
rect 216790 123086 216854 123150
rect 217470 123086 217534 123150
rect 21766 122678 21830 122742
rect 22310 122814 22374 122878
rect 22446 122814 22510 122878
rect 22310 122678 22374 122742
rect 22582 122678 22646 122742
rect 22990 122814 23054 122878
rect 22990 122678 23054 122742
rect 23398 122814 23462 122878
rect 23534 122678 23598 122742
rect 21766 122406 21830 122470
rect 22310 122406 22374 122470
rect 22582 122406 22646 122470
rect 22718 122270 22782 122334
rect 22990 122406 23054 122470
rect 23126 122270 23190 122334
rect 23534 122406 23598 122470
rect 23398 122270 23462 122334
rect 195166 122814 195230 122878
rect 195166 122678 195230 122742
rect 195438 122814 195502 122878
rect 195574 122678 195638 122742
rect 196254 122814 196318 122878
rect 195846 122678 195910 122742
rect 196662 122678 196726 122742
rect 216790 122678 216854 122742
rect 195166 122406 195230 122470
rect 195030 122270 195094 122334
rect 195574 122406 195638 122470
rect 195438 122270 195502 122334
rect 195846 122406 195910 122470
rect 196118 122270 196182 122334
rect 196662 122406 196726 122470
rect 21766 121998 21830 122062
rect 22446 121998 22510 122062
rect 22718 121998 22782 122062
rect 23126 121998 23190 122062
rect 21766 121726 21830 121790
rect 21766 121590 21830 121654
rect 22446 121726 22510 121790
rect 22174 121590 22238 121654
rect 23398 121998 23462 122062
rect 28294 121726 28358 121790
rect 195030 121998 195094 122062
rect 190134 121726 190198 121790
rect 1230 121318 1294 121382
rect 21766 121318 21830 121382
rect 21902 121182 21966 121246
rect 22174 121318 22238 121382
rect 21902 120910 21966 120974
rect 21766 120774 21830 120838
rect 22446 120774 22510 120838
rect 23126 120774 23190 120838
rect 28294 121454 28358 121518
rect 28294 121318 28358 121382
rect 28294 121046 28358 121110
rect 28430 120910 28494 120974
rect 190134 121454 190198 121518
rect 190270 121318 190334 121382
rect 190270 121046 190334 121110
rect 190270 120910 190334 120974
rect 195438 121998 195502 122062
rect 196118 121998 196182 122062
rect 196798 121998 196862 122062
rect 196118 121590 196182 121654
rect 196798 121726 196862 121790
rect 196662 121590 196726 121654
rect 217470 121454 217534 121518
rect 23398 120774 23462 120838
rect 21766 120502 21830 120566
rect 21766 120366 21830 120430
rect 22446 120502 22510 120566
rect 22174 120366 22238 120430
rect 22718 120366 22782 120430
rect 23126 120502 23190 120566
rect 23126 120366 23190 120430
rect 23398 120502 23462 120566
rect 23398 120366 23462 120430
rect 28294 120502 28358 120566
rect 28430 120502 28494 120566
rect 28294 120230 28358 120294
rect 21766 120094 21830 120158
rect 21902 119958 21966 120022
rect 22174 120094 22238 120158
rect 22718 120094 22782 120158
rect 22310 119958 22374 120022
rect 23126 120094 23190 120158
rect 23126 119958 23190 120022
rect 23398 120094 23462 120158
rect 195166 120774 195230 120838
rect 195438 120774 195502 120838
rect 196118 121318 196182 121382
rect 196662 121318 196726 121382
rect 196798 121182 196862 121246
rect 218150 121046 218214 121110
rect 195846 120774 195910 120838
rect 196798 120910 196862 120974
rect 196662 120774 196726 120838
rect 190134 120502 190198 120566
rect 190270 120502 190334 120566
rect 195166 120502 195230 120566
rect 195166 120366 195230 120430
rect 195438 120502 195502 120566
rect 195574 120366 195638 120430
rect 195846 120502 195910 120566
rect 195982 120366 196046 120430
rect 196662 120502 196726 120566
rect 196798 120366 196862 120430
rect 190134 120230 190198 120294
rect 23398 119958 23462 120022
rect 195166 120094 195230 120158
rect 195030 119958 195094 120022
rect 195574 120094 195638 120158
rect 195574 119958 195638 120022
rect 195982 120094 196046 120158
rect 195982 119958 196046 120022
rect 196798 120094 196862 120158
rect 196798 119958 196862 120022
rect 217470 119822 217534 119886
rect 1230 119686 1294 119750
rect 21902 119686 21966 119750
rect 21766 119550 21830 119614
rect 22310 119686 22374 119750
rect 22446 119550 22510 119614
rect 23126 119686 23190 119750
rect 23126 119550 23190 119614
rect 23398 119686 23462 119750
rect 23534 119550 23598 119614
rect 195030 119686 195094 119750
rect 195166 119550 195230 119614
rect 195574 119686 195638 119750
rect 195438 119550 195502 119614
rect 195982 119686 196046 119750
rect 195846 119550 195910 119614
rect 196254 119550 196318 119614
rect 196798 119686 196862 119750
rect 196662 119550 196726 119614
rect 21766 119278 21830 119342
rect 22446 119278 22510 119342
rect 22310 119142 22374 119206
rect 23126 119278 23190 119342
rect 23126 119142 23190 119206
rect 23534 119278 23598 119342
rect 195166 119278 195230 119342
rect 23534 119142 23598 119206
rect 195030 119142 195094 119206
rect 195438 119278 195502 119342
rect 195438 119142 195502 119206
rect 195846 119278 195910 119342
rect 196254 119278 196318 119342
rect 195846 119142 195910 119206
rect 196118 119142 196182 119206
rect 196662 119278 196726 119342
rect 21902 118734 21966 118798
rect 22310 118870 22374 118934
rect 22718 118734 22782 118798
rect 23126 118870 23190 118934
rect 22990 118734 23054 118798
rect 23534 118870 23598 118934
rect 23398 118734 23462 118798
rect 195030 118870 195094 118934
rect 195030 118734 195094 118798
rect 195438 118870 195502 118934
rect 195438 118734 195502 118798
rect 195846 118870 195910 118934
rect 196118 118870 196182 118934
rect 195846 118734 195910 118798
rect 196798 118734 196862 118798
rect 21902 118462 21966 118526
rect 22174 118326 22238 118390
rect 22718 118462 22782 118526
rect 22582 118326 22646 118390
rect 22990 118462 23054 118526
rect 23126 118326 23190 118390
rect 23398 118462 23462 118526
rect 23534 118326 23598 118390
rect 195030 118462 195094 118526
rect 1230 118054 1294 118118
rect 195166 118326 195230 118390
rect 195438 118462 195502 118526
rect 195438 118326 195502 118390
rect 195846 118462 195910 118526
rect 195846 118326 195910 118390
rect 196118 118326 196182 118390
rect 196798 118462 196862 118526
rect 218150 118462 218214 118526
rect 21766 118054 21830 118118
rect 22174 118054 22238 118118
rect 22582 118054 22646 118118
rect 22446 117918 22510 117982
rect 23126 118054 23190 118118
rect 23126 117918 23190 117982
rect 23534 118054 23598 118118
rect 23398 117918 23462 117982
rect 21766 117782 21830 117846
rect 22446 117646 22510 117710
rect 22582 117510 22646 117574
rect 23126 117646 23190 117710
rect 23398 117646 23462 117710
rect 28294 117646 28358 117710
rect 195166 118054 195230 118118
rect 195030 117918 195094 117982
rect 195438 118054 195502 118118
rect 195438 117918 195502 117982
rect 195846 118054 195910 118118
rect 196118 118054 196182 118118
rect 196662 118054 196726 118118
rect 217470 118190 217534 118254
rect 195030 117646 195094 117710
rect 21766 117238 21830 117302
rect 22582 117238 22646 117302
rect 21766 116966 21830 117030
rect 21902 116830 21966 116894
rect 22310 116830 22374 116894
rect 22446 116830 22510 116894
rect 28294 117374 28358 117438
rect 28430 117374 28494 117438
rect 28430 117102 28494 117166
rect 28566 116966 28630 117030
rect 190134 117374 190198 117438
rect 190134 117102 190198 117166
rect 190270 116966 190334 117030
rect 195438 117646 195502 117710
rect 195846 117510 195910 117574
rect 196662 117782 196726 117846
rect 216493 117670 216557 117674
rect 216493 117614 216497 117670
rect 216497 117614 216553 117670
rect 216553 117614 216557 117670
rect 216493 117610 216557 117614
rect 21902 116558 21966 116622
rect 1230 116422 1294 116486
rect 21902 116422 21966 116486
rect 22310 116558 22374 116622
rect 22446 116558 22510 116622
rect 23126 116422 23190 116486
rect 23534 116422 23598 116486
rect 28566 116694 28630 116758
rect 28430 116558 28494 116622
rect 190270 116694 190334 116758
rect 190270 116558 190334 116622
rect 195846 117238 195910 117302
rect 196662 117238 196726 117302
rect 195846 116830 195910 116894
rect 196118 116830 196182 116894
rect 196662 116966 196726 117030
rect 196798 116830 196862 116894
rect 216790 116830 216854 116894
rect 195166 116422 195230 116486
rect 195438 116422 195502 116486
rect 195846 116558 195910 116622
rect 196118 116558 196182 116622
rect 196798 116558 196862 116622
rect 196798 116422 196862 116486
rect 216790 116422 216854 116486
rect 28430 116286 28494 116350
rect 21902 116150 21966 116214
rect 21902 116014 21966 116078
rect 22174 116014 22238 116078
rect 22582 116014 22646 116078
rect 23126 116150 23190 116214
rect 22990 116014 23054 116078
rect 23534 116150 23598 116214
rect 23398 116014 23462 116078
rect 190270 116286 190334 116350
rect 217470 116286 217534 116350
rect 195166 116150 195230 116214
rect 21902 115742 21966 115806
rect 21902 115606 21966 115670
rect 22174 115742 22238 115806
rect 22582 115742 22646 115806
rect 22310 115606 22374 115670
rect 22446 115606 22510 115670
rect 22990 115742 23054 115806
rect 22990 115606 23054 115670
rect 23398 115742 23462 115806
rect 23398 115606 23462 115670
rect 195166 116014 195230 116078
rect 195438 116150 195502 116214
rect 195438 116014 195502 116078
rect 195982 116014 196046 116078
rect 196118 116014 196182 116078
rect 196798 116150 196862 116214
rect 196798 116014 196862 116078
rect 195166 115742 195230 115806
rect 195030 115606 195094 115670
rect 195438 115742 195502 115806
rect 195438 115606 195502 115670
rect 195982 115742 196046 115806
rect 196118 115742 196182 115806
rect 196390 115606 196454 115670
rect 196798 115742 196862 115806
rect 196798 115606 196862 115670
rect 21902 115334 21966 115398
rect 21766 115198 21830 115262
rect 22310 115334 22374 115398
rect 22446 115334 22510 115398
rect 22174 115198 22238 115262
rect 22446 115198 22510 115262
rect 22990 115334 23054 115398
rect 23126 115198 23190 115262
rect 23398 115334 23462 115398
rect 23534 115198 23598 115262
rect 195030 115334 195094 115398
rect 195166 115198 195230 115262
rect 195438 115334 195502 115398
rect 195438 115198 195502 115262
rect 195846 115198 195910 115262
rect 196390 115334 196454 115398
rect 196254 115198 196318 115262
rect 196798 115334 196862 115398
rect 196662 115198 196726 115262
rect 21766 114926 21830 114990
rect 21766 114790 21830 114854
rect 22174 114926 22238 114990
rect 22446 114926 22510 114990
rect 22446 114790 22510 114854
rect 23126 114926 23190 114990
rect 23126 114790 23190 114854
rect 23534 114926 23598 114990
rect 23398 114790 23462 114854
rect 195166 114926 195230 114990
rect 195030 114790 195094 114854
rect 195438 114926 195502 114990
rect 195574 114790 195638 114854
rect 195846 114926 195910 114990
rect 195982 114790 196046 114854
rect 196254 114926 196318 114990
rect 196662 114926 196726 114990
rect 196798 114790 196862 114854
rect 217470 114790 217534 114854
rect 1230 114654 1294 114718
rect 21766 114518 21830 114582
rect 22446 114518 22510 114582
rect 22174 114382 22238 114446
rect 23126 114518 23190 114582
rect 22990 114382 23054 114446
rect 23398 114518 23462 114582
rect 23534 114382 23598 114446
rect 28566 114246 28630 114310
rect 195030 114518 195094 114582
rect 195030 114382 195094 114446
rect 195574 114518 195638 114582
rect 195438 114382 195502 114446
rect 195982 114518 196046 114582
rect 196390 114382 196454 114446
rect 196798 114518 196862 114582
rect 190270 114246 190334 114310
rect 22174 114110 22238 114174
rect 22990 114110 23054 114174
rect 23126 113974 23190 114038
rect 23534 114110 23598 114174
rect 23534 113974 23598 114038
rect 28566 113974 28630 114038
rect 22174 113566 22238 113630
rect 23126 113702 23190 113766
rect 23534 113702 23598 113766
rect 28294 113702 28358 113766
rect 190270 113974 190334 114038
rect 195030 114110 195094 114174
rect 195166 113974 195230 114038
rect 195438 114110 195502 114174
rect 195574 113974 195638 114038
rect 196390 114110 196454 114174
rect 21766 113294 21830 113358
rect 22174 113294 22238 113358
rect 28294 113430 28358 113494
rect 1230 113022 1294 113086
rect 21766 113022 21830 113086
rect 21766 112886 21830 112950
rect 22582 112886 22646 112950
rect 28430 113022 28494 113086
rect 190134 113430 190198 113494
rect 190134 113158 190198 113222
rect 190270 113158 190334 113222
rect 195166 113702 195230 113766
rect 195574 113702 195638 113766
rect 195982 113566 196046 113630
rect 196118 113566 196182 113630
rect 190134 113022 190198 113086
rect 21766 112614 21830 112678
rect 21902 112478 21966 112542
rect 22582 112614 22646 112678
rect 23126 112478 23190 112542
rect 23398 112478 23462 112542
rect 28430 112750 28494 112814
rect 190270 112750 190334 112814
rect 190134 112614 190198 112678
rect 195982 113294 196046 113358
rect 196118 113294 196182 113358
rect 196662 113294 196726 113358
rect 195982 112886 196046 112950
rect 196662 113022 196726 113086
rect 196662 112886 196726 112950
rect 217470 112886 217534 112950
rect 195030 112478 195094 112542
rect 195574 112478 195638 112542
rect 195982 112614 196046 112678
rect 21902 112206 21966 112270
rect 21902 112070 21966 112134
rect 22310 112070 22374 112134
rect 22446 112070 22510 112134
rect 23126 112206 23190 112270
rect 22990 112070 23054 112134
rect 23398 112206 23462 112270
rect 196662 112614 196726 112678
rect 196798 112478 196862 112542
rect 23398 112070 23462 112134
rect 21902 111798 21966 111862
rect 21902 111662 21966 111726
rect 22310 111798 22374 111862
rect 22446 111798 22510 111862
rect 22174 111662 22238 111726
rect 22582 111662 22646 111726
rect 22990 111798 23054 111862
rect 23126 111662 23190 111726
rect 23398 111798 23462 111862
rect 23534 111662 23598 111726
rect 28294 111798 28358 111862
rect 28294 111526 28358 111590
rect 1230 111254 1294 111318
rect 21902 111390 21966 111454
rect 21902 111254 21966 111318
rect 22174 111390 22238 111454
rect 22582 111390 22646 111454
rect 22446 111254 22510 111318
rect 23126 111390 23190 111454
rect 23126 111254 23190 111318
rect 23534 111390 23598 111454
rect 195030 112206 195094 112270
rect 195030 112070 195094 112134
rect 195574 112206 195638 112270
rect 195438 112070 195502 112134
rect 196798 112206 196862 112270
rect 196662 112070 196726 112134
rect 195030 111798 195094 111862
rect 195030 111662 195094 111726
rect 195438 111798 195502 111862
rect 195574 111662 195638 111726
rect 195982 111662 196046 111726
rect 196662 111798 196726 111862
rect 196662 111662 196726 111726
rect 23398 111254 23462 111318
rect 195030 111390 195094 111454
rect 195030 111254 195094 111318
rect 195574 111390 195638 111454
rect 195438 111254 195502 111318
rect 195982 111390 196046 111454
rect 196390 111254 196454 111318
rect 196662 111390 196726 111454
rect 196798 111254 196862 111318
rect 217470 111390 217534 111454
rect 21902 110982 21966 111046
rect 21766 110846 21830 110910
rect 22446 110982 22510 111046
rect 22174 110846 22238 110910
rect 22582 110846 22646 110910
rect 23126 110982 23190 111046
rect 23126 110846 23190 110910
rect 23398 110982 23462 111046
rect 23534 110846 23598 110910
rect 195030 110982 195094 111046
rect 195166 110846 195230 110910
rect 195438 110982 195502 111046
rect 195574 110846 195638 110910
rect 196390 110982 196454 111046
rect 196254 110846 196318 110910
rect 196798 110982 196862 111046
rect 196662 110846 196726 110910
rect 21766 110574 21830 110638
rect 22174 110574 22238 110638
rect 22582 110574 22646 110638
rect 22174 110438 22238 110502
rect 22446 110438 22510 110502
rect 23126 110574 23190 110638
rect 23126 110438 23190 110502
rect 23534 110574 23598 110638
rect 195166 110574 195230 110638
rect 23534 110438 23598 110502
rect 195166 110438 195230 110502
rect 195574 110574 195638 110638
rect 195438 110438 195502 110502
rect 195846 110438 195910 110502
rect 196254 110574 196318 110638
rect 196662 110574 196726 110638
rect 190270 110302 190334 110366
rect 22174 110166 22238 110230
rect 22446 110166 22510 110230
rect 22446 110030 22510 110094
rect 23126 110166 23190 110230
rect 22990 110030 23054 110094
rect 23534 110166 23598 110230
rect 23398 110030 23462 110094
rect 1230 109622 1294 109686
rect 22446 109758 22510 109822
rect 22582 109622 22646 109686
rect 22990 109758 23054 109822
rect 22990 109622 23054 109686
rect 23398 109758 23462 109822
rect 23534 109622 23598 109686
rect 190134 110030 190198 110094
rect 190270 110030 190334 110094
rect 195166 110166 195230 110230
rect 195030 110030 195094 110094
rect 195438 110166 195502 110230
rect 195574 110030 195638 110094
rect 195846 110166 195910 110230
rect 195030 109758 195094 109822
rect 190134 109622 190198 109686
rect 195166 109622 195230 109686
rect 195574 109758 195638 109822
rect 195574 109622 195638 109686
rect 196118 109622 196182 109686
rect 217470 109758 217534 109822
rect 190270 109486 190334 109550
rect 21766 109350 21830 109414
rect 22582 109350 22646 109414
rect 22990 109350 23054 109414
rect 23534 109350 23598 109414
rect 21766 109078 21830 109142
rect 21766 108942 21830 109006
rect 22446 108942 22510 109006
rect 21766 108670 21830 108734
rect 21766 108534 21830 108598
rect 22446 108670 22510 108734
rect 28430 109078 28494 109142
rect 190270 109214 190334 109278
rect 190270 109078 190334 109142
rect 195166 109350 195230 109414
rect 195574 109350 195638 109414
rect 196118 109350 196182 109414
rect 196798 109350 196862 109414
rect 28430 108806 28494 108870
rect 28294 108670 28358 108734
rect 190270 108806 190334 108870
rect 190134 108670 190198 108734
rect 21766 108262 21830 108326
rect 1230 108126 1294 108190
rect 21902 108126 21966 108190
rect 22718 108126 22782 108190
rect 23126 108126 23190 108190
rect 23398 108126 23462 108190
rect 28294 108398 28358 108462
rect 190134 108398 190198 108462
rect 196118 108942 196182 109006
rect 196798 109078 196862 109142
rect 196798 108942 196862 109006
rect 196118 108670 196182 108734
rect 196798 108670 196862 108734
rect 196662 108534 196726 108598
rect 196254 108398 196318 108462
rect 190134 108262 190198 108326
rect 21902 107854 21966 107918
rect 21902 107718 21966 107782
rect 22718 107854 22782 107918
rect 22446 107718 22510 107782
rect 23126 107854 23190 107918
rect 22990 107718 23054 107782
rect 23398 107854 23462 107918
rect 23398 107718 23462 107782
rect 28430 107854 28494 107918
rect 195030 108126 195094 108190
rect 195438 108126 195502 108190
rect 196118 108262 196182 108326
rect 196118 108126 196182 108190
rect 196662 108262 196726 108326
rect 196798 108126 196862 108190
rect 217470 108126 217534 108190
rect 190134 107854 190198 107918
rect 190270 107854 190334 107918
rect 195030 107854 195094 107918
rect 195166 107718 195230 107782
rect 195438 107854 195502 107918
rect 195574 107718 195638 107782
rect 196118 107854 196182 107918
rect 196390 107718 196454 107782
rect 196798 107854 196862 107918
rect 196798 107718 196862 107782
rect 28430 107582 28494 107646
rect 21902 107446 21966 107510
rect 21902 107310 21966 107374
rect 22446 107446 22510 107510
rect 22174 107310 22238 107374
rect 22582 107310 22646 107374
rect 22990 107446 23054 107510
rect 22990 107310 23054 107374
rect 23398 107446 23462 107510
rect 23398 107310 23462 107374
rect 190270 107582 190334 107646
rect 195166 107446 195230 107510
rect 195030 107310 195094 107374
rect 195574 107446 195638 107510
rect 195438 107310 195502 107374
rect 195982 107310 196046 107374
rect 196390 107446 196454 107510
rect 196254 107310 196318 107374
rect 196798 107446 196862 107510
rect 196798 107310 196862 107374
rect 21902 107038 21966 107102
rect 21902 106902 21966 106966
rect 22174 107038 22238 107102
rect 22582 107038 22646 107102
rect 22310 106902 22374 106966
rect 22990 107038 23054 107102
rect 23126 106902 23190 106966
rect 23398 107038 23462 107102
rect 23398 106902 23462 106966
rect 195030 107038 195094 107102
rect 195030 106902 195094 106966
rect 195438 107038 195502 107102
rect 195438 106902 195502 106966
rect 195982 107038 196046 107102
rect 196254 107038 196318 107102
rect 196118 106902 196182 106966
rect 196798 107038 196862 107102
rect 196798 106902 196862 106966
rect 21902 106630 21966 106694
rect 22310 106630 22374 106694
rect 22174 106494 22238 106558
rect 23126 106630 23190 106694
rect 23126 106494 23190 106558
rect 23398 106630 23462 106694
rect 23534 106494 23598 106558
rect 1230 106358 1294 106422
rect 195030 106630 195094 106694
rect 195166 106494 195230 106558
rect 195438 106630 195502 106694
rect 195574 106494 195638 106558
rect 196118 106630 196182 106694
rect 195846 106494 195910 106558
rect 196254 106494 196318 106558
rect 196798 106630 196862 106694
rect 22174 106222 22238 106286
rect 23126 106222 23190 106286
rect 23126 106086 23190 106150
rect 23534 106222 23598 106286
rect 23534 106086 23598 106150
rect 195166 106222 195230 106286
rect 195166 106086 195230 106150
rect 195574 106222 195638 106286
rect 195574 106086 195638 106150
rect 195846 106222 195910 106286
rect 196254 106222 196318 106286
rect 217470 106222 217534 106286
rect 22174 105678 22238 105742
rect 22582 105678 22646 105742
rect 23126 105814 23190 105878
rect 23126 105678 23190 105742
rect 23534 105814 23598 105878
rect 23534 105678 23598 105742
rect 28566 105542 28630 105606
rect 195166 105814 195230 105878
rect 195166 105678 195230 105742
rect 195574 105814 195638 105878
rect 195438 105678 195502 105742
rect 196254 105678 196318 105742
rect 190270 105542 190334 105606
rect 21766 105406 21830 105470
rect 22174 105406 22238 105470
rect 22582 105406 22646 105470
rect 23126 105406 23190 105470
rect 23534 105406 23598 105470
rect 21766 105134 21830 105198
rect 21766 104998 21830 105062
rect 22446 104998 22510 105062
rect 22582 104998 22646 105062
rect 1230 104726 1294 104790
rect 21766 104726 21830 104790
rect 21766 104590 21830 104654
rect 22446 104726 22510 104790
rect 22582 104726 22646 104790
rect 28566 105270 28630 105334
rect 28430 105134 28494 105198
rect 190270 105270 190334 105334
rect 195166 105406 195230 105470
rect 195438 105406 195502 105470
rect 190270 105134 190334 105198
rect 28430 104862 28494 104926
rect 21766 104318 21830 104382
rect 21766 104182 21830 104246
rect 22582 104182 22646 104246
rect 22990 104182 23054 104246
rect 190270 104862 190334 104926
rect 190270 104454 190334 104518
rect 196254 105406 196318 105470
rect 196662 105406 196726 105470
rect 195846 104998 195910 105062
rect 196118 104998 196182 105062
rect 196662 105134 196726 105198
rect 196798 104998 196862 105062
rect 23534 104182 23598 104246
rect 21766 103910 21830 103974
rect 21902 103774 21966 103838
rect 22582 103910 22646 103974
rect 22990 103910 23054 103974
rect 22990 103774 23054 103838
rect 23534 103910 23598 103974
rect 23398 103774 23462 103838
rect 190270 104182 190334 104246
rect 195166 104182 195230 104246
rect 195574 104182 195638 104246
rect 195846 104726 195910 104790
rect 196118 104726 196182 104790
rect 196798 104726 196862 104790
rect 196662 104590 196726 104654
rect 217470 104590 217534 104654
rect 195846 104182 195910 104246
rect 196662 104318 196726 104382
rect 196662 104182 196726 104246
rect 195166 103910 195230 103974
rect 195030 103774 195094 103838
rect 195574 103910 195638 103974
rect 195438 103774 195502 103838
rect 195846 103910 195910 103974
rect 196662 103910 196726 103974
rect 196798 103774 196862 103838
rect 21902 103502 21966 103566
rect 21766 103366 21830 103430
rect 22446 103366 22510 103430
rect 22990 103502 23054 103566
rect 23126 103366 23190 103430
rect 23398 103502 23462 103566
rect 23398 103366 23462 103430
rect 195030 103502 195094 103566
rect 195166 103366 195230 103430
rect 195438 103502 195502 103566
rect 195574 103366 195638 103430
rect 195846 103366 195910 103430
rect 196798 103502 196862 103566
rect 196798 103366 196862 103430
rect 1230 103094 1294 103158
rect 21766 103094 21830 103158
rect 21902 102958 21966 103022
rect 22446 103094 22510 103158
rect 22310 102958 22374 103022
rect 22718 102958 22782 103022
rect 23126 103094 23190 103158
rect 22990 102958 23054 103022
rect 23398 103094 23462 103158
rect 23398 102958 23462 103022
rect 21902 102686 21966 102750
rect 22310 102686 22374 102750
rect 22718 102686 22782 102750
rect 22446 102550 22510 102614
rect 22990 102686 23054 102750
rect 22990 102550 23054 102614
rect 23398 102686 23462 102750
rect 195166 103094 195230 103158
rect 195166 102958 195230 103022
rect 195574 103094 195638 103158
rect 195438 102958 195502 103022
rect 195846 103094 195910 103158
rect 196798 103094 196862 103158
rect 196798 102958 196862 103022
rect 217470 102958 217534 103022
rect 23398 102550 23462 102614
rect 195166 102686 195230 102750
rect 195030 102550 195094 102614
rect 195438 102686 195502 102750
rect 195574 102550 195638 102614
rect 195982 102550 196046 102614
rect 196390 102550 196454 102614
rect 196798 102686 196862 102750
rect 21902 102142 21966 102206
rect 22446 102278 22510 102342
rect 22990 102278 23054 102342
rect 23126 102142 23190 102206
rect 23398 102278 23462 102342
rect 23534 102142 23598 102206
rect 195030 102278 195094 102342
rect 195166 102142 195230 102206
rect 195574 102278 195638 102342
rect 195438 102142 195502 102206
rect 195982 102278 196046 102342
rect 196390 102278 196454 102342
rect 196118 102142 196182 102206
rect 196662 102142 196726 102206
rect 21902 101870 21966 101934
rect 22310 101734 22374 101798
rect 22446 101734 22510 101798
rect 23126 101870 23190 101934
rect 23126 101734 23190 101798
rect 23534 101870 23598 101934
rect 195166 101870 195230 101934
rect 23534 101734 23598 101798
rect 28430 101598 28494 101662
rect 195030 101734 195094 101798
rect 195438 101870 195502 101934
rect 195438 101734 195502 101798
rect 196118 101870 196182 101934
rect 195846 101734 195910 101798
rect 196662 101870 196726 101934
rect 21902 101462 21966 101526
rect 22310 101462 22374 101526
rect 22446 101462 22510 101526
rect 23126 101462 23190 101526
rect 22990 101326 23054 101390
rect 23534 101462 23598 101526
rect 23534 101326 23598 101390
rect 28430 101326 28494 101390
rect 1230 101190 1294 101254
rect 21902 101190 21966 101254
rect 22174 100918 22238 100982
rect 22582 100918 22646 100982
rect 22990 101054 23054 101118
rect 23534 101054 23598 101118
rect 21766 100646 21830 100710
rect 22174 100646 22238 100710
rect 22582 100646 22646 100710
rect 21766 100374 21830 100438
rect 21766 100238 21830 100302
rect 22446 100238 22510 100302
rect 23126 100238 23190 100302
rect 23398 100238 23462 100302
rect 21766 99966 21830 100030
rect 21766 99830 21830 99894
rect 1230 99558 1294 99622
rect 22446 99966 22510 100030
rect 23126 99966 23190 100030
rect 23126 99830 23190 99894
rect 23398 99966 23462 100030
rect 23534 99830 23598 99894
rect 190270 101326 190334 101390
rect 195030 101462 195094 101526
rect 195030 101326 195094 101390
rect 195438 101462 195502 101526
rect 195438 101326 195502 101390
rect 195846 101462 195910 101526
rect 196798 101462 196862 101526
rect 217470 101326 217534 101390
rect 195030 101054 195094 101118
rect 190270 100918 190334 100982
rect 195438 101054 195502 101118
rect 195846 100918 195910 100982
rect 196254 100918 196318 100982
rect 196798 101190 196862 101254
rect 195846 100646 195910 100710
rect 196254 100646 196318 100710
rect 196662 100646 196726 100710
rect 195030 100238 195094 100302
rect 195574 100238 195638 100302
rect 195846 100238 195910 100302
rect 196662 100374 196726 100438
rect 196798 100238 196862 100302
rect 195030 99966 195094 100030
rect 195166 99830 195230 99894
rect 195574 99966 195638 100030
rect 195574 99830 195638 99894
rect 195846 99966 195910 100030
rect 21766 99558 21830 99622
rect 21902 99422 21966 99486
rect 22718 99422 22782 99486
rect 23126 99558 23190 99622
rect 23126 99422 23190 99486
rect 23534 99558 23598 99622
rect 23398 99422 23462 99486
rect 196798 99966 196862 100030
rect 196662 99830 196726 99894
rect 217470 99694 217534 99758
rect 195166 99558 195230 99622
rect 195030 99422 195094 99486
rect 195574 99558 195638 99622
rect 195574 99422 195638 99486
rect 196662 99558 196726 99622
rect 196798 99422 196862 99486
rect 21902 99150 21966 99214
rect 21766 99014 21830 99078
rect 22718 99150 22782 99214
rect 23126 99150 23190 99214
rect 23126 99014 23190 99078
rect 23398 99150 23462 99214
rect 23534 99014 23598 99078
rect 195030 99150 195094 99214
rect 195030 99014 195094 99078
rect 195574 99150 195638 99214
rect 195574 99014 195638 99078
rect 196118 99014 196182 99078
rect 196798 99150 196862 99214
rect 196798 99014 196862 99078
rect 21766 98742 21830 98806
rect 21766 98606 21830 98670
rect 22174 98606 22238 98670
rect 22718 98606 22782 98670
rect 23126 98742 23190 98806
rect 22990 98606 23054 98670
rect 23534 98742 23598 98806
rect 23534 98606 23598 98670
rect 195030 98742 195094 98806
rect 195030 98606 195094 98670
rect 195574 98742 195638 98806
rect 195574 98606 195638 98670
rect 196118 98742 196182 98806
rect 195982 98606 196046 98670
rect 196798 98742 196862 98806
rect 196662 98606 196726 98670
rect 21766 98334 21830 98398
rect 21902 98198 21966 98262
rect 22174 98334 22238 98398
rect 22718 98334 22782 98398
rect 22310 98198 22374 98262
rect 22446 98198 22510 98262
rect 22990 98334 23054 98398
rect 23126 98198 23190 98262
rect 23534 98334 23598 98398
rect 23398 98198 23462 98262
rect 195030 98334 195094 98398
rect 195030 98198 195094 98262
rect 195574 98334 195638 98398
rect 195574 98198 195638 98262
rect 195982 98334 196046 98398
rect 196390 98198 196454 98262
rect 196662 98334 196726 98398
rect 196798 98198 196862 98262
rect 1230 97926 1294 97990
rect 21902 97926 21966 97990
rect 22310 97926 22374 97990
rect 22446 97926 22510 97990
rect 22174 97790 22238 97854
rect 23126 97926 23190 97990
rect 22990 97790 23054 97854
rect 23398 97926 23462 97990
rect 23534 97790 23598 97854
rect 195030 97926 195094 97990
rect 195166 97790 195230 97854
rect 195574 97926 195638 97990
rect 195438 97790 195502 97854
rect 195846 97790 195910 97854
rect 196390 97926 196454 97990
rect 196254 97790 196318 97854
rect 196798 97926 196862 97990
rect 217470 97790 217534 97854
rect 22174 97518 22238 97582
rect 22990 97518 23054 97582
rect 22990 97382 23054 97446
rect 23534 97518 23598 97582
rect 23534 97382 23598 97446
rect 22718 96974 22782 97038
rect 22990 97110 23054 97174
rect 23534 97110 23598 97174
rect 21766 96702 21830 96766
rect 22718 96702 22782 96766
rect 21766 96430 21830 96494
rect 21766 96294 21830 96358
rect 22310 96294 22374 96358
rect 1230 96158 1294 96222
rect 195166 97518 195230 97582
rect 195030 97382 195094 97446
rect 195438 97518 195502 97582
rect 195574 97382 195638 97446
rect 195846 97518 195910 97582
rect 196254 97518 196318 97582
rect 195030 97110 195094 97174
rect 28566 96838 28630 96902
rect 28566 96566 28630 96630
rect 28430 96430 28494 96494
rect 190134 96430 190198 96494
rect 195574 97110 195638 97174
rect 196254 96974 196318 97038
rect 196254 96702 196318 96766
rect 196662 96702 196726 96766
rect 28430 96158 28494 96222
rect 21766 96022 21830 96086
rect 21766 95886 21830 95950
rect 22310 96022 22374 96086
rect 22990 95886 23054 95950
rect 23398 95886 23462 95950
rect 28430 96022 28494 96086
rect 190134 96158 190198 96222
rect 195982 96294 196046 96358
rect 196118 96294 196182 96358
rect 196662 96430 196726 96494
rect 196662 96294 196726 96358
rect 217470 96294 217534 96358
rect 195030 95886 195094 95950
rect 195574 95886 195638 95950
rect 195982 96022 196046 96086
rect 196118 96022 196182 96086
rect 28430 95750 28494 95814
rect 21766 95614 21830 95678
rect 21766 95478 21830 95542
rect 22582 95478 22646 95542
rect 22990 95614 23054 95678
rect 22990 95478 23054 95542
rect 23398 95614 23462 95678
rect 196662 96022 196726 96086
rect 196798 95886 196862 95950
rect 196254 95750 196318 95814
rect 23534 95478 23598 95542
rect 21766 95206 21830 95270
rect 21902 95070 21966 95134
rect 22582 95206 22646 95270
rect 22718 95070 22782 95134
rect 22990 95206 23054 95270
rect 23126 95070 23190 95134
rect 23534 95206 23598 95270
rect 23398 95070 23462 95134
rect 195030 95614 195094 95678
rect 195166 95478 195230 95542
rect 195574 95614 195638 95678
rect 195574 95478 195638 95542
rect 196118 95614 196182 95678
rect 196118 95478 196182 95542
rect 196798 95614 196862 95678
rect 196662 95478 196726 95542
rect 190270 95206 190334 95270
rect 195166 95206 195230 95270
rect 195030 95070 195094 95134
rect 195574 95206 195638 95270
rect 195574 95070 195638 95134
rect 196118 95206 196182 95270
rect 195982 95070 196046 95134
rect 196662 95206 196726 95270
rect 196798 95070 196862 95134
rect 21902 94798 21966 94862
rect 1230 94662 1294 94726
rect 21766 94662 21830 94726
rect 22718 94798 22782 94862
rect 22310 94662 22374 94726
rect 22446 94662 22510 94726
rect 23126 94798 23190 94862
rect 22990 94662 23054 94726
rect 23398 94798 23462 94862
rect 190270 94934 190334 94998
rect 23534 94662 23598 94726
rect 195030 94798 195094 94862
rect 195030 94662 195094 94726
rect 195574 94798 195638 94862
rect 195574 94662 195638 94726
rect 195982 94798 196046 94862
rect 196118 94662 196182 94726
rect 196798 94798 196862 94862
rect 196662 94662 196726 94726
rect 217470 94526 217534 94590
rect 21766 94390 21830 94454
rect 21766 94254 21830 94318
rect 22310 94390 22374 94454
rect 22446 94390 22510 94454
rect 22718 94254 22782 94318
rect 22990 94390 23054 94454
rect 22990 94254 23054 94318
rect 23534 94390 23598 94454
rect 23534 94254 23598 94318
rect 21766 93982 21830 94046
rect 22718 93982 22782 94046
rect 22310 93846 22374 93910
rect 22990 93982 23054 94046
rect 22990 93846 23054 93910
rect 23534 93982 23598 94046
rect 195030 94390 195094 94454
rect 195030 94254 195094 94318
rect 195574 94390 195638 94454
rect 195438 94254 195502 94318
rect 196118 94390 196182 94454
rect 195982 94254 196046 94318
rect 196118 94254 196182 94318
rect 196254 94254 196318 94318
rect 196662 94390 196726 94454
rect 196662 94254 196726 94318
rect 23398 93846 23462 93910
rect 28294 93710 28358 93774
rect 195030 93982 195094 94046
rect 195030 93846 195094 93910
rect 195438 93982 195502 94046
rect 195438 93846 195502 93910
rect 195982 93982 196046 94046
rect 196118 93982 196182 94046
rect 196254 93982 196318 94046
rect 195982 93846 196046 93910
rect 196662 93982 196726 94046
rect 22310 93574 22374 93638
rect 22990 93574 23054 93638
rect 22990 93438 23054 93502
rect 23398 93574 23462 93638
rect 23534 93438 23598 93502
rect 28294 93438 28358 93502
rect 22990 93166 23054 93230
rect 23126 93030 23190 93094
rect 23534 93166 23598 93230
rect 195030 93574 195094 93638
rect 195166 93438 195230 93502
rect 195438 93574 195502 93638
rect 195574 93438 195638 93502
rect 195982 93574 196046 93638
rect 195166 93166 195230 93230
rect 23398 93030 23462 93094
rect 1230 92758 1294 92822
rect 195030 93030 195094 93094
rect 195574 93166 195638 93230
rect 195574 93030 195638 93094
rect 190270 92894 190334 92958
rect 21902 92758 21966 92822
rect 21902 92486 21966 92550
rect 21766 92350 21830 92414
rect 22446 92350 22510 92414
rect 23126 92758 23190 92822
rect 23398 92758 23462 92822
rect 28566 92486 28630 92550
rect 190270 92622 190334 92686
rect 190134 92486 190198 92550
rect 195030 92758 195094 92822
rect 195574 92758 195638 92822
rect 196798 92758 196862 92822
rect 217470 92894 217534 92958
rect 21766 92078 21830 92142
rect 21766 91942 21830 92006
rect 22446 92078 22510 92142
rect 22990 91942 23054 92006
rect 23534 91942 23598 92006
rect 28566 92214 28630 92278
rect 190134 92214 190198 92278
rect 196118 92350 196182 92414
rect 196798 92486 196862 92550
rect 196662 92350 196726 92414
rect 195166 91942 195230 92006
rect 195438 91942 195502 92006
rect 22446 91806 22510 91870
rect 21766 91670 21830 91734
rect 21902 91534 21966 91598
rect 22446 91534 22510 91598
rect 22718 91534 22782 91598
rect 22990 91670 23054 91734
rect 23126 91534 23190 91598
rect 23534 91670 23598 91734
rect 196118 92078 196182 92142
rect 196662 92078 196726 92142
rect 196798 91942 196862 92006
rect 23534 91534 23598 91598
rect 1230 91126 1294 91190
rect 21902 91262 21966 91326
rect 21766 91126 21830 91190
rect 22718 91262 22782 91326
rect 22174 91126 22238 91190
rect 22582 91126 22646 91190
rect 23126 91262 23190 91326
rect 22990 91126 23054 91190
rect 23534 91262 23598 91326
rect 23534 91126 23598 91190
rect 195166 91670 195230 91734
rect 195030 91534 195094 91598
rect 195438 91670 195502 91734
rect 195438 91534 195502 91598
rect 196254 91534 196318 91598
rect 196798 91670 196862 91734
rect 196662 91534 196726 91598
rect 195030 91262 195094 91326
rect 195166 91126 195230 91190
rect 195438 91262 195502 91326
rect 195574 91126 195638 91190
rect 196254 91262 196318 91326
rect 195846 91126 195910 91190
rect 196662 91262 196726 91326
rect 196662 91126 196726 91190
rect 217470 91262 217534 91326
rect 21766 90854 21830 90918
rect 21902 90718 21966 90782
rect 22174 90854 22238 90918
rect 22582 90854 22646 90918
rect 22718 90718 22782 90782
rect 22990 90854 23054 90918
rect 23126 90718 23190 90782
rect 23534 90854 23598 90918
rect 23398 90718 23462 90782
rect 195166 90854 195230 90918
rect 195030 90718 195094 90782
rect 195574 90854 195638 90918
rect 195574 90718 195638 90782
rect 195846 90854 195910 90918
rect 196118 90718 196182 90782
rect 196662 90854 196726 90918
rect 196798 90718 196862 90782
rect 21902 90446 21966 90510
rect 21902 90310 21966 90374
rect 22718 90446 22782 90510
rect 22310 90310 22374 90374
rect 23126 90446 23190 90510
rect 22990 90310 23054 90374
rect 23398 90446 23462 90510
rect 23534 90310 23598 90374
rect 195030 90446 195094 90510
rect 195030 90310 195094 90374
rect 195574 90446 195638 90510
rect 195574 90310 195638 90374
rect 196118 90446 196182 90510
rect 195846 90310 195910 90374
rect 196798 90446 196862 90510
rect 196798 90310 196862 90374
rect 21902 90038 21966 90102
rect 22310 90038 22374 90102
rect 22174 89902 22238 89966
rect 22718 89902 22782 89966
rect 22990 90038 23054 90102
rect 22990 89902 23054 89966
rect 23534 90038 23598 90102
rect 23534 89902 23598 89966
rect 195030 90038 195094 90102
rect 1230 89494 1294 89558
rect 28566 89766 28630 89830
rect 22174 89630 22238 89694
rect 22718 89630 22782 89694
rect 22990 89630 23054 89694
rect 23126 89494 23190 89558
rect 23534 89630 23598 89694
rect 23398 89494 23462 89558
rect 28566 89494 28630 89558
rect 22174 89086 22238 89150
rect 23126 89222 23190 89286
rect 23126 89086 23190 89150
rect 23398 89222 23462 89286
rect 23534 89086 23598 89150
rect 195030 89902 195094 89966
rect 195574 90038 195638 90102
rect 195438 89902 195502 89966
rect 195846 90038 195910 90102
rect 195982 89902 196046 89966
rect 196118 89902 196182 89966
rect 196798 90038 196862 90102
rect 195030 89630 195094 89694
rect 195030 89494 195094 89558
rect 195438 89630 195502 89694
rect 195438 89494 195502 89558
rect 195982 89630 196046 89694
rect 196118 89630 196182 89694
rect 217470 89630 217534 89694
rect 195030 89222 195094 89286
rect 195166 89086 195230 89150
rect 195438 89222 195502 89286
rect 195438 89086 195502 89150
rect 195982 89086 196046 89150
rect 196254 89086 196318 89150
rect 190134 88950 190198 89014
rect 21902 88814 21966 88878
rect 22174 88814 22238 88878
rect 23126 88814 23190 88878
rect 23534 88814 23598 88878
rect 21902 88542 21966 88606
rect 21902 88406 21966 88470
rect 22174 88406 22238 88470
rect 22446 88406 22510 88470
rect 28430 88542 28494 88606
rect 190134 88678 190198 88742
rect 190270 88678 190334 88742
rect 195166 88814 195230 88878
rect 195438 88814 195502 88878
rect 195982 88814 196046 88878
rect 196254 88814 196318 88878
rect 196662 88814 196726 88878
rect 21902 88134 21966 88198
rect 21766 87998 21830 88062
rect 22174 88134 22238 88198
rect 22446 88134 22510 88198
rect 1230 87862 1294 87926
rect 21766 87726 21830 87790
rect 21766 87590 21830 87654
rect 22310 87590 22374 87654
rect 22446 87590 22510 87654
rect 22582 87590 22646 87654
rect 23126 87590 23190 87654
rect 28430 88270 28494 88334
rect 28566 88134 28630 88198
rect 28566 87862 28630 87926
rect 190270 88270 190334 88334
rect 190134 87862 190198 87926
rect 196118 88406 196182 88470
rect 196662 88542 196726 88606
rect 196798 88406 196862 88470
rect 23534 87590 23598 87654
rect 21766 87318 21830 87382
rect 21766 87182 21830 87246
rect 22310 87318 22374 87382
rect 22446 87318 22510 87382
rect 22582 87318 22646 87382
rect 22174 87182 22238 87246
rect 22446 87182 22510 87246
rect 23126 87318 23190 87382
rect 22990 87182 23054 87246
rect 23534 87318 23598 87382
rect 23398 87182 23462 87246
rect 28430 87318 28494 87382
rect 190134 87590 190198 87654
rect 195030 87590 195094 87654
rect 195574 87590 195638 87654
rect 196118 88134 196182 88198
rect 196798 88134 196862 88198
rect 196662 87998 196726 88062
rect 195982 87590 196046 87654
rect 196390 87590 196454 87654
rect 196662 87726 196726 87790
rect 217470 87726 217534 87790
rect 196662 87590 196726 87654
rect 190270 87318 190334 87382
rect 195030 87318 195094 87382
rect 195030 87182 195094 87246
rect 195574 87318 195638 87382
rect 195438 87182 195502 87246
rect 195982 87318 196046 87382
rect 196390 87318 196454 87382
rect 196254 87182 196318 87246
rect 196662 87318 196726 87382
rect 196662 87182 196726 87246
rect 28430 87046 28494 87110
rect 21766 86910 21830 86974
rect 21766 86774 21830 86838
rect 22174 86910 22238 86974
rect 22446 86910 22510 86974
rect 22582 86774 22646 86838
rect 22990 86910 23054 86974
rect 23126 86774 23190 86838
rect 23398 86910 23462 86974
rect 190270 87046 190334 87110
rect 195030 86910 195094 86974
rect 23534 86774 23598 86838
rect 195166 86774 195230 86838
rect 195438 86910 195502 86974
rect 195574 86774 195638 86838
rect 196254 86910 196318 86974
rect 195846 86774 195910 86838
rect 196118 86774 196182 86838
rect 196662 86910 196726 86974
rect 196662 86774 196726 86838
rect 21766 86502 21830 86566
rect 21902 86366 21966 86430
rect 22582 86502 22646 86566
rect 22310 86366 22374 86430
rect 23126 86502 23190 86566
rect 23126 86366 23190 86430
rect 23534 86502 23598 86566
rect 23398 86366 23462 86430
rect 195166 86502 195230 86566
rect 195030 86366 195094 86430
rect 195574 86502 195638 86566
rect 195438 86366 195502 86430
rect 195846 86502 195910 86566
rect 196118 86502 196182 86566
rect 195982 86366 196046 86430
rect 196118 86366 196182 86430
rect 196662 86502 196726 86566
rect 196798 86366 196862 86430
rect 1230 86230 1294 86294
rect 21902 86094 21966 86158
rect 22310 86094 22374 86158
rect 23126 86094 23190 86158
rect 23126 85958 23190 86022
rect 23398 86094 23462 86158
rect 23398 85958 23462 86022
rect 195030 86094 195094 86158
rect 195030 85958 195094 86022
rect 195438 86094 195502 86158
rect 195574 85958 195638 86022
rect 195982 86094 196046 86158
rect 196118 86094 196182 86158
rect 195846 85958 195910 86022
rect 196798 86094 196862 86158
rect 217470 86094 217534 86158
rect 21902 85550 21966 85614
rect 22174 85550 22238 85614
rect 22582 85550 22646 85614
rect 23126 85686 23190 85750
rect 23126 85550 23190 85614
rect 23398 85686 23462 85750
rect 23398 85550 23462 85614
rect 195030 85686 195094 85750
rect 195030 85550 195094 85614
rect 195574 85686 195638 85750
rect 195438 85550 195502 85614
rect 195846 85686 195910 85750
rect 195982 85550 196046 85614
rect 196798 85550 196862 85614
rect 21902 85278 21966 85342
rect 22174 85278 22238 85342
rect 22582 85278 22646 85342
rect 22310 85142 22374 85206
rect 23126 85278 23190 85342
rect 23126 85142 23190 85206
rect 23398 85278 23462 85342
rect 23398 85142 23462 85206
rect 28294 85006 28358 85070
rect 195030 85278 195094 85342
rect 195030 85142 195094 85206
rect 195438 85278 195502 85342
rect 195574 85142 195638 85206
rect 195982 85278 196046 85342
rect 196390 85142 196454 85206
rect 196798 85278 196862 85342
rect 21902 84870 21966 84934
rect 22310 84870 22374 84934
rect 23126 84870 23190 84934
rect 23126 84734 23190 84798
rect 23398 84870 23462 84934
rect 23534 84734 23598 84798
rect 28294 84734 28358 84798
rect 1230 84462 1294 84526
rect 21902 84598 21966 84662
rect 22310 84326 22374 84390
rect 22446 84326 22510 84390
rect 23126 84462 23190 84526
rect 21902 84054 21966 84118
rect 22310 84054 22374 84118
rect 22446 84054 22510 84118
rect 21902 83782 21966 83846
rect 21766 83646 21830 83710
rect 22310 83646 22374 83710
rect 22582 83646 22646 83710
rect 23126 83646 23190 83710
rect 23534 84462 23598 84526
rect 28430 84462 28494 84526
rect 195030 84870 195094 84934
rect 195166 84734 195230 84798
rect 195574 84870 195638 84934
rect 195438 84734 195502 84798
rect 196390 84870 196454 84934
rect 196798 84870 196862 84934
rect 195166 84462 195230 84526
rect 28430 84190 28494 84254
rect 28566 84190 28630 84254
rect 28566 83918 28630 83982
rect 28566 83782 28630 83846
rect 190270 84190 190334 84254
rect 190270 83918 190334 83982
rect 23534 83646 23598 83710
rect 21766 83374 21830 83438
rect 21766 83238 21830 83302
rect 22310 83374 22374 83438
rect 22582 83374 22646 83438
rect 23126 83374 23190 83438
rect 23126 83238 23190 83302
rect 23534 83374 23598 83438
rect 23534 83238 23598 83302
rect 28430 83374 28494 83438
rect 28566 83374 28630 83438
rect 28430 83102 28494 83166
rect 21766 82966 21830 83030
rect 21766 82830 21830 82894
rect 22718 82830 22782 82894
rect 23126 82966 23190 83030
rect 23126 82830 23190 82894
rect 23534 82966 23598 83030
rect 195438 84462 195502 84526
rect 195846 84326 195910 84390
rect 196118 84326 196182 84390
rect 196798 84598 196862 84662
rect 217470 84326 217534 84390
rect 195846 84054 195910 84118
rect 196118 84054 196182 84118
rect 196798 84054 196862 84118
rect 195166 83646 195230 83710
rect 195438 83646 195502 83710
rect 195846 83646 195910 83710
rect 196798 83782 196862 83846
rect 196662 83646 196726 83710
rect 195166 83374 195230 83438
rect 195166 83238 195230 83302
rect 195438 83374 195502 83438
rect 195574 83238 195638 83302
rect 195846 83374 195910 83438
rect 195982 83238 196046 83302
rect 196390 83238 196454 83302
rect 196662 83374 196726 83438
rect 196662 83238 196726 83302
rect 23534 82830 23598 82894
rect 1230 82694 1294 82758
rect 195166 82966 195230 83030
rect 195166 82830 195230 82894
rect 195574 82966 195638 83030
rect 195438 82830 195502 82894
rect 195982 82966 196046 83030
rect 196390 82966 196454 83030
rect 196254 82830 196318 82894
rect 196662 82966 196726 83030
rect 196798 82830 196862 82894
rect 217470 82830 217534 82894
rect 21766 82558 21830 82622
rect 21766 82422 21830 82486
rect 22718 82558 22782 82622
rect 22174 82422 22238 82486
rect 22582 82422 22646 82486
rect 23126 82558 23190 82622
rect 23126 82422 23190 82486
rect 23534 82558 23598 82622
rect 23534 82422 23598 82486
rect 195166 82558 195230 82622
rect 195166 82422 195230 82486
rect 195438 82558 195502 82622
rect 195438 82422 195502 82486
rect 195846 82422 195910 82486
rect 196254 82558 196318 82622
rect 196254 82422 196318 82486
rect 196798 82558 196862 82622
rect 196662 82422 196726 82486
rect 21766 82150 21830 82214
rect 21902 82014 21966 82078
rect 22174 82150 22238 82214
rect 22582 82150 22646 82214
rect 22718 82014 22782 82078
rect 23126 82150 23190 82214
rect 23126 82014 23190 82078
rect 23534 82150 23598 82214
rect 23398 82014 23462 82078
rect 195166 82150 195230 82214
rect 195030 82014 195094 82078
rect 195438 82150 195502 82214
rect 195438 82014 195502 82078
rect 195846 82150 195910 82214
rect 196254 82150 196318 82214
rect 195982 82014 196046 82078
rect 196662 82150 196726 82214
rect 196798 82014 196862 82078
rect 21902 81742 21966 81806
rect 21766 81606 21830 81670
rect 22718 81742 22782 81806
rect 22310 81606 22374 81670
rect 22446 81606 22510 81670
rect 23126 81742 23190 81806
rect 23126 81606 23190 81670
rect 23398 81742 23462 81806
rect 23534 81606 23598 81670
rect 195030 81742 195094 81806
rect 195166 81606 195230 81670
rect 195438 81742 195502 81806
rect 195438 81606 195502 81670
rect 195982 81742 196046 81806
rect 196118 81606 196182 81670
rect 196798 81742 196862 81806
rect 196662 81606 196726 81670
rect 21766 81334 21830 81398
rect 1230 81062 1294 81126
rect 22310 81334 22374 81398
rect 22446 81334 22510 81398
rect 22582 81198 22646 81262
rect 23126 81334 23190 81398
rect 22990 81198 23054 81262
rect 23534 81334 23598 81398
rect 23534 81198 23598 81262
rect 195166 81334 195230 81398
rect 28566 81062 28630 81126
rect 195166 81198 195230 81262
rect 195438 81334 195502 81398
rect 195438 81198 195502 81262
rect 196118 81334 196182 81398
rect 195982 81198 196046 81262
rect 196118 81198 196182 81262
rect 196662 81334 196726 81398
rect 217470 81198 217534 81262
rect 21902 80926 21966 80990
rect 22446 80926 22510 80990
rect 22582 80926 22646 80990
rect 22990 80926 23054 80990
rect 22990 80790 23054 80854
rect 23534 80926 23598 80990
rect 23398 80790 23462 80854
rect 28430 80790 28494 80854
rect 28566 80790 28630 80854
rect 21902 80654 21966 80718
rect 22446 80654 22510 80718
rect 22446 80382 22510 80446
rect 22990 80518 23054 80582
rect 23398 80518 23462 80582
rect 195166 80926 195230 80990
rect 195030 80790 195094 80854
rect 195438 80926 195502 80990
rect 195574 80790 195638 80854
rect 195982 80926 196046 80990
rect 196118 80926 196182 80990
rect 196662 80926 196726 80990
rect 21766 80110 21830 80174
rect 22446 80110 22510 80174
rect 21766 79838 21830 79902
rect 21902 79702 21966 79766
rect 22310 79702 22374 79766
rect 22446 79702 22510 79766
rect 1230 79566 1294 79630
rect 28430 80382 28494 80446
rect 28294 80246 28358 80310
rect 28294 79974 28358 80038
rect 28430 79974 28494 80038
rect 195030 80518 195094 80582
rect 195574 80518 195638 80582
rect 195982 80382 196046 80446
rect 196662 80654 196726 80718
rect 190134 80246 190198 80310
rect 190134 79974 190198 80038
rect 195982 80110 196046 80174
rect 196798 80110 196862 80174
rect 190270 79838 190334 79902
rect 28430 79566 28494 79630
rect 21902 79430 21966 79494
rect 21766 79294 21830 79358
rect 22310 79430 22374 79494
rect 22446 79430 22510 79494
rect 23126 79294 23190 79358
rect 23534 79294 23598 79358
rect 28566 79430 28630 79494
rect 28566 79158 28630 79222
rect 21766 79022 21830 79086
rect 21902 78886 21966 78950
rect 22582 78886 22646 78950
rect 23126 79022 23190 79086
rect 22990 78886 23054 78950
rect 23534 79022 23598 79086
rect 23398 78886 23462 78950
rect 190270 79566 190334 79630
rect 190270 79430 190334 79494
rect 196390 79702 196454 79766
rect 196798 79838 196862 79902
rect 196798 79702 196862 79766
rect 195166 79294 195230 79358
rect 195574 79294 195638 79358
rect 190270 79158 190334 79222
rect 196390 79430 196454 79494
rect 196798 79430 196862 79494
rect 196662 79294 196726 79358
rect 217470 79294 217534 79358
rect 195166 79022 195230 79086
rect 195166 78886 195230 78950
rect 195574 79022 195638 79086
rect 195438 78886 195502 78950
rect 195846 78886 195910 78950
rect 196118 78886 196182 78950
rect 196662 79022 196726 79086
rect 196798 78886 196862 78950
rect 21902 78614 21966 78678
rect 21902 78478 21966 78542
rect 22582 78614 22646 78678
rect 22174 78478 22238 78542
rect 22718 78478 22782 78542
rect 22990 78614 23054 78678
rect 22990 78478 23054 78542
rect 23398 78614 23462 78678
rect 23398 78478 23462 78542
rect 195166 78614 195230 78678
rect 195166 78478 195230 78542
rect 195438 78614 195502 78678
rect 195574 78478 195638 78542
rect 195846 78614 195910 78678
rect 196118 78614 196182 78678
rect 195846 78478 195910 78542
rect 196798 78614 196862 78678
rect 196798 78478 196862 78542
rect 21902 78206 21966 78270
rect 21766 78070 21830 78134
rect 22174 78206 22238 78270
rect 22718 78206 22782 78270
rect 22582 78070 22646 78134
rect 22990 78206 23054 78270
rect 22990 78070 23054 78134
rect 23398 78206 23462 78270
rect 195166 78206 195230 78270
rect 23534 78070 23598 78134
rect 195166 78070 195230 78134
rect 195574 78206 195638 78270
rect 195438 78070 195502 78134
rect 195846 78206 195910 78270
rect 195846 78070 195910 78134
rect 196798 78206 196862 78270
rect 196662 78070 196726 78134
rect 1230 77662 1294 77726
rect 21766 77798 21830 77862
rect 21902 77662 21966 77726
rect 22582 77798 22646 77862
rect 22446 77662 22510 77726
rect 22990 77798 23054 77862
rect 22990 77662 23054 77726
rect 23534 77798 23598 77862
rect 23398 77662 23462 77726
rect 195166 77798 195230 77862
rect 195030 77662 195094 77726
rect 195438 77798 195502 77862
rect 195438 77662 195502 77726
rect 195846 77798 195910 77862
rect 195982 77662 196046 77726
rect 196390 77662 196454 77726
rect 196662 77798 196726 77862
rect 196798 77662 196862 77726
rect 217470 77798 217534 77862
rect 21902 77390 21966 77454
rect 22446 77390 22510 77454
rect 22310 77254 22374 77318
rect 22990 77390 23054 77454
rect 22990 77254 23054 77318
rect 23398 77390 23462 77454
rect 23534 77254 23598 77318
rect 195030 77390 195094 77454
rect 195166 77254 195230 77318
rect 195438 77390 195502 77454
rect 195438 77254 195502 77318
rect 195982 77390 196046 77454
rect 196390 77390 196454 77454
rect 195846 77254 195910 77318
rect 196390 77254 196454 77318
rect 196798 77390 196862 77454
rect 190134 77118 190198 77182
rect 22310 76982 22374 77046
rect 22990 76982 23054 77046
rect 22990 76846 23054 76910
rect 23534 76982 23598 77046
rect 23534 76846 23598 76910
rect 22310 76438 22374 76502
rect 22446 76438 22510 76502
rect 22990 76574 23054 76638
rect 23534 76574 23598 76638
rect 190134 76846 190198 76910
rect 195166 76982 195230 77046
rect 195166 76846 195230 76910
rect 195438 76982 195502 77046
rect 195438 76846 195502 76910
rect 195846 76982 195910 77046
rect 196390 76982 196454 77046
rect 1230 76166 1294 76230
rect 21766 76166 21830 76230
rect 22310 76166 22374 76230
rect 22446 76166 22510 76230
rect 28566 76302 28630 76366
rect 190270 76302 190334 76366
rect 21766 75894 21830 75958
rect 21766 75758 21830 75822
rect 22174 75758 22238 75822
rect 22446 75758 22510 75822
rect 28566 76030 28630 76094
rect 28430 75894 28494 75958
rect 190270 76030 190334 76094
rect 195166 76574 195230 76638
rect 195438 76574 195502 76638
rect 195846 76438 195910 76502
rect 196118 76438 196182 76502
rect 190134 75894 190198 75958
rect 23262 75622 23326 75686
rect 21766 75486 21830 75550
rect 21902 75350 21966 75414
rect 22174 75486 22238 75550
rect 22446 75486 22510 75550
rect 23126 75350 23190 75414
rect 28430 75622 28494 75686
rect 23398 75350 23462 75414
rect 25302 75350 25366 75414
rect 28430 75486 28494 75550
rect 190134 75622 190198 75686
rect 195846 76166 195910 76230
rect 196118 76166 196182 76230
rect 196798 76166 196862 76230
rect 217470 76030 217534 76094
rect 196118 75758 196182 75822
rect 196390 75758 196454 75822
rect 196798 75894 196862 75958
rect 196662 75758 196726 75822
rect 190270 75486 190334 75550
rect 193126 75350 193190 75414
rect 23262 75214 23326 75278
rect 28430 75214 28494 75278
rect 21902 75078 21966 75142
rect 21766 74942 21830 75006
rect 22174 74942 22238 75006
rect 23126 75078 23190 75142
rect 22990 74942 23054 75006
rect 23398 75078 23462 75142
rect 25302 75078 25366 75142
rect 190270 75214 190334 75278
rect 195030 75350 195094 75414
rect 195438 75350 195502 75414
rect 196118 75486 196182 75550
rect 196390 75486 196454 75550
rect 196662 75486 196726 75550
rect 196798 75350 196862 75414
rect 193126 75078 193190 75142
rect 195030 75078 195094 75142
rect 23534 74942 23598 75006
rect 21766 74670 21830 74734
rect 1230 74534 1294 74598
rect 21766 74534 21830 74598
rect 22174 74670 22238 74734
rect 22990 74670 23054 74734
rect 22990 74534 23054 74598
rect 23534 74670 23598 74734
rect 23534 74534 23598 74598
rect 195166 74942 195230 75006
rect 195438 75078 195502 75142
rect 195438 74942 195502 75006
rect 196254 74942 196318 75006
rect 196798 75078 196862 75142
rect 196662 74942 196726 75006
rect 195166 74670 195230 74734
rect 195166 74534 195230 74598
rect 195438 74670 195502 74734
rect 195438 74534 195502 74598
rect 195846 74534 195910 74598
rect 196254 74670 196318 74734
rect 196390 74534 196454 74598
rect 196662 74670 196726 74734
rect 196798 74534 196862 74598
rect 217470 74534 217534 74598
rect 21766 74262 21830 74326
rect 21766 74126 21830 74190
rect 22174 74126 22238 74190
rect 22718 74126 22782 74190
rect 22990 74262 23054 74326
rect 22990 74126 23054 74190
rect 23534 74262 23598 74326
rect 23534 74126 23598 74190
rect 195166 74262 195230 74326
rect 195166 74126 195230 74190
rect 195438 74262 195502 74326
rect 195438 74126 195502 74190
rect 195846 74262 195910 74326
rect 196390 74262 196454 74326
rect 196118 74126 196182 74190
rect 196798 74262 196862 74326
rect 196662 74126 196726 74190
rect 21766 73854 21830 73918
rect 21766 73718 21830 73782
rect 22174 73854 22238 73918
rect 22718 73854 22782 73918
rect 22582 73718 22646 73782
rect 22990 73854 23054 73918
rect 23126 73718 23190 73782
rect 23534 73854 23598 73918
rect 23534 73718 23598 73782
rect 195166 73854 195230 73918
rect 195166 73718 195230 73782
rect 195438 73854 195502 73918
rect 195574 73718 195638 73782
rect 196118 73854 196182 73918
rect 195846 73718 195910 73782
rect 196254 73718 196318 73782
rect 196662 73854 196726 73918
rect 196662 73718 196726 73782
rect 21766 73446 21830 73510
rect 22174 73310 22238 73374
rect 22582 73446 22646 73510
rect 22718 73310 22782 73374
rect 23126 73446 23190 73510
rect 23126 73310 23190 73374
rect 23534 73446 23598 73510
rect 23398 73310 23462 73374
rect 195166 73446 195230 73510
rect 195030 73310 195094 73374
rect 195574 73446 195638 73510
rect 195438 73310 195502 73374
rect 195846 73446 195910 73510
rect 196254 73446 196318 73510
rect 195982 73310 196046 73374
rect 196118 73310 196182 73374
rect 196662 73446 196726 73510
rect 22174 73038 22238 73102
rect 22718 73038 22782 73102
rect 23126 73038 23190 73102
rect 23126 72902 23190 72966
rect 23398 73038 23462 73102
rect 23534 72902 23598 72966
rect 28294 72902 28358 72966
rect 1230 72630 1294 72694
rect 22718 72494 22782 72558
rect 23126 72630 23190 72694
rect 22990 72494 23054 72558
rect 23534 72630 23598 72694
rect 23398 72494 23462 72558
rect 195030 73038 195094 73102
rect 195030 72902 195094 72966
rect 195438 73038 195502 73102
rect 195574 72902 195638 72966
rect 195982 73038 196046 73102
rect 196118 73038 196182 73102
rect 195030 72630 195094 72694
rect 28294 72494 28358 72558
rect 28566 72358 28630 72422
rect 195030 72494 195094 72558
rect 195574 72630 195638 72694
rect 195438 72494 195502 72558
rect 196118 72494 196182 72558
rect 217470 72766 217534 72830
rect 21902 72222 21966 72286
rect 22718 72222 22782 72286
rect 21902 71950 21966 72014
rect 21902 71814 21966 71878
rect 22310 71814 22374 71878
rect 22446 71814 22510 71878
rect 22990 72222 23054 72286
rect 23398 72222 23462 72286
rect 28566 72086 28630 72150
rect 28566 71950 28630 72014
rect 190134 71950 190198 72014
rect 195030 72222 195094 72286
rect 195438 72222 195502 72286
rect 196118 72222 196182 72286
rect 196798 72222 196862 72286
rect 21902 71542 21966 71606
rect 21902 71406 21966 71470
rect 22310 71542 22374 71606
rect 22446 71542 22510 71606
rect 1230 70998 1294 71062
rect 21902 71134 21966 71198
rect 21902 70998 21966 71062
rect 22990 70998 23054 71062
rect 28566 71678 28630 71742
rect 28430 71270 28494 71334
rect 28294 71134 28358 71198
rect 190134 71678 190198 71742
rect 190134 71542 190198 71606
rect 190134 71270 190198 71334
rect 190270 71270 190334 71334
rect 196390 71814 196454 71878
rect 196798 71950 196862 72014
rect 196798 71814 196862 71878
rect 23398 70998 23462 71062
rect 28430 70998 28494 71062
rect 21902 70726 21966 70790
rect 21766 70590 21830 70654
rect 22446 70590 22510 70654
rect 22990 70726 23054 70790
rect 22990 70590 23054 70654
rect 23398 70726 23462 70790
rect 23534 70590 23598 70654
rect 28294 70726 28358 70790
rect 28566 70726 28630 70790
rect 28566 70454 28630 70518
rect 21766 70318 21830 70382
rect 21902 70182 21966 70246
rect 22446 70318 22510 70382
rect 22310 70182 22374 70246
rect 22582 70182 22646 70246
rect 22990 70318 23054 70382
rect 22990 70182 23054 70246
rect 23534 70318 23598 70382
rect 23534 70182 23598 70246
rect 190270 70998 190334 71062
rect 195030 70998 195094 71062
rect 195574 70998 195638 71062
rect 196390 71542 196454 71606
rect 196798 71542 196862 71606
rect 196662 71406 196726 71470
rect 196390 70998 196454 71062
rect 196662 71134 196726 71198
rect 196798 70998 196862 71062
rect 217470 71134 217534 71198
rect 190134 70726 190198 70790
rect 195030 70726 195094 70790
rect 195166 70590 195230 70654
rect 195574 70726 195638 70790
rect 195438 70590 195502 70654
rect 196390 70726 196454 70790
rect 196118 70590 196182 70654
rect 196254 70590 196318 70654
rect 196798 70726 196862 70790
rect 196662 70590 196726 70654
rect 190134 70454 190198 70518
rect 195166 70318 195230 70382
rect 195030 70182 195094 70246
rect 195438 70318 195502 70382
rect 195438 70182 195502 70246
rect 196118 70318 196182 70382
rect 196254 70318 196318 70382
rect 195982 70182 196046 70246
rect 196118 70182 196182 70246
rect 196662 70318 196726 70382
rect 196662 70182 196726 70246
rect 21902 69910 21966 69974
rect 21766 69774 21830 69838
rect 22310 69910 22374 69974
rect 22582 69910 22646 69974
rect 22310 69774 22374 69838
rect 22582 69774 22646 69838
rect 22990 69910 23054 69974
rect 22990 69774 23054 69838
rect 23534 69910 23598 69974
rect 23534 69774 23598 69838
rect 195030 69910 195094 69974
rect 195030 69774 195094 69838
rect 195438 69910 195502 69974
rect 195438 69774 195502 69838
rect 195982 69910 196046 69974
rect 196118 69910 196182 69974
rect 196254 69774 196318 69838
rect 196662 69910 196726 69974
rect 196798 69774 196862 69838
rect 21766 69502 21830 69566
rect 1230 69366 1294 69430
rect 22310 69502 22374 69566
rect 22582 69502 22646 69566
rect 22582 69366 22646 69430
rect 22990 69502 23054 69566
rect 22990 69366 23054 69430
rect 23534 69502 23598 69566
rect 195030 69502 195094 69566
rect 23534 69366 23598 69430
rect 195166 69366 195230 69430
rect 195438 69502 195502 69566
rect 195574 69366 195638 69430
rect 196254 69502 196318 69566
rect 195846 69366 195910 69430
rect 196118 69366 196182 69430
rect 196798 69502 196862 69566
rect 21902 68958 21966 69022
rect 22582 69094 22646 69158
rect 22718 68958 22782 69022
rect 22990 69094 23054 69158
rect 23126 68958 23190 69022
rect 23534 69094 23598 69158
rect 23398 68958 23462 69022
rect 195166 69094 195230 69158
rect 195030 68958 195094 69022
rect 195574 69094 195638 69158
rect 195438 68958 195502 69022
rect 195846 69094 195910 69158
rect 196118 69094 196182 69158
rect 217470 69230 217534 69294
rect 196798 68958 196862 69022
rect 21902 68686 21966 68750
rect 22718 68686 22782 68750
rect 22310 68550 22374 68614
rect 23126 68686 23190 68750
rect 22990 68550 23054 68614
rect 23398 68686 23462 68750
rect 23534 68550 23598 68614
rect 195030 68686 195094 68750
rect 195030 68550 195094 68614
rect 195438 68686 195502 68750
rect 195574 68550 195638 68614
rect 195846 68550 195910 68614
rect 196798 68686 196862 68750
rect 190134 68414 190198 68478
rect 21766 68278 21830 68342
rect 22310 68278 22374 68342
rect 22990 68278 23054 68342
rect 23534 68278 23598 68342
rect 21766 68006 21830 68070
rect 21902 67870 21966 67934
rect 22446 67870 22510 67934
rect 1230 67734 1294 67798
rect 28430 68006 28494 68070
rect 190134 68142 190198 68206
rect 195030 68278 195094 68342
rect 190134 68006 190198 68070
rect 28430 67734 28494 67798
rect 21902 67598 21966 67662
rect 21902 67462 21966 67526
rect 22446 67598 22510 67662
rect 21902 67190 21966 67254
rect 21902 67054 21966 67118
rect 22582 67054 22646 67118
rect 23126 67054 23190 67118
rect 23398 67054 23462 67118
rect 28294 67598 28358 67662
rect 28294 67326 28358 67390
rect 190134 67734 190198 67798
rect 195574 68278 195638 68342
rect 195846 68278 195910 68342
rect 196662 68278 196726 68342
rect 196662 68006 196726 68070
rect 196798 67870 196862 67934
rect 196798 67598 196862 67662
rect 217470 67598 217534 67662
rect 196662 67462 196726 67526
rect 21902 66782 21966 66846
rect 21902 66646 21966 66710
rect 22582 66782 22646 66846
rect 22310 66646 22374 66710
rect 22718 66646 22782 66710
rect 23126 66782 23190 66846
rect 22990 66646 23054 66710
rect 23398 66782 23462 66846
rect 23398 66646 23462 66710
rect 28294 66782 28358 66846
rect 195030 67054 195094 67118
rect 195438 67054 195502 67118
rect 196662 67190 196726 67254
rect 196798 67054 196862 67118
rect 190270 66782 190334 66846
rect 195030 66782 195094 66846
rect 195030 66646 195094 66710
rect 195438 66782 195502 66846
rect 195438 66646 195502 66710
rect 196390 66646 196454 66710
rect 196798 66782 196862 66846
rect 196798 66646 196862 66710
rect 28294 66510 28358 66574
rect 21902 66374 21966 66438
rect 21766 66238 21830 66302
rect 22310 66374 22374 66438
rect 22718 66374 22782 66438
rect 22174 66238 22238 66302
rect 22446 66238 22510 66302
rect 22990 66374 23054 66438
rect 23126 66238 23190 66302
rect 23398 66374 23462 66438
rect 190270 66510 190334 66574
rect 23534 66238 23598 66302
rect 1230 66102 1294 66166
rect 195030 66374 195094 66438
rect 195166 66238 195230 66302
rect 195438 66374 195502 66438
rect 195438 66238 195502 66302
rect 195846 66238 195910 66302
rect 196390 66374 196454 66438
rect 196254 66238 196318 66302
rect 196798 66374 196862 66438
rect 196662 66238 196726 66302
rect 21766 65966 21830 66030
rect 21766 65830 21830 65894
rect 22174 65966 22238 66030
rect 22446 65966 22510 66030
rect 22582 65830 22646 65894
rect 23126 65966 23190 66030
rect 23126 65830 23190 65894
rect 23534 65966 23598 66030
rect 23398 65830 23462 65894
rect 21766 65558 21830 65622
rect 22582 65558 22646 65622
rect 22174 65422 22238 65486
rect 22446 65422 22510 65486
rect 23126 65558 23190 65622
rect 22990 65422 23054 65486
rect 23398 65558 23462 65622
rect 195166 65966 195230 66030
rect 195166 65830 195230 65894
rect 195438 65966 195502 66030
rect 195574 65830 195638 65894
rect 195846 65966 195910 66030
rect 196254 65966 196318 66030
rect 195982 65830 196046 65894
rect 196118 65830 196182 65894
rect 196662 65966 196726 66030
rect 217470 65966 217534 66030
rect 196662 65830 196726 65894
rect 23398 65422 23462 65486
rect 195166 65558 195230 65622
rect 195030 65422 195094 65486
rect 195574 65558 195638 65622
rect 195438 65422 195502 65486
rect 195982 65558 196046 65622
rect 196118 65558 196182 65622
rect 196254 65422 196318 65486
rect 196662 65558 196726 65622
rect 21766 65014 21830 65078
rect 22174 65150 22238 65214
rect 22446 65150 22510 65214
rect 22582 65014 22646 65078
rect 22990 65150 23054 65214
rect 23126 65014 23190 65078
rect 23398 65150 23462 65214
rect 23534 65014 23598 65078
rect 195030 65150 195094 65214
rect 195166 65014 195230 65078
rect 195438 65150 195502 65214
rect 195574 65014 195638 65078
rect 196254 65150 196318 65214
rect 195846 65014 195910 65078
rect 196118 65014 196182 65078
rect 196662 65014 196726 65078
rect 21766 64742 21830 64806
rect 22582 64742 22646 64806
rect 22446 64606 22510 64670
rect 22718 64606 22782 64670
rect 23126 64742 23190 64806
rect 23126 64606 23190 64670
rect 23534 64742 23598 64806
rect 23398 64606 23462 64670
rect 28566 64470 28630 64534
rect 195166 64742 195230 64806
rect 195030 64606 195094 64670
rect 195574 64742 195638 64806
rect 195574 64606 195638 64670
rect 195846 64742 195910 64806
rect 196118 64742 196182 64806
rect 195982 64606 196046 64670
rect 196662 64742 196726 64806
rect 21902 64334 21966 64398
rect 1230 64198 1294 64262
rect 22446 64334 22510 64398
rect 22718 64334 22782 64398
rect 23126 64334 23190 64398
rect 23126 64198 23190 64262
rect 23398 64334 23462 64398
rect 23398 64198 23462 64262
rect 28566 64198 28630 64262
rect 21902 64062 21966 64126
rect 22718 63790 22782 63854
rect 23126 63926 23190 63990
rect 23398 63926 23462 63990
rect 21902 63518 21966 63582
rect 22718 63518 22782 63582
rect 21902 63246 21966 63310
rect 21902 63110 21966 63174
rect 22310 63110 22374 63174
rect 22446 63110 22510 63174
rect 195030 64334 195094 64398
rect 195166 64198 195230 64262
rect 195574 64334 195638 64398
rect 195574 64198 195638 64262
rect 195982 64334 196046 64398
rect 196798 64334 196862 64398
rect 217470 64334 217534 64398
rect 195166 63926 195230 63990
rect 28430 63654 28494 63718
rect 28294 63382 28358 63446
rect 28430 63382 28494 63446
rect 195574 63926 195638 63990
rect 195982 63790 196046 63854
rect 196798 64062 196862 64126
rect 190134 63654 190198 63718
rect 190134 63382 190198 63446
rect 190134 63246 190198 63310
rect 21902 62838 21966 62902
rect 21766 62702 21830 62766
rect 22310 62838 22374 62902
rect 22446 62838 22510 62902
rect 1230 62566 1294 62630
rect 22990 62702 23054 62766
rect 23398 62702 23462 62766
rect 28294 62974 28358 63038
rect 190134 62974 190198 63038
rect 190134 62838 190198 62902
rect 195982 63518 196046 63582
rect 196798 63518 196862 63582
rect 196118 63110 196182 63174
rect 196798 63246 196862 63310
rect 196662 63110 196726 63174
rect 195030 62702 195094 62766
rect 195438 62702 195502 62766
rect 21766 62430 21830 62494
rect 21902 62294 21966 62358
rect 22718 62294 22782 62358
rect 22990 62430 23054 62494
rect 23126 62294 23190 62358
rect 23398 62430 23462 62494
rect 23398 62294 23462 62358
rect 190134 62566 190198 62630
rect 196118 62838 196182 62902
rect 196662 62838 196726 62902
rect 196798 62702 196862 62766
rect 217470 62702 217534 62766
rect 195030 62430 195094 62494
rect 195030 62294 195094 62358
rect 195438 62430 195502 62494
rect 195438 62294 195502 62358
rect 195982 62294 196046 62358
rect 196798 62430 196862 62494
rect 196798 62294 196862 62358
rect 21902 62022 21966 62086
rect 21766 61886 21830 61950
rect 22174 61886 22238 61950
rect 22718 62022 22782 62086
rect 22582 61886 22646 61950
rect 23126 62022 23190 62086
rect 22990 61886 23054 61950
rect 23398 62022 23462 62086
rect 23534 61886 23598 61950
rect 195030 62022 195094 62086
rect 195166 61886 195230 61950
rect 195438 62022 195502 62086
rect 195574 61886 195638 61950
rect 195982 62022 196046 62086
rect 196118 61886 196182 61950
rect 196254 61886 196318 61950
rect 196798 62022 196862 62086
rect 196662 61886 196726 61950
rect 21766 61614 21830 61678
rect 21902 61478 21966 61542
rect 22174 61614 22238 61678
rect 22582 61614 22646 61678
rect 22990 61614 23054 61678
rect 23126 61478 23190 61542
rect 23534 61614 23598 61678
rect 195166 61614 195230 61678
rect 23534 61478 23598 61542
rect 195166 61478 195230 61542
rect 195574 61614 195638 61678
rect 195574 61478 195638 61542
rect 196118 61614 196182 61678
rect 196254 61614 196318 61678
rect 195982 61478 196046 61542
rect 196662 61614 196726 61678
rect 196662 61478 196726 61542
rect 21902 61206 21966 61270
rect 21902 61070 21966 61134
rect 22174 61070 22238 61134
rect 23126 61206 23190 61270
rect 22718 61070 22782 61134
rect 22990 61070 23054 61134
rect 23534 61206 23598 61270
rect 23534 61070 23598 61134
rect 195166 61206 195230 61270
rect 195030 61070 195094 61134
rect 195574 61206 195638 61270
rect 195438 61070 195502 61134
rect 195982 61206 196046 61270
rect 196118 61070 196182 61134
rect 196662 61206 196726 61270
rect 196662 61070 196726 61134
rect 217470 61070 217534 61134
rect 1230 60934 1294 60998
rect 21902 60798 21966 60862
rect 22174 60798 22238 60862
rect 22718 60798 22782 60862
rect 22582 60662 22646 60726
rect 22990 60798 23054 60862
rect 22990 60662 23054 60726
rect 23534 60798 23598 60862
rect 195030 60798 195094 60862
rect 23534 60662 23598 60726
rect 195166 60662 195230 60726
rect 195438 60798 195502 60862
rect 195438 60662 195502 60726
rect 196118 60798 196182 60862
rect 195846 60662 195910 60726
rect 196254 60662 196318 60726
rect 196662 60798 196726 60862
rect 22582 60390 22646 60454
rect 22990 60390 23054 60454
rect 23126 60254 23190 60318
rect 23534 60390 23598 60454
rect 23398 60254 23462 60318
rect 28294 60254 28358 60318
rect 22582 59846 22646 59910
rect 23126 59982 23190 60046
rect 23398 59982 23462 60046
rect 195166 60390 195230 60454
rect 195030 60254 195094 60318
rect 195438 60390 195502 60454
rect 195438 60254 195502 60318
rect 195846 60390 195910 60454
rect 196254 60390 196318 60454
rect 21766 59574 21830 59638
rect 22582 59574 22646 59638
rect 1230 59166 1294 59230
rect 21766 59302 21830 59366
rect 21902 59166 21966 59230
rect 22582 59166 22646 59230
rect 21902 58894 21966 58958
rect 21766 58758 21830 58822
rect 22582 58894 22646 58958
rect 22990 58758 23054 58822
rect 28294 59846 28358 59910
rect 28566 59302 28630 59366
rect 195030 59982 195094 60046
rect 195438 59982 195502 60046
rect 190270 59302 190334 59366
rect 28566 59030 28630 59094
rect 23534 58758 23598 58822
rect 28566 58894 28630 58958
rect 28566 58622 28630 58686
rect 21766 58486 21830 58550
rect 21902 58350 21966 58414
rect 22582 58350 22646 58414
rect 22990 58486 23054 58550
rect 22990 58350 23054 58414
rect 23534 58486 23598 58550
rect 190270 59030 190334 59094
rect 196662 59574 196726 59638
rect 195982 59166 196046 59230
rect 196662 59302 196726 59366
rect 196798 59166 196862 59230
rect 217470 59302 217534 59366
rect 190134 58894 190198 58958
rect 195166 58758 195230 58822
rect 195438 58758 195502 58822
rect 195982 58894 196046 58958
rect 190134 58622 190198 58686
rect 196798 58894 196862 58958
rect 196798 58758 196862 58822
rect 195166 58486 195230 58550
rect 23534 58350 23598 58414
rect 21902 58078 21966 58142
rect 21902 57942 21966 58006
rect 22582 58078 22646 58142
rect 22990 58078 23054 58142
rect 22990 57942 23054 58006
rect 23534 58078 23598 58142
rect 23398 57942 23462 58006
rect 28430 58078 28494 58142
rect 195030 58350 195094 58414
rect 195438 58486 195502 58550
rect 195438 58350 195502 58414
rect 195982 58350 196046 58414
rect 196118 58350 196182 58414
rect 196798 58486 196862 58550
rect 196662 58350 196726 58414
rect 195030 58078 195094 58142
rect 195030 57942 195094 58006
rect 195438 58078 195502 58142
rect 195574 57942 195638 58006
rect 195982 58078 196046 58142
rect 196118 58078 196182 58142
rect 196390 57942 196454 58006
rect 196662 58078 196726 58142
rect 196798 57942 196862 58006
rect 28430 57806 28494 57870
rect 1230 57670 1294 57734
rect 21902 57670 21966 57734
rect 21766 57534 21830 57598
rect 22174 57534 22238 57598
rect 22582 57534 22646 57598
rect 22990 57670 23054 57734
rect 22990 57534 23054 57598
rect 23398 57670 23462 57734
rect 23534 57534 23598 57598
rect 195030 57670 195094 57734
rect 195166 57534 195230 57598
rect 195574 57670 195638 57734
rect 195438 57534 195502 57598
rect 196390 57670 196454 57734
rect 196118 57534 196182 57598
rect 196254 57534 196318 57598
rect 196798 57670 196862 57734
rect 196662 57534 196726 57598
rect 217470 57534 217534 57598
rect 21766 57262 21830 57326
rect 21766 57126 21830 57190
rect 22174 57262 22238 57326
rect 22582 57262 22646 57326
rect 22990 57262 23054 57326
rect 23126 57126 23190 57190
rect 23534 57262 23598 57326
rect 23534 57126 23598 57190
rect 195166 57262 195230 57326
rect 195166 57126 195230 57190
rect 195438 57262 195502 57326
rect 195438 57126 195502 57190
rect 196118 57262 196182 57326
rect 196254 57262 196318 57326
rect 195846 57126 195910 57190
rect 196118 57126 196182 57190
rect 196662 57262 196726 57326
rect 196798 57126 196862 57190
rect 21766 56854 21830 56918
rect 22174 56718 22238 56782
rect 22718 56718 22782 56782
rect 23126 56854 23190 56918
rect 22990 56718 23054 56782
rect 23534 56854 23598 56918
rect 23534 56718 23598 56782
rect 195166 56854 195230 56918
rect 195166 56718 195230 56782
rect 195438 56854 195502 56918
rect 195438 56718 195502 56782
rect 195846 56854 195910 56918
rect 196118 56854 196182 56918
rect 196254 56718 196318 56782
rect 196798 56854 196862 56918
rect 190270 56582 190334 56646
rect 1230 55902 1294 55966
rect 22174 56446 22238 56510
rect 22718 56446 22782 56510
rect 22990 56446 23054 56510
rect 22990 56310 23054 56374
rect 23534 56446 23598 56510
rect 23534 56310 23598 56374
rect 22718 55902 22782 55966
rect 22990 56038 23054 56102
rect 22990 55902 23054 55966
rect 23534 56038 23598 56102
rect 23398 55902 23462 55966
rect 190270 56310 190334 56374
rect 195166 56446 195230 56510
rect 195166 56310 195230 56374
rect 195438 56446 195502 56510
rect 195574 56310 195638 56374
rect 196254 56446 196318 56510
rect 28294 55766 28358 55830
rect 195166 56038 195230 56102
rect 195030 55902 195094 55966
rect 195574 56038 195638 56102
rect 195438 55902 195502 55966
rect 195982 55902 196046 55966
rect 196118 55902 196182 55966
rect 21766 55630 21830 55694
rect 22718 55630 22782 55694
rect 21766 55358 21830 55422
rect 21766 55222 21830 55286
rect 22582 55222 22646 55286
rect 22990 55630 23054 55694
rect 23398 55630 23462 55694
rect 21766 54950 21830 55014
rect 21902 54814 21966 54878
rect 22582 54950 22646 55014
rect 21902 54542 21966 54606
rect 21766 54406 21830 54470
rect 22446 54406 22510 54470
rect 23126 54406 23190 54470
rect 28294 55494 28358 55558
rect 28294 55358 28358 55422
rect 190134 55358 190198 55422
rect 195030 55630 195094 55694
rect 195438 55630 195502 55694
rect 195982 55630 196046 55694
rect 196118 55630 196182 55694
rect 217470 55902 217534 55966
rect 196662 55630 196726 55694
rect 28294 55086 28358 55150
rect 28566 54950 28630 55014
rect 190134 55086 190198 55150
rect 190270 54950 190334 55014
rect 28294 54678 28358 54742
rect 28566 54678 28630 54742
rect 190270 54678 190334 54742
rect 23398 54406 23462 54470
rect 28294 54406 28358 54470
rect 1230 54134 1294 54198
rect 21766 54134 21830 54198
rect 21902 53998 21966 54062
rect 22446 54134 22510 54198
rect 22310 53998 22374 54062
rect 22718 53998 22782 54062
rect 23126 54134 23190 54198
rect 22990 53998 23054 54062
rect 23398 54134 23462 54198
rect 23398 53998 23462 54062
rect 196118 55222 196182 55286
rect 196662 55358 196726 55422
rect 196662 55222 196726 55286
rect 195166 54406 195230 54470
rect 195574 54406 195638 54470
rect 196118 54950 196182 55014
rect 196662 54950 196726 55014
rect 196798 54814 196862 54878
rect 195846 54406 195910 54470
rect 196390 54406 196454 54470
rect 196798 54542 196862 54606
rect 196798 54406 196862 54470
rect 217470 54270 217534 54334
rect 195166 54134 195230 54198
rect 195166 53998 195230 54062
rect 195574 54134 195638 54198
rect 195574 53998 195638 54062
rect 195846 54134 195910 54198
rect 196390 54134 196454 54198
rect 196798 54134 196862 54198
rect 196798 53998 196862 54062
rect 21902 53726 21966 53790
rect 21902 53590 21966 53654
rect 22310 53726 22374 53790
rect 22718 53726 22782 53790
rect 22990 53726 23054 53790
rect 23126 53590 23190 53654
rect 23398 53726 23462 53790
rect 23398 53590 23462 53654
rect 195166 53726 195230 53790
rect 195030 53590 195094 53654
rect 195574 53726 195638 53790
rect 195574 53590 195638 53654
rect 196390 53590 196454 53654
rect 196798 53726 196862 53790
rect 196798 53590 196862 53654
rect 21902 53318 21966 53382
rect 21766 53182 21830 53246
rect 22446 53182 22510 53246
rect 23126 53318 23190 53382
rect 22990 53182 23054 53246
rect 23398 53318 23462 53382
rect 23534 53182 23598 53246
rect 21766 52910 21830 52974
rect 22446 52910 22510 52974
rect 22310 52774 22374 52838
rect 22990 52910 23054 52974
rect 22990 52774 23054 52838
rect 23534 52910 23598 52974
rect 195030 53318 195094 53382
rect 195166 53182 195230 53246
rect 195574 53318 195638 53382
rect 195438 53182 195502 53246
rect 195846 53182 195910 53246
rect 196390 53318 196454 53382
rect 196390 53182 196454 53246
rect 196798 53318 196862 53382
rect 196662 53182 196726 53246
rect 195166 52910 195230 52974
rect 23398 52774 23462 52838
rect 1230 52502 1294 52566
rect 195166 52774 195230 52838
rect 195438 52910 195502 52974
rect 195438 52774 195502 52838
rect 195846 52910 195910 52974
rect 196390 52910 196454 52974
rect 195982 52774 196046 52838
rect 196118 52774 196182 52838
rect 196390 52774 196454 52838
rect 196662 52910 196726 52974
rect 22310 52502 22374 52566
rect 22990 52502 23054 52566
rect 22990 52366 23054 52430
rect 23398 52502 23462 52566
rect 23398 52366 23462 52430
rect 195166 52502 195230 52566
rect 195166 52366 195230 52430
rect 195438 52502 195502 52566
rect 195438 52366 195502 52430
rect 195982 52502 196046 52566
rect 196118 52502 196182 52566
rect 196390 52502 196454 52566
rect 22446 51958 22510 52022
rect 22990 52094 23054 52158
rect 23126 51958 23190 52022
rect 23398 52094 23462 52158
rect 195166 52094 195230 52158
rect 23534 51958 23598 52022
rect 28294 51822 28358 51886
rect 195166 51958 195230 52022
rect 195438 52094 195502 52158
rect 195438 51958 195502 52022
rect 195846 51958 195910 52022
rect 217470 52638 217534 52702
rect 21902 51686 21966 51750
rect 22446 51686 22510 51750
rect 21902 51414 21966 51478
rect 21766 51278 21830 51342
rect 22718 51278 22782 51342
rect 23126 51686 23190 51750
rect 23534 51686 23598 51750
rect 28294 51550 28358 51614
rect 28294 51414 28358 51478
rect 190270 51414 190334 51478
rect 195166 51686 195230 51750
rect 195438 51686 195502 51750
rect 195846 51686 195910 51750
rect 196662 51686 196726 51750
rect 1230 50870 1294 50934
rect 21766 51006 21830 51070
rect 21766 50870 21830 50934
rect 22718 51006 22782 51070
rect 21766 50598 21830 50662
rect 21902 50462 21966 50526
rect 22718 50462 22782 50526
rect 22990 50462 23054 50526
rect 28294 51142 28358 51206
rect 23398 50462 23462 50526
rect 21902 50190 21966 50254
rect 21766 50054 21830 50118
rect 22718 50190 22782 50254
rect 22310 50054 22374 50118
rect 22990 50190 23054 50254
rect 22990 50054 23054 50118
rect 23398 50190 23462 50254
rect 23398 50054 23462 50118
rect 28294 50190 28358 50254
rect 28294 49918 28358 49982
rect 21766 49782 21830 49846
rect 21766 49646 21830 49710
rect 22310 49782 22374 49846
rect 22174 49646 22238 49710
rect 22718 49646 22782 49710
rect 22990 49782 23054 49846
rect 22990 49646 23054 49710
rect 23398 49782 23462 49846
rect 23398 49646 23462 49710
rect 190270 51142 190334 51206
rect 195982 51278 196046 51342
rect 196662 51414 196726 51478
rect 196662 51278 196726 51342
rect 195030 50462 195094 50526
rect 195438 50462 195502 50526
rect 195982 51006 196046 51070
rect 196662 51006 196726 51070
rect 196662 50870 196726 50934
rect 217470 50734 217534 50798
rect 195982 50462 196046 50526
rect 196662 50598 196726 50662
rect 196798 50462 196862 50526
rect 195030 50190 195094 50254
rect 195030 50054 195094 50118
rect 195438 50190 195502 50254
rect 195438 50054 195502 50118
rect 195982 50190 196046 50254
rect 196390 50054 196454 50118
rect 196798 50190 196862 50254
rect 196798 50054 196862 50118
rect 195030 49782 195094 49846
rect 195438 49782 195502 49846
rect 195030 49646 195094 49710
rect 195438 49646 195502 49710
rect 195846 49646 195910 49710
rect 196390 49782 196454 49846
rect 196798 49782 196862 49846
rect 196662 49646 196726 49710
rect 21766 49374 21830 49438
rect 1230 49238 1294 49302
rect 21902 49238 21966 49302
rect 22174 49374 22238 49438
rect 22718 49374 22782 49438
rect 22310 49238 22374 49302
rect 22990 49374 23054 49438
rect 23126 49238 23190 49302
rect 23398 49374 23462 49438
rect 23398 49238 23462 49302
rect 195030 49374 195094 49438
rect 195030 49238 195094 49302
rect 195438 49374 195502 49438
rect 195574 49238 195638 49302
rect 195846 49374 195910 49438
rect 196390 49238 196454 49302
rect 196662 49374 196726 49438
rect 196798 49238 196862 49302
rect 21902 48966 21966 49030
rect 22310 48966 22374 49030
rect 22174 48830 22238 48894
rect 23126 48966 23190 49030
rect 22990 48830 23054 48894
rect 23398 48966 23462 49030
rect 23534 48830 23598 48894
rect 217470 49102 217534 49166
rect 195030 48966 195094 49030
rect 195166 48830 195230 48894
rect 195574 48966 195638 49030
rect 195438 48830 195502 48894
rect 195846 48830 195910 48894
rect 196390 48966 196454 49030
rect 196254 48830 196318 48894
rect 196798 48966 196862 49030
rect 21902 48422 21966 48486
rect 22174 48558 22238 48622
rect 22310 48422 22374 48486
rect 22582 48422 22646 48486
rect 22990 48558 23054 48622
rect 23126 48422 23190 48486
rect 23534 48558 23598 48622
rect 23534 48422 23598 48486
rect 21902 48150 21966 48214
rect 22310 48150 22374 48214
rect 22582 48150 22646 48214
rect 22718 48014 22782 48078
rect 23126 48150 23190 48214
rect 22990 48014 23054 48078
rect 23534 48150 23598 48214
rect 195166 48558 195230 48622
rect 195030 48422 195094 48486
rect 195438 48558 195502 48622
rect 195574 48422 195638 48486
rect 195846 48558 195910 48622
rect 196254 48558 196318 48622
rect 195846 48422 195910 48486
rect 196118 48422 196182 48486
rect 196798 48422 196862 48486
rect 23534 48014 23598 48078
rect 195030 48150 195094 48214
rect 195166 48014 195230 48078
rect 195574 48150 195638 48214
rect 195438 48014 195502 48078
rect 195846 48150 195910 48214
rect 196118 48150 196182 48214
rect 196254 48014 196318 48078
rect 196798 48150 196862 48214
rect 21902 47742 21966 47806
rect 22718 47742 22782 47806
rect 1230 47606 1294 47670
rect 22990 47742 23054 47806
rect 22990 47606 23054 47670
rect 23534 47742 23598 47806
rect 23534 47606 23598 47670
rect 21902 47470 21966 47534
rect 22446 47198 22510 47262
rect 22990 47334 23054 47398
rect 23534 47334 23598 47398
rect 195166 47742 195230 47806
rect 195166 47606 195230 47670
rect 195438 47742 195502 47806
rect 195438 47606 195502 47670
rect 21902 46926 21966 46990
rect 22446 46926 22510 46990
rect 22310 46790 22374 46854
rect 28294 47062 28358 47126
rect 28294 46790 28358 46854
rect 21902 46654 21966 46718
rect 21766 46518 21830 46582
rect 22446 46654 22510 46718
rect 22582 46518 22646 46582
rect 22990 46518 23054 46582
rect 195166 47334 195230 47398
rect 195438 47334 195502 47398
rect 196254 47742 196318 47806
rect 196662 47742 196726 47806
rect 196662 47470 196726 47534
rect 217470 47470 217534 47534
rect 23534 46518 23598 46582
rect 21766 46246 21830 46310
rect 21902 46110 21966 46174
rect 1230 45974 1294 46038
rect 22582 46246 22646 46310
rect 22990 46246 23054 46310
rect 23126 46110 23190 46174
rect 23534 46246 23598 46310
rect 23398 46110 23462 46174
rect 195166 46518 195230 46582
rect 196798 46926 196862 46990
rect 195438 46518 195502 46582
rect 196254 46518 196318 46582
rect 196798 46654 196862 46718
rect 196662 46518 196726 46582
rect 190134 46246 190198 46310
rect 195166 46246 195230 46310
rect 195030 46110 195094 46174
rect 195438 46246 195502 46310
rect 195574 46110 195638 46174
rect 21902 45838 21966 45902
rect 21902 45702 21966 45766
rect 22174 45702 22238 45766
rect 23126 45838 23190 45902
rect 23126 45702 23190 45766
rect 23398 45838 23462 45902
rect 190134 45974 190198 46038
rect 196254 46246 196318 46310
rect 196662 46246 196726 46310
rect 196798 46110 196862 46174
rect 217470 45974 217534 46038
rect 23534 45702 23598 45766
rect 14694 45566 14758 45630
rect 195030 45838 195094 45902
rect 195166 45702 195230 45766
rect 195574 45838 195638 45902
rect 195574 45702 195638 45766
rect 195846 45702 195910 45766
rect 196798 45838 196862 45902
rect 196662 45702 196726 45766
rect 21902 45430 21966 45494
rect 21902 45294 21966 45358
rect 22174 45430 22238 45494
rect 22718 45294 22782 45358
rect 23126 45430 23190 45494
rect 22990 45294 23054 45358
rect 23534 45430 23598 45494
rect 23534 45294 23598 45358
rect 195166 45430 195230 45494
rect 195166 45294 195230 45358
rect 195574 45430 195638 45494
rect 195438 45294 195502 45358
rect 195846 45430 195910 45494
rect 195846 45294 195910 45358
rect 196118 45294 196182 45358
rect 196662 45430 196726 45494
rect 196662 45294 196726 45358
rect 21902 45022 21966 45086
rect 21902 44886 21966 44950
rect 22718 45022 22782 45086
rect 22310 44886 22374 44950
rect 22990 45022 23054 45086
rect 23126 44886 23190 44950
rect 23534 45022 23598 45086
rect 23398 44886 23462 44950
rect 195166 45022 195230 45086
rect 195030 44886 195094 44950
rect 195438 45022 195502 45086
rect 195438 44886 195502 44950
rect 195846 45022 195910 45086
rect 196118 45022 196182 45086
rect 196390 44886 196454 44950
rect 196662 45022 196726 45086
rect 196798 44886 196862 44950
rect 21902 44614 21966 44678
rect 21766 44478 21830 44542
rect 22310 44614 22374 44678
rect 22174 44478 22238 44542
rect 22582 44478 22646 44542
rect 23126 44614 23190 44678
rect 22990 44478 23054 44542
rect 23398 44614 23462 44678
rect 23534 44478 23598 44542
rect 1230 44070 1294 44134
rect 14558 44070 14622 44134
rect 21766 44206 21830 44270
rect 22174 44206 22238 44270
rect 22582 44206 22646 44270
rect 22446 44070 22510 44134
rect 22990 44206 23054 44270
rect 23126 44070 23190 44134
rect 23534 44206 23598 44270
rect 195030 44614 195094 44678
rect 195166 44478 195230 44542
rect 195438 44614 195502 44678
rect 195574 44478 195638 44542
rect 196390 44614 196454 44678
rect 196254 44478 196318 44542
rect 196798 44614 196862 44678
rect 196662 44478 196726 44542
rect 195166 44206 195230 44270
rect 23534 44070 23598 44134
rect 195030 44070 195094 44134
rect 195574 44206 195638 44270
rect 195574 44070 195638 44134
rect 195982 44070 196046 44134
rect 196254 44206 196318 44270
rect 196390 44070 196454 44134
rect 196662 44206 196726 44270
rect 217470 44206 217534 44270
rect 22446 43798 22510 43862
rect 23126 43798 23190 43862
rect 22990 43662 23054 43726
rect 23534 43798 23598 43862
rect 23398 43662 23462 43726
rect 22446 43254 22510 43318
rect 22990 43390 23054 43454
rect 23398 43390 23462 43454
rect 195030 43798 195094 43862
rect 195030 43662 195094 43726
rect 195574 43798 195638 43862
rect 195574 43662 195638 43726
rect 195982 43798 196046 43862
rect 196390 43798 196454 43862
rect 190134 43390 190198 43454
rect 195030 43390 195094 43454
rect 21766 42982 21830 43046
rect 22446 42982 22510 43046
rect 14694 42846 14758 42910
rect 22446 42846 22510 42910
rect 14694 42710 14758 42774
rect 21766 42710 21830 42774
rect 21766 42574 21830 42638
rect 22446 42574 22510 42638
rect 22718 42574 22782 42638
rect 1230 42438 1294 42502
rect 28294 43118 28358 43182
rect 28294 42846 28358 42910
rect 28566 42846 28630 42910
rect 28294 42710 28358 42774
rect 190134 43118 190198 43182
rect 190270 43118 190334 43182
rect 190270 42846 190334 42910
rect 190270 42710 190334 42774
rect 195574 43390 195638 43454
rect 196390 43254 196454 43318
rect 196390 42982 196454 43046
rect 196662 42982 196726 43046
rect 21766 42302 21830 42366
rect 21766 42166 21830 42230
rect 22718 42302 22782 42366
rect 23126 42166 23190 42230
rect 23534 42166 23598 42230
rect 28294 42438 28358 42502
rect 28566 42438 28630 42502
rect 190270 42438 190334 42502
rect 195166 42166 195230 42230
rect 196390 42574 196454 42638
rect 196662 42710 196726 42774
rect 196662 42574 196726 42638
rect 217470 42574 217534 42638
rect 195574 42166 195638 42230
rect 21766 41894 21830 41958
rect 21902 41758 21966 41822
rect 22446 41758 22510 41822
rect 22718 41758 22782 41822
rect 23126 41894 23190 41958
rect 22990 41758 23054 41822
rect 23534 41894 23598 41958
rect 23398 41758 23462 41822
rect 14558 41486 14622 41550
rect 21902 41486 21966 41550
rect 21902 41350 21966 41414
rect 22446 41486 22510 41550
rect 22718 41486 22782 41550
rect 22310 41350 22374 41414
rect 22990 41486 23054 41550
rect 23126 41350 23190 41414
rect 23398 41486 23462 41550
rect 23398 41350 23462 41414
rect 28294 41486 28358 41550
rect 196390 42302 196454 42366
rect 196662 42302 196726 42366
rect 196662 42166 196726 42230
rect 195166 41894 195230 41958
rect 195030 41758 195094 41822
rect 195574 41894 195638 41958
rect 195438 41758 195502 41822
rect 196662 41894 196726 41958
rect 196798 41758 196862 41822
rect 190134 41486 190198 41550
rect 195030 41486 195094 41550
rect 195166 41350 195230 41414
rect 195438 41486 195502 41550
rect 195574 41350 195638 41414
rect 195846 41350 195910 41414
rect 196390 41350 196454 41414
rect 196798 41486 196862 41550
rect 196798 41350 196862 41414
rect 14558 41214 14622 41278
rect 28294 41214 28358 41278
rect 21902 41078 21966 41142
rect 21902 40942 21966 41006
rect 22310 41078 22374 41142
rect 22582 40942 22646 41006
rect 23126 41078 23190 41142
rect 22990 40942 23054 41006
rect 23398 41078 23462 41142
rect 23534 40942 23598 41006
rect 190134 41214 190198 41278
rect 195166 41078 195230 41142
rect 1230 40806 1294 40870
rect 195166 40942 195230 41006
rect 195574 41078 195638 41142
rect 195438 40942 195502 41006
rect 195846 41078 195910 41142
rect 196390 41078 196454 41142
rect 196798 41078 196862 41142
rect 196662 40942 196726 41006
rect 217470 40806 217534 40870
rect 21902 40670 21966 40734
rect 21902 40534 21966 40598
rect 22582 40670 22646 40734
rect 22310 40534 22374 40598
rect 22990 40670 23054 40734
rect 23126 40534 23190 40598
rect 23534 40670 23598 40734
rect 23398 40534 23462 40598
rect 195166 40670 195230 40734
rect 195030 40534 195094 40598
rect 195438 40670 195502 40734
rect 195438 40534 195502 40598
rect 196390 40534 196454 40598
rect 196662 40670 196726 40734
rect 196798 40534 196862 40598
rect 21902 40262 21966 40326
rect 22310 40262 22374 40326
rect 22174 40126 22238 40190
rect 22446 40126 22510 40190
rect 23126 40262 23190 40326
rect 22990 40126 23054 40190
rect 23398 40262 23462 40326
rect 23534 40126 23598 40190
rect 14694 39990 14758 40054
rect 14694 39854 14758 39918
rect 28294 39990 28358 40054
rect 195030 40262 195094 40326
rect 195166 40126 195230 40190
rect 195438 40262 195502 40326
rect 195574 40126 195638 40190
rect 195846 40126 195910 40190
rect 196390 40262 196454 40326
rect 196254 40126 196318 40190
rect 196798 40262 196862 40326
rect 190134 39990 190198 40054
rect 22174 39854 22238 39918
rect 22446 39854 22510 39918
rect 22990 39854 23054 39918
rect 22990 39718 23054 39782
rect 23534 39854 23598 39918
rect 23398 39718 23462 39782
rect 28294 39718 28358 39782
rect 22174 39310 22238 39374
rect 22446 39310 22510 39374
rect 22990 39446 23054 39510
rect 22990 39310 23054 39374
rect 23398 39446 23462 39510
rect 190134 39718 190198 39782
rect 195166 39854 195230 39918
rect 195166 39718 195230 39782
rect 195574 39854 195638 39918
rect 195574 39718 195638 39782
rect 195846 39854 195910 39918
rect 196254 39854 196318 39918
rect 23398 39310 23462 39374
rect 1230 39174 1294 39238
rect 195166 39446 195230 39510
rect 195166 39310 195230 39374
rect 195574 39446 195638 39510
rect 195438 39310 195502 39374
rect 196254 39310 196318 39374
rect 21766 39038 21830 39102
rect 22174 39038 22238 39102
rect 22446 39038 22510 39102
rect 22990 39038 23054 39102
rect 23398 39038 23462 39102
rect 21766 38766 21830 38830
rect 14558 38630 14622 38694
rect 21902 38630 21966 38694
rect 22582 38630 22646 38694
rect 14558 38494 14622 38558
rect 21902 38358 21966 38422
rect 21902 38222 21966 38286
rect 22582 38358 22646 38422
rect 22990 38222 23054 38286
rect 28294 38766 28358 38830
rect 190134 38902 190198 38966
rect 195166 39038 195230 39102
rect 190270 38766 190334 38830
rect 28294 38494 28358 38558
rect 23398 38222 23462 38286
rect 190134 38494 190198 38558
rect 190270 38494 190334 38558
rect 195438 39038 195502 39102
rect 196254 39038 196318 39102
rect 196662 39038 196726 39102
rect 217470 39038 217534 39102
rect 195846 38630 195910 38694
rect 196662 38766 196726 38830
rect 196662 38630 196726 38694
rect 195166 38222 195230 38286
rect 195438 38222 195502 38286
rect 195846 38358 195910 38422
rect 21902 37950 21966 38014
rect 21766 37814 21830 37878
rect 22174 37814 22238 37878
rect 22582 37814 22646 37878
rect 22990 37950 23054 38014
rect 22990 37814 23054 37878
rect 23398 37950 23462 38014
rect 23534 37814 23598 37878
rect 196662 38358 196726 38422
rect 196798 38222 196862 38286
rect 195166 37950 195230 38014
rect 21766 37542 21830 37606
rect 1230 37406 1294 37470
rect 21902 37406 21966 37470
rect 22174 37542 22238 37606
rect 22582 37542 22646 37606
rect 22718 37406 22782 37470
rect 22990 37542 23054 37606
rect 22990 37406 23054 37470
rect 23534 37542 23598 37606
rect 23398 37406 23462 37470
rect 195166 37814 195230 37878
rect 195438 37950 195502 38014
rect 195438 37814 195502 37878
rect 196254 37814 196318 37878
rect 196798 37950 196862 38014
rect 196662 37814 196726 37878
rect 190134 37542 190198 37606
rect 195166 37542 195230 37606
rect 195030 37406 195094 37470
rect 195438 37542 195502 37606
rect 195574 37406 195638 37470
rect 196254 37542 196318 37606
rect 196662 37542 196726 37606
rect 196798 37406 196862 37470
rect 217470 37542 217534 37606
rect 14694 37134 14758 37198
rect 14694 36998 14758 37062
rect 21902 37134 21966 37198
rect 21902 36998 21966 37062
rect 22718 37134 22782 37198
rect 22310 36998 22374 37062
rect 22990 37134 23054 37198
rect 22990 36998 23054 37062
rect 23398 37134 23462 37198
rect 190134 37270 190198 37334
rect 23534 36998 23598 37062
rect 195030 37134 195094 37198
rect 195166 36998 195230 37062
rect 195574 37134 195638 37198
rect 195574 36998 195638 37062
rect 196798 37134 196862 37198
rect 196798 36998 196862 37062
rect 21902 36726 21966 36790
rect 21902 36590 21966 36654
rect 22310 36726 22374 36790
rect 22582 36590 22646 36654
rect 22990 36726 23054 36790
rect 22990 36590 23054 36654
rect 23534 36726 23598 36790
rect 23534 36590 23598 36654
rect 195166 36726 195230 36790
rect 195166 36590 195230 36654
rect 195574 36726 195638 36790
rect 195438 36590 195502 36654
rect 196798 36726 196862 36790
rect 196798 36590 196862 36654
rect 21902 36318 21966 36382
rect 22582 36318 22646 36382
rect 22446 36182 22510 36246
rect 22718 36182 22782 36246
rect 22990 36318 23054 36382
rect 23126 36182 23190 36246
rect 23534 36318 23598 36382
rect 23398 36182 23462 36246
rect 1230 35638 1294 35702
rect 14558 35774 14622 35838
rect 28294 36046 28358 36110
rect 195166 36318 195230 36382
rect 195030 36182 195094 36246
rect 195438 36318 195502 36382
rect 195438 36182 195502 36246
rect 196390 36182 196454 36246
rect 196798 36318 196862 36382
rect 18502 35638 18566 35702
rect 22446 35910 22510 35974
rect 22718 35910 22782 35974
rect 23126 35910 23190 35974
rect 22990 35774 23054 35838
rect 23398 35910 23462 35974
rect 23534 35774 23598 35838
rect 28294 35774 28358 35838
rect 22310 35366 22374 35430
rect 22446 35366 22510 35430
rect 22990 35502 23054 35566
rect 22990 35366 23054 35430
rect 23534 35502 23598 35566
rect 195030 35910 195094 35974
rect 195166 35774 195230 35838
rect 195438 35910 195502 35974
rect 195438 35774 195502 35838
rect 196390 35910 196454 35974
rect 195166 35502 195230 35566
rect 23398 35366 23462 35430
rect 195166 35366 195230 35430
rect 195438 35502 195502 35566
rect 195438 35366 195502 35430
rect 195982 35366 196046 35430
rect 196118 35366 196182 35430
rect 217470 35774 217534 35838
rect 190270 35230 190334 35294
rect 21902 35094 21966 35158
rect 22310 35094 22374 35158
rect 22446 35094 22510 35158
rect 22990 35094 23054 35158
rect 21902 34822 21966 34886
rect 21766 34686 21830 34750
rect 22174 34686 22238 34750
rect 22582 34686 22646 34750
rect 23398 35094 23462 35158
rect 28430 34822 28494 34886
rect 190270 34958 190334 35022
rect 190134 34822 190198 34886
rect 195166 35094 195230 35158
rect 195438 35094 195502 35158
rect 195982 35094 196046 35158
rect 196118 35094 196182 35158
rect 196798 35094 196862 35158
rect 14694 34414 14758 34478
rect 21766 34414 21830 34478
rect 21766 34278 21830 34342
rect 22174 34414 22238 34478
rect 16598 34142 16662 34206
rect 22582 34414 22646 34478
rect 1230 34006 1294 34070
rect 18502 34006 18566 34070
rect 18230 33870 18294 33934
rect 18910 33870 18974 33934
rect 19318 33870 19382 33934
rect 21766 34006 21830 34070
rect 21766 33870 21830 33934
rect 22174 33870 22238 33934
rect 22582 33870 22646 33934
rect 28430 34550 28494 34614
rect 28294 34414 28358 34478
rect 28294 34142 28358 34206
rect 28430 34142 28494 34206
rect 22990 33870 23054 33934
rect 190134 34550 190198 34614
rect 190134 34414 190198 34478
rect 190134 34142 190198 34206
rect 23534 33870 23598 33934
rect 28430 33870 28494 33934
rect 21766 33598 21830 33662
rect 21766 33462 21830 33526
rect 22174 33598 22238 33662
rect 22582 33598 22646 33662
rect 22582 33462 22646 33526
rect 22990 33598 23054 33662
rect 23126 33462 23190 33526
rect 23534 33598 23598 33662
rect 23534 33462 23598 33526
rect 195846 34686 195910 34750
rect 196798 34822 196862 34886
rect 196662 34686 196726 34750
rect 195846 34414 195910 34478
rect 196662 34414 196726 34478
rect 196662 34278 196726 34342
rect 195166 33870 195230 33934
rect 195438 33870 195502 33934
rect 217470 34142 217534 34206
rect 196390 33870 196454 33934
rect 196662 34006 196726 34070
rect 196662 33870 196726 33934
rect 198838 33870 198902 33934
rect 199110 33870 199174 33934
rect 200470 33870 200534 33934
rect 195166 33598 195230 33662
rect 195166 33462 195230 33526
rect 195438 33598 195502 33662
rect 195574 33462 195638 33526
rect 196390 33598 196454 33662
rect 196118 33462 196182 33526
rect 196390 33462 196454 33526
rect 196662 33598 196726 33662
rect 196662 33462 196726 33526
rect 18230 33190 18294 33254
rect 18094 33054 18158 33118
rect 18910 33190 18974 33254
rect 19318 33190 19382 33254
rect 18774 33054 18838 33118
rect 19454 33054 19518 33118
rect 21766 33190 21830 33254
rect 21902 33054 21966 33118
rect 22582 33190 22646 33254
rect 22446 33054 22510 33118
rect 23126 33190 23190 33254
rect 22990 33054 23054 33118
rect 23534 33190 23598 33254
rect 23398 33054 23462 33118
rect 195166 33190 195230 33254
rect 195030 33054 195094 33118
rect 195574 33190 195638 33254
rect 195574 33054 195638 33118
rect 196118 33190 196182 33254
rect 196390 33190 196454 33254
rect 195982 33054 196046 33118
rect 196118 33054 196182 33118
rect 196662 33190 196726 33254
rect 196798 33054 196862 33118
rect 198838 33190 198902 33254
rect 199110 33190 199174 33254
rect 199110 33054 199174 33118
rect 199790 33054 199854 33118
rect 200470 33190 200534 33254
rect 200470 33054 200534 33118
rect 21902 32782 21966 32846
rect 21902 32646 21966 32710
rect 22446 32782 22510 32846
rect 22990 32782 23054 32846
rect 23126 32646 23190 32710
rect 23398 32782 23462 32846
rect 23398 32646 23462 32710
rect 195030 32782 195094 32846
rect 195166 32646 195230 32710
rect 195574 32782 195638 32846
rect 195438 32646 195502 32710
rect 195982 32782 196046 32846
rect 196118 32782 196182 32846
rect 195982 32646 196046 32710
rect 196390 32646 196454 32710
rect 196798 32782 196862 32846
rect 196798 32646 196862 32710
rect 1230 32374 1294 32438
rect 18094 32374 18158 32438
rect 18094 32238 18158 32302
rect 18910 32374 18974 32438
rect 18910 32238 18974 32302
rect 19454 32374 19518 32438
rect 19454 32238 19518 32302
rect 19862 32238 19926 32302
rect 21902 32374 21966 32438
rect 22174 32238 22238 32302
rect 22718 32238 22782 32302
rect 23126 32374 23190 32438
rect 22990 32238 23054 32302
rect 23398 32374 23462 32438
rect 23534 32238 23598 32302
rect 217470 32510 217534 32574
rect 195166 32374 195230 32438
rect 195166 32238 195230 32302
rect 195438 32374 195502 32438
rect 195438 32238 195502 32302
rect 195982 32374 196046 32438
rect 196390 32374 196454 32438
rect 196118 32238 196182 32302
rect 196798 32374 196862 32438
rect 198974 32238 199038 32302
rect 199110 32374 199174 32438
rect 199246 32238 199310 32302
rect 199926 32374 199990 32438
rect 200470 32374 200534 32438
rect 200470 32238 200534 32302
rect 201830 32238 201894 32302
rect 21902 31830 21966 31894
rect 22174 31966 22238 32030
rect 22718 31966 22782 32030
rect 22310 31830 22374 31894
rect 22446 31830 22510 31894
rect 22990 31966 23054 32030
rect 23126 31830 23190 31894
rect 23534 31966 23598 32030
rect 23398 31830 23462 31894
rect 195166 31966 195230 32030
rect 195030 31830 195094 31894
rect 195438 31966 195502 32030
rect 195438 31830 195502 31894
rect 196118 31966 196182 32030
rect 196390 31830 196454 31894
rect 196662 31830 196726 31894
rect 16598 31558 16662 31622
rect 18094 31558 18158 31622
rect 18910 31558 18974 31622
rect 19454 31558 19518 31622
rect 18910 31422 18974 31486
rect 19318 31422 19382 31486
rect 19862 31558 19926 31622
rect 21902 31558 21966 31622
rect 22310 31558 22374 31622
rect 22446 31558 22510 31622
rect 22582 31422 22646 31486
rect 23126 31558 23190 31622
rect 22990 31422 23054 31486
rect 23398 31558 23462 31622
rect 23534 31422 23598 31486
rect 195030 31558 195094 31622
rect 28566 31286 28630 31350
rect 21766 31150 21830 31214
rect 22582 31150 22646 31214
rect 22990 31150 23054 31214
rect 22990 31014 23054 31078
rect 23534 31150 23598 31214
rect 23534 31014 23598 31078
rect 28566 31014 28630 31078
rect 21766 30878 21830 30942
rect 1230 30742 1294 30806
rect 22038 30606 22102 30670
rect 22174 30606 22238 30670
rect 22582 30606 22646 30670
rect 22990 30742 23054 30806
rect 2109 30352 2173 30356
rect 2109 30296 2113 30352
rect 2113 30296 2169 30352
rect 2169 30296 2173 30352
rect 2109 30292 2173 30296
rect 21766 30334 21830 30398
rect 22174 30334 22238 30398
rect 22038 30198 22102 30262
rect 22582 30334 22646 30398
rect 23534 30742 23598 30806
rect 195166 31422 195230 31486
rect 195438 31558 195502 31622
rect 195438 31422 195502 31486
rect 195846 31422 195910 31486
rect 196390 31558 196454 31622
rect 196254 31422 196318 31486
rect 196662 31558 196726 31622
rect 198974 31558 199038 31622
rect 198838 31422 198902 31486
rect 199246 31558 199310 31622
rect 199110 31422 199174 31486
rect 200470 31558 200534 31622
rect 199790 31422 199854 31486
rect 201830 31558 201894 31622
rect 190134 31286 190198 31350
rect 190134 31014 190198 31078
rect 195166 31150 195230 31214
rect 195030 31014 195094 31078
rect 195438 31150 195502 31214
rect 195574 31014 195638 31078
rect 195846 31150 195910 31214
rect 196254 31150 196318 31214
rect 196662 31150 196726 31214
rect 198838 31014 198902 31078
rect 196662 30878 196726 30942
rect 18230 29926 18294 29990
rect 18910 30062 18974 30126
rect 18774 29926 18838 29990
rect 19318 30062 19382 30126
rect 19318 29926 19382 29990
rect 21766 30062 21830 30126
rect 19862 29926 19926 29990
rect 21902 29926 21966 29990
rect 22446 29926 22510 29990
rect 23126 29926 23190 29990
rect 23398 29926 23462 29990
rect 190134 30470 190198 30534
rect 190134 30198 190198 30262
rect 195030 30742 195094 30806
rect 195574 30742 195638 30806
rect 196254 30606 196318 30670
rect 217470 30606 217534 30670
rect 550 29654 614 29718
rect 21902 29654 21966 29718
rect 21902 29518 21966 29582
rect 22446 29654 22510 29718
rect 22310 29518 22374 29582
rect 22718 29518 22782 29582
rect 23126 29654 23190 29718
rect 22990 29518 23054 29582
rect 23398 29654 23462 29718
rect 23398 29518 23462 29582
rect 195166 29926 195230 29990
rect 195438 29926 195502 29990
rect 196254 30334 196318 30398
rect 196662 30334 196726 30398
rect 195846 29926 195910 29990
rect 196662 30062 196726 30126
rect 196798 29926 196862 29990
rect 199110 30062 199174 30126
rect 199110 29926 199174 29990
rect 199382 29926 199446 29990
rect 199790 30062 199854 30126
rect 199926 29926 199990 29990
rect 200606 29926 200670 29990
rect 195166 29654 195230 29718
rect 195166 29518 195230 29582
rect 195438 29654 195502 29718
rect 195438 29518 195502 29582
rect 195846 29654 195910 29718
rect 195846 29518 195910 29582
rect 196798 29654 196862 29718
rect 199110 29654 199174 29718
rect 196662 29518 196726 29582
rect 18230 29246 18294 29310
rect 1230 29110 1294 29174
rect 18230 29110 18294 29174
rect 18910 29246 18974 29310
rect 19318 29246 19382 29310
rect 18910 29110 18974 29174
rect 19454 29110 19518 29174
rect 19862 29246 19926 29310
rect 21902 29246 21966 29310
rect 21766 29110 21830 29174
rect 22310 29246 22374 29310
rect 22718 29246 22782 29310
rect 22582 29110 22646 29174
rect 22990 29246 23054 29310
rect 23126 29110 23190 29174
rect 23398 29246 23462 29310
rect 23534 29110 23598 29174
rect 195166 29246 195230 29310
rect 195166 29110 195230 29174
rect 195438 29246 195502 29310
rect 195438 29110 195502 29174
rect 195846 29246 195910 29310
rect 195846 29110 195910 29174
rect 196254 29110 196318 29174
rect 196662 29246 196726 29310
rect 196662 29110 196726 29174
rect 198838 29110 198902 29174
rect 199382 29246 199446 29310
rect 199246 29110 199310 29174
rect 199790 29246 199854 29310
rect 200606 29246 200670 29310
rect 200470 29110 200534 29174
rect 217470 28974 217534 29038
rect 21766 28838 21830 28902
rect 21902 28702 21966 28766
rect 22310 28702 22374 28766
rect 22582 28838 22646 28902
rect 22718 28702 22782 28766
rect 23126 28838 23190 28902
rect 22990 28702 23054 28766
rect 23534 28838 23598 28902
rect 23398 28702 23462 28766
rect 195166 28838 195230 28902
rect 195030 28702 195094 28766
rect 195438 28838 195502 28902
rect 195438 28702 195502 28766
rect 195846 28838 195910 28902
rect 196254 28838 196318 28902
rect 196662 28838 196726 28902
rect 196798 28702 196862 28766
rect 18910 28566 18974 28630
rect 18230 28430 18294 28494
rect 18094 28294 18158 28358
rect 18366 28294 18430 28358
rect 19454 28430 19518 28494
rect 19046 28294 19110 28358
rect 19318 28294 19382 28358
rect 19454 28294 19518 28358
rect 19862 28294 19926 28358
rect 21902 28430 21966 28494
rect 21902 28294 21966 28358
rect 22310 28430 22374 28494
rect 22718 28430 22782 28494
rect 22446 28294 22510 28358
rect 22990 28430 23054 28494
rect 22990 28294 23054 28358
rect 23398 28430 23462 28494
rect 23398 28294 23462 28358
rect 195030 28430 195094 28494
rect 195166 28294 195230 28358
rect 195438 28430 195502 28494
rect 195438 28294 195502 28358
rect 196390 28294 196454 28358
rect 196798 28430 196862 28494
rect 196798 28294 196862 28358
rect 198838 28430 198902 28494
rect 198974 28294 199038 28358
rect 199246 28430 199310 28494
rect 199382 28294 199446 28358
rect 200470 28430 200534 28494
rect 200470 28294 200534 28358
rect 1910 28022 1974 28086
rect 18366 28022 18430 28086
rect 19318 28022 19382 28086
rect 21902 28022 21966 28086
rect 21766 27886 21830 27950
rect 22446 28022 22510 28086
rect 22174 27886 22238 27950
rect 22582 27886 22646 27950
rect 22990 28022 23054 28086
rect 23126 27886 23190 27950
rect 23398 28022 23462 28086
rect 23398 27886 23462 27950
rect 195166 28022 195230 28086
rect 195166 27886 195230 27950
rect 195438 28022 195502 28086
rect 195438 27886 195502 27950
rect 195982 27886 196046 27950
rect 196390 28022 196454 28086
rect 196798 28022 196862 28086
rect 196798 27886 196862 27950
rect 1230 27478 1294 27542
rect 1910 27478 1974 27542
rect 18094 27614 18158 27678
rect 19046 27614 19110 27678
rect 19454 27614 19518 27678
rect 19862 27614 19926 27678
rect 19454 27478 19518 27542
rect 19726 27478 19790 27542
rect 21766 27614 21830 27678
rect 22174 27614 22238 27678
rect 22582 27614 22646 27678
rect 22310 27478 22374 27542
rect 23126 27614 23190 27678
rect 23126 27478 23190 27542
rect 23398 27614 23462 27678
rect 23398 27478 23462 27542
rect 195166 27614 195230 27678
rect 195030 27478 195094 27542
rect 195438 27614 195502 27678
rect 195438 27478 195502 27542
rect 195982 27614 196046 27678
rect 196390 27478 196454 27542
rect 196798 27614 196862 27678
rect 198974 27614 199038 27678
rect 199382 27614 199446 27678
rect 200470 27614 200534 27678
rect 200470 27478 200534 27542
rect 21902 27206 21966 27270
rect 22310 27206 22374 27270
rect 23126 27206 23190 27270
rect 23126 27070 23190 27134
rect 23398 27206 23462 27270
rect 23534 27070 23598 27134
rect 21902 26934 21966 26998
rect 550 26662 614 26726
rect 22174 26662 22238 26726
rect 22446 26662 22510 26726
rect 23126 26798 23190 26862
rect 23534 26798 23598 26862
rect 195030 27206 195094 27270
rect 195166 27070 195230 27134
rect 195438 27206 195502 27270
rect 195574 27070 195638 27134
rect 196390 27206 196454 27270
rect 198974 27342 199038 27406
rect 217470 27342 217534 27406
rect 196798 27206 196862 27270
rect 21902 26390 21966 26454
rect 22174 26390 22238 26454
rect 22446 26390 22510 26454
rect 18638 25982 18702 26046
rect 19454 26118 19518 26182
rect 19454 25846 19518 25910
rect 19726 26118 19790 26182
rect 21902 26118 21966 26182
rect 21766 25982 21830 26046
rect 22174 25982 22238 26046
rect 22582 25982 22646 26046
rect 28566 26526 28630 26590
rect 28566 26254 28630 26318
rect 19726 25846 19790 25910
rect 28430 26118 28494 26182
rect 195166 26798 195230 26862
rect 190270 26526 190334 26590
rect 190270 26254 190334 26318
rect 190270 26118 190334 26182
rect 21766 25710 21830 25774
rect 1230 25574 1294 25638
rect 18774 25574 18838 25638
rect 19318 25574 19382 25638
rect 21902 25574 21966 25638
rect 22174 25710 22238 25774
rect 19726 25438 19790 25502
rect 22582 25710 22646 25774
rect 23126 25574 23190 25638
rect 23398 25574 23462 25638
rect 28430 25846 28494 25910
rect 28294 25710 28358 25774
rect 190270 25846 190334 25910
rect 195574 26798 195638 26862
rect 196390 26662 196454 26726
rect 196798 26934 196862 26998
rect 196390 26390 196454 26454
rect 196798 26390 196862 26454
rect 196254 25982 196318 26046
rect 196798 26118 196862 26182
rect 196662 25982 196726 26046
rect 198974 26118 199038 26182
rect 199654 25982 199718 26046
rect 200470 26118 200534 26182
rect 200198 25982 200262 26046
rect 201286 25982 201350 26046
rect 199382 25846 199446 25910
rect 195030 25574 195094 25638
rect 195438 25574 195502 25638
rect 28294 25438 28358 25502
rect 17142 25166 17206 25230
rect 18638 25302 18702 25366
rect 18774 25302 18838 25366
rect 19318 25302 19382 25366
rect 19454 25302 19518 25366
rect 17550 25166 17614 25230
rect 21902 25302 21966 25366
rect 21902 25166 21966 25230
rect 23126 25302 23190 25366
rect 23398 25302 23462 25366
rect 196254 25710 196318 25774
rect 196662 25710 196726 25774
rect 196662 25574 196726 25638
rect 217470 25710 217534 25774
rect 23398 25166 23462 25230
rect 195030 25302 195094 25366
rect 195030 25166 195094 25230
rect 195438 25302 195502 25366
rect 196662 25302 196726 25366
rect 199382 25302 199446 25366
rect 199382 25166 199446 25230
rect 199654 25302 199718 25366
rect 200198 25302 200262 25366
rect 199926 25166 199990 25230
rect 201286 25302 201350 25366
rect 201150 25166 201214 25230
rect 204006 25166 204070 25230
rect 23398 24758 23462 24822
rect 23126 24486 23190 24550
rect 199382 24894 199446 24958
rect 199926 24894 199990 24958
rect 204006 24894 204070 24958
rect 204142 24758 204206 24822
rect 29926 24622 29990 24686
rect 29382 24350 29446 24414
rect 30606 24350 30670 24414
rect 32238 24214 32302 24278
rect 32918 24214 32982 24278
rect 33462 24214 33526 24278
rect 34142 24214 34206 24278
rect 35502 24214 35566 24278
rect 39310 24350 39374 24414
rect 37134 24214 37198 24278
rect 38494 24214 38558 24278
rect 40942 24214 41006 24278
rect 41622 24214 41686 24278
rect 42846 24214 42910 24278
rect 44614 24214 44678 24278
rect 45430 24214 45494 24278
rect 47198 24214 47262 24278
rect 48014 24214 48078 24278
rect 49646 24214 49710 24278
rect 50462 24214 50526 24278
rect 50870 24214 50934 24278
rect 51686 24214 51750 24278
rect 52910 24214 52974 24278
rect 54678 24214 54742 24278
rect 55358 24214 55422 24278
rect 58078 24350 58142 24414
rect 56582 24214 56646 24278
rect 59710 24214 59774 24278
rect 60390 24214 60454 24278
rect 61614 24214 61678 24278
rect 62158 24214 62222 24278
rect 62838 24214 62902 24278
rect 64062 24214 64126 24278
rect 66646 24214 66710 24278
rect 67870 24214 67934 24278
rect 68414 24214 68478 24278
rect 69094 24214 69158 24278
rect 69638 24214 69702 24278
rect 70318 24214 70382 24278
rect 70862 24214 70926 24278
rect 71678 24214 71742 24278
rect 73446 24214 73510 24278
rect 74670 24214 74734 24278
rect 75214 24214 75278 24278
rect 75894 24214 75958 24278
rect 76574 24214 76638 24278
rect 78342 24214 78406 24278
rect 79566 24214 79630 24278
rect 80518 24214 80582 24278
rect 82014 24214 82078 24278
rect 83374 24214 83438 24278
rect 84598 24214 84662 24278
rect 85686 24214 85750 24278
rect 86502 24214 86566 24278
rect 88406 24214 88470 24278
rect 89086 24214 89150 24278
rect 89766 24214 89830 24278
rect 92078 24214 92142 24278
rect 94662 24214 94726 24278
rect 95342 24214 95406 24278
rect 95750 24214 95814 24278
rect 97110 24214 97174 24278
rect 97790 24214 97854 24278
rect 100782 24214 100846 24278
rect 101598 24214 101662 24278
rect 102142 24214 102206 24278
rect 103366 24214 103430 24278
rect 104046 24214 104110 24278
rect 104590 24214 104654 24278
rect 105270 24214 105334 24278
rect 109622 24214 109686 24278
rect 110302 24214 110366 24278
rect 110846 24214 110910 24278
rect 111526 24214 111590 24278
rect 112750 24214 112814 24278
rect 114246 24350 114310 24414
rect 113294 24214 113358 24278
rect 115334 24214 115398 24278
rect 117102 24214 117166 24278
rect 117646 24214 117710 24278
rect 119006 24214 119070 24278
rect 120230 24214 120294 24278
rect 121998 24214 122062 24278
rect 122950 24214 123014 24278
rect 123902 24214 123966 24278
rect 124446 24214 124510 24278
rect 125806 24214 125870 24278
rect 127030 24214 127094 24278
rect 128934 24214 128998 24278
rect 130294 24214 130358 24278
rect 131654 24214 131718 24278
rect 133286 24214 133350 24278
rect 134510 24214 134574 24278
rect 135190 24214 135254 24278
rect 136686 24350 136750 24414
rect 135734 24214 135798 24278
rect 138182 24214 138246 24278
rect 139542 24214 139606 24278
rect 140222 24214 140286 24278
rect 141854 24214 141918 24278
rect 145390 24350 145454 24414
rect 143214 24214 143278 24278
rect 144030 24214 144094 24278
rect 146478 24214 146542 24278
rect 147022 24214 147086 24278
rect 147702 24214 147766 24278
rect 149062 24214 149126 24278
rect 150422 24214 150486 24278
rect 152054 24214 152118 24278
rect 152734 24214 152798 24278
rect 153278 24214 153342 24278
rect 154502 24214 154566 24278
rect 155182 24214 155246 24278
rect 155726 24214 155790 24278
rect 156950 24214 157014 24278
rect 158174 24214 158238 24278
rect 159534 24214 159598 24278
rect 160214 24214 160278 24278
rect 160758 24214 160822 24278
rect 161438 24214 161502 24278
rect 163206 24214 163270 24278
rect 164430 24214 164494 24278
rect 165382 24214 165446 24278
rect 166878 24214 166942 24278
rect 168238 24214 168302 24278
rect 169462 24214 169526 24278
rect 170550 24214 170614 24278
rect 171366 24214 171430 24278
rect 171910 24214 171974 24278
rect 173270 24214 173334 24278
rect 175174 24214 175238 24278
rect 179118 24350 179182 24414
rect 176942 24214 177006 24278
rect 178166 24214 178230 24278
rect 180206 24214 180270 24278
rect 181430 24214 181494 24278
rect 183198 24214 183262 24278
rect 185646 24214 185710 24278
rect 186462 24214 186526 24278
rect 195030 24350 195094 24414
rect 187686 24214 187750 24278
rect 188910 24214 188974 24278
rect 1230 23942 1294 24006
rect 217470 24078 217534 24142
rect 550 23806 614 23870
rect 17142 23942 17206 24006
rect 15238 23806 15302 23870
rect 29382 23670 29446 23734
rect 29654 23534 29718 23598
rect 30606 23670 30670 23734
rect 32238 23670 32302 23734
rect 32918 23670 32982 23734
rect 33462 23670 33526 23734
rect 34142 23670 34206 23734
rect 34686 23534 34750 23598
rect 35502 23670 35566 23734
rect 37134 23670 37198 23734
rect 38494 23670 38558 23734
rect 39310 23670 39374 23734
rect 39718 23534 39782 23598
rect 40942 23670 41006 23734
rect 41622 23670 41686 23734
rect 42846 23670 42910 23734
rect 44614 23670 44678 23734
rect 45430 23670 45494 23734
rect 45430 23534 45494 23598
rect 47198 23670 47262 23734
rect 48014 23670 48078 23734
rect 49646 23670 49710 23734
rect 49374 23534 49438 23598
rect 50462 23670 50526 23734
rect 50870 23670 50934 23734
rect 51686 23670 51750 23734
rect 52910 23670 52974 23734
rect 54678 23670 54742 23734
rect 54270 23534 54334 23598
rect 55358 23670 55422 23734
rect 56582 23670 56646 23734
rect 58078 23670 58142 23734
rect 59710 23670 59774 23734
rect 60390 23670 60454 23734
rect 60798 23534 60862 23598
rect 61614 23670 61678 23734
rect 62158 23670 62222 23734
rect 62838 23670 62902 23734
rect 64062 23670 64126 23734
rect 64606 23534 64670 23598
rect 66646 23670 66710 23734
rect 67870 23670 67934 23734
rect 68414 23670 68478 23734
rect 69094 23670 69158 23734
rect 69638 23670 69702 23734
rect 70318 23670 70382 23734
rect 70862 23670 70926 23734
rect 70318 23534 70382 23598
rect 71678 23670 71742 23734
rect 73446 23670 73510 23734
rect 74670 23670 74734 23734
rect 75214 23670 75278 23734
rect 75894 23670 75958 23734
rect 75350 23534 75414 23598
rect 76574 23670 76638 23734
rect 78342 23670 78406 23734
rect 79566 23670 79630 23734
rect 80518 23670 80582 23734
rect 82014 23670 82078 23734
rect 83374 23670 83438 23734
rect 84598 23670 84662 23734
rect 84190 23534 84254 23598
rect 85686 23670 85750 23734
rect 86502 23670 86566 23734
rect 88406 23670 88470 23734
rect 89086 23670 89150 23734
rect 89766 23670 89830 23734
rect 89630 23534 89694 23598
rect 92078 23670 92142 23734
rect 94662 23670 94726 23734
rect 95342 23670 95406 23734
rect 95750 23670 95814 23734
rect 95342 23534 95406 23598
rect 97110 23670 97174 23734
rect 97790 23670 97854 23734
rect 99558 23534 99622 23598
rect 100782 23670 100846 23734
rect 101598 23670 101662 23734
rect 102142 23670 102206 23734
rect 103366 23670 103430 23734
rect 104046 23670 104110 23734
rect 104590 23670 104654 23734
rect 105270 23670 105334 23734
rect 105270 23534 105334 23598
rect 109622 23670 109686 23734
rect 110302 23670 110366 23734
rect 110846 23670 110910 23734
rect 110302 23534 110366 23598
rect 111526 23670 111590 23734
rect 112750 23670 112814 23734
rect 113294 23670 113358 23734
rect 114246 23670 114310 23734
rect 114518 23534 114582 23598
rect 115334 23670 115398 23734
rect 117102 23670 117166 23734
rect 117646 23670 117710 23734
rect 119006 23670 119070 23734
rect 119278 23534 119342 23598
rect 120230 23670 120294 23734
rect 121998 23670 122062 23734
rect 122950 23670 123014 23734
rect 123902 23670 123966 23734
rect 124446 23670 124510 23734
rect 124582 23534 124646 23598
rect 125806 23670 125870 23734
rect 127030 23670 127094 23734
rect 128934 23670 128998 23734
rect 130294 23670 130358 23734
rect 130294 23534 130358 23598
rect 131654 23670 131718 23734
rect 133286 23670 133350 23734
rect 134510 23670 134574 23734
rect 134102 23534 134166 23598
rect 135190 23670 135254 23734
rect 135734 23670 135798 23734
rect 136686 23670 136750 23734
rect 138182 23670 138246 23734
rect 139542 23670 139606 23734
rect 139134 23534 139198 23598
rect 140222 23670 140286 23734
rect 141854 23670 141918 23734
rect 143214 23670 143278 23734
rect 144030 23670 144094 23734
rect 145390 23670 145454 23734
rect 145662 23534 145726 23598
rect 146478 23670 146542 23734
rect 147022 23670 147086 23734
rect 147702 23670 147766 23734
rect 149062 23670 149126 23734
rect 149470 23534 149534 23598
rect 150422 23670 150486 23734
rect 152054 23670 152118 23734
rect 152734 23670 152798 23734
rect 153278 23670 153342 23734
rect 154502 23670 154566 23734
rect 155182 23670 155246 23734
rect 155726 23670 155790 23734
rect 155182 23534 155246 23598
rect 156950 23670 157014 23734
rect 158174 23670 158238 23734
rect 159534 23670 159598 23734
rect 160214 23670 160278 23734
rect 160758 23670 160822 23734
rect 160214 23534 160278 23598
rect 161438 23670 161502 23734
rect 163206 23670 163270 23734
rect 164430 23670 164494 23734
rect 164158 23534 164222 23598
rect 165382 23670 165446 23734
rect 166878 23670 166942 23734
rect 168238 23670 168302 23734
rect 169462 23670 169526 23734
rect 170550 23670 170614 23734
rect 170142 23534 170206 23598
rect 171366 23670 171430 23734
rect 171910 23670 171974 23734
rect 173270 23670 173334 23734
rect 175174 23670 175238 23734
rect 174494 23534 174558 23598
rect 176942 23670 177006 23734
rect 178166 23670 178230 23734
rect 179118 23670 179182 23734
rect 180206 23670 180270 23734
rect 180206 23534 180270 23598
rect 181430 23670 181494 23734
rect 183198 23670 183262 23734
rect 184422 23534 184486 23598
rect 185646 23670 185710 23734
rect 186462 23670 186526 23734
rect 187686 23670 187750 23734
rect 188910 23670 188974 23734
rect 201150 23534 201214 23598
rect 204006 23262 204070 23326
rect 2109 22885 2173 22949
rect 17550 22582 17614 22646
rect 15102 22446 15166 22510
rect 1230 22310 1294 22374
rect 21902 22310 21966 22374
rect 217470 22310 217534 22374
rect 21766 22174 21830 22238
rect 29926 22174 29990 22238
rect 29926 22038 29990 22102
rect 35094 22038 35158 22102
rect 39990 22038 40054 22102
rect 44886 22038 44950 22102
rect 50054 22038 50118 22102
rect 55086 22038 55150 22102
rect 59710 22038 59774 22102
rect 64878 22038 64942 22102
rect 70046 22038 70110 22102
rect 75078 22038 75142 22102
rect 79838 22038 79902 22102
rect 85006 22038 85070 22102
rect 90038 22038 90102 22102
rect 94798 22038 94862 22102
rect 99966 22038 100030 22102
rect 104998 22038 105062 22102
rect 110030 22038 110094 22102
rect 114790 22038 114854 22102
rect 119958 22038 120022 22102
rect 124990 22038 125054 22102
rect 129750 22038 129814 22102
rect 134918 22038 134982 22102
rect 139950 22038 140014 22102
rect 144846 22038 144910 22102
rect 149742 22038 149806 22102
rect 154910 22038 154974 22102
rect 159942 22038 160006 22102
rect 164838 22038 164902 22102
rect 169870 22038 169934 22102
rect 174902 22038 174966 22102
rect 179662 22038 179726 22102
rect 184694 22038 184758 22102
rect 204142 22038 204206 22102
rect 204142 21902 204206 21966
rect 550 20950 614 21014
rect 15238 21086 15302 21150
rect 15238 20950 15302 21014
rect 23126 20950 23190 21014
rect 20542 20814 20606 20878
rect 1230 20678 1294 20742
rect 204006 20678 204070 20742
rect 2726 20542 2790 20606
rect 204006 20542 204070 20606
rect 217470 20542 217534 20606
rect 2726 19726 2790 19790
rect 15102 19726 15166 19790
rect 15102 19590 15166 19654
rect 29926 19590 29990 19654
rect 30062 19590 30126 19654
rect 34958 19590 35022 19654
rect 35094 19590 35158 19654
rect 39854 19590 39918 19654
rect 39990 19590 40054 19654
rect 44886 19590 44950 19654
rect 45022 19590 45086 19654
rect 49918 19590 49982 19654
rect 50054 19590 50118 19654
rect 54950 19590 55014 19654
rect 55086 19590 55150 19654
rect 59710 19590 59774 19654
rect 59982 19590 60046 19654
rect 64878 19590 64942 19654
rect 65014 19590 65078 19654
rect 69910 19590 69974 19654
rect 70046 19590 70110 19654
rect 74942 19590 75006 19654
rect 75078 19590 75142 19654
rect 79838 19590 79902 19654
rect 79974 19590 80038 19654
rect 84870 19590 84934 19654
rect 85006 19590 85070 19654
rect 89902 19590 89966 19654
rect 90038 19590 90102 19654
rect 94798 19590 94862 19654
rect 94934 19590 94998 19654
rect 99830 19590 99894 19654
rect 99966 19590 100030 19654
rect 104862 19590 104926 19654
rect 104998 19590 105062 19654
rect 109894 19590 109958 19654
rect 110030 19590 110094 19654
rect 114790 19590 114854 19654
rect 114926 19590 114990 19654
rect 119822 19590 119886 19654
rect 119958 19590 120022 19654
rect 124854 19590 124918 19654
rect 124990 19590 125054 19654
rect 129750 19590 129814 19654
rect 129886 19590 129950 19654
rect 134782 19590 134846 19654
rect 134918 19590 134982 19654
rect 139814 19590 139878 19654
rect 139950 19590 140014 19654
rect 144710 19590 144774 19654
rect 144846 19590 144910 19654
rect 149742 19590 149806 19654
rect 149878 19590 149942 19654
rect 154774 19590 154838 19654
rect 154910 19590 154974 19654
rect 159806 19590 159870 19654
rect 159942 19590 160006 19654
rect 164702 19590 164766 19654
rect 164838 19590 164902 19654
rect 169734 19590 169798 19654
rect 169870 19590 169934 19654
rect 174766 19590 174830 19654
rect 174902 19590 174966 19654
rect 179662 19590 179726 19654
rect 179798 19590 179862 19654
rect 184558 19590 184622 19654
rect 184694 19590 184758 19654
rect 21766 19454 21830 19518
rect 21766 19318 21830 19382
rect 204142 19182 204206 19246
rect 204278 19046 204342 19110
rect 217470 19046 217534 19110
rect 1230 18910 1294 18974
rect 29654 18910 29718 18974
rect 29790 18774 29854 18838
rect 34686 18910 34750 18974
rect 34686 18774 34750 18838
rect 39718 18910 39782 18974
rect 39718 18774 39782 18838
rect 45430 18910 45494 18974
rect 49374 18910 49438 18974
rect 54270 18910 54334 18974
rect 44750 18774 44814 18838
rect 49646 18774 49710 18838
rect 54678 18774 54742 18838
rect 60798 18910 60862 18974
rect 64606 18910 64670 18974
rect 59710 18774 59774 18838
rect 64878 18774 64942 18838
rect 70318 18910 70382 18974
rect 75350 18910 75414 18974
rect 69774 18774 69838 18838
rect 74670 18774 74734 18838
rect 84190 18910 84254 18974
rect 79702 18774 79766 18838
rect 84734 18774 84798 18838
rect 89630 18910 89694 18974
rect 89766 18774 89830 18838
rect 95342 18910 95406 18974
rect 99558 18910 99622 18974
rect 94798 18774 94862 18838
rect 99694 18774 99758 18838
rect 105270 18910 105334 18974
rect 110302 18910 110366 18974
rect 114518 18910 114582 18974
rect 119278 18910 119342 18974
rect 104590 18774 104654 18838
rect 109758 18774 109822 18838
rect 114790 18774 114854 18838
rect 119550 18774 119614 18838
rect 124582 18910 124646 18974
rect 124582 18774 124646 18838
rect 130294 18910 130358 18974
rect 134102 18910 134166 18974
rect 139134 18910 139198 18974
rect 129614 18774 129678 18838
rect 134510 18774 134574 18838
rect 139542 18774 139606 18838
rect 145662 18910 145726 18974
rect 149470 18910 149534 18974
rect 144574 18774 144638 18838
rect 149606 18774 149670 18838
rect 155182 18910 155246 18974
rect 160214 18910 160278 18974
rect 164158 18910 164222 18974
rect 154638 18774 154702 18838
rect 159534 18774 159598 18838
rect 164566 18774 164630 18838
rect 170142 18910 170206 18974
rect 174494 18910 174558 18974
rect 169598 18774 169662 18838
rect 174630 18774 174694 18838
rect 180206 18910 180270 18974
rect 184422 18910 184486 18974
rect 179662 18774 179726 18838
rect 184422 18774 184486 18838
rect 550 18366 614 18430
rect 15238 18366 15302 18430
rect 15238 18094 15302 18158
rect 20542 18094 20606 18158
rect 29790 18094 29854 18158
rect 34686 18094 34750 18158
rect 20406 17958 20470 18022
rect 29926 17958 29990 18022
rect 34822 17958 34886 18022
rect 39718 18094 39782 18158
rect 44750 18094 44814 18158
rect 49646 18094 49710 18158
rect 54678 18094 54742 18158
rect 59710 18094 59774 18158
rect 39718 17958 39782 18022
rect 44886 17958 44950 18022
rect 49782 17958 49846 18022
rect 54814 17958 54878 18022
rect 59846 17958 59910 18022
rect 64878 18094 64942 18158
rect 69774 18094 69838 18158
rect 74670 18094 74734 18158
rect 79702 18094 79766 18158
rect 84734 18094 84798 18158
rect 89766 18094 89830 18158
rect 94798 18094 94862 18158
rect 64742 17958 64806 18022
rect 69774 17958 69838 18022
rect 74806 17958 74870 18022
rect 79838 17958 79902 18022
rect 84734 17958 84798 18022
rect 89766 17958 89830 18022
rect 94798 17958 94862 18022
rect 99694 18094 99758 18158
rect 104590 18094 104654 18158
rect 109758 18094 109822 18158
rect 114790 18094 114854 18158
rect 119550 18094 119614 18158
rect 124582 18094 124646 18158
rect 129614 18094 129678 18158
rect 134510 18094 134574 18158
rect 139542 18094 139606 18158
rect 144574 18094 144638 18158
rect 149606 18094 149670 18158
rect 154638 18094 154702 18158
rect 159534 18094 159598 18158
rect 99558 17958 99622 18022
rect 104726 17958 104790 18022
rect 109758 17958 109822 18022
rect 114790 17958 114854 18022
rect 119686 17958 119750 18022
rect 124718 17958 124782 18022
rect 129750 17958 129814 18022
rect 134646 17958 134710 18022
rect 139678 17958 139742 18022
rect 144710 17958 144774 18022
rect 149742 17958 149806 18022
rect 154638 17958 154702 18022
rect 159670 17958 159734 18022
rect 164566 18094 164630 18158
rect 169598 18094 169662 18158
rect 174630 18094 174694 18158
rect 179662 18094 179726 18158
rect 164566 17958 164630 18022
rect 169598 17958 169662 18022
rect 174630 17958 174694 18022
rect 179662 17958 179726 18022
rect 184422 18094 184486 18158
rect 184422 17958 184486 18022
rect 30062 17822 30126 17886
rect 28974 17550 29038 17614
rect 34958 17822 35022 17886
rect 34550 17550 34614 17614
rect 34958 17550 35022 17614
rect 39446 17550 39510 17614
rect 39854 17822 39918 17886
rect 45022 17822 45086 17886
rect 39854 17550 39918 17614
rect 44206 17550 44270 17614
rect 49918 17822 49982 17886
rect 49510 17550 49574 17614
rect 49918 17550 49982 17614
rect 54950 17822 55014 17886
rect 54542 17550 54606 17614
rect 59982 17822 60046 17886
rect 54950 17550 55014 17614
rect 59302 17550 59366 17614
rect 64470 17550 64534 17614
rect 65014 17822 65078 17886
rect 64878 17550 64942 17614
rect 69910 17822 69974 17886
rect 69502 17550 69566 17614
rect 74942 17822 75006 17886
rect 69910 17550 69974 17614
rect 74398 17550 74462 17614
rect 79974 17822 80038 17886
rect 79430 17550 79494 17614
rect 84870 17822 84934 17886
rect 84326 17550 84390 17614
rect 89902 17822 89966 17886
rect 84870 17550 84934 17614
rect 89358 17550 89422 17614
rect 94934 17822 94998 17886
rect 94390 17550 94454 17614
rect 99830 17822 99894 17886
rect 99422 17550 99486 17614
rect 99694 17550 99758 17614
rect 104862 17822 104926 17886
rect 104318 17550 104382 17614
rect 109894 17822 109958 17886
rect 109078 17550 109142 17614
rect 114926 17822 114990 17886
rect 114382 17550 114446 17614
rect 119822 17822 119886 17886
rect 119278 17550 119342 17614
rect 124854 17822 124918 17886
rect 119822 17550 119886 17614
rect 124310 17550 124374 17614
rect 129886 17822 129950 17886
rect 129342 17550 129406 17614
rect 134782 17822 134846 17886
rect 134374 17550 134438 17614
rect 134782 17550 134846 17614
rect 139814 17822 139878 17886
rect 139270 17550 139334 17614
rect 144846 17822 144910 17886
rect 144302 17550 144366 17614
rect 149878 17822 149942 17886
rect 149062 17550 149126 17614
rect 154774 17822 154838 17886
rect 154230 17550 154294 17614
rect 159806 17822 159870 17886
rect 154774 17550 154838 17614
rect 159262 17550 159326 17614
rect 164294 17550 164358 17614
rect 164702 17822 164766 17886
rect 164702 17550 164766 17614
rect 169734 17822 169798 17886
rect 169190 17550 169254 17614
rect 174766 17822 174830 17886
rect 169734 17550 169798 17614
rect 174222 17550 174286 17614
rect 179798 17822 179862 17886
rect 179254 17550 179318 17614
rect 184558 17822 184622 17886
rect 204006 17822 204070 17886
rect 204142 17686 204206 17750
rect 184286 17550 184350 17614
rect 184558 17550 184622 17614
rect 29790 17414 29854 17478
rect 44750 17414 44814 17478
rect 59710 17414 59774 17478
rect 74670 17414 74734 17478
rect 79702 17414 79766 17478
rect 89630 17414 89694 17478
rect 94662 17414 94726 17478
rect 104590 17414 104654 17478
rect 109622 17414 109686 17478
rect 114654 17414 114718 17478
rect 124582 17414 124646 17478
rect 129614 17414 129678 17478
rect 139542 17414 139606 17478
rect 144574 17414 144638 17478
rect 149606 17414 149670 17478
rect 159534 17414 159598 17478
rect 174494 17414 174558 17478
rect 179526 17414 179590 17478
rect 1230 17278 1294 17342
rect 49918 17142 49982 17206
rect 134782 17142 134846 17206
rect 217470 17142 217534 17206
rect 29790 17006 29854 17070
rect 15102 16870 15166 16934
rect 29790 16870 29854 16934
rect 34958 17006 35022 17070
rect 39854 17006 39918 17070
rect 44750 17006 44814 17070
rect 34958 16870 35022 16934
rect 39854 16870 39918 16934
rect 44614 16870 44678 16934
rect 50054 17006 50118 17070
rect 54950 17006 55014 17070
rect 59710 17006 59774 17070
rect 49918 16870 49982 16934
rect 54950 16870 55014 16934
rect 59574 16870 59638 16934
rect 64878 17006 64942 17070
rect 69910 17006 69974 17070
rect 74670 17006 74734 17070
rect 64878 16870 64942 16934
rect 69910 16870 69974 16934
rect 79702 17006 79766 17070
rect 84870 17006 84934 17070
rect 89630 17006 89694 17070
rect 74670 16870 74734 16934
rect 79294 16870 79358 16934
rect 79974 16870 80038 16934
rect 84870 16870 84934 16934
rect 89630 16870 89694 16934
rect 94662 17006 94726 17070
rect 99694 17006 99758 17070
rect 104590 17006 104654 17070
rect 94934 16870 94998 16934
rect 99694 16870 99758 16934
rect 99830 16870 99894 16934
rect 104454 16870 104518 16934
rect 109622 17006 109686 17070
rect 109486 16870 109550 16934
rect 114654 17006 114718 17070
rect 114654 16870 114718 16934
rect 119822 17006 119886 17070
rect 124582 17006 124646 17070
rect 129614 17006 129678 17070
rect 134918 17006 134982 17070
rect 139542 17006 139606 17070
rect 144574 17006 144638 17070
rect 149606 17006 149670 17070
rect 119550 16870 119614 16934
rect 119822 16870 119886 16934
rect 124854 16870 124918 16934
rect 129886 16870 129950 16934
rect 134782 16870 134846 16934
rect 139814 16870 139878 16934
rect 144846 16870 144910 16934
rect 149470 16870 149534 16934
rect 154774 17006 154838 17070
rect 159534 17006 159598 17070
rect 154774 16870 154838 16934
rect 159534 16870 159598 16934
rect 164702 17006 164766 17070
rect 169734 17006 169798 17070
rect 174494 17006 174558 17070
rect 164702 16870 164766 16934
rect 169462 16870 169526 16934
rect 179526 17006 179590 17070
rect 184558 17006 184622 17070
rect 174766 16870 174830 16934
rect 179798 16870 179862 16934
rect 184558 16870 184622 16934
rect 184694 16870 184758 16934
rect 15102 16734 15166 16798
rect 21766 16734 21830 16798
rect 21766 16462 21830 16526
rect 29926 16462 29990 16526
rect 34822 16462 34886 16526
rect 29654 16326 29718 16390
rect 34822 16326 34886 16390
rect 39718 16462 39782 16526
rect 39718 16326 39782 16390
rect 44886 16462 44950 16526
rect 49782 16462 49846 16526
rect 44750 16326 44814 16390
rect 49782 16326 49846 16390
rect 54814 16462 54878 16526
rect 59846 16462 59910 16526
rect 64742 16462 64806 16526
rect 54814 16326 54878 16390
rect 59710 16326 59774 16390
rect 64742 16326 64806 16390
rect 69774 16462 69838 16526
rect 74806 16462 74870 16526
rect 79838 16462 79902 16526
rect 84734 16462 84798 16526
rect 69774 16326 69838 16390
rect 74534 16326 74598 16390
rect 79702 16326 79766 16390
rect 84598 16326 84662 16390
rect 89766 16462 89830 16526
rect 94798 16462 94862 16526
rect 99558 16462 99622 16526
rect 89494 16326 89558 16390
rect 94662 16326 94726 16390
rect 99558 16326 99622 16390
rect 104726 16462 104790 16526
rect 109758 16462 109822 16526
rect 114790 16462 114854 16526
rect 119686 16462 119750 16526
rect 104590 16326 104654 16390
rect 109622 16326 109686 16390
rect 114518 16326 114582 16390
rect 119686 16326 119750 16390
rect 124718 16462 124782 16526
rect 129750 16462 129814 16526
rect 134646 16462 134710 16526
rect 124582 16326 124646 16390
rect 129614 16326 129678 16390
rect 134646 16326 134710 16390
rect 139678 16462 139742 16526
rect 144710 16462 144774 16526
rect 149742 16462 149806 16526
rect 154638 16462 154702 16526
rect 159670 16462 159734 16526
rect 164566 16462 164630 16526
rect 139542 16326 139606 16390
rect 144574 16326 144638 16390
rect 149606 16326 149670 16390
rect 154502 16326 154566 16390
rect 159398 16326 159462 16390
rect 164566 16326 164630 16390
rect 169598 16462 169662 16526
rect 169598 16326 169662 16390
rect 174630 16462 174694 16526
rect 179662 16462 179726 16526
rect 184422 16462 184486 16526
rect 174494 16326 174558 16390
rect 179526 16326 179590 16390
rect 184422 16326 184486 16390
rect 204278 16462 204342 16526
rect 29790 16190 29854 16254
rect 34958 16190 35022 16254
rect 39854 16190 39918 16254
rect 44614 16190 44678 16254
rect 29246 15782 29310 15846
rect 50054 16190 50118 16254
rect 54950 16190 55014 16254
rect 59574 16190 59638 16254
rect 64878 16190 64942 16254
rect 69910 16190 69974 16254
rect 74670 16190 74734 16254
rect 49918 15918 49982 15982
rect 79974 16190 80038 16254
rect 84870 16190 84934 16254
rect 89630 16190 89694 16254
rect 94934 16190 94998 16254
rect 99830 16190 99894 16254
rect 104454 16190 104518 16254
rect 109486 16190 109550 16254
rect 79294 16054 79358 16118
rect 114654 16190 114718 16254
rect 119822 16190 119886 16254
rect 124854 16190 124918 16254
rect 129886 16190 129950 16254
rect 134918 16190 134982 16254
rect 139814 16190 139878 16254
rect 144846 16190 144910 16254
rect 149470 16190 149534 16254
rect 99694 16054 99758 16118
rect 119550 16054 119614 16118
rect 154774 16190 154838 16254
rect 159534 16190 159598 16254
rect 134782 15918 134846 15982
rect 164702 16190 164766 16254
rect 169462 16190 169526 16254
rect 174766 16190 174830 16254
rect 179798 16190 179862 16254
rect 184694 16190 184758 16254
rect 204006 16190 204070 16254
rect 184558 16054 184622 16118
rect 189182 15782 189246 15846
rect 217470 15646 217534 15710
rect 1230 15510 1294 15574
rect 15238 15510 15302 15574
rect 29518 15510 29582 15574
rect 29654 15510 29718 15574
rect 34822 15510 34886 15574
rect 39718 15510 39782 15574
rect 44750 15510 44814 15574
rect 49782 15510 49846 15574
rect 54814 15510 54878 15574
rect 59710 15510 59774 15574
rect 64742 15510 64806 15574
rect 69774 15510 69838 15574
rect 74534 15510 74598 15574
rect 79702 15510 79766 15574
rect 84598 15510 84662 15574
rect 89494 15510 89558 15574
rect 94662 15510 94726 15574
rect 99558 15510 99622 15574
rect 104590 15510 104654 15574
rect 109622 15510 109686 15574
rect 114518 15510 114582 15574
rect 119686 15510 119750 15574
rect 124582 15510 124646 15574
rect 129614 15510 129678 15574
rect 134646 15510 134710 15574
rect 139542 15510 139606 15574
rect 144574 15510 144638 15574
rect 149606 15510 149670 15574
rect 154502 15510 154566 15574
rect 159398 15510 159462 15574
rect 164566 15510 164630 15574
rect 169598 15510 169662 15574
rect 174494 15510 174558 15574
rect 179526 15510 179590 15574
rect 184422 15510 184486 15574
rect 189046 15510 189110 15574
rect 15238 15374 15302 15438
rect 20406 15238 20470 15302
rect 21902 15102 21966 15166
rect 29518 15102 29582 15166
rect 189046 15102 189110 15166
rect 204142 14966 204206 15030
rect 550 14150 614 14214
rect 1230 13878 1294 13942
rect 15102 14014 15166 14078
rect 29246 14014 29310 14078
rect 189182 14014 189246 14078
rect 21766 13878 21830 13942
rect 217470 14014 217534 14078
rect 20406 13742 20470 13806
rect 204006 13606 204070 13670
rect 2046 12518 2110 12582
rect 15238 12654 15302 12718
rect 21902 12382 21966 12446
rect 1230 12246 1294 12310
rect 2046 12246 2110 12310
rect 217470 12110 217534 12174
rect 20406 11022 20470 11086
rect 1230 10614 1294 10678
rect 217470 10478 217534 10542
rect 1230 8982 1294 9046
rect 217470 8846 217534 8910
rect 1230 7078 1294 7142
rect 217470 7214 217534 7278
rect 1230 5446 1294 5510
rect 217470 5582 217534 5646
rect 1230 3814 1294 3878
rect 217470 3950 217534 4014
rect 16870 3542 16934 3606
rect 16462 2590 16526 2654
rect 17686 2590 17750 2654
rect 18774 2590 18838 2654
rect 19998 2590 20062 2654
rect 21086 2590 21150 2654
rect 22310 2590 22374 2654
rect 23534 2590 23598 2654
rect 24622 2590 24686 2654
rect 25982 2590 26046 2654
rect 27070 2590 27134 2654
rect 28294 2590 28358 2654
rect 29246 2590 29310 2654
rect 30606 2590 30670 2654
rect 31694 2590 31758 2654
rect 32782 2590 32846 2654
rect 34006 2590 34070 2654
rect 35094 2590 35158 2654
rect 36454 2590 36518 2654
rect 37542 2590 37606 2654
rect 38630 2590 38694 2654
rect 39854 2590 39918 2654
rect 40942 2590 41006 2654
rect 42302 2590 42366 2654
rect 43390 2590 43454 2654
rect 44614 2590 44678 2654
rect 45838 2590 45902 2654
rect 46926 2590 46990 2654
rect 48014 2590 48078 2654
rect 49102 2590 49166 2654
rect 50326 2590 50390 2654
rect 51550 2590 51614 2654
rect 52774 2590 52838 2654
rect 53862 2590 53926 2654
rect 54950 2590 55014 2654
rect 56174 2590 56238 2654
rect 57398 2590 57462 2654
rect 58622 2590 58686 2654
rect 59846 2590 59910 2654
rect 60798 2590 60862 2654
rect 1230 2182 1294 2246
rect 3678 1820 3718 1838
rect 3718 1820 3742 1838
rect 3678 1774 3742 1820
rect 5446 1820 5454 1838
rect 5454 1820 5510 1838
rect 5446 1774 5510 1820
rect 6942 1774 7006 1838
rect 8710 1820 8758 1838
rect 8758 1820 8774 1838
rect 8710 1774 8774 1820
rect 10478 1820 10494 1838
rect 10494 1820 10542 1838
rect 10478 1774 10542 1820
rect 12110 1820 12118 1838
rect 12118 1820 12174 1838
rect 12110 1774 12174 1820
rect 13742 1820 13798 1838
rect 13798 1820 13806 1838
rect 13742 1774 13806 1820
rect 15510 1820 15534 1838
rect 15534 1820 15574 1838
rect 15510 1774 15574 1820
rect 17142 1820 17158 1838
rect 17158 1820 17206 1838
rect 17142 1774 17206 1820
rect 19046 1774 19110 1838
rect 20406 1774 20470 1838
rect 22174 1820 22198 1838
rect 22198 1820 22238 1838
rect 22174 1774 22238 1820
rect 23942 1774 24006 1838
rect 25438 1774 25502 1838
rect 27206 1820 27238 1838
rect 27238 1820 27270 1838
rect 27206 1774 27270 1820
rect 28838 1774 28902 1838
rect 30470 1774 30534 1838
rect 32374 1774 32438 1838
rect 33870 1774 33934 1838
rect 35502 1774 35566 1838
rect 37270 1820 37318 1838
rect 37318 1820 37334 1838
rect 37270 1774 37334 1820
rect 38902 1774 38966 1838
rect 40806 1774 40870 1838
rect 42438 1774 42502 1838
rect 43934 1774 43998 1838
rect 45702 1820 45718 1838
rect 45718 1820 45766 1838
rect 45702 1774 45766 1820
rect 47470 1774 47534 1838
rect 48966 1774 49030 1838
rect 50734 1820 50758 1838
rect 50758 1820 50798 1838
rect 50734 1774 50798 1820
rect 217470 2046 217534 2110
rect 52366 1774 52430 1838
rect 54134 1820 54174 1838
rect 54174 1820 54198 1838
rect 54134 1774 54198 1820
rect 55902 1774 55966 1838
rect 57670 1774 57734 1838
rect 59166 1820 59214 1838
rect 59214 1820 59230 1838
rect 59166 1774 59230 1820
rect 61070 1774 61134 1838
rect 62430 1774 62494 1838
rect 64062 1774 64126 1838
rect 65966 1774 66030 1838
rect 67462 1774 67526 1838
rect 69230 1820 69238 1838
rect 69238 1820 69294 1838
rect 69230 1774 69294 1820
rect 70862 1820 70918 1838
rect 70918 1820 70926 1838
rect 70862 1774 70926 1820
rect 72494 1774 72558 1838
rect 74262 1820 74278 1838
rect 74278 1820 74326 1838
rect 74262 1774 74326 1820
rect 75894 1774 75958 1838
rect 77662 1820 77694 1838
rect 77694 1820 77726 1838
rect 77662 1774 77726 1820
rect 79294 1820 79318 1838
rect 79318 1820 79358 1838
rect 79294 1774 79358 1820
rect 80926 1774 80990 1838
rect 82694 1820 82734 1838
rect 82734 1820 82758 1838
rect 82694 1774 82758 1820
rect 84598 1774 84662 1838
rect 85958 1774 86022 1838
rect 87726 1820 87774 1838
rect 87774 1820 87790 1838
rect 87726 1774 87790 1820
rect 89494 1774 89558 1838
rect 91126 1820 91134 1838
rect 91134 1820 91190 1838
rect 91126 1774 91190 1820
rect 92622 1774 92686 1838
rect 94662 1774 94726 1838
rect 96158 1820 96174 1838
rect 96174 1820 96222 1838
rect 96158 1774 96222 1820
rect 97790 1820 97798 1838
rect 97798 1820 97854 1838
rect 97790 1774 97854 1820
rect 99558 1774 99622 1838
rect 101190 1820 101214 1838
rect 101214 1820 101254 1838
rect 101190 1774 101254 1820
rect 102958 1774 103022 1838
rect 104454 1774 104518 1838
rect 106222 1820 106254 1838
rect 106254 1820 106286 1838
rect 106222 1774 106286 1820
rect 107854 1820 107878 1838
rect 107878 1820 107918 1838
rect 107854 1774 107918 1820
rect 109486 1774 109550 1838
rect 111118 1774 111182 1838
rect 112886 1820 112918 1838
rect 112918 1820 112950 1838
rect 112886 1774 112950 1820
rect 114654 1774 114718 1838
rect 116150 1774 116214 1838
rect 117918 1820 117958 1838
rect 117958 1820 117982 1838
rect 117918 1774 117982 1820
rect 119686 1820 119694 1838
rect 119694 1820 119750 1838
rect 119686 1774 119750 1820
rect 121454 1774 121518 1838
rect 122950 1820 122998 1838
rect 122998 1820 123014 1838
rect 122950 1774 123014 1820
rect 124718 1820 124734 1838
rect 124734 1820 124782 1838
rect 124718 1774 124782 1820
rect 126214 1774 126278 1838
rect 127982 1820 128038 1838
rect 128038 1820 128046 1838
rect 127982 1774 128046 1820
rect 129614 1774 129678 1838
rect 131382 1820 131398 1838
rect 131398 1820 131446 1838
rect 131382 1774 131446 1820
rect 133150 1774 133214 1838
rect 134646 1774 134710 1838
rect 136414 1820 136438 1838
rect 136438 1820 136478 1838
rect 136414 1774 136478 1820
rect 138182 1774 138246 1838
rect 139678 1774 139742 1838
rect 141446 1820 141478 1838
rect 141478 1820 141510 1838
rect 141446 1774 141510 1820
rect 143214 1774 143278 1838
rect 144710 1774 144774 1838
rect 146478 1820 146518 1838
rect 146518 1820 146542 1838
rect 146478 1774 146542 1820
rect 148110 1774 148174 1838
rect 150014 1774 150078 1838
rect 151646 1774 151710 1838
rect 153142 1774 153206 1838
rect 154910 1820 154918 1838
rect 154918 1820 154974 1838
rect 154910 1774 154974 1820
rect 156678 1774 156742 1838
rect 158174 1774 158238 1838
rect 159942 1820 159958 1838
rect 159958 1820 160006 1838
rect 159942 1774 160006 1820
rect 161710 1774 161774 1838
rect 163206 1774 163270 1838
rect 164974 1820 164998 1838
rect 164998 1820 165038 1838
rect 164974 1774 165038 1820
rect 166606 1774 166670 1838
rect 168374 1820 168414 1838
rect 168414 1820 168438 1838
rect 168374 1774 168438 1820
rect 170142 1774 170206 1838
rect 171638 1774 171702 1838
rect 173406 1820 173454 1838
rect 173454 1820 173470 1838
rect 173406 1774 173470 1820
rect 175174 1774 175238 1838
rect 176670 1774 176734 1838
rect 178438 1820 178494 1838
rect 178494 1820 178502 1838
rect 178438 1774 178502 1820
rect 180206 1774 180270 1838
rect 181702 1774 181766 1838
rect 183470 1820 183478 1838
rect 183478 1820 183534 1838
rect 183470 1774 183534 1820
rect 185102 1820 185158 1838
rect 185158 1820 185166 1838
rect 185102 1774 185166 1820
rect 186870 1820 186894 1838
rect 186894 1820 186934 1838
rect 186870 1774 186934 1820
rect 188638 1774 188702 1838
rect 190134 1774 190198 1838
rect 191902 1820 191934 1838
rect 191934 1820 191966 1838
rect 191902 1774 191966 1820
rect 193670 1774 193734 1838
rect 195166 1774 195230 1838
rect 196934 1820 196974 1838
rect 196974 1820 196998 1838
rect 196934 1774 196998 1820
rect 198702 1774 198766 1838
rect 200198 1774 200262 1838
rect 201966 1820 202014 1838
rect 202014 1820 202030 1838
rect 201966 1774 202030 1820
rect 203598 1820 203638 1838
rect 203638 1820 203662 1838
rect 203598 1774 203662 1820
rect 205230 1774 205294 1838
rect 207134 1774 207198 1838
rect 208630 1820 208678 1838
rect 208678 1820 208694 1838
rect 208630 1774 208694 1820
rect 210398 1820 210414 1838
rect 210414 1820 210462 1838
rect 210398 1774 210462 1820
rect 211894 1774 211958 1838
rect 213662 1820 213718 1838
rect 213718 1820 213726 1838
rect 213662 1774 213726 1820
rect 215430 1820 215454 1838
rect 215454 1820 215494 1838
rect 215430 1774 215494 1820
rect 958 1230 1022 1294
rect 1094 1230 1158 1294
rect 1230 1230 1294 1294
rect 3678 1230 3742 1294
rect 5446 1230 5510 1294
rect 6942 1230 7006 1294
rect 8710 1230 8774 1294
rect 10478 1230 10542 1294
rect 12110 1230 12174 1294
rect 13742 1230 13806 1294
rect 15510 1230 15574 1294
rect 17142 1230 17206 1294
rect 19046 1230 19110 1294
rect 20406 1230 20470 1294
rect 22174 1230 22238 1294
rect 23942 1230 24006 1294
rect 25438 1230 25502 1294
rect 27206 1230 27270 1294
rect 28838 1230 28902 1294
rect 30470 1230 30534 1294
rect 32374 1230 32438 1294
rect 33870 1230 33934 1294
rect 35502 1230 35566 1294
rect 37270 1230 37334 1294
rect 38902 1230 38966 1294
rect 40806 1230 40870 1294
rect 42438 1230 42502 1294
rect 43934 1230 43998 1294
rect 45702 1230 45766 1294
rect 47470 1230 47534 1294
rect 48966 1230 49030 1294
rect 50734 1230 50798 1294
rect 52366 1230 52430 1294
rect 54134 1230 54198 1294
rect 55902 1230 55966 1294
rect 57670 1230 57734 1294
rect 59166 1230 59230 1294
rect 61070 1230 61134 1294
rect 62430 1230 62494 1294
rect 64062 1230 64126 1294
rect 65966 1230 66030 1294
rect 67462 1230 67526 1294
rect 69230 1230 69294 1294
rect 70862 1230 70926 1294
rect 72494 1230 72558 1294
rect 74262 1230 74326 1294
rect 75894 1230 75958 1294
rect 77662 1230 77726 1294
rect 79294 1230 79358 1294
rect 80926 1230 80990 1294
rect 82694 1230 82758 1294
rect 84598 1230 84662 1294
rect 85958 1230 86022 1294
rect 87726 1230 87790 1294
rect 89494 1230 89558 1294
rect 91126 1230 91190 1294
rect 92622 1230 92686 1294
rect 94662 1230 94726 1294
rect 96158 1230 96222 1294
rect 97790 1230 97854 1294
rect 99558 1230 99622 1294
rect 101190 1230 101254 1294
rect 102958 1230 103022 1294
rect 104454 1230 104518 1294
rect 106222 1230 106286 1294
rect 107854 1230 107918 1294
rect 109486 1230 109550 1294
rect 111118 1230 111182 1294
rect 112886 1230 112950 1294
rect 114654 1230 114718 1294
rect 116150 1230 116214 1294
rect 117918 1230 117982 1294
rect 119686 1230 119750 1294
rect 121454 1230 121518 1294
rect 122950 1230 123014 1294
rect 124718 1230 124782 1294
rect 126214 1230 126278 1294
rect 127982 1230 128046 1294
rect 129614 1230 129678 1294
rect 131382 1230 131446 1294
rect 133150 1230 133214 1294
rect 134646 1230 134710 1294
rect 136414 1230 136478 1294
rect 138182 1230 138246 1294
rect 139678 1230 139742 1294
rect 141446 1230 141510 1294
rect 143214 1230 143278 1294
rect 144710 1230 144774 1294
rect 146478 1230 146542 1294
rect 148110 1230 148174 1294
rect 150014 1230 150078 1294
rect 151646 1230 151710 1294
rect 153142 1230 153206 1294
rect 154910 1230 154974 1294
rect 156678 1230 156742 1294
rect 158174 1230 158238 1294
rect 159942 1230 160006 1294
rect 161710 1230 161774 1294
rect 163206 1230 163270 1294
rect 164974 1230 165038 1294
rect 166606 1230 166670 1294
rect 168374 1230 168438 1294
rect 170142 1230 170206 1294
rect 171638 1230 171702 1294
rect 173406 1230 173470 1294
rect 175174 1230 175238 1294
rect 176670 1230 176734 1294
rect 178438 1230 178502 1294
rect 180206 1230 180270 1294
rect 181702 1230 181766 1294
rect 183470 1230 183534 1294
rect 185102 1230 185166 1294
rect 186870 1230 186934 1294
rect 188638 1230 188702 1294
rect 190134 1230 190198 1294
rect 191902 1230 191966 1294
rect 193670 1230 193734 1294
rect 195166 1230 195230 1294
rect 196934 1230 196998 1294
rect 198702 1230 198766 1294
rect 200198 1230 200262 1294
rect 201966 1230 202030 1294
rect 203598 1230 203662 1294
rect 205230 1230 205294 1294
rect 207134 1230 207198 1294
rect 208630 1230 208694 1294
rect 210398 1230 210462 1294
rect 211894 1230 211958 1294
rect 213662 1230 213726 1294
rect 215430 1230 215494 1294
rect 217470 1230 217534 1294
rect 217606 1230 217670 1294
rect 217742 1230 217806 1294
rect 958 1094 1022 1158
rect 1094 1094 1158 1158
rect 1230 1094 1294 1158
rect 217470 1094 217534 1158
rect 217606 1094 217670 1158
rect 217742 1094 217806 1158
rect 958 958 1022 1022
rect 1094 958 1158 1022
rect 1230 958 1294 1022
rect 217470 958 217534 1022
rect 217606 958 217670 1022
rect 217742 958 217806 1022
rect 278 550 342 614
rect 414 550 478 614
rect 550 550 614 614
rect 16870 550 16934 614
rect 218150 550 218214 614
rect 218286 550 218350 614
rect 218422 550 218486 614
rect 278 414 342 478
rect 414 414 478 478
rect 550 414 614 478
rect 218150 414 218214 478
rect 218286 414 218350 478
rect 218422 414 218486 478
rect 278 278 342 342
rect 414 278 478 342
rect 550 278 614 342
rect 218150 278 218214 342
rect 218286 278 218350 342
rect 218422 278 218486 342
<< metal4 >>
rect 272 143822 620 143828
rect 272 143758 278 143822
rect 342 143758 414 143822
rect 478 143758 550 143822
rect 614 143758 620 143822
rect 272 143686 620 143758
rect 272 143622 278 143686
rect 342 143622 414 143686
rect 478 143622 550 143686
rect 614 143622 620 143686
rect 272 143550 620 143622
rect 272 143486 278 143550
rect 342 143486 414 143550
rect 478 143486 550 143550
rect 614 143486 620 143550
rect 272 29718 620 143486
rect 272 29654 550 29718
rect 614 29654 620 29718
rect 272 26726 620 29654
rect 272 26662 550 26726
rect 614 26662 620 26726
rect 272 23870 620 26662
rect 272 23806 550 23870
rect 614 23806 620 23870
rect 272 21014 620 23806
rect 272 20950 550 21014
rect 614 20950 620 21014
rect 272 18430 620 20950
rect 272 18366 550 18430
rect 614 18366 620 18430
rect 272 14214 620 18366
rect 272 14150 550 14214
rect 614 14150 620 14214
rect 272 614 620 14150
rect 952 143142 1300 143148
rect 952 143078 958 143142
rect 1022 143078 1094 143142
rect 1158 143078 1230 143142
rect 1294 143078 1300 143142
rect 952 143006 1300 143078
rect 952 142942 958 143006
rect 1022 142942 1094 143006
rect 1158 142942 1230 143006
rect 1294 142942 1300 143006
rect 952 142870 1300 142942
rect 952 142806 958 142870
rect 1022 142806 1094 142870
rect 1158 142806 1230 142870
rect 1294 142806 1300 142870
rect 952 141782 1300 142806
rect 1904 142870 1980 142876
rect 1904 142806 1910 142870
rect 1974 142806 1980 142870
rect 1904 142462 1980 142806
rect 1904 142430 1910 142462
rect 1909 142398 1910 142430
rect 1974 142430 1980 142462
rect 3672 142870 3748 142876
rect 3672 142806 3678 142870
rect 3742 142806 3748 142870
rect 3672 142462 3748 142806
rect 3672 142430 3678 142462
rect 1974 142398 1975 142430
rect 1909 142397 1975 142398
rect 3677 142398 3678 142430
rect 3742 142430 3748 142462
rect 5440 142870 5516 142876
rect 5440 142806 5446 142870
rect 5510 142806 5516 142870
rect 5440 142462 5516 142806
rect 5440 142430 5446 142462
rect 3742 142398 3743 142430
rect 3677 142397 3743 142398
rect 5445 142398 5446 142430
rect 5510 142430 5516 142462
rect 7208 142870 7284 142876
rect 7208 142806 7214 142870
rect 7278 142806 7284 142870
rect 7208 142462 7284 142806
rect 7208 142430 7214 142462
rect 5510 142398 5511 142430
rect 5445 142397 5511 142398
rect 7213 142398 7214 142430
rect 7278 142430 7284 142462
rect 8704 142870 8780 142876
rect 8704 142806 8710 142870
rect 8774 142806 8780 142870
rect 8704 142462 8780 142806
rect 8704 142430 8710 142462
rect 7278 142398 7279 142430
rect 7213 142397 7279 142398
rect 8709 142398 8710 142430
rect 8774 142430 8780 142462
rect 10472 142870 10548 142876
rect 10472 142806 10478 142870
rect 10542 142806 10548 142870
rect 10472 142462 10548 142806
rect 10472 142430 10478 142462
rect 8774 142398 8775 142430
rect 8709 142397 8775 142398
rect 10477 142398 10478 142430
rect 10542 142430 10548 142462
rect 12240 142870 12316 142876
rect 12240 142806 12246 142870
rect 12310 142806 12316 142870
rect 12240 142462 12316 142806
rect 12240 142430 12246 142462
rect 10542 142398 10543 142430
rect 10477 142397 10543 142398
rect 12245 142398 12246 142430
rect 12310 142430 12316 142462
rect 13736 142870 13812 142876
rect 13736 142806 13742 142870
rect 13806 142806 13812 142870
rect 13736 142462 13812 142806
rect 13736 142430 13742 142462
rect 12310 142398 12311 142430
rect 12245 142397 12311 142398
rect 13741 142398 13742 142430
rect 13806 142430 13812 142462
rect 15368 142870 15444 142876
rect 15368 142806 15374 142870
rect 15438 142806 15444 142870
rect 15368 142462 15444 142806
rect 15368 142430 15374 142462
rect 13806 142398 13807 142430
rect 13741 142397 13807 142398
rect 15373 142398 15374 142430
rect 15438 142430 15444 142462
rect 17136 142870 17212 142876
rect 17136 142806 17142 142870
rect 17206 142806 17212 142870
rect 17136 142462 17212 142806
rect 17136 142430 17142 142462
rect 15438 142398 15439 142430
rect 15373 142397 15439 142398
rect 17141 142398 17142 142430
rect 17206 142430 17212 142462
rect 18904 142870 18980 142876
rect 18904 142806 18910 142870
rect 18974 142806 18980 142870
rect 18904 142462 18980 142806
rect 18904 142430 18910 142462
rect 17206 142398 17207 142430
rect 17141 142397 17207 142398
rect 18909 142398 18910 142430
rect 18974 142430 18980 142462
rect 20400 142870 20476 142876
rect 20400 142806 20406 142870
rect 20470 142806 20476 142870
rect 20400 142462 20476 142806
rect 20400 142430 20406 142462
rect 18974 142398 18975 142430
rect 18909 142397 18975 142398
rect 20405 142398 20406 142430
rect 20470 142430 20476 142462
rect 22168 142870 22244 142876
rect 22168 142806 22174 142870
rect 22238 142806 22244 142870
rect 22168 142462 22244 142806
rect 22168 142430 22174 142462
rect 20470 142398 20471 142430
rect 20405 142397 20471 142398
rect 22173 142398 22174 142430
rect 22238 142430 22244 142462
rect 23936 142870 24012 142876
rect 23936 142806 23942 142870
rect 24006 142806 24012 142870
rect 23936 142462 24012 142806
rect 23936 142430 23942 142462
rect 22238 142398 22239 142430
rect 22173 142397 22239 142398
rect 23941 142398 23942 142430
rect 24006 142430 24012 142462
rect 25432 142870 25508 142876
rect 25432 142806 25438 142870
rect 25502 142806 25508 142870
rect 25432 142462 25508 142806
rect 25432 142430 25438 142462
rect 24006 142398 24007 142430
rect 23941 142397 24007 142398
rect 25437 142398 25438 142430
rect 25502 142430 25508 142462
rect 27200 142870 27276 142876
rect 27200 142806 27206 142870
rect 27270 142806 27276 142870
rect 27200 142462 27276 142806
rect 27200 142430 27206 142462
rect 25502 142398 25503 142430
rect 25437 142397 25503 142398
rect 27205 142398 27206 142430
rect 27270 142430 27276 142462
rect 28968 142870 29044 142876
rect 28968 142806 28974 142870
rect 29038 142806 29044 142870
rect 28968 142462 29044 142806
rect 28968 142430 28974 142462
rect 27270 142398 27271 142430
rect 27205 142397 27271 142398
rect 28973 142398 28974 142430
rect 29038 142430 29044 142462
rect 29038 142398 29039 142430
rect 28973 142397 29039 142398
rect 952 141718 1230 141782
rect 1294 141718 1300 141782
rect 952 139878 1300 141718
rect 952 139814 1230 139878
rect 1294 139814 1300 139878
rect 952 138246 1300 139814
rect 952 138182 1230 138246
rect 1294 138182 1300 138246
rect 952 136750 1300 138182
rect 952 136686 1230 136750
rect 1294 136686 1300 136750
rect 952 134982 1300 136686
rect 952 134918 1230 134982
rect 1294 134918 1300 134982
rect 952 133214 1300 134918
rect 952 133150 1230 133214
rect 1294 133150 1300 133214
rect 29512 133214 29588 144100
rect 30464 142870 30540 142876
rect 30464 142806 30470 142870
rect 30534 142806 30540 142870
rect 30464 142462 30540 142806
rect 30464 142430 30470 142462
rect 30469 142398 30470 142430
rect 30534 142430 30540 142462
rect 32232 142870 32308 142876
rect 32232 142806 32238 142870
rect 32302 142806 32308 142870
rect 32232 142462 32308 142806
rect 32232 142430 32238 142462
rect 30534 142398 30535 142430
rect 30469 142397 30535 142398
rect 32237 142398 32238 142430
rect 32302 142430 32308 142462
rect 33864 142870 33940 142876
rect 33864 142806 33870 142870
rect 33934 142806 33940 142870
rect 33864 142462 33940 142806
rect 33864 142430 33870 142462
rect 32302 142398 32303 142430
rect 32237 142397 32303 142398
rect 33869 142398 33870 142430
rect 33934 142430 33940 142462
rect 33934 142398 33935 142430
rect 33869 142397 33935 142398
rect 29512 133182 29518 133214
rect 952 131582 1300 133150
rect 29517 133150 29518 133182
rect 29582 133182 29588 133214
rect 34408 133214 34484 144100
rect 35496 142870 35572 142876
rect 35496 142806 35502 142870
rect 35566 142806 35572 142870
rect 35496 142462 35572 142806
rect 35496 142430 35502 142462
rect 35501 142398 35502 142430
rect 35566 142430 35572 142462
rect 37400 142870 37476 142876
rect 37400 142806 37406 142870
rect 37470 142806 37476 142870
rect 37400 142462 37476 142806
rect 37400 142430 37406 142462
rect 35566 142398 35567 142430
rect 35501 142397 35567 142398
rect 37405 142398 37406 142430
rect 37470 142430 37476 142462
rect 38896 142870 38972 142876
rect 38896 142806 38902 142870
rect 38966 142806 38972 142870
rect 38896 142462 38972 142806
rect 38896 142430 38902 142462
rect 37470 142398 37471 142430
rect 37405 142397 37471 142398
rect 38901 142398 38902 142430
rect 38966 142430 38972 142462
rect 38966 142398 38967 142430
rect 38901 142397 38967 142398
rect 34408 133182 34414 133214
rect 29582 133150 29583 133182
rect 29517 133149 29583 133150
rect 34413 133150 34414 133182
rect 34478 133182 34484 133214
rect 39440 133214 39516 144100
rect 40664 142870 40740 142876
rect 40664 142806 40670 142870
rect 40734 142806 40740 142870
rect 40664 142462 40740 142806
rect 40664 142430 40670 142462
rect 40669 142398 40670 142430
rect 40734 142430 40740 142462
rect 42432 142870 42508 142876
rect 42432 142806 42438 142870
rect 42502 142806 42508 142870
rect 42432 142462 42508 142806
rect 42432 142430 42438 142462
rect 40734 142398 40735 142430
rect 40669 142397 40735 142398
rect 42437 142398 42438 142430
rect 42502 142430 42508 142462
rect 43928 142870 44004 142876
rect 43928 142806 43934 142870
rect 43998 142806 44004 142870
rect 43928 142462 44004 142806
rect 43928 142430 43934 142462
rect 42502 142398 42503 142430
rect 42437 142397 42503 142398
rect 43933 142398 43934 142430
rect 43998 142430 44004 142462
rect 43998 142398 43999 142430
rect 43933 142397 43999 142398
rect 39440 133182 39446 133214
rect 34478 133150 34479 133182
rect 34413 133149 34479 133150
rect 39445 133150 39446 133182
rect 39510 133182 39516 133214
rect 44472 133214 44548 144100
rect 45696 142870 45772 142876
rect 45696 142806 45702 142870
rect 45766 142806 45772 142870
rect 45696 142462 45772 142806
rect 45696 142430 45702 142462
rect 45701 142398 45702 142430
rect 45766 142430 45772 142462
rect 47464 142870 47540 142876
rect 47464 142806 47470 142870
rect 47534 142806 47540 142870
rect 47464 142462 47540 142806
rect 47464 142430 47470 142462
rect 45766 142398 45767 142430
rect 45701 142397 45767 142398
rect 47469 142398 47470 142430
rect 47534 142430 47540 142462
rect 48960 142870 49036 142876
rect 48960 142806 48966 142870
rect 49030 142806 49036 142870
rect 48960 142462 49036 142806
rect 48960 142430 48966 142462
rect 47534 142398 47535 142430
rect 47469 142397 47535 142398
rect 48965 142398 48966 142430
rect 49030 142430 49036 142462
rect 49030 142398 49031 142430
rect 48965 142397 49031 142398
rect 44472 133182 44478 133214
rect 39510 133150 39511 133182
rect 39445 133149 39511 133150
rect 44477 133150 44478 133182
rect 44542 133182 44548 133214
rect 49504 133214 49580 144100
rect 50728 142870 50804 142876
rect 50728 142806 50734 142870
rect 50798 142806 50804 142870
rect 50728 142462 50804 142806
rect 50728 142430 50734 142462
rect 50733 142398 50734 142430
rect 50798 142430 50804 142462
rect 52360 142870 52436 142876
rect 52360 142806 52366 142870
rect 52430 142806 52436 142870
rect 52360 142462 52436 142806
rect 52360 142430 52366 142462
rect 50798 142398 50799 142430
rect 50733 142397 50799 142398
rect 52365 142398 52366 142430
rect 52430 142430 52436 142462
rect 53992 142870 54068 142876
rect 53992 142806 53998 142870
rect 54062 142806 54068 142870
rect 53992 142462 54068 142806
rect 53992 142430 53998 142462
rect 52430 142398 52431 142430
rect 52365 142397 52431 142398
rect 53997 142398 53998 142430
rect 54062 142430 54068 142462
rect 54062 142398 54063 142430
rect 53997 142397 54063 142398
rect 49504 133182 49510 133214
rect 44542 133150 44543 133182
rect 44477 133149 44543 133150
rect 49509 133150 49510 133182
rect 49574 133182 49580 133214
rect 54536 133214 54612 144100
rect 55896 142870 55972 142876
rect 55896 142806 55902 142870
rect 55966 142806 55972 142870
rect 55896 142462 55972 142806
rect 55896 142430 55902 142462
rect 55901 142398 55902 142430
rect 55966 142430 55972 142462
rect 57392 142870 57468 142876
rect 57392 142806 57398 142870
rect 57462 142806 57468 142870
rect 57392 142462 57468 142806
rect 57392 142430 57398 142462
rect 55966 142398 55967 142430
rect 55901 142397 55967 142398
rect 57397 142398 57398 142430
rect 57462 142430 57468 142462
rect 59160 142870 59236 142876
rect 59160 142806 59166 142870
rect 59230 142806 59236 142870
rect 59160 142462 59236 142806
rect 59160 142430 59166 142462
rect 57462 142398 57463 142430
rect 57397 142397 57463 142398
rect 59165 142398 59166 142430
rect 59230 142430 59236 142462
rect 59230 142398 59231 142430
rect 59165 142397 59231 142398
rect 54536 133182 54542 133214
rect 49574 133150 49575 133182
rect 49509 133149 49575 133150
rect 54541 133150 54542 133182
rect 54606 133182 54612 133214
rect 59432 133214 59508 144100
rect 60928 142870 61004 142876
rect 60928 142806 60934 142870
rect 60998 142806 61004 142870
rect 60928 142462 61004 142806
rect 60928 142430 60934 142462
rect 60933 142398 60934 142430
rect 60998 142430 61004 142462
rect 62424 142870 62500 142876
rect 62424 142806 62430 142870
rect 62494 142806 62500 142870
rect 62424 142462 62500 142806
rect 62424 142430 62430 142462
rect 60998 142398 60999 142430
rect 60933 142397 60999 142398
rect 62429 142398 62430 142430
rect 62494 142430 62500 142462
rect 64056 142870 64132 142876
rect 64056 142806 64062 142870
rect 64126 142806 64132 142870
rect 64056 142462 64132 142806
rect 64056 142430 64062 142462
rect 62494 142398 62495 142430
rect 62429 142397 62495 142398
rect 64061 142398 64062 142430
rect 64126 142430 64132 142462
rect 64126 142398 64127 142430
rect 64061 142397 64127 142398
rect 59432 133182 59438 133214
rect 54606 133150 54607 133182
rect 54541 133149 54607 133150
rect 59437 133150 59438 133182
rect 59502 133182 59508 133214
rect 64464 133214 64540 144100
rect 65960 142870 66036 142876
rect 65960 142806 65966 142870
rect 66030 142806 66036 142870
rect 65960 142462 66036 142806
rect 65960 142430 65966 142462
rect 65965 142398 65966 142430
rect 66030 142430 66036 142462
rect 67456 142870 67532 142876
rect 67456 142806 67462 142870
rect 67526 142806 67532 142870
rect 67456 142462 67532 142806
rect 67456 142430 67462 142462
rect 66030 142398 66031 142430
rect 65965 142397 66031 142398
rect 67461 142398 67462 142430
rect 67526 142430 67532 142462
rect 69360 142870 69436 142876
rect 69360 142806 69366 142870
rect 69430 142806 69436 142870
rect 69360 142462 69436 142806
rect 69360 142430 69366 142462
rect 67526 142398 67527 142430
rect 67461 142397 67527 142398
rect 69365 142398 69366 142430
rect 69430 142430 69436 142462
rect 69430 142398 69431 142430
rect 69365 142397 69431 142398
rect 64464 133182 64470 133214
rect 59502 133150 59503 133182
rect 59437 133149 59503 133150
rect 64469 133150 64470 133182
rect 64534 133182 64540 133214
rect 69496 133214 69572 144100
rect 70856 142870 70932 142876
rect 70856 142806 70862 142870
rect 70926 142806 70932 142870
rect 70856 142462 70932 142806
rect 70856 142430 70862 142462
rect 70861 142398 70862 142430
rect 70926 142430 70932 142462
rect 72488 142870 72564 142876
rect 72488 142806 72494 142870
rect 72558 142806 72564 142870
rect 72488 142462 72564 142806
rect 72488 142430 72494 142462
rect 70926 142398 70927 142430
rect 70861 142397 70927 142398
rect 72493 142398 72494 142430
rect 72558 142430 72564 142462
rect 74256 142870 74332 142876
rect 74256 142806 74262 142870
rect 74326 142806 74332 142870
rect 74256 142462 74332 142806
rect 74256 142430 74262 142462
rect 72558 142398 72559 142430
rect 72493 142397 72559 142398
rect 74261 142398 74262 142430
rect 74326 142430 74332 142462
rect 74326 142398 74327 142430
rect 74261 142397 74327 142398
rect 69496 133182 69502 133214
rect 64534 133150 64535 133182
rect 64469 133149 64535 133150
rect 69501 133150 69502 133182
rect 69566 133182 69572 133214
rect 74528 133214 74604 144100
rect 75888 142870 75964 142876
rect 75888 142806 75894 142870
rect 75958 142806 75964 142870
rect 75888 142462 75964 142806
rect 75888 142430 75894 142462
rect 75893 142398 75894 142430
rect 75958 142430 75964 142462
rect 77656 142870 77732 142876
rect 77656 142806 77662 142870
rect 77726 142806 77732 142870
rect 77656 142462 77732 142806
rect 77656 142430 77662 142462
rect 75958 142398 75959 142430
rect 75893 142397 75959 142398
rect 77661 142398 77662 142430
rect 77726 142430 77732 142462
rect 79424 142870 79500 142876
rect 79424 142806 79430 142870
rect 79494 142806 79500 142870
rect 79424 142462 79500 142806
rect 79424 142430 79430 142462
rect 77726 142398 77727 142430
rect 77661 142397 77727 142398
rect 79429 142398 79430 142430
rect 79494 142430 79500 142462
rect 79494 142398 79495 142430
rect 79429 142397 79495 142398
rect 74528 133182 74534 133214
rect 69566 133150 69567 133182
rect 69501 133149 69567 133150
rect 74533 133150 74534 133182
rect 74598 133182 74604 133214
rect 79560 133214 79636 144100
rect 80920 142870 80996 142876
rect 80920 142806 80926 142870
rect 80990 142806 80996 142870
rect 80920 142462 80996 142806
rect 80920 142430 80926 142462
rect 80925 142398 80926 142430
rect 80990 142430 80996 142462
rect 82688 142870 82764 142876
rect 82688 142806 82694 142870
rect 82758 142806 82764 142870
rect 82688 142462 82764 142806
rect 82688 142430 82694 142462
rect 80990 142398 80991 142430
rect 80925 142397 80991 142398
rect 82693 142398 82694 142430
rect 82758 142430 82764 142462
rect 82758 142398 82759 142430
rect 82693 142397 82759 142398
rect 79560 133182 79566 133214
rect 74598 133150 74599 133182
rect 74533 133149 74599 133150
rect 79565 133150 79566 133182
rect 79630 133182 79636 133214
rect 84320 133214 84396 144100
rect 84592 142870 84668 142876
rect 84592 142806 84598 142870
rect 84662 142806 84668 142870
rect 84592 142462 84668 142806
rect 84592 142430 84598 142462
rect 84597 142398 84598 142430
rect 84662 142430 84668 142462
rect 85952 142870 86028 142876
rect 85952 142806 85958 142870
rect 86022 142806 86028 142870
rect 85952 142462 86028 142806
rect 85952 142430 85958 142462
rect 84662 142398 84663 142430
rect 84597 142397 84663 142398
rect 85957 142398 85958 142430
rect 86022 142430 86028 142462
rect 87720 142870 87796 142876
rect 87720 142806 87726 142870
rect 87790 142806 87796 142870
rect 87720 142462 87796 142806
rect 87720 142430 87726 142462
rect 86022 142398 86023 142430
rect 85957 142397 86023 142398
rect 87725 142398 87726 142430
rect 87790 142430 87796 142462
rect 87790 142398 87791 142430
rect 87725 142397 87791 142398
rect 84320 133182 84326 133214
rect 79630 133150 79631 133182
rect 79565 133149 79631 133150
rect 84325 133150 84326 133182
rect 84390 133182 84396 133214
rect 89352 133214 89428 144100
rect 89488 142870 89564 142876
rect 89488 142806 89494 142870
rect 89558 142806 89564 142870
rect 89488 142462 89564 142806
rect 89488 142430 89494 142462
rect 89493 142398 89494 142430
rect 89558 142430 89564 142462
rect 90984 142870 91060 142876
rect 90984 142806 90990 142870
rect 91054 142806 91060 142870
rect 90984 142462 91060 142806
rect 90984 142430 90990 142462
rect 89558 142398 89559 142430
rect 89493 142397 89559 142398
rect 90989 142398 90990 142430
rect 91054 142430 91060 142462
rect 92888 142870 92964 142876
rect 92888 142806 92894 142870
rect 92958 142806 92964 142870
rect 92888 142462 92964 142806
rect 92888 142430 92894 142462
rect 91054 142398 91055 142430
rect 90989 142397 91055 142398
rect 92893 142398 92894 142430
rect 92958 142430 92964 142462
rect 94384 142870 94460 142876
rect 94384 142806 94390 142870
rect 94454 142806 94460 142870
rect 94384 142462 94460 142806
rect 94384 142430 94390 142462
rect 92958 142398 92959 142430
rect 92893 142397 92959 142398
rect 94389 142398 94390 142430
rect 94454 142430 94460 142462
rect 94454 142398 94455 142430
rect 94389 142397 94455 142398
rect 89352 133182 89358 133214
rect 84390 133150 84391 133182
rect 84325 133149 84391 133150
rect 89357 133150 89358 133182
rect 89422 133182 89428 133214
rect 94520 133214 94596 144100
rect 96152 142870 96228 142876
rect 96152 142806 96158 142870
rect 96222 142806 96228 142870
rect 96152 142462 96228 142806
rect 96152 142430 96158 142462
rect 96157 142398 96158 142430
rect 96222 142430 96228 142462
rect 97784 142870 97860 142876
rect 97784 142806 97790 142870
rect 97854 142806 97860 142870
rect 97784 142462 97860 142806
rect 97784 142430 97790 142462
rect 96222 142398 96223 142430
rect 96157 142397 96223 142398
rect 97789 142398 97790 142430
rect 97854 142430 97860 142462
rect 97854 142398 97855 142430
rect 97789 142397 97855 142398
rect 94520 133182 94526 133214
rect 89422 133150 89423 133182
rect 89357 133149 89423 133150
rect 94525 133150 94526 133182
rect 94590 133182 94596 133214
rect 99416 133214 99492 144100
rect 99552 142870 99628 142876
rect 99552 142806 99558 142870
rect 99622 142806 99628 142870
rect 99552 142462 99628 142806
rect 99552 142430 99558 142462
rect 99557 142398 99558 142430
rect 99622 142430 99628 142462
rect 101184 142870 101260 142876
rect 101184 142806 101190 142870
rect 101254 142806 101260 142870
rect 101184 142462 101260 142806
rect 101184 142430 101190 142462
rect 99622 142398 99623 142430
rect 99557 142397 99623 142398
rect 101189 142398 101190 142430
rect 101254 142430 101260 142462
rect 102952 142870 103028 142876
rect 102952 142806 102958 142870
rect 103022 142806 103028 142870
rect 102952 142462 103028 142806
rect 102952 142430 102958 142462
rect 101254 142398 101255 142430
rect 101189 142397 101255 142398
rect 102957 142398 102958 142430
rect 103022 142430 103028 142462
rect 103022 142398 103023 142430
rect 102957 142397 103023 142398
rect 99416 133182 99422 133214
rect 94590 133150 94591 133182
rect 94525 133149 94591 133150
rect 99421 133150 99422 133182
rect 99486 133182 99492 133214
rect 104312 133214 104388 144100
rect 104448 142870 104524 142876
rect 104448 142806 104454 142870
rect 104518 142806 104524 142870
rect 104448 142462 104524 142806
rect 104448 142430 104454 142462
rect 104453 142398 104454 142430
rect 104518 142430 104524 142462
rect 106216 142870 106292 142876
rect 106216 142806 106222 142870
rect 106286 142806 106292 142870
rect 106216 142462 106292 142806
rect 106216 142430 106222 142462
rect 104518 142398 104519 142430
rect 104453 142397 104519 142398
rect 106221 142398 106222 142430
rect 106286 142430 106292 142462
rect 107848 142870 107924 142876
rect 107848 142806 107854 142870
rect 107918 142806 107924 142870
rect 107848 142462 107924 142806
rect 107848 142430 107854 142462
rect 106286 142398 106287 142430
rect 106221 142397 106287 142398
rect 107853 142398 107854 142430
rect 107918 142430 107924 142462
rect 107918 142398 107919 142430
rect 107853 142397 107919 142398
rect 104312 133182 104318 133214
rect 99486 133150 99487 133182
rect 99421 133149 99487 133150
rect 104317 133150 104318 133182
rect 104382 133182 104388 133214
rect 109344 133214 109420 144100
rect 109616 142870 109692 142876
rect 109616 142806 109622 142870
rect 109686 142806 109692 142870
rect 109616 142462 109692 142806
rect 109616 142430 109622 142462
rect 109621 142398 109622 142430
rect 109686 142430 109692 142462
rect 111112 142870 111188 142876
rect 111112 142806 111118 142870
rect 111182 142806 111188 142870
rect 111112 142462 111188 142806
rect 111112 142430 111118 142462
rect 109686 142398 109687 142430
rect 109621 142397 109687 142398
rect 111117 142398 111118 142430
rect 111182 142430 111188 142462
rect 112880 142870 112956 142876
rect 112880 142806 112886 142870
rect 112950 142806 112956 142870
rect 112880 142462 112956 142806
rect 112880 142430 112886 142462
rect 111182 142398 111183 142430
rect 111117 142397 111183 142398
rect 112885 142398 112886 142430
rect 112950 142430 112956 142462
rect 112950 142398 112951 142430
rect 112885 142397 112951 142398
rect 109344 133182 109350 133214
rect 104382 133150 104383 133182
rect 104317 133149 104383 133150
rect 109349 133150 109350 133182
rect 109414 133182 109420 133214
rect 114376 133214 114452 144100
rect 114648 142870 114724 142876
rect 114648 142806 114654 142870
rect 114718 142806 114724 142870
rect 114648 142462 114724 142806
rect 114648 142430 114654 142462
rect 114653 142398 114654 142430
rect 114718 142430 114724 142462
rect 116144 142870 116220 142876
rect 116144 142806 116150 142870
rect 116214 142806 116220 142870
rect 116144 142462 116220 142806
rect 116144 142430 116150 142462
rect 114718 142398 114719 142430
rect 114653 142397 114719 142398
rect 116149 142398 116150 142430
rect 116214 142430 116220 142462
rect 117912 142870 117988 142876
rect 117912 142806 117918 142870
rect 117982 142806 117988 142870
rect 117912 142462 117988 142806
rect 117912 142430 117918 142462
rect 116214 142398 116215 142430
rect 116149 142397 116215 142398
rect 117917 142398 117918 142430
rect 117982 142430 117988 142462
rect 117982 142398 117983 142430
rect 117917 142397 117983 142398
rect 114376 133182 114382 133214
rect 109414 133150 109415 133182
rect 109349 133149 109415 133150
rect 114381 133150 114382 133182
rect 114446 133182 114452 133214
rect 119272 133214 119348 144100
rect 119680 142870 119756 142876
rect 119680 142806 119686 142870
rect 119750 142806 119756 142870
rect 119680 142462 119756 142806
rect 119680 142430 119686 142462
rect 119685 142398 119686 142430
rect 119750 142430 119756 142462
rect 121312 142870 121388 142876
rect 121312 142806 121318 142870
rect 121382 142806 121388 142870
rect 121312 142462 121388 142806
rect 121312 142430 121318 142462
rect 119750 142398 119751 142430
rect 119685 142397 119751 142398
rect 121317 142398 121318 142430
rect 121382 142430 121388 142462
rect 122944 142870 123020 142876
rect 122944 142806 122950 142870
rect 123014 142806 123020 142870
rect 122944 142462 123020 142806
rect 122944 142430 122950 142462
rect 121382 142398 121383 142430
rect 121317 142397 121383 142398
rect 122949 142398 122950 142430
rect 123014 142430 123020 142462
rect 123014 142398 123015 142430
rect 122949 142397 123015 142398
rect 119272 133182 119278 133214
rect 114446 133150 114447 133182
rect 114381 133149 114447 133150
rect 119277 133150 119278 133182
rect 119342 133182 119348 133214
rect 124304 133214 124380 144100
rect 124712 142870 124788 142876
rect 124712 142806 124718 142870
rect 124782 142806 124788 142870
rect 124712 142462 124788 142806
rect 124712 142430 124718 142462
rect 124717 142398 124718 142430
rect 124782 142430 124788 142462
rect 126208 142870 126284 142876
rect 126208 142806 126214 142870
rect 126278 142806 126284 142870
rect 126208 142462 126284 142806
rect 126208 142430 126214 142462
rect 124782 142398 124783 142430
rect 124717 142397 124783 142398
rect 126213 142398 126214 142430
rect 126278 142430 126284 142462
rect 127976 142870 128052 142876
rect 127976 142806 127982 142870
rect 128046 142806 128052 142870
rect 127976 142462 128052 142806
rect 127976 142430 127982 142462
rect 126278 142398 126279 142430
rect 126213 142397 126279 142398
rect 127981 142398 127982 142430
rect 128046 142430 128052 142462
rect 128046 142398 128047 142430
rect 127981 142397 128047 142398
rect 124304 133182 124310 133214
rect 119342 133150 119343 133182
rect 119277 133149 119343 133150
rect 124309 133150 124310 133182
rect 124374 133182 124380 133214
rect 129336 133214 129412 144100
rect 129608 142870 129684 142876
rect 129608 142806 129614 142870
rect 129678 142806 129684 142870
rect 129608 142462 129684 142806
rect 129608 142430 129614 142462
rect 129613 142398 129614 142430
rect 129678 142430 129684 142462
rect 131376 142870 131452 142876
rect 131376 142806 131382 142870
rect 131446 142806 131452 142870
rect 131376 142462 131452 142806
rect 131376 142430 131382 142462
rect 129678 142398 129679 142430
rect 129613 142397 129679 142398
rect 131381 142398 131382 142430
rect 131446 142430 131452 142462
rect 133144 142870 133220 142876
rect 133144 142806 133150 142870
rect 133214 142806 133220 142870
rect 133144 142462 133220 142806
rect 133144 142430 133150 142462
rect 131446 142398 131447 142430
rect 131381 142397 131447 142398
rect 133149 142398 133150 142430
rect 133214 142430 133220 142462
rect 133214 142398 133215 142430
rect 133149 142397 133215 142398
rect 129336 133182 129342 133214
rect 124374 133150 124375 133182
rect 124309 133149 124375 133150
rect 129341 133150 129342 133182
rect 129406 133182 129412 133214
rect 134368 133214 134444 144100
rect 134640 142870 134716 142876
rect 134640 142806 134646 142870
rect 134710 142806 134716 142870
rect 134640 142462 134716 142806
rect 134640 142430 134646 142462
rect 134645 142398 134646 142430
rect 134710 142430 134716 142462
rect 136408 142870 136484 142876
rect 136408 142806 136414 142870
rect 136478 142806 136484 142870
rect 136408 142462 136484 142806
rect 136408 142430 136414 142462
rect 134710 142398 134711 142430
rect 134645 142397 134711 142398
rect 136413 142398 136414 142430
rect 136478 142430 136484 142462
rect 138176 142870 138252 142876
rect 138176 142806 138182 142870
rect 138246 142806 138252 142870
rect 138176 142462 138252 142806
rect 138176 142430 138182 142462
rect 136478 142398 136479 142430
rect 136413 142397 136479 142398
rect 138181 142398 138182 142430
rect 138246 142430 138252 142462
rect 138246 142398 138247 142430
rect 138181 142397 138247 142398
rect 134368 133182 134374 133214
rect 129406 133150 129407 133182
rect 129341 133149 129407 133150
rect 134373 133150 134374 133182
rect 134438 133182 134444 133214
rect 139400 133214 139476 144100
rect 139672 142870 139748 142876
rect 139672 142806 139678 142870
rect 139742 142806 139748 142870
rect 139672 142462 139748 142806
rect 139672 142430 139678 142462
rect 139677 142398 139678 142430
rect 139742 142430 139748 142462
rect 141440 142870 141516 142876
rect 141440 142806 141446 142870
rect 141510 142806 141516 142870
rect 141440 142462 141516 142806
rect 141440 142430 141446 142462
rect 139742 142398 139743 142430
rect 139677 142397 139743 142398
rect 141445 142398 141446 142430
rect 141510 142430 141516 142462
rect 143208 142870 143284 142876
rect 143208 142806 143214 142870
rect 143278 142806 143284 142870
rect 143208 142462 143284 142806
rect 143208 142430 143214 142462
rect 141510 142398 141511 142430
rect 141445 142397 141511 142398
rect 143213 142398 143214 142430
rect 143278 142430 143284 142462
rect 143278 142398 143279 142430
rect 143213 142397 143279 142398
rect 139400 133182 139406 133214
rect 134438 133150 134439 133182
rect 134373 133149 134439 133150
rect 139405 133150 139406 133182
rect 139470 133182 139476 133214
rect 144296 133214 144372 144100
rect 144704 142870 144780 142876
rect 144704 142806 144710 142870
rect 144774 142806 144780 142870
rect 144704 142462 144780 142806
rect 144704 142430 144710 142462
rect 144709 142398 144710 142430
rect 144774 142430 144780 142462
rect 146472 142870 146548 142876
rect 146472 142806 146478 142870
rect 146542 142806 146548 142870
rect 146472 142462 146548 142806
rect 146472 142430 146478 142462
rect 144774 142398 144775 142430
rect 144709 142397 144775 142398
rect 146477 142398 146478 142430
rect 146542 142430 146548 142462
rect 148104 142870 148180 142876
rect 148104 142806 148110 142870
rect 148174 142806 148180 142870
rect 148104 142462 148180 142806
rect 148104 142430 148110 142462
rect 146542 142398 146543 142430
rect 146477 142397 146543 142398
rect 148109 142398 148110 142430
rect 148174 142430 148180 142462
rect 148174 142398 148175 142430
rect 148109 142397 148175 142398
rect 144296 133182 144302 133214
rect 139470 133150 139471 133182
rect 139405 133149 139471 133150
rect 144301 133150 144302 133182
rect 144366 133182 144372 133214
rect 149328 133214 149404 144100
rect 149736 142870 149812 142876
rect 149736 142806 149742 142870
rect 149806 142806 149812 142870
rect 149736 142462 149812 142806
rect 149736 142430 149742 142462
rect 149741 142398 149742 142430
rect 149806 142430 149812 142462
rect 151640 142870 151716 142876
rect 151640 142806 151646 142870
rect 151710 142806 151716 142870
rect 151640 142462 151716 142806
rect 151640 142430 151646 142462
rect 149806 142398 149807 142430
rect 149741 142397 149807 142398
rect 151645 142398 151646 142430
rect 151710 142430 151716 142462
rect 153136 142870 153212 142876
rect 153136 142806 153142 142870
rect 153206 142806 153212 142870
rect 153136 142462 153212 142806
rect 153136 142430 153142 142462
rect 151710 142398 151711 142430
rect 151645 142397 151711 142398
rect 153141 142398 153142 142430
rect 153206 142430 153212 142462
rect 153206 142398 153207 142430
rect 153141 142397 153207 142398
rect 149328 133182 149334 133214
rect 144366 133150 144367 133182
rect 144301 133149 144367 133150
rect 149333 133150 149334 133182
rect 149398 133182 149404 133214
rect 154360 133214 154436 144100
rect 154768 142870 154844 142876
rect 154768 142806 154774 142870
rect 154838 142806 154844 142870
rect 154768 142462 154844 142806
rect 154768 142430 154774 142462
rect 154773 142398 154774 142430
rect 154838 142430 154844 142462
rect 156672 142870 156748 142876
rect 156672 142806 156678 142870
rect 156742 142806 156748 142870
rect 156672 142462 156748 142806
rect 156672 142430 156678 142462
rect 154838 142398 154839 142430
rect 154773 142397 154839 142398
rect 156677 142398 156678 142430
rect 156742 142430 156748 142462
rect 158168 142870 158244 142876
rect 158168 142806 158174 142870
rect 158238 142806 158244 142870
rect 158168 142462 158244 142806
rect 158168 142430 158174 142462
rect 156742 142398 156743 142430
rect 156677 142397 156743 142398
rect 158173 142398 158174 142430
rect 158238 142430 158244 142462
rect 158238 142398 158239 142430
rect 158173 142397 158239 142398
rect 154360 133182 154366 133214
rect 149398 133150 149399 133182
rect 149333 133149 149399 133150
rect 154365 133150 154366 133182
rect 154430 133182 154436 133214
rect 159392 133214 159468 144100
rect 159936 142870 160012 142876
rect 159936 142806 159942 142870
rect 160006 142806 160012 142870
rect 159936 142462 160012 142806
rect 159936 142430 159942 142462
rect 159941 142398 159942 142430
rect 160006 142430 160012 142462
rect 161704 142870 161780 142876
rect 161704 142806 161710 142870
rect 161774 142806 161780 142870
rect 161704 142462 161780 142806
rect 161704 142430 161710 142462
rect 160006 142398 160007 142430
rect 159941 142397 160007 142398
rect 161709 142398 161710 142430
rect 161774 142430 161780 142462
rect 163200 142870 163276 142876
rect 163200 142806 163206 142870
rect 163270 142806 163276 142870
rect 163200 142462 163276 142806
rect 163200 142430 163206 142462
rect 161774 142398 161775 142430
rect 161709 142397 161775 142398
rect 163205 142398 163206 142430
rect 163270 142430 163276 142462
rect 163270 142398 163271 142430
rect 163205 142397 163271 142398
rect 159392 133182 159398 133214
rect 154430 133150 154431 133182
rect 154365 133149 154431 133150
rect 159397 133150 159398 133182
rect 159462 133182 159468 133214
rect 164424 133214 164500 144100
rect 164968 142870 165044 142876
rect 164968 142806 164974 142870
rect 165038 142806 165044 142870
rect 164968 142462 165044 142806
rect 164968 142430 164974 142462
rect 164973 142398 164974 142430
rect 165038 142430 165044 142462
rect 166600 142870 166676 142876
rect 166600 142806 166606 142870
rect 166670 142806 166676 142870
rect 166600 142462 166676 142806
rect 166600 142430 166606 142462
rect 165038 142398 165039 142430
rect 164973 142397 165039 142398
rect 166605 142398 166606 142430
rect 166670 142430 166676 142462
rect 168232 142870 168308 142876
rect 168232 142806 168238 142870
rect 168302 142806 168308 142870
rect 168232 142462 168308 142806
rect 168232 142430 168238 142462
rect 166670 142398 166671 142430
rect 166605 142397 166671 142398
rect 168237 142398 168238 142430
rect 168302 142430 168308 142462
rect 168302 142398 168303 142430
rect 168237 142397 168303 142398
rect 164424 133182 164430 133214
rect 159462 133150 159463 133182
rect 159397 133149 159463 133150
rect 164429 133150 164430 133182
rect 164494 133182 164500 133214
rect 169184 133214 169260 144100
rect 170136 142870 170212 142876
rect 170136 142806 170142 142870
rect 170206 142806 170212 142870
rect 170136 142462 170212 142806
rect 170136 142430 170142 142462
rect 170141 142398 170142 142430
rect 170206 142430 170212 142462
rect 171632 142870 171708 142876
rect 171632 142806 171638 142870
rect 171702 142806 171708 142870
rect 171632 142462 171708 142806
rect 171632 142430 171638 142462
rect 170206 142398 170207 142430
rect 170141 142397 170207 142398
rect 171637 142398 171638 142430
rect 171702 142430 171708 142462
rect 173400 142870 173476 142876
rect 173400 142806 173406 142870
rect 173470 142806 173476 142870
rect 173400 142462 173476 142806
rect 173400 142430 173406 142462
rect 171702 142398 171703 142430
rect 171637 142397 171703 142398
rect 173405 142398 173406 142430
rect 173470 142430 173476 142462
rect 173470 142398 173471 142430
rect 173405 142397 173471 142398
rect 169184 133182 169190 133214
rect 164494 133150 164495 133182
rect 164429 133149 164495 133150
rect 169189 133150 169190 133182
rect 169254 133182 169260 133214
rect 174216 133214 174292 144100
rect 175168 142870 175244 142876
rect 175168 142806 175174 142870
rect 175238 142806 175244 142870
rect 175168 142462 175244 142806
rect 175168 142430 175174 142462
rect 175173 142398 175174 142430
rect 175238 142430 175244 142462
rect 176664 142870 176740 142876
rect 176664 142806 176670 142870
rect 176734 142806 176740 142870
rect 176664 142462 176740 142806
rect 176664 142430 176670 142462
rect 175238 142398 175239 142430
rect 175173 142397 175239 142398
rect 176669 142398 176670 142430
rect 176734 142430 176740 142462
rect 178432 142870 178508 142876
rect 178432 142806 178438 142870
rect 178502 142806 178508 142870
rect 178432 142462 178508 142806
rect 178432 142430 178438 142462
rect 176734 142398 176735 142430
rect 176669 142397 176735 142398
rect 178437 142398 178438 142430
rect 178502 142430 178508 142462
rect 178502 142398 178503 142430
rect 178437 142397 178503 142398
rect 174216 133182 174222 133214
rect 169254 133150 169255 133182
rect 169189 133149 169255 133150
rect 174221 133150 174222 133182
rect 174286 133182 174292 133214
rect 179384 133214 179460 144100
rect 180200 142870 180276 142876
rect 180200 142806 180206 142870
rect 180270 142806 180276 142870
rect 180200 142462 180276 142806
rect 180200 142430 180206 142462
rect 180205 142398 180206 142430
rect 180270 142430 180276 142462
rect 181696 142870 181772 142876
rect 181696 142806 181702 142870
rect 181766 142806 181772 142870
rect 181696 142462 181772 142806
rect 181696 142430 181702 142462
rect 180270 142398 180271 142430
rect 180205 142397 180271 142398
rect 181701 142398 181702 142430
rect 181766 142430 181772 142462
rect 183328 142870 183404 142876
rect 183328 142806 183334 142870
rect 183398 142806 183404 142870
rect 183328 142462 183404 142806
rect 183328 142430 183334 142462
rect 181766 142398 181767 142430
rect 181701 142397 181767 142398
rect 183333 142398 183334 142430
rect 183398 142430 183404 142462
rect 183398 142398 183399 142430
rect 183333 142397 183399 142398
rect 179384 133182 179390 133214
rect 174286 133150 174287 133182
rect 174221 133149 174287 133150
rect 179389 133150 179390 133182
rect 179454 133182 179460 133214
rect 184280 133214 184356 144100
rect 198152 143550 198228 143556
rect 198152 143486 198158 143550
rect 198222 143486 198228 143550
rect 185096 142870 185172 142876
rect 185096 142806 185102 142870
rect 185166 142806 185172 142870
rect 185096 142462 185172 142806
rect 185096 142430 185102 142462
rect 185101 142398 185102 142430
rect 185166 142430 185172 142462
rect 186728 142870 186804 142876
rect 186728 142806 186734 142870
rect 186798 142806 186804 142870
rect 186728 142462 186804 142806
rect 186728 142430 186734 142462
rect 185166 142398 185167 142430
rect 185101 142397 185167 142398
rect 186733 142398 186734 142430
rect 186798 142430 186804 142462
rect 188632 142870 188708 142876
rect 188632 142806 188638 142870
rect 188702 142806 188708 142870
rect 188632 142462 188708 142806
rect 188632 142430 188638 142462
rect 186798 142398 186799 142430
rect 186733 142397 186799 142398
rect 188637 142398 188638 142430
rect 188702 142430 188708 142462
rect 190128 142870 190204 142876
rect 190128 142806 190134 142870
rect 190198 142806 190204 142870
rect 190128 142462 190204 142806
rect 190128 142430 190134 142462
rect 188702 142398 188703 142430
rect 188637 142397 188703 142398
rect 190133 142398 190134 142430
rect 190198 142430 190204 142462
rect 191896 142870 191972 142876
rect 191896 142806 191902 142870
rect 191966 142806 191972 142870
rect 191896 142462 191972 142806
rect 191896 142430 191902 142462
rect 190198 142398 190199 142430
rect 190133 142397 190199 142398
rect 191901 142398 191902 142430
rect 191966 142430 191972 142462
rect 193664 142870 193740 142876
rect 193664 142806 193670 142870
rect 193734 142806 193740 142870
rect 193664 142462 193740 142806
rect 193664 142430 193670 142462
rect 191966 142398 191967 142430
rect 191901 142397 191967 142398
rect 193669 142398 193670 142430
rect 193734 142430 193740 142462
rect 195160 142870 195236 142876
rect 195160 142806 195166 142870
rect 195230 142806 195236 142870
rect 195160 142462 195236 142806
rect 195160 142430 195166 142462
rect 193734 142398 193735 142430
rect 193669 142397 193735 142398
rect 195165 142398 195166 142430
rect 195230 142430 195236 142462
rect 196928 142870 197004 142876
rect 196928 142806 196934 142870
rect 196998 142806 197004 142870
rect 196928 142462 197004 142806
rect 196928 142430 196934 142462
rect 195230 142398 195231 142430
rect 195165 142397 195231 142398
rect 196933 142398 196934 142430
rect 196998 142430 197004 142462
rect 196998 142398 196999 142430
rect 196933 142397 196999 142398
rect 198152 140694 198228 143486
rect 198152 140662 198158 140694
rect 198157 140630 198158 140662
rect 198222 140662 198228 140694
rect 198288 141918 198364 141924
rect 198288 141854 198294 141918
rect 198358 141854 198364 141918
rect 198222 140630 198223 140662
rect 198157 140629 198223 140630
rect 198152 140558 198228 140564
rect 198152 140494 198158 140558
rect 198222 140494 198228 140558
rect 197885 139742 197951 139743
rect 197885 139710 197886 139742
rect 197880 139678 197886 139710
rect 197950 139710 197951 139742
rect 197950 139678 197956 139710
rect 196661 138382 196727 138383
rect 196661 138350 196662 138382
rect 196656 138318 196662 138350
rect 196726 138350 196727 138382
rect 196726 138318 196732 138350
rect 196656 135662 196732 138318
rect 197880 137158 197956 139678
rect 198152 138518 198228 140494
rect 198288 139878 198364 141854
rect 198560 141510 198636 144100
rect 198832 142870 198908 142876
rect 198832 142806 198838 142870
rect 198902 142806 198908 142870
rect 198832 142462 198908 142806
rect 198832 142430 198838 142462
rect 198837 142398 198838 142430
rect 198902 142430 198908 142462
rect 198902 142398 198903 142430
rect 198837 142397 198903 142398
rect 199245 142326 199311 142327
rect 199245 142294 199246 142326
rect 199240 142262 199246 142294
rect 199310 142294 199311 142326
rect 199310 142262 199316 142294
rect 199240 142054 199316 142262
rect 199240 141990 199246 142054
rect 199310 141990 199316 142054
rect 199240 141984 199316 141990
rect 198560 141478 198566 141510
rect 198565 141446 198566 141478
rect 198630 141478 198636 141510
rect 199920 141510 199996 144100
rect 200192 142870 200268 142876
rect 200192 142806 200198 142870
rect 200262 142806 200268 142870
rect 200192 142462 200268 142806
rect 200192 142430 200198 142462
rect 200197 142398 200198 142430
rect 200262 142430 200268 142462
rect 200262 142398 200263 142430
rect 200197 142397 200263 142398
rect 200469 142326 200535 142327
rect 200469 142294 200470 142326
rect 200464 142262 200470 142294
rect 200534 142294 200535 142326
rect 200534 142262 200540 142294
rect 200464 142054 200540 142262
rect 200464 141990 200470 142054
rect 200534 141990 200540 142054
rect 200464 141984 200540 141990
rect 199920 141478 199926 141510
rect 198630 141446 198631 141478
rect 198565 141445 198631 141446
rect 199925 141446 199926 141478
rect 199990 141478 199996 141510
rect 201008 141510 201084 144100
rect 218144 143822 218492 143828
rect 218144 143758 218150 143822
rect 218214 143758 218286 143822
rect 218350 143758 218422 143822
rect 218486 143758 218492 143822
rect 218144 143686 218492 143758
rect 218144 143622 218150 143686
rect 218214 143622 218286 143686
rect 218350 143622 218422 143686
rect 218486 143622 218492 143686
rect 218144 143550 218492 143622
rect 218144 143486 218150 143550
rect 218214 143486 218286 143550
rect 218350 143486 218422 143550
rect 218486 143486 218492 143550
rect 217464 143142 217812 143148
rect 217464 143078 217470 143142
rect 217534 143078 217606 143142
rect 217670 143078 217742 143142
rect 217806 143078 217812 143142
rect 217464 143006 217812 143078
rect 217464 142942 217470 143006
rect 217534 142942 217606 143006
rect 217670 142942 217742 143006
rect 217806 142942 217812 143006
rect 201960 142870 202036 142876
rect 201960 142806 201966 142870
rect 202030 142806 202036 142870
rect 201960 142462 202036 142806
rect 201960 142430 201966 142462
rect 201965 142398 201966 142430
rect 202030 142430 202036 142462
rect 203592 142870 203668 142876
rect 203592 142806 203598 142870
rect 203662 142806 203668 142870
rect 203592 142462 203668 142806
rect 203592 142430 203598 142462
rect 202030 142398 202031 142430
rect 201965 142397 202031 142398
rect 203597 142398 203598 142430
rect 203662 142430 203668 142462
rect 205224 142870 205300 142876
rect 205224 142806 205230 142870
rect 205294 142806 205300 142870
rect 205224 142462 205300 142806
rect 205224 142430 205230 142462
rect 203662 142398 203663 142430
rect 203597 142397 203663 142398
rect 205229 142398 205230 142430
rect 205294 142430 205300 142462
rect 206856 142870 206932 142876
rect 206856 142806 206862 142870
rect 206926 142806 206932 142870
rect 206856 142462 206932 142806
rect 206856 142430 206862 142462
rect 205294 142398 205295 142430
rect 205229 142397 205295 142398
rect 206861 142398 206862 142430
rect 206926 142430 206932 142462
rect 208624 142870 208700 142876
rect 208624 142806 208630 142870
rect 208694 142806 208700 142870
rect 208624 142462 208700 142806
rect 208624 142430 208630 142462
rect 206926 142398 206927 142430
rect 206861 142397 206927 142398
rect 208629 142398 208630 142430
rect 208694 142430 208700 142462
rect 210392 142870 210468 142876
rect 210392 142806 210398 142870
rect 210462 142806 210468 142870
rect 210392 142462 210468 142806
rect 210392 142430 210398 142462
rect 208694 142398 208695 142430
rect 208629 142397 208695 142398
rect 210397 142398 210398 142430
rect 210462 142430 210468 142462
rect 212024 142870 212100 142876
rect 212024 142806 212030 142870
rect 212094 142806 212100 142870
rect 212024 142462 212100 142806
rect 212024 142430 212030 142462
rect 210462 142398 210463 142430
rect 210397 142397 210463 142398
rect 212029 142398 212030 142430
rect 212094 142430 212100 142462
rect 213656 142870 213732 142876
rect 213656 142806 213662 142870
rect 213726 142806 213732 142870
rect 213656 142462 213732 142806
rect 213656 142430 213662 142462
rect 212094 142398 212095 142430
rect 212029 142397 212095 142398
rect 213661 142398 213662 142430
rect 213726 142430 213732 142462
rect 215424 142870 215500 142876
rect 215424 142806 215430 142870
rect 215494 142806 215500 142870
rect 215424 142462 215500 142806
rect 215424 142430 215430 142462
rect 213726 142398 213727 142430
rect 213661 142397 213727 142398
rect 215429 142398 215430 142430
rect 215494 142430 215500 142462
rect 217464 142870 217812 142942
rect 217464 142806 217470 142870
rect 217534 142806 217606 142870
rect 217670 142806 217742 142870
rect 217806 142806 217812 142870
rect 215494 142398 215495 142430
rect 215429 142397 215495 142398
rect 201008 141478 201014 141510
rect 199990 141446 199991 141478
rect 199925 141445 199991 141446
rect 201013 141446 201014 141478
rect 201078 141478 201084 141510
rect 217464 141782 217812 142806
rect 217464 141718 217470 141782
rect 217534 141718 217812 141782
rect 201078 141446 201079 141478
rect 201013 141445 201079 141446
rect 198288 139846 198294 139878
rect 198293 139814 198294 139846
rect 198358 139846 198364 139878
rect 217464 140014 217812 141718
rect 217464 139950 217470 140014
rect 217534 139950 217812 140014
rect 198358 139814 198359 139846
rect 198293 139813 198359 139814
rect 198152 138486 198158 138518
rect 198157 138454 198158 138486
rect 198222 138486 198228 138518
rect 198222 138454 198223 138486
rect 198157 138453 198223 138454
rect 197880 137094 197886 137158
rect 197950 137094 197956 137158
rect 197880 137088 197956 137094
rect 217464 138382 217812 139950
rect 217464 138318 217470 138382
rect 217534 138318 217812 138382
rect 196656 135598 196662 135662
rect 196726 135598 196732 135662
rect 196656 135592 196732 135598
rect 197880 136886 197956 136892
rect 197880 136822 197886 136886
rect 197950 136822 197956 136886
rect 197880 134302 197956 136822
rect 217464 136614 217812 138318
rect 217464 136550 217470 136614
rect 217534 136550 217812 136614
rect 198021 135526 198087 135527
rect 198021 135494 198022 135526
rect 197880 134270 197886 134302
rect 197885 134238 197886 134270
rect 197950 134270 197956 134302
rect 198016 135462 198022 135494
rect 198086 135494 198087 135526
rect 198086 135462 198092 135494
rect 197950 134238 197951 134270
rect 197885 134237 197951 134238
rect 184280 133182 184286 133214
rect 179454 133150 179455 133182
rect 179389 133149 179455 133150
rect 184285 133150 184286 133182
rect 184350 133182 184356 133214
rect 196656 134166 196732 134172
rect 196656 134102 196662 134166
rect 196726 134102 196732 134166
rect 184350 133150 184351 133182
rect 184285 133149 184351 133150
rect 29925 133078 29991 133079
rect 29925 133046 29926 133078
rect 29920 133014 29926 133046
rect 29990 133046 29991 133078
rect 34821 133078 34887 133079
rect 34821 133046 34822 133078
rect 29990 133014 29996 133046
rect 29784 132670 29860 132676
rect 29784 132606 29790 132670
rect 29854 132606 29860 132670
rect 29784 131990 29860 132606
rect 29784 131958 29790 131990
rect 29789 131926 29790 131958
rect 29854 131958 29860 131990
rect 29854 131926 29855 131958
rect 29789 131925 29855 131926
rect 952 131518 1230 131582
rect 1294 131518 1300 131582
rect 952 129814 1300 131518
rect 952 129750 1230 129814
rect 1294 129750 1300 129814
rect 952 128182 1300 129750
rect 29648 131854 29724 131860
rect 29648 131790 29654 131854
rect 29718 131790 29724 131854
rect 952 128118 1230 128182
rect 1294 128118 1300 128182
rect 952 126550 1300 128118
rect 952 126486 1230 126550
rect 1294 126486 1300 126550
rect 952 124918 1300 126486
rect 28832 128590 28908 128596
rect 28832 128526 28838 128590
rect 28902 128526 28908 128590
rect 28832 126414 28908 128526
rect 29648 127230 29724 131790
rect 29920 131310 29996 133014
rect 34816 133014 34822 133046
rect 34886 133046 34887 133078
rect 39853 133078 39919 133079
rect 39853 133046 39854 133078
rect 34886 133014 34892 133046
rect 34680 132670 34756 132676
rect 34680 132606 34686 132670
rect 34750 132606 34756 132670
rect 34680 131990 34756 132606
rect 34680 131958 34686 131990
rect 34685 131926 34686 131958
rect 34750 131958 34756 131990
rect 34750 131926 34751 131958
rect 34685 131925 34751 131926
rect 29920 131246 29926 131310
rect 29990 131246 29996 131310
rect 29920 131240 29996 131246
rect 34816 131310 34892 133014
rect 39848 133014 39854 133046
rect 39918 133046 39919 133078
rect 44885 133078 44951 133079
rect 44885 133046 44886 133078
rect 39918 133014 39924 133046
rect 39712 132670 39788 132676
rect 39712 132606 39718 132670
rect 39782 132606 39788 132670
rect 39712 131990 39788 132606
rect 39712 131958 39718 131990
rect 39717 131926 39718 131958
rect 39782 131958 39788 131990
rect 39782 131926 39783 131958
rect 39717 131925 39783 131926
rect 35773 131854 35839 131855
rect 35773 131822 35774 131854
rect 34816 131246 34822 131310
rect 34886 131246 34892 131310
rect 34816 131240 34892 131246
rect 35768 131790 35774 131822
rect 35838 131822 35839 131854
rect 39712 131854 39788 131860
rect 35838 131790 35844 131822
rect 29925 131174 29991 131175
rect 29925 131142 29926 131174
rect 29920 131110 29926 131142
rect 29990 131142 29991 131174
rect 34957 131174 35023 131175
rect 34957 131142 34958 131174
rect 29990 131110 29996 131142
rect 29920 128726 29996 131110
rect 29920 128662 29926 128726
rect 29990 128662 29996 128726
rect 29920 128656 29996 128662
rect 34952 131110 34958 131142
rect 35022 131142 35023 131174
rect 35022 131110 35028 131142
rect 34952 128726 35028 131110
rect 34952 128662 34958 128726
rect 35022 128662 35028 128726
rect 34952 128656 35028 128662
rect 29648 127198 29654 127230
rect 29653 127166 29654 127198
rect 29718 127198 29724 127230
rect 35768 127230 35844 131790
rect 29718 127166 29719 127198
rect 29653 127165 29719 127166
rect 35768 127166 35774 127230
rect 35838 127166 35844 127230
rect 39712 131790 39718 131854
rect 39782 131790 39788 131854
rect 39712 127230 39788 131790
rect 39848 131310 39924 133014
rect 44880 133014 44886 133046
rect 44950 133046 44951 133078
rect 49917 133078 49983 133079
rect 49917 133046 49918 133078
rect 44950 133014 44956 133046
rect 44744 132670 44820 132676
rect 44744 132606 44750 132670
rect 44814 132606 44820 132670
rect 44744 131990 44820 132606
rect 44744 131958 44750 131990
rect 44749 131926 44750 131958
rect 44814 131958 44820 131990
rect 44814 131926 44815 131958
rect 44749 131925 44815 131926
rect 39848 131246 39854 131310
rect 39918 131246 39924 131310
rect 39848 131240 39924 131246
rect 44336 131854 44412 131860
rect 44336 131790 44342 131854
rect 44406 131790 44412 131854
rect 39989 131174 40055 131175
rect 39989 131142 39990 131174
rect 39984 131110 39990 131142
rect 40054 131142 40055 131174
rect 40054 131110 40060 131142
rect 39984 128726 40060 131110
rect 39984 128662 39990 128726
rect 40054 128662 40060 128726
rect 39984 128656 40060 128662
rect 39712 127198 39718 127230
rect 35768 127160 35844 127166
rect 39717 127166 39718 127198
rect 39782 127198 39788 127230
rect 44336 127230 44412 131790
rect 44880 131310 44956 133014
rect 49912 133014 49918 133046
rect 49982 133046 49983 133078
rect 54813 133078 54879 133079
rect 54813 133046 54814 133078
rect 49982 133014 49988 133046
rect 49640 132670 49716 132676
rect 49640 132606 49646 132670
rect 49710 132606 49716 132670
rect 49640 131990 49716 132606
rect 49640 131958 49646 131990
rect 49645 131926 49646 131958
rect 49710 131958 49716 131990
rect 49710 131926 49711 131958
rect 49645 131925 49711 131926
rect 44880 131246 44886 131310
rect 44950 131246 44956 131310
rect 44880 131240 44956 131246
rect 49912 131310 49988 133014
rect 54808 133014 54814 133046
rect 54878 133046 54879 133078
rect 59845 133078 59911 133079
rect 59845 133046 59846 133078
rect 54878 133014 54884 133046
rect 54672 132670 54748 132676
rect 54672 132606 54678 132670
rect 54742 132606 54748 132670
rect 54672 131990 54748 132606
rect 54672 131958 54678 131990
rect 54677 131926 54678 131958
rect 54742 131958 54748 131990
rect 54742 131926 54743 131958
rect 54677 131925 54743 131926
rect 50733 131854 50799 131855
rect 50733 131822 50734 131854
rect 49912 131246 49918 131310
rect 49982 131246 49988 131310
rect 49912 131240 49988 131246
rect 50728 131790 50734 131822
rect 50798 131822 50799 131854
rect 54672 131854 54748 131860
rect 50798 131790 50804 131822
rect 44885 131174 44951 131175
rect 44885 131142 44886 131174
rect 44880 131110 44886 131142
rect 44950 131142 44951 131174
rect 49917 131174 49983 131175
rect 49917 131142 49918 131174
rect 44950 131110 44956 131142
rect 44880 128726 44956 131110
rect 44880 128662 44886 128726
rect 44950 128662 44956 128726
rect 44880 128656 44956 128662
rect 49912 131110 49918 131142
rect 49982 131142 49983 131174
rect 49982 131110 49988 131142
rect 49912 128726 49988 131110
rect 49912 128662 49918 128726
rect 49982 128662 49988 128726
rect 49912 128656 49988 128662
rect 44336 127198 44342 127230
rect 39782 127166 39783 127198
rect 39717 127165 39783 127166
rect 44341 127166 44342 127198
rect 44406 127198 44412 127230
rect 50728 127230 50804 131790
rect 44406 127166 44407 127198
rect 44341 127165 44407 127166
rect 50728 127166 50734 127230
rect 50798 127166 50804 127230
rect 54672 131790 54678 131854
rect 54742 131790 54748 131854
rect 54672 127230 54748 131790
rect 54808 131310 54884 133014
rect 59840 133014 59846 133046
rect 59910 133046 59911 133078
rect 64741 133078 64807 133079
rect 64741 133046 64742 133078
rect 59910 133014 59916 133046
rect 59704 132670 59780 132676
rect 59704 132606 59710 132670
rect 59774 132606 59780 132670
rect 59704 131990 59780 132606
rect 59704 131958 59710 131990
rect 59709 131926 59710 131958
rect 59774 131958 59780 131990
rect 59774 131926 59775 131958
rect 59709 131925 59775 131926
rect 54808 131246 54814 131310
rect 54878 131246 54884 131310
rect 54808 131240 54884 131246
rect 59840 131310 59916 133014
rect 64736 133014 64742 133046
rect 64806 133046 64807 133078
rect 69909 133078 69975 133079
rect 69909 133046 69910 133078
rect 64806 133014 64812 133046
rect 60797 131854 60863 131855
rect 60797 131822 60798 131854
rect 59840 131246 59846 131310
rect 59910 131246 59916 131310
rect 59840 131240 59916 131246
rect 60792 131790 60798 131822
rect 60862 131822 60863 131854
rect 64600 131854 64676 131860
rect 60862 131790 60868 131822
rect 54808 131174 54884 131180
rect 54808 131110 54814 131174
rect 54878 131110 54884 131174
rect 59981 131174 60047 131175
rect 59981 131142 59982 131174
rect 54808 128726 54884 131110
rect 54808 128694 54814 128726
rect 54813 128662 54814 128694
rect 54878 128694 54884 128726
rect 59976 131110 59982 131142
rect 60046 131142 60047 131174
rect 60046 131110 60052 131142
rect 59976 128726 60052 131110
rect 54878 128662 54879 128694
rect 54813 128661 54879 128662
rect 59976 128662 59982 128726
rect 60046 128662 60052 128726
rect 59976 128656 60052 128662
rect 54672 127198 54678 127230
rect 50728 127160 50804 127166
rect 54677 127166 54678 127198
rect 54742 127198 54748 127230
rect 60792 127230 60868 131790
rect 54742 127166 54743 127198
rect 54677 127165 54743 127166
rect 60792 127166 60798 127230
rect 60862 127166 60868 127230
rect 64600 131790 64606 131854
rect 64670 131790 64676 131854
rect 64600 127230 64676 131790
rect 64736 131310 64812 133014
rect 69904 133014 69910 133046
rect 69974 133046 69975 133078
rect 74805 133078 74871 133079
rect 74805 133046 74806 133078
rect 69974 133014 69980 133046
rect 64872 132670 64948 132676
rect 64872 132606 64878 132670
rect 64942 132606 64948 132670
rect 64872 131990 64948 132606
rect 64872 131958 64878 131990
rect 64877 131926 64878 131958
rect 64942 131958 64948 131990
rect 69768 132670 69844 132676
rect 69768 132606 69774 132670
rect 69838 132606 69844 132670
rect 69768 131990 69844 132606
rect 69768 131958 69774 131990
rect 64942 131926 64943 131958
rect 64877 131925 64943 131926
rect 69773 131926 69774 131958
rect 69838 131958 69844 131990
rect 69838 131926 69839 131958
rect 69773 131925 69839 131926
rect 64736 131246 64742 131310
rect 64806 131246 64812 131310
rect 64736 131240 64812 131246
rect 69224 131854 69300 131860
rect 69224 131790 69230 131854
rect 69294 131790 69300 131854
rect 64877 131174 64943 131175
rect 64877 131142 64878 131174
rect 64872 131110 64878 131142
rect 64942 131142 64943 131174
rect 64942 131110 64948 131142
rect 64872 128726 64948 131110
rect 64872 128662 64878 128726
rect 64942 128662 64948 128726
rect 64872 128656 64948 128662
rect 64600 127198 64606 127230
rect 60792 127160 60868 127166
rect 64605 127166 64606 127198
rect 64670 127198 64676 127230
rect 69224 127230 69300 131790
rect 69904 131310 69980 133014
rect 74800 133014 74806 133046
rect 74870 133046 74871 133078
rect 79837 133078 79903 133079
rect 79837 133046 79838 133078
rect 74870 133014 74876 133046
rect 74664 132670 74740 132676
rect 74664 132606 74670 132670
rect 74734 132606 74740 132670
rect 74664 131990 74740 132606
rect 74664 131958 74670 131990
rect 74669 131926 74670 131958
rect 74734 131958 74740 131990
rect 74734 131926 74735 131958
rect 74669 131925 74735 131926
rect 69904 131246 69910 131310
rect 69974 131246 69980 131310
rect 69904 131240 69980 131246
rect 74664 131854 74740 131860
rect 74664 131790 74670 131854
rect 74734 131790 74740 131854
rect 69909 131174 69975 131175
rect 69909 131142 69910 131174
rect 69904 131110 69910 131142
rect 69974 131142 69975 131174
rect 69974 131110 69980 131142
rect 69904 128726 69980 131110
rect 69904 128662 69910 128726
rect 69974 128662 69980 128726
rect 69904 128656 69980 128662
rect 69224 127198 69230 127230
rect 64670 127166 64671 127198
rect 64605 127165 64671 127166
rect 69229 127166 69230 127198
rect 69294 127198 69300 127230
rect 74664 127230 74740 131790
rect 74800 131310 74876 133014
rect 79832 133014 79838 133046
rect 79902 133046 79903 133078
rect 84869 133078 84935 133079
rect 84869 133046 84870 133078
rect 79902 133014 79908 133046
rect 79696 132670 79772 132676
rect 79696 132606 79702 132670
rect 79766 132606 79772 132670
rect 79696 131990 79772 132606
rect 79696 131958 79702 131990
rect 79701 131926 79702 131958
rect 79766 131958 79772 131990
rect 79766 131926 79767 131958
rect 79701 131925 79767 131926
rect 74800 131246 74806 131310
rect 74870 131246 74876 131310
rect 74800 131240 74876 131246
rect 79288 131854 79364 131860
rect 79288 131790 79294 131854
rect 79358 131790 79364 131854
rect 74941 131174 75007 131175
rect 74941 131142 74942 131174
rect 74936 131110 74942 131142
rect 75006 131142 75007 131174
rect 75006 131110 75012 131142
rect 74936 128726 75012 131110
rect 74936 128662 74942 128726
rect 75006 128662 75012 128726
rect 74936 128656 75012 128662
rect 74664 127198 74670 127230
rect 69294 127166 69295 127198
rect 69229 127165 69295 127166
rect 74669 127166 74670 127198
rect 74734 127198 74740 127230
rect 79288 127230 79364 131790
rect 79832 131310 79908 133014
rect 84864 133014 84870 133046
rect 84934 133046 84935 133078
rect 89901 133078 89967 133079
rect 89901 133046 89902 133078
rect 84934 133014 84940 133046
rect 84728 132670 84804 132676
rect 84728 132606 84734 132670
rect 84798 132606 84804 132670
rect 84728 131990 84804 132606
rect 84728 131958 84734 131990
rect 84733 131926 84734 131958
rect 84798 131958 84804 131990
rect 84798 131926 84799 131958
rect 84733 131925 84799 131926
rect 79832 131246 79838 131310
rect 79902 131246 79908 131310
rect 79832 131240 79908 131246
rect 84184 131854 84260 131860
rect 84184 131790 84190 131854
rect 84254 131790 84260 131854
rect 79837 131174 79903 131175
rect 79837 131142 79838 131174
rect 79832 131110 79838 131142
rect 79902 131142 79903 131174
rect 79902 131110 79908 131142
rect 79832 128726 79908 131110
rect 79832 128662 79838 128726
rect 79902 128662 79908 128726
rect 79832 128656 79908 128662
rect 79288 127198 79294 127230
rect 74734 127166 74735 127198
rect 74669 127165 74735 127166
rect 79293 127166 79294 127198
rect 79358 127198 79364 127230
rect 84184 127230 84260 131790
rect 84864 131310 84940 133014
rect 89896 133014 89902 133046
rect 89966 133046 89967 133078
rect 94933 133078 94999 133079
rect 94933 133046 94934 133078
rect 89966 133014 89972 133046
rect 89760 132670 89836 132676
rect 89760 132606 89766 132670
rect 89830 132606 89836 132670
rect 89760 131990 89836 132606
rect 89760 131958 89766 131990
rect 89765 131926 89766 131958
rect 89830 131958 89836 131990
rect 89830 131926 89831 131958
rect 89765 131925 89831 131926
rect 84864 131246 84870 131310
rect 84934 131246 84940 131310
rect 84864 131240 84940 131246
rect 89624 131854 89700 131860
rect 89624 131790 89630 131854
rect 89694 131790 89700 131854
rect 84869 131174 84935 131175
rect 84869 131142 84870 131174
rect 84864 131110 84870 131142
rect 84934 131142 84935 131174
rect 84934 131110 84940 131142
rect 84864 128726 84940 131110
rect 84864 128662 84870 128726
rect 84934 128662 84940 128726
rect 84864 128656 84940 128662
rect 84184 127198 84190 127230
rect 79358 127166 79359 127198
rect 79293 127165 79359 127166
rect 84189 127166 84190 127198
rect 84254 127198 84260 127230
rect 89624 127230 89700 131790
rect 89896 131310 89972 133014
rect 94928 133014 94934 133046
rect 94998 133046 94999 133078
rect 99829 133078 99895 133079
rect 99829 133046 99830 133078
rect 94998 133014 95004 133046
rect 94792 132670 94868 132676
rect 94792 132606 94798 132670
rect 94862 132606 94868 132670
rect 94792 131990 94868 132606
rect 94792 131958 94798 131990
rect 94797 131926 94798 131958
rect 94862 131958 94868 131990
rect 94862 131926 94863 131958
rect 94797 131925 94863 131926
rect 89896 131246 89902 131310
rect 89966 131246 89972 131310
rect 89896 131240 89972 131246
rect 94656 131854 94732 131860
rect 94656 131790 94662 131854
rect 94726 131790 94732 131854
rect 89901 131174 89967 131175
rect 89901 131142 89902 131174
rect 89896 131110 89902 131142
rect 89966 131142 89967 131174
rect 89966 131110 89972 131142
rect 89896 128726 89972 131110
rect 89896 128662 89902 128726
rect 89966 128662 89972 128726
rect 89896 128656 89972 128662
rect 89624 127198 89630 127230
rect 84254 127166 84255 127198
rect 84189 127165 84255 127166
rect 89629 127166 89630 127198
rect 89694 127198 89700 127230
rect 94656 127230 94732 131790
rect 94928 131310 95004 133014
rect 99824 133014 99830 133046
rect 99894 133046 99895 133078
rect 104725 133078 104791 133079
rect 104725 133046 104726 133078
rect 99894 133014 99900 133046
rect 99688 132670 99764 132676
rect 99688 132606 99694 132670
rect 99758 132606 99764 132670
rect 99688 131990 99764 132606
rect 99688 131958 99694 131990
rect 99693 131926 99694 131958
rect 99758 131958 99764 131990
rect 99758 131926 99759 131958
rect 99693 131925 99759 131926
rect 94928 131246 94934 131310
rect 94998 131246 95004 131310
rect 94928 131240 95004 131246
rect 99552 131854 99628 131860
rect 99552 131790 99558 131854
rect 99622 131790 99628 131854
rect 94933 131174 94999 131175
rect 94933 131142 94934 131174
rect 94928 131110 94934 131142
rect 94998 131142 94999 131174
rect 94998 131110 95004 131142
rect 94928 128726 95004 131110
rect 94928 128662 94934 128726
rect 94998 128662 95004 128726
rect 94928 128656 95004 128662
rect 94656 127198 94662 127230
rect 89694 127166 89695 127198
rect 89629 127165 89695 127166
rect 94661 127166 94662 127198
rect 94726 127198 94732 127230
rect 99552 127230 99628 131790
rect 99824 131310 99900 133014
rect 104720 133014 104726 133046
rect 104790 133046 104791 133078
rect 109893 133078 109959 133079
rect 109893 133046 109894 133078
rect 104790 133014 104796 133046
rect 104584 132670 104660 132676
rect 104584 132606 104590 132670
rect 104654 132606 104660 132670
rect 104584 131990 104660 132606
rect 104584 131958 104590 131990
rect 104589 131926 104590 131958
rect 104654 131958 104660 131990
rect 104654 131926 104655 131958
rect 104589 131925 104655 131926
rect 99824 131246 99830 131310
rect 99894 131246 99900 131310
rect 99824 131240 99900 131246
rect 104312 131854 104388 131860
rect 104312 131790 104318 131854
rect 104382 131790 104388 131854
rect 99829 131174 99895 131175
rect 99829 131142 99830 131174
rect 99824 131110 99830 131142
rect 99894 131142 99895 131174
rect 99894 131110 99900 131142
rect 99824 128726 99900 131110
rect 99824 128662 99830 128726
rect 99894 128662 99900 128726
rect 99824 128656 99900 128662
rect 99552 127198 99558 127230
rect 94726 127166 94727 127198
rect 94661 127165 94727 127166
rect 99557 127166 99558 127198
rect 99622 127198 99628 127230
rect 104312 127230 104388 131790
rect 104720 131310 104796 133014
rect 109888 133014 109894 133046
rect 109958 133046 109959 133078
rect 114789 133078 114855 133079
rect 114789 133046 114790 133078
rect 109958 133014 109964 133046
rect 109752 132670 109828 132676
rect 109752 132606 109758 132670
rect 109822 132606 109828 132670
rect 109752 131990 109828 132606
rect 109752 131958 109758 131990
rect 109757 131926 109758 131958
rect 109822 131958 109828 131990
rect 109822 131926 109823 131958
rect 109757 131925 109823 131926
rect 104720 131246 104726 131310
rect 104790 131246 104796 131310
rect 104720 131240 104796 131246
rect 109616 131854 109692 131860
rect 109616 131790 109622 131854
rect 109686 131790 109692 131854
rect 104861 131174 104927 131175
rect 104861 131142 104862 131174
rect 104856 131110 104862 131142
rect 104926 131142 104927 131174
rect 104926 131110 104932 131142
rect 104856 128726 104932 131110
rect 104856 128662 104862 128726
rect 104926 128662 104932 128726
rect 104856 128656 104932 128662
rect 104312 127198 104318 127230
rect 99622 127166 99623 127198
rect 99557 127165 99623 127166
rect 104317 127166 104318 127198
rect 104382 127198 104388 127230
rect 109616 127230 109692 131790
rect 109888 131310 109964 133014
rect 114784 133014 114790 133046
rect 114854 133046 114855 133078
rect 119685 133078 119751 133079
rect 119685 133046 119686 133078
rect 114854 133014 114860 133046
rect 114784 132812 114860 133014
rect 114648 132736 114860 132812
rect 119680 133014 119686 133046
rect 119750 133046 119751 133078
rect 124717 133078 124783 133079
rect 124717 133046 124718 133078
rect 119750 133014 119756 133046
rect 109888 131246 109894 131310
rect 109958 131246 109964 131310
rect 109888 131240 109964 131246
rect 114240 131854 114316 131860
rect 114240 131790 114246 131854
rect 114310 131790 114316 131854
rect 109893 131174 109959 131175
rect 109893 131142 109894 131174
rect 109888 131110 109894 131142
rect 109958 131142 109959 131174
rect 109958 131110 109964 131142
rect 109888 128726 109964 131110
rect 109888 128662 109894 128726
rect 109958 128662 109964 128726
rect 109888 128656 109964 128662
rect 109616 127198 109622 127230
rect 104382 127166 104383 127198
rect 104317 127165 104383 127166
rect 109621 127166 109622 127198
rect 109686 127198 109692 127230
rect 114240 127230 114316 131790
rect 114648 131310 114724 132736
rect 114784 132670 114860 132676
rect 114784 132606 114790 132670
rect 114854 132606 114860 132670
rect 114784 131990 114860 132606
rect 114784 131958 114790 131990
rect 114789 131926 114790 131958
rect 114854 131958 114860 131990
rect 119544 132670 119620 132676
rect 119544 132606 119550 132670
rect 119614 132606 119620 132670
rect 119544 131990 119620 132606
rect 119544 131958 119550 131990
rect 114854 131926 114855 131958
rect 114789 131925 114855 131926
rect 119549 131926 119550 131958
rect 119614 131958 119620 131990
rect 119614 131926 119615 131958
rect 119549 131925 119615 131926
rect 114648 131246 114654 131310
rect 114718 131246 114724 131310
rect 114648 131240 114724 131246
rect 119680 131310 119756 133014
rect 124712 133014 124718 133046
rect 124782 133046 124783 133078
rect 129749 133078 129815 133079
rect 129749 133046 129750 133078
rect 124782 133014 124788 133046
rect 124576 132670 124652 132676
rect 124576 132606 124582 132670
rect 124646 132606 124652 132670
rect 124576 131990 124652 132606
rect 124576 131958 124582 131990
rect 124581 131926 124582 131958
rect 124646 131958 124652 131990
rect 124646 131926 124647 131958
rect 124581 131925 124647 131926
rect 120229 131854 120295 131855
rect 120229 131822 120230 131854
rect 119680 131246 119686 131310
rect 119750 131246 119756 131310
rect 119680 131240 119756 131246
rect 120224 131790 120230 131822
rect 120294 131822 120295 131854
rect 124576 131854 124652 131860
rect 120294 131790 120300 131822
rect 114648 131174 114724 131180
rect 114648 131110 114654 131174
rect 114718 131110 114724 131174
rect 119821 131174 119887 131175
rect 119821 131142 119822 131174
rect 114648 128726 114724 131110
rect 114648 128694 114654 128726
rect 114653 128662 114654 128694
rect 114718 128694 114724 128726
rect 119816 131110 119822 131142
rect 119886 131142 119887 131174
rect 119886 131110 119892 131142
rect 119816 128726 119892 131110
rect 114718 128662 114719 128694
rect 114653 128661 114719 128662
rect 119816 128662 119822 128726
rect 119886 128662 119892 128726
rect 119816 128656 119892 128662
rect 114240 127198 114246 127230
rect 109686 127166 109687 127198
rect 109621 127165 109687 127166
rect 114245 127166 114246 127198
rect 114310 127198 114316 127230
rect 120224 127230 120300 131790
rect 114310 127166 114311 127198
rect 114245 127165 114311 127166
rect 120224 127166 120230 127230
rect 120294 127166 120300 127230
rect 124576 131790 124582 131854
rect 124646 131790 124652 131854
rect 124576 127230 124652 131790
rect 124712 131310 124788 133014
rect 129744 133014 129750 133046
rect 129814 133046 129815 133078
rect 134781 133078 134847 133079
rect 134781 133046 134782 133078
rect 129814 133014 129820 133046
rect 129608 132670 129684 132676
rect 129608 132606 129614 132670
rect 129678 132606 129684 132670
rect 129608 131990 129684 132606
rect 129608 131958 129614 131990
rect 129613 131926 129614 131958
rect 129678 131958 129684 131990
rect 129678 131926 129679 131958
rect 129613 131925 129679 131926
rect 124712 131246 124718 131310
rect 124782 131246 124788 131310
rect 124712 131240 124788 131246
rect 129200 131854 129276 131860
rect 129200 131790 129206 131854
rect 129270 131790 129276 131854
rect 124853 131174 124919 131175
rect 124853 131142 124854 131174
rect 124848 131110 124854 131142
rect 124918 131142 124919 131174
rect 124918 131110 124924 131142
rect 124848 128726 124924 131110
rect 124848 128662 124854 128726
rect 124918 128662 124924 128726
rect 124848 128656 124924 128662
rect 124576 127198 124582 127230
rect 120224 127160 120300 127166
rect 124581 127166 124582 127198
rect 124646 127198 124652 127230
rect 129200 127230 129276 131790
rect 129744 131310 129820 133014
rect 134776 133014 134782 133046
rect 134846 133046 134847 133078
rect 139677 133078 139743 133079
rect 139677 133046 139678 133078
rect 134846 133014 134852 133046
rect 134640 132670 134716 132676
rect 134640 132606 134646 132670
rect 134710 132606 134716 132670
rect 134640 131990 134716 132606
rect 134640 131958 134646 131990
rect 134645 131926 134646 131958
rect 134710 131958 134716 131990
rect 134710 131926 134711 131958
rect 134645 131925 134711 131926
rect 129744 131246 129750 131310
rect 129814 131246 129820 131310
rect 129744 131240 129820 131246
rect 134776 131310 134852 133014
rect 139672 133014 139678 133046
rect 139742 133046 139743 133078
rect 144709 133078 144775 133079
rect 144709 133046 144710 133078
rect 139742 133014 139748 133046
rect 139536 132670 139612 132676
rect 139536 132606 139542 132670
rect 139606 132606 139612 132670
rect 139536 131990 139612 132606
rect 139536 131958 139542 131990
rect 139541 131926 139542 131958
rect 139606 131958 139612 131990
rect 139606 131926 139607 131958
rect 139541 131925 139607 131926
rect 135597 131854 135663 131855
rect 135597 131822 135598 131854
rect 134776 131246 134782 131310
rect 134846 131246 134852 131310
rect 134776 131240 134852 131246
rect 135592 131790 135598 131822
rect 135662 131822 135663 131854
rect 139536 131854 139612 131860
rect 135662 131790 135668 131822
rect 129749 131174 129815 131175
rect 129749 131142 129750 131174
rect 129744 131110 129750 131142
rect 129814 131142 129815 131174
rect 134781 131174 134847 131175
rect 134781 131142 134782 131174
rect 129814 131110 129820 131142
rect 129744 128726 129820 131110
rect 129744 128662 129750 128726
rect 129814 128662 129820 128726
rect 129744 128656 129820 128662
rect 134776 131110 134782 131142
rect 134846 131142 134847 131174
rect 134846 131110 134852 131142
rect 134776 128726 134852 131110
rect 134776 128662 134782 128726
rect 134846 128662 134852 128726
rect 134776 128656 134852 128662
rect 129200 127198 129206 127230
rect 124646 127166 124647 127198
rect 124581 127165 124647 127166
rect 129205 127166 129206 127198
rect 129270 127198 129276 127230
rect 135592 127230 135668 131790
rect 129270 127166 129271 127198
rect 129205 127165 129271 127166
rect 135592 127166 135598 127230
rect 135662 127166 135668 127230
rect 139536 131790 139542 131854
rect 139606 131790 139612 131854
rect 139536 127230 139612 131790
rect 139672 131310 139748 133014
rect 144704 133014 144710 133046
rect 144774 133046 144775 133078
rect 149741 133078 149807 133079
rect 149741 133046 149742 133078
rect 144774 133014 144780 133046
rect 144568 132670 144644 132676
rect 144568 132606 144574 132670
rect 144638 132606 144644 132670
rect 144568 131990 144644 132606
rect 144568 131958 144574 131990
rect 144573 131926 144574 131958
rect 144638 131958 144644 131990
rect 144638 131926 144639 131958
rect 144573 131925 144639 131926
rect 139672 131246 139678 131310
rect 139742 131246 139748 131310
rect 139672 131240 139748 131246
rect 144704 131310 144780 133014
rect 149736 133014 149742 133046
rect 149806 133046 149807 133078
rect 154773 133078 154839 133079
rect 154773 133046 154774 133078
rect 149806 133014 149812 133046
rect 149600 132670 149676 132676
rect 149600 132606 149606 132670
rect 149670 132606 149676 132670
rect 149600 131990 149676 132606
rect 149600 131958 149606 131990
rect 149605 131926 149606 131958
rect 149670 131958 149676 131990
rect 149670 131926 149671 131958
rect 149605 131925 149671 131926
rect 145253 131854 145319 131855
rect 145253 131822 145254 131854
rect 144704 131246 144710 131310
rect 144774 131246 144780 131310
rect 144704 131240 144780 131246
rect 145248 131790 145254 131822
rect 145318 131822 145319 131854
rect 149464 131854 149540 131860
rect 145318 131790 145324 131822
rect 139813 131174 139879 131175
rect 139813 131142 139814 131174
rect 139808 131110 139814 131142
rect 139878 131142 139879 131174
rect 144845 131174 144911 131175
rect 144845 131142 144846 131174
rect 139878 131110 139884 131142
rect 139808 128726 139884 131110
rect 139808 128662 139814 128726
rect 139878 128662 139884 128726
rect 139808 128656 139884 128662
rect 144840 131110 144846 131142
rect 144910 131142 144911 131174
rect 144910 131110 144916 131142
rect 144840 128726 144916 131110
rect 144840 128662 144846 128726
rect 144910 128662 144916 128726
rect 144840 128656 144916 128662
rect 139536 127198 139542 127230
rect 135592 127160 135668 127166
rect 139541 127166 139542 127198
rect 139606 127198 139612 127230
rect 145248 127230 145324 131790
rect 139606 127166 139607 127198
rect 139541 127165 139607 127166
rect 145248 127166 145254 127230
rect 145318 127166 145324 127230
rect 149464 131790 149470 131854
rect 149534 131790 149540 131854
rect 149464 127230 149540 131790
rect 149736 131310 149812 133014
rect 154768 133014 154774 133046
rect 154838 133046 154839 133078
rect 159805 133078 159871 133079
rect 159805 133046 159806 133078
rect 154838 133014 154844 133046
rect 154632 132670 154708 132676
rect 154632 132606 154638 132670
rect 154702 132606 154708 132670
rect 154632 131990 154708 132606
rect 154632 131958 154638 131990
rect 154637 131926 154638 131958
rect 154702 131958 154708 131990
rect 154702 131926 154703 131958
rect 154637 131925 154703 131926
rect 149736 131246 149742 131310
rect 149806 131246 149812 131310
rect 149736 131240 149812 131246
rect 154088 131854 154164 131860
rect 154088 131790 154094 131854
rect 154158 131790 154164 131854
rect 149600 131174 149676 131180
rect 149600 131110 149606 131174
rect 149670 131110 149676 131174
rect 149600 128726 149676 131110
rect 149600 128694 149606 128726
rect 149605 128662 149606 128694
rect 149670 128694 149676 128726
rect 149670 128662 149671 128694
rect 149605 128661 149671 128662
rect 149464 127198 149470 127230
rect 145248 127160 145324 127166
rect 149469 127166 149470 127198
rect 149534 127198 149540 127230
rect 154088 127230 154164 131790
rect 154768 131310 154844 133014
rect 159800 133014 159806 133046
rect 159870 133046 159871 133078
rect 164701 133078 164767 133079
rect 164701 133046 164702 133078
rect 159870 133014 159876 133046
rect 159664 132670 159740 132676
rect 159664 132606 159670 132670
rect 159734 132606 159740 132670
rect 159664 131990 159740 132606
rect 159664 131958 159670 131990
rect 159669 131926 159670 131958
rect 159734 131958 159740 131990
rect 159734 131926 159735 131958
rect 159669 131925 159735 131926
rect 154768 131246 154774 131310
rect 154838 131246 154844 131310
rect 154768 131240 154844 131246
rect 159800 131310 159876 133014
rect 164696 133014 164702 133046
rect 164766 133046 164767 133078
rect 169733 133078 169799 133079
rect 169733 133046 169734 133078
rect 164766 133014 164772 133046
rect 164560 132670 164636 132676
rect 164560 132606 164566 132670
rect 164630 132606 164636 132670
rect 164560 131990 164636 132606
rect 164560 131958 164566 131990
rect 164565 131926 164566 131958
rect 164630 131958 164636 131990
rect 164630 131926 164631 131958
rect 164565 131925 164631 131926
rect 160213 131854 160279 131855
rect 160213 131822 160214 131854
rect 159800 131246 159806 131310
rect 159870 131246 159876 131310
rect 159800 131240 159876 131246
rect 160208 131790 160214 131822
rect 160278 131822 160279 131854
rect 160278 131790 160284 131822
rect 154773 131174 154839 131175
rect 154773 131142 154774 131174
rect 154768 131110 154774 131142
rect 154838 131142 154839 131174
rect 159805 131174 159871 131175
rect 159805 131142 159806 131174
rect 154838 131110 154844 131142
rect 154768 128726 154844 131110
rect 154768 128662 154774 128726
rect 154838 128662 154844 128726
rect 154768 128656 154844 128662
rect 159800 131110 159806 131142
rect 159870 131142 159871 131174
rect 159870 131110 159876 131142
rect 159800 128726 159876 131110
rect 159800 128662 159806 128726
rect 159870 128662 159876 128726
rect 159800 128656 159876 128662
rect 154088 127198 154094 127230
rect 149534 127166 149535 127198
rect 149469 127165 149535 127166
rect 154093 127166 154094 127198
rect 154158 127198 154164 127230
rect 160208 127230 160284 131790
rect 164696 131310 164772 133014
rect 169728 133014 169734 133046
rect 169798 133046 169799 133078
rect 174765 133078 174831 133079
rect 174765 133046 174766 133078
rect 169798 133014 169804 133046
rect 169592 132670 169668 132676
rect 169592 132606 169598 132670
rect 169662 132606 169668 132670
rect 169592 131990 169668 132606
rect 169592 131958 169598 131990
rect 169597 131926 169598 131958
rect 169662 131958 169668 131990
rect 169662 131926 169663 131958
rect 169597 131925 169663 131926
rect 165517 131854 165583 131855
rect 165517 131822 165518 131854
rect 164696 131246 164702 131310
rect 164766 131246 164772 131310
rect 164696 131240 164772 131246
rect 165512 131790 165518 131822
rect 165582 131822 165583 131854
rect 165582 131790 165588 131822
rect 164701 131174 164767 131175
rect 164701 131142 164702 131174
rect 164696 131110 164702 131142
rect 164766 131142 164767 131174
rect 164766 131110 164772 131142
rect 164696 128726 164772 131110
rect 164696 128662 164702 128726
rect 164766 128662 164772 128726
rect 164696 128656 164772 128662
rect 154158 127166 154159 127198
rect 154093 127165 154159 127166
rect 160208 127166 160214 127230
rect 160278 127166 160284 127230
rect 160208 127160 160284 127166
rect 165512 127230 165588 131790
rect 169728 131310 169804 133014
rect 174760 133014 174766 133046
rect 174830 133046 174831 133078
rect 179797 133078 179863 133079
rect 179797 133046 179798 133078
rect 174830 133014 174836 133046
rect 174624 132670 174700 132676
rect 174624 132606 174630 132670
rect 174694 132606 174700 132670
rect 174624 131990 174700 132606
rect 174624 131958 174630 131990
rect 174629 131926 174630 131958
rect 174694 131958 174700 131990
rect 174694 131926 174695 131958
rect 174629 131925 174695 131926
rect 170141 131854 170207 131855
rect 170141 131822 170142 131854
rect 169728 131246 169734 131310
rect 169798 131246 169804 131310
rect 169728 131240 169804 131246
rect 170136 131790 170142 131822
rect 170206 131822 170207 131854
rect 174488 131854 174564 131860
rect 170206 131790 170212 131822
rect 169733 131174 169799 131175
rect 169733 131142 169734 131174
rect 169728 131110 169734 131142
rect 169798 131142 169799 131174
rect 169798 131110 169804 131142
rect 169728 128726 169804 131110
rect 169728 128662 169734 128726
rect 169798 128662 169804 128726
rect 169728 128656 169804 128662
rect 165512 127166 165518 127230
rect 165582 127166 165588 127230
rect 165512 127160 165588 127166
rect 170136 127230 170212 131790
rect 170136 127166 170142 127230
rect 170206 127166 170212 127230
rect 174488 131790 174494 131854
rect 174558 131790 174564 131854
rect 174488 127230 174564 131790
rect 174760 131310 174836 133014
rect 179792 133014 179798 133046
rect 179862 133046 179863 133078
rect 184557 133078 184623 133079
rect 184557 133046 184558 133078
rect 179862 133014 179868 133046
rect 179656 132670 179732 132676
rect 179656 132606 179662 132670
rect 179726 132606 179732 132670
rect 179656 131990 179732 132606
rect 179656 131958 179662 131990
rect 179661 131926 179662 131958
rect 179726 131958 179732 131990
rect 179726 131926 179727 131958
rect 179661 131925 179727 131926
rect 174760 131246 174766 131310
rect 174830 131246 174836 131310
rect 174760 131240 174836 131246
rect 179520 131854 179596 131860
rect 179520 131790 179526 131854
rect 179590 131790 179596 131854
rect 174624 131174 174700 131180
rect 174624 131110 174630 131174
rect 174694 131110 174700 131174
rect 174624 128726 174700 131110
rect 174624 128694 174630 128726
rect 174629 128662 174630 128694
rect 174694 128694 174700 128726
rect 174694 128662 174695 128694
rect 174629 128661 174695 128662
rect 174488 127198 174494 127230
rect 170136 127160 170212 127166
rect 174493 127166 174494 127198
rect 174558 127198 174564 127230
rect 179520 127230 179596 131790
rect 179792 131310 179868 133014
rect 184552 133014 184558 133046
rect 184622 133046 184623 133078
rect 184622 133014 184628 133046
rect 184416 132670 184492 132676
rect 184416 132606 184422 132670
rect 184486 132606 184492 132670
rect 184416 131990 184492 132606
rect 184416 131958 184422 131990
rect 184421 131926 184422 131958
rect 184486 131958 184492 131990
rect 184486 131926 184487 131958
rect 184421 131925 184487 131926
rect 179792 131246 179798 131310
rect 179862 131246 179868 131310
rect 179792 131240 179868 131246
rect 184416 131854 184492 131860
rect 184416 131790 184422 131854
rect 184486 131790 184492 131854
rect 179797 131174 179863 131175
rect 179797 131142 179798 131174
rect 179792 131110 179798 131142
rect 179862 131142 179863 131174
rect 179862 131110 179868 131142
rect 179792 128726 179868 131110
rect 179792 128662 179798 128726
rect 179862 128662 179868 128726
rect 179792 128656 179868 128662
rect 179520 127198 179526 127230
rect 174558 127166 174559 127198
rect 174493 127165 174559 127166
rect 179525 127166 179526 127198
rect 179590 127198 179596 127230
rect 184416 127230 184492 131790
rect 184552 131310 184628 133014
rect 196525 132670 196591 132671
rect 196525 132638 196526 132670
rect 184552 131246 184558 131310
rect 184622 131246 184628 131310
rect 184552 131240 184628 131246
rect 196520 132606 196526 132638
rect 196590 132638 196591 132670
rect 196590 132606 196596 132638
rect 184693 131174 184759 131175
rect 184693 131142 184694 131174
rect 184688 131110 184694 131142
rect 184758 131142 184759 131174
rect 184758 131110 184764 131142
rect 184688 128726 184764 131110
rect 196520 130086 196596 132606
rect 196656 131446 196732 134102
rect 198016 132806 198092 135462
rect 198016 132742 198022 132806
rect 198086 132742 198092 132806
rect 198016 132736 198092 132742
rect 203320 135254 203396 135260
rect 203320 135190 203326 135254
rect 203390 135190 203396 135254
rect 216789 135254 216855 135255
rect 216789 135222 216790 135254
rect 203320 132670 203396 135190
rect 216784 135190 216790 135222
rect 216854 135222 216855 135254
rect 216854 135190 216860 135222
rect 216784 134982 216860 135190
rect 216784 134918 216790 134982
rect 216854 134918 216860 134982
rect 216784 134912 216860 134918
rect 217464 134846 217812 136550
rect 217464 134782 217470 134846
rect 217534 134782 217812 134846
rect 203456 133894 203532 133900
rect 203456 133830 203462 133894
rect 203526 133830 203532 133894
rect 203597 133894 203663 133895
rect 203597 133862 203598 133894
rect 203456 132806 203532 133830
rect 203456 132774 203462 132806
rect 203461 132742 203462 132774
rect 203526 132774 203532 132806
rect 203592 133830 203598 133862
rect 203662 133862 203663 133894
rect 203662 133830 203668 133862
rect 203526 132742 203527 132774
rect 203461 132741 203527 132742
rect 203320 132638 203326 132670
rect 203325 132606 203326 132638
rect 203390 132638 203396 132670
rect 203390 132606 203391 132638
rect 203325 132605 203391 132606
rect 203325 132534 203391 132535
rect 203325 132502 203326 132534
rect 196656 131414 196662 131446
rect 196661 131382 196662 131414
rect 196726 131414 196732 131446
rect 203320 132470 203326 132502
rect 203390 132502 203391 132534
rect 203456 132534 203532 132540
rect 203390 132470 203396 132502
rect 196726 131382 196727 131414
rect 196661 131381 196727 131382
rect 196520 130022 196526 130086
rect 196590 130022 196596 130086
rect 196520 130016 196596 130022
rect 197880 131310 197956 131316
rect 197880 131246 197886 131310
rect 197950 131246 197956 131310
rect 184688 128662 184694 128726
rect 184758 128662 184764 128726
rect 184688 128656 184764 128662
rect 196520 129814 196596 129820
rect 196520 129750 196526 129814
rect 196590 129750 196596 129814
rect 190405 128590 190471 128591
rect 190405 128558 190406 128590
rect 184416 127198 184422 127230
rect 179590 127166 179591 127198
rect 179525 127165 179591 127166
rect 184421 127166 184422 127198
rect 184486 127198 184492 127230
rect 190400 128526 190406 128558
rect 190470 128558 190471 128590
rect 190470 128526 190476 128558
rect 184486 127166 184487 127198
rect 184421 127165 184487 127166
rect 29653 127094 29719 127095
rect 29653 127062 29654 127094
rect 29648 127030 29654 127062
rect 29718 127062 29719 127094
rect 30877 127094 30943 127095
rect 30877 127062 30878 127094
rect 29718 127030 29724 127062
rect 29648 126686 29724 127030
rect 29648 126622 29654 126686
rect 29718 126622 29724 126686
rect 29648 126616 29724 126622
rect 30872 127030 30878 127062
rect 30942 127062 30943 127094
rect 31688 127094 31764 127100
rect 30942 127030 30948 127062
rect 30872 126686 30948 127030
rect 30872 126622 30878 126686
rect 30942 126622 30948 126686
rect 31688 127030 31694 127094
rect 31758 127030 31764 127094
rect 31688 126686 31764 127030
rect 31688 126654 31694 126686
rect 30872 126616 30948 126622
rect 31693 126622 31694 126654
rect 31758 126654 31764 126686
rect 32912 127094 32988 127100
rect 32912 127030 32918 127094
rect 32982 127030 32988 127094
rect 33461 127094 33527 127095
rect 33461 127062 33462 127094
rect 32912 126686 32988 127030
rect 32912 126654 32918 126686
rect 31758 126622 31759 126654
rect 31693 126621 31759 126622
rect 32917 126622 32918 126654
rect 32982 126654 32988 126686
rect 33456 127030 33462 127062
rect 33526 127062 33527 127094
rect 34136 127094 34212 127100
rect 33526 127030 33532 127062
rect 33456 126686 33532 127030
rect 32982 126622 32983 126654
rect 32917 126621 32983 126622
rect 33456 126622 33462 126686
rect 33526 126622 33532 126686
rect 34136 127030 34142 127094
rect 34206 127030 34212 127094
rect 34685 127094 34751 127095
rect 34685 127062 34686 127094
rect 34136 126686 34212 127030
rect 34136 126654 34142 126686
rect 33456 126616 33532 126622
rect 34141 126622 34142 126654
rect 34206 126654 34212 126686
rect 34680 127030 34686 127062
rect 34750 127062 34751 127094
rect 35909 127094 35975 127095
rect 35909 127062 35910 127094
rect 34750 127030 34756 127062
rect 34680 126686 34756 127030
rect 34206 126622 34207 126654
rect 34141 126621 34207 126622
rect 34680 126622 34686 126686
rect 34750 126622 34756 126686
rect 34680 126616 34756 126622
rect 35904 127030 35910 127062
rect 35974 127062 35975 127094
rect 36584 127094 36660 127100
rect 35974 127030 35980 127062
rect 35904 126686 35980 127030
rect 35904 126622 35910 126686
rect 35974 126622 35980 126686
rect 36584 127030 36590 127094
rect 36654 127030 36660 127094
rect 37133 127094 37199 127095
rect 37133 127062 37134 127094
rect 36584 126686 36660 127030
rect 36584 126654 36590 126686
rect 35904 126616 35980 126622
rect 36589 126622 36590 126654
rect 36654 126654 36660 126686
rect 37128 127030 37134 127062
rect 37198 127062 37199 127094
rect 38085 127094 38151 127095
rect 38085 127062 38086 127094
rect 37198 127030 37204 127062
rect 37128 126686 37204 127030
rect 36654 126622 36655 126654
rect 36589 126621 36655 126622
rect 37128 126622 37134 126686
rect 37198 126622 37204 126686
rect 37128 126616 37204 126622
rect 38080 127030 38086 127062
rect 38150 127062 38151 127094
rect 39445 127094 39511 127095
rect 39445 127062 39446 127094
rect 38150 127030 38156 127062
rect 38080 126686 38156 127030
rect 38080 126622 38086 126686
rect 38150 126622 38156 126686
rect 38080 126616 38156 126622
rect 39440 127030 39446 127062
rect 39510 127062 39511 127094
rect 40392 127094 40468 127100
rect 39510 127030 39516 127062
rect 39440 126686 39516 127030
rect 39440 126622 39446 126686
rect 39510 126622 39516 126686
rect 40392 127030 40398 127094
rect 40462 127030 40468 127094
rect 40392 126686 40468 127030
rect 40392 126654 40398 126686
rect 39440 126616 39516 126622
rect 40397 126622 40398 126654
rect 40462 126654 40468 126686
rect 41616 127094 41692 127100
rect 41616 127030 41622 127094
rect 41686 127030 41692 127094
rect 42165 127094 42231 127095
rect 42165 127062 42166 127094
rect 41616 126686 41692 127030
rect 41616 126654 41622 126686
rect 40462 126622 40463 126654
rect 40397 126621 40463 126622
rect 41621 126622 41622 126654
rect 41686 126654 41692 126686
rect 42160 127030 42166 127062
rect 42230 127062 42231 127094
rect 42976 127094 43052 127100
rect 42230 127030 42236 127062
rect 42160 126686 42236 127030
rect 41686 126622 41687 126654
rect 41621 126621 41687 126622
rect 42160 126622 42166 126686
rect 42230 126622 42236 126686
rect 42976 127030 42982 127094
rect 43046 127030 43052 127094
rect 42976 126686 43052 127030
rect 42976 126654 42982 126686
rect 42160 126616 42236 126622
rect 42981 126622 42982 126654
rect 43046 126654 43052 126686
rect 43248 127094 43324 127100
rect 43248 127030 43254 127094
rect 43318 127030 43324 127094
rect 44613 127094 44679 127095
rect 44613 127062 44614 127094
rect 43248 126686 43324 127030
rect 43248 126654 43254 126686
rect 43046 126622 43047 126654
rect 42981 126621 43047 126622
rect 43253 126622 43254 126654
rect 43318 126654 43324 126686
rect 44608 127030 44614 127062
rect 44678 127062 44679 127094
rect 45424 127094 45500 127100
rect 44678 127030 44684 127062
rect 44608 126686 44684 127030
rect 43318 126622 43319 126654
rect 43253 126621 43319 126622
rect 44608 126622 44614 126686
rect 44678 126622 44684 126686
rect 45424 127030 45430 127094
rect 45494 127030 45500 127094
rect 45973 127094 46039 127095
rect 45973 127062 45974 127094
rect 45424 126686 45500 127030
rect 45424 126654 45430 126686
rect 44608 126616 44684 126622
rect 45429 126622 45430 126654
rect 45494 126654 45500 126686
rect 45968 127030 45974 127062
rect 46038 127062 46039 127094
rect 46648 127094 46724 127100
rect 46038 127030 46044 127062
rect 45968 126686 46044 127030
rect 45494 126622 45495 126654
rect 45429 126621 45495 126622
rect 45968 126622 45974 126686
rect 46038 126622 46044 126686
rect 46648 127030 46654 127094
rect 46718 127030 46724 127094
rect 46789 127094 46855 127095
rect 46789 127062 46790 127094
rect 46648 126686 46724 127030
rect 46648 126654 46654 126686
rect 45968 126616 46044 126622
rect 46653 126622 46654 126654
rect 46718 126654 46724 126686
rect 46784 127030 46790 127062
rect 46854 127062 46855 127094
rect 48421 127094 48487 127095
rect 48421 127062 48422 127094
rect 46854 127030 46860 127062
rect 46784 126686 46860 127030
rect 46718 126622 46719 126654
rect 46653 126621 46719 126622
rect 46784 126622 46790 126686
rect 46854 126622 46860 126686
rect 46784 126616 46860 126622
rect 48416 127030 48422 127062
rect 48486 127062 48487 127094
rect 49096 127094 49172 127100
rect 48486 127030 48492 127062
rect 48416 126686 48492 127030
rect 48416 126622 48422 126686
rect 48486 126622 48492 126686
rect 49096 127030 49102 127094
rect 49166 127030 49172 127094
rect 49096 126686 49172 127030
rect 49096 126654 49102 126686
rect 48416 126616 48492 126622
rect 49101 126622 49102 126654
rect 49166 126654 49172 126686
rect 50320 127094 50396 127100
rect 50320 127030 50326 127094
rect 50390 127030 50396 127094
rect 50869 127094 50935 127095
rect 50869 127062 50870 127094
rect 50320 126686 50396 127030
rect 50320 126654 50326 126686
rect 49166 126622 49167 126654
rect 49101 126621 49167 126622
rect 50325 126622 50326 126654
rect 50390 126654 50396 126686
rect 50864 127030 50870 127062
rect 50934 127062 50935 127094
rect 52229 127094 52295 127095
rect 52229 127062 52230 127094
rect 50934 127030 50940 127062
rect 50864 126686 50940 127030
rect 50390 126622 50391 126654
rect 50325 126621 50391 126622
rect 50864 126622 50870 126686
rect 50934 126622 50940 126686
rect 50864 126616 50940 126622
rect 52224 127030 52230 127062
rect 52294 127062 52295 127094
rect 52773 127094 52839 127095
rect 52773 127062 52774 127094
rect 52294 127030 52300 127062
rect 52224 126686 52300 127030
rect 52224 126622 52230 126686
rect 52294 126622 52300 126686
rect 52224 126616 52300 126622
rect 52768 127030 52774 127062
rect 52838 127062 52839 127094
rect 53317 127094 53383 127095
rect 53317 127062 53318 127094
rect 52838 127030 52844 127062
rect 52768 126686 52844 127030
rect 52768 126622 52774 126686
rect 52838 126622 52844 126686
rect 52768 126616 52844 126622
rect 53312 127030 53318 127062
rect 53382 127062 53383 127094
rect 54128 127094 54204 127100
rect 53382 127030 53388 127062
rect 53312 126686 53388 127030
rect 53312 126622 53318 126686
rect 53382 126622 53388 126686
rect 54128 127030 54134 127094
rect 54198 127030 54204 127094
rect 54677 127094 54743 127095
rect 54677 127062 54678 127094
rect 54128 126686 54204 127030
rect 54128 126654 54134 126686
rect 53312 126616 53388 126622
rect 54133 126622 54134 126654
rect 54198 126654 54204 126686
rect 54672 127030 54678 127062
rect 54742 127062 54743 127094
rect 55352 127094 55428 127100
rect 54742 127030 54748 127062
rect 54672 126686 54748 127030
rect 54198 126622 54199 126654
rect 54133 126621 54199 126622
rect 54672 126622 54678 126686
rect 54742 126622 54748 126686
rect 55352 127030 55358 127094
rect 55422 127030 55428 127094
rect 55901 127094 55967 127095
rect 55901 127062 55902 127094
rect 55352 126686 55428 127030
rect 55352 126654 55358 126686
rect 54672 126616 54748 126622
rect 55357 126622 55358 126654
rect 55422 126654 55428 126686
rect 55896 127030 55902 127062
rect 55966 127062 55967 127094
rect 57125 127094 57191 127095
rect 57125 127062 57126 127094
rect 55966 127030 55972 127062
rect 55896 126686 55972 127030
rect 55422 126622 55423 126654
rect 55357 126621 55423 126622
rect 55896 126622 55902 126686
rect 55966 126622 55972 126686
rect 55896 126616 55972 126622
rect 57120 127030 57126 127062
rect 57190 127062 57191 127094
rect 57800 127094 57876 127100
rect 57190 127030 57196 127062
rect 57120 126686 57196 127030
rect 57120 126622 57126 126686
rect 57190 126622 57196 126686
rect 57800 127030 57806 127094
rect 57870 127030 57876 127094
rect 59573 127094 59639 127095
rect 59573 127062 59574 127094
rect 57800 126686 57876 127030
rect 57800 126654 57806 126686
rect 57120 126616 57196 126622
rect 57805 126622 57806 126654
rect 57870 126654 57876 126686
rect 59568 127030 59574 127062
rect 59638 127062 59639 127094
rect 60933 127094 60999 127095
rect 60933 127062 60934 127094
rect 59638 127030 59644 127062
rect 59568 126686 59644 127030
rect 57870 126622 57871 126654
rect 57805 126621 57871 126622
rect 59568 126622 59574 126686
rect 59638 126622 59644 126686
rect 59568 126616 59644 126622
rect 60928 127030 60934 127062
rect 60998 127062 60999 127094
rect 61477 127094 61543 127095
rect 61477 127062 61478 127094
rect 60998 127030 61004 127062
rect 60928 126686 61004 127030
rect 60928 126622 60934 126686
rect 60998 126622 61004 126686
rect 60928 126616 61004 126622
rect 61472 127030 61478 127062
rect 61542 127062 61543 127094
rect 61608 127094 61684 127100
rect 61542 127030 61548 127062
rect 61472 126686 61548 127030
rect 61472 126622 61478 126686
rect 61542 126622 61548 126686
rect 61608 127030 61614 127094
rect 61678 127030 61684 127094
rect 62157 127094 62223 127095
rect 62157 127062 62158 127094
rect 61608 126686 61684 127030
rect 61608 126654 61614 126686
rect 61472 126616 61548 126622
rect 61613 126622 61614 126654
rect 61678 126654 61684 126686
rect 62152 127030 62158 127062
rect 62222 127062 62223 127094
rect 62832 127094 62908 127100
rect 62222 127030 62228 127062
rect 62152 126686 62228 127030
rect 61678 126622 61679 126654
rect 61613 126621 61679 126622
rect 62152 126622 62158 126686
rect 62222 126622 62228 126686
rect 62832 127030 62838 127094
rect 62902 127030 62908 127094
rect 63381 127094 63447 127095
rect 63381 127062 63382 127094
rect 62832 126686 62908 127030
rect 62832 126654 62838 126686
rect 62152 126616 62228 126622
rect 62837 126622 62838 126654
rect 62902 126654 62908 126686
rect 63376 127030 63382 127062
rect 63446 127062 63447 127094
rect 64056 127094 64132 127100
rect 63446 127030 63452 127062
rect 63376 126686 63452 127030
rect 62902 126622 62903 126654
rect 62837 126621 62903 126622
rect 63376 126622 63382 126686
rect 63446 126622 63452 126686
rect 64056 127030 64062 127094
rect 64126 127030 64132 127094
rect 64056 126686 64132 127030
rect 64056 126654 64062 126686
rect 63376 126616 63452 126622
rect 64061 126622 64062 126654
rect 64126 126654 64132 126686
rect 65688 127094 65764 127100
rect 65688 127030 65694 127094
rect 65758 127030 65764 127094
rect 65688 126686 65764 127030
rect 65688 126654 65694 126686
rect 64126 126622 64127 126654
rect 64061 126621 64127 126622
rect 65693 126622 65694 126654
rect 65758 126654 65764 126686
rect 66640 127094 66716 127100
rect 66640 127030 66646 127094
rect 66710 127030 66716 127094
rect 67189 127094 67255 127095
rect 67189 127062 67190 127094
rect 66640 126686 66716 127030
rect 66640 126654 66646 126686
rect 65758 126622 65759 126654
rect 65693 126621 65759 126622
rect 66645 126622 66646 126654
rect 66710 126654 66716 126686
rect 67184 127030 67190 127062
rect 67254 127062 67255 127094
rect 67320 127094 67396 127100
rect 67254 127030 67260 127062
rect 67184 126686 67260 127030
rect 66710 126622 66711 126654
rect 66645 126621 66711 126622
rect 67184 126622 67190 126686
rect 67254 126622 67260 126686
rect 67320 127030 67326 127094
rect 67390 127030 67396 127094
rect 68413 127094 68479 127095
rect 68413 127062 68414 127094
rect 67320 126686 67396 127030
rect 67320 126654 67326 126686
rect 67184 126616 67260 126622
rect 67325 126622 67326 126654
rect 67390 126654 67396 126686
rect 68408 127030 68414 127062
rect 68478 127062 68479 127094
rect 69088 127094 69164 127100
rect 68478 127030 68484 127062
rect 68408 126686 68484 127030
rect 67390 126622 67391 126654
rect 67325 126621 67391 126622
rect 68408 126622 68414 126686
rect 68478 126622 68484 126686
rect 69088 127030 69094 127094
rect 69158 127030 69164 127094
rect 69637 127094 69703 127095
rect 69637 127062 69638 127094
rect 69088 126686 69164 127030
rect 69088 126654 69094 126686
rect 68408 126616 68484 126622
rect 69093 126622 69094 126654
rect 69158 126654 69164 126686
rect 69632 127030 69638 127062
rect 69702 127062 69703 127094
rect 70312 127094 70388 127100
rect 69702 127030 69708 127062
rect 69632 126686 69708 127030
rect 69158 126622 69159 126654
rect 69093 126621 69159 126622
rect 69632 126622 69638 126686
rect 69702 126622 69708 126686
rect 70312 127030 70318 127094
rect 70382 127030 70388 127094
rect 70861 127094 70927 127095
rect 70861 127062 70862 127094
rect 70312 126686 70388 127030
rect 70312 126654 70318 126686
rect 69632 126616 69708 126622
rect 70317 126622 70318 126654
rect 70382 126654 70388 126686
rect 70856 127030 70862 127062
rect 70926 127062 70927 127094
rect 71944 127094 72020 127100
rect 70926 127030 70932 127062
rect 70856 126686 70932 127030
rect 70382 126622 70383 126654
rect 70317 126621 70383 126622
rect 70856 126622 70862 126686
rect 70926 126622 70932 126686
rect 71944 127030 71950 127094
rect 72014 127030 72020 127094
rect 71944 126686 72020 127030
rect 71944 126654 71950 126686
rect 70856 126616 70932 126622
rect 71949 126622 71950 126654
rect 72014 126654 72020 126686
rect 72896 127094 72972 127100
rect 72896 127030 72902 127094
rect 72966 127030 72972 127094
rect 72896 126686 72972 127030
rect 72896 126654 72902 126686
rect 72014 126622 72015 126654
rect 71949 126621 72015 126622
rect 72901 126622 72902 126654
rect 72966 126654 72972 126686
rect 74120 127094 74196 127100
rect 74120 127030 74126 127094
rect 74190 127030 74196 127094
rect 75213 127094 75279 127095
rect 75213 127062 75214 127094
rect 74120 126686 74196 127030
rect 74120 126654 74126 126686
rect 72966 126622 72967 126654
rect 72901 126621 72967 126622
rect 74125 126622 74126 126654
rect 74190 126654 74196 126686
rect 75208 127030 75214 127062
rect 75278 127062 75279 127094
rect 75344 127094 75420 127100
rect 75278 127030 75284 127062
rect 75208 126686 75284 127030
rect 74190 126622 74191 126654
rect 74125 126621 74191 126622
rect 75208 126622 75214 126686
rect 75278 126622 75284 126686
rect 75344 127030 75350 127094
rect 75414 127030 75420 127094
rect 75893 127094 75959 127095
rect 75893 127062 75894 127094
rect 75344 126686 75420 127030
rect 75344 126654 75350 126686
rect 75208 126616 75284 126622
rect 75349 126622 75350 126654
rect 75414 126654 75420 126686
rect 75888 127030 75894 127062
rect 75958 127062 75959 127094
rect 76568 127094 76644 127100
rect 75958 127030 75964 127062
rect 75888 126686 75964 127030
rect 75414 126622 75415 126654
rect 75349 126621 75415 126622
rect 75888 126622 75894 126686
rect 75958 126622 75964 126686
rect 76568 127030 76574 127094
rect 76638 127030 76644 127094
rect 77117 127094 77183 127095
rect 77117 127062 77118 127094
rect 76568 126686 76644 127030
rect 76568 126654 76574 126686
rect 75888 126616 75964 126622
rect 76573 126622 76574 126654
rect 76638 126654 76644 126686
rect 77112 127030 77118 127062
rect 77182 127062 77183 127094
rect 77792 127094 77868 127100
rect 77182 127030 77188 127062
rect 77112 126686 77188 127030
rect 76638 126622 76639 126654
rect 76573 126621 76639 126622
rect 77112 126622 77118 126686
rect 77182 126622 77188 126686
rect 77792 127030 77798 127094
rect 77862 127030 77868 127094
rect 78341 127094 78407 127095
rect 78341 127062 78342 127094
rect 77792 126686 77868 127030
rect 77792 126654 77798 126686
rect 77112 126616 77188 126622
rect 77797 126622 77798 126654
rect 77862 126654 77868 126686
rect 78336 127030 78342 127062
rect 78406 127062 78407 127094
rect 79565 127094 79631 127095
rect 79565 127062 79566 127094
rect 78406 127030 78412 127062
rect 78336 126686 78412 127030
rect 77862 126622 77863 126654
rect 77797 126621 77863 126622
rect 78336 126622 78342 126686
rect 78406 126622 78412 126686
rect 78336 126616 78412 126622
rect 79560 127030 79566 127062
rect 79630 127062 79631 127094
rect 80925 127094 80991 127095
rect 80925 127062 80926 127094
rect 79630 127030 79636 127062
rect 79560 126686 79636 127030
rect 79560 126622 79566 126686
rect 79630 126622 79636 126686
rect 79560 126616 79636 126622
rect 80920 127030 80926 127062
rect 80990 127062 80991 127094
rect 81469 127094 81535 127095
rect 81469 127062 81470 127094
rect 80990 127030 80996 127062
rect 80920 126686 80996 127030
rect 80920 126622 80926 126686
rect 80990 126622 80996 126686
rect 80920 126616 80996 126622
rect 81464 127030 81470 127062
rect 81534 127062 81535 127094
rect 81600 127094 81676 127100
rect 81534 127030 81540 127062
rect 81464 126686 81540 127030
rect 81464 126622 81470 126686
rect 81534 126622 81540 126686
rect 81600 127030 81606 127094
rect 81670 127030 81676 127094
rect 82013 127094 82079 127095
rect 82013 127062 82014 127094
rect 81600 126686 81676 127030
rect 81600 126654 81606 126686
rect 81464 126616 81540 126622
rect 81605 126622 81606 126654
rect 81670 126654 81676 126686
rect 82008 127030 82014 127062
rect 82078 127062 82079 127094
rect 82824 127094 82900 127100
rect 82078 127030 82084 127062
rect 82008 126686 82084 127030
rect 81670 126622 81671 126654
rect 81605 126621 81671 126622
rect 82008 126622 82014 126686
rect 82078 126622 82084 126686
rect 82824 127030 82830 127094
rect 82894 127030 82900 127094
rect 82824 126686 82900 127030
rect 82824 126654 82830 126686
rect 82008 126616 82084 126622
rect 82829 126622 82830 126654
rect 82894 126654 82900 126686
rect 84048 127094 84124 127100
rect 84048 127030 84054 127094
rect 84118 127030 84124 127094
rect 84597 127094 84663 127095
rect 84597 127062 84598 127094
rect 84048 126686 84124 127030
rect 84048 126654 84054 126686
rect 82894 126622 82895 126654
rect 82829 126621 82895 126622
rect 84053 126622 84054 126654
rect 84118 126654 84124 126686
rect 84592 127030 84598 127062
rect 84662 127062 84663 127094
rect 85272 127094 85348 127100
rect 84662 127030 84668 127062
rect 84592 126686 84668 127030
rect 84118 126622 84119 126654
rect 84053 126621 84119 126622
rect 84592 126622 84598 126686
rect 84662 126622 84668 126686
rect 85272 127030 85278 127094
rect 85342 127030 85348 127094
rect 85821 127094 85887 127095
rect 85821 127062 85822 127094
rect 85272 126686 85348 127030
rect 85272 126654 85278 126686
rect 84592 126616 84668 126622
rect 85277 126622 85278 126654
rect 85342 126654 85348 126686
rect 85816 127030 85822 127062
rect 85886 127062 85887 127094
rect 86496 127094 86572 127100
rect 85886 127030 85892 127062
rect 85816 126686 85892 127030
rect 85342 126622 85343 126654
rect 85277 126621 85343 126622
rect 85816 126622 85822 126686
rect 85886 126622 85892 126686
rect 86496 127030 86502 127094
rect 86566 127030 86572 127094
rect 87045 127094 87111 127095
rect 87045 127062 87046 127094
rect 86496 126686 86572 127030
rect 86496 126654 86502 126686
rect 85816 126616 85892 126622
rect 86501 126622 86502 126654
rect 86566 126654 86572 126686
rect 87040 127030 87046 127062
rect 87110 127062 87111 127094
rect 88405 127094 88471 127095
rect 88405 127062 88406 127094
rect 87110 127030 87116 127062
rect 87040 126686 87116 127030
rect 86566 126622 86567 126654
rect 86501 126621 86567 126622
rect 87040 126622 87046 126686
rect 87110 126622 87116 126686
rect 87040 126616 87116 126622
rect 88400 127030 88406 127062
rect 88470 127062 88471 127094
rect 89221 127094 89287 127095
rect 89221 127062 89222 127094
rect 88470 127030 88476 127062
rect 88400 126686 88476 127030
rect 88400 126622 88406 126686
rect 88470 126622 88476 126686
rect 88400 126616 88476 126622
rect 89216 127030 89222 127062
rect 89286 127062 89287 127094
rect 90304 127094 90380 127100
rect 89286 127030 89292 127062
rect 89216 126550 89292 127030
rect 90304 127030 90310 127094
rect 90374 127030 90380 127094
rect 90853 127094 90919 127095
rect 90853 127062 90854 127094
rect 90304 126686 90380 127030
rect 90304 126654 90310 126686
rect 90309 126622 90310 126654
rect 90374 126654 90380 126686
rect 90848 127030 90854 127062
rect 90918 127062 90919 127094
rect 91528 127094 91604 127100
rect 90918 127030 90924 127062
rect 90848 126686 90924 127030
rect 90374 126622 90375 126654
rect 90309 126621 90375 126622
rect 90848 126622 90854 126686
rect 90918 126622 90924 126686
rect 91528 127030 91534 127094
rect 91598 127030 91604 127094
rect 91528 126686 91604 127030
rect 91528 126654 91534 126686
rect 90848 126616 90924 126622
rect 91533 126622 91534 126654
rect 91598 126654 91604 126686
rect 92752 127094 92828 127100
rect 92752 127030 92758 127094
rect 92822 127030 92828 127094
rect 93301 127094 93367 127095
rect 93301 127062 93302 127094
rect 92752 126686 92828 127030
rect 92752 126654 92758 126686
rect 91598 126622 91599 126654
rect 91533 126621 91599 126622
rect 92757 126622 92758 126654
rect 92822 126654 92828 126686
rect 93296 127030 93302 127062
rect 93366 127062 93367 127094
rect 94661 127094 94727 127095
rect 94661 127062 94662 127094
rect 93366 127030 93372 127062
rect 93296 126686 93372 127030
rect 92822 126622 92823 126654
rect 92757 126621 92823 126622
rect 93296 126622 93302 126686
rect 93366 126622 93372 126686
rect 93296 126616 93372 126622
rect 94656 127030 94662 127062
rect 94726 127062 94727 127094
rect 95336 127094 95412 127100
rect 94726 127030 94732 127062
rect 94656 126686 94732 127030
rect 94656 126622 94662 126686
rect 94726 126622 94732 126686
rect 95336 127030 95342 127094
rect 95406 127030 95412 127094
rect 95749 127094 95815 127095
rect 95749 127062 95750 127094
rect 95336 126686 95412 127030
rect 95336 126654 95342 126686
rect 94656 126616 94732 126622
rect 95341 126622 95342 126654
rect 95406 126654 95412 126686
rect 95744 127030 95750 127062
rect 95814 127062 95815 127094
rect 96560 127094 96636 127100
rect 95814 127030 95820 127062
rect 95744 126686 95820 127030
rect 95406 126622 95407 126654
rect 95341 126621 95407 126622
rect 95744 126622 95750 126686
rect 95814 126622 95820 126686
rect 96560 127030 96566 127094
rect 96630 127030 96636 127094
rect 97109 127094 97175 127095
rect 97109 127062 97110 127094
rect 96560 126686 96636 127030
rect 96560 126654 96566 126686
rect 95744 126616 95820 126622
rect 96565 126622 96566 126654
rect 96630 126654 96636 126686
rect 97104 127030 97110 127062
rect 97174 127062 97175 127094
rect 97925 127094 97991 127095
rect 97925 127062 97926 127094
rect 97174 127030 97180 127062
rect 97104 126686 97180 127030
rect 96630 126622 96631 126654
rect 96565 126621 96631 126622
rect 97104 126622 97110 126686
rect 97174 126622 97180 126686
rect 97104 126616 97180 126622
rect 97920 127030 97926 127062
rect 97990 127062 97991 127094
rect 99557 127094 99623 127095
rect 99557 127062 99558 127094
rect 97990 127030 97996 127062
rect 89216 126486 89222 126550
rect 89286 126486 89292 126550
rect 89216 126480 89292 126486
rect 97920 126550 97996 127030
rect 99552 127030 99558 127062
rect 99622 127062 99623 127094
rect 100232 127094 100308 127100
rect 99622 127030 99628 127062
rect 99552 126686 99628 127030
rect 99552 126622 99558 126686
rect 99622 126622 99628 126686
rect 100232 127030 100238 127094
rect 100302 127030 100308 127094
rect 100509 127094 100575 127095
rect 100509 127062 100510 127094
rect 100232 126686 100308 127030
rect 100232 126654 100238 126686
rect 99552 126616 99628 126622
rect 100237 126622 100238 126654
rect 100302 126654 100308 126686
rect 100504 127030 100510 127062
rect 100574 127062 100575 127094
rect 102005 127094 102071 127095
rect 102005 127062 102006 127094
rect 100574 127030 100580 127062
rect 100504 126686 100580 127030
rect 100302 126622 100303 126654
rect 100237 126621 100303 126622
rect 100504 126622 100510 126686
rect 100574 126622 100580 126686
rect 100504 126616 100580 126622
rect 102000 127030 102006 127062
rect 102070 127062 102071 127094
rect 103365 127094 103431 127095
rect 103365 127062 103366 127094
rect 102070 127030 102076 127062
rect 102000 126686 102076 127030
rect 102000 126622 102006 126686
rect 102070 126622 102076 126686
rect 102000 126616 102076 126622
rect 103360 127030 103366 127062
rect 103430 127062 103431 127094
rect 104040 127094 104116 127100
rect 103430 127030 103436 127062
rect 103360 126686 103436 127030
rect 103360 126622 103366 126686
rect 103430 126622 103436 126686
rect 104040 127030 104046 127094
rect 104110 127030 104116 127094
rect 104589 127094 104655 127095
rect 104589 127062 104590 127094
rect 104040 126686 104116 127030
rect 104040 126654 104046 126686
rect 103360 126616 103436 126622
rect 104045 126622 104046 126654
rect 104110 126654 104116 126686
rect 104584 127030 104590 127062
rect 104654 127062 104655 127094
rect 105264 127094 105340 127100
rect 104654 127030 104660 127062
rect 104584 126686 104660 127030
rect 104110 126622 104111 126654
rect 104045 126621 104111 126622
rect 104584 126622 104590 126686
rect 104654 126622 104660 126686
rect 105264 127030 105270 127094
rect 105334 127030 105340 127094
rect 105813 127094 105879 127095
rect 105813 127062 105814 127094
rect 105264 126686 105340 127030
rect 105264 126654 105270 126686
rect 104584 126616 104660 126622
rect 105269 126622 105270 126654
rect 105334 126654 105340 126686
rect 105808 127030 105814 127062
rect 105878 127062 105879 127094
rect 106488 127094 106564 127100
rect 105878 127030 105884 127062
rect 105808 126686 105884 127030
rect 105334 126622 105335 126654
rect 105269 126621 105335 126622
rect 105808 126622 105814 126686
rect 105878 126622 105884 126686
rect 106488 127030 106494 127094
rect 106558 127030 106564 127094
rect 106488 126686 106564 127030
rect 106488 126654 106494 126686
rect 105808 126616 105884 126622
rect 106493 126622 106494 126654
rect 106558 126654 106564 126686
rect 108120 127094 108196 127100
rect 108120 127030 108126 127094
rect 108190 127030 108196 127094
rect 109213 127094 109279 127095
rect 109213 127062 109214 127094
rect 108120 126686 108196 127030
rect 108120 126654 108126 126686
rect 106558 126622 106559 126654
rect 106493 126621 106559 126622
rect 108125 126622 108126 126654
rect 108190 126654 108196 126686
rect 109208 127030 109214 127062
rect 109278 127062 109279 127094
rect 110296 127094 110372 127100
rect 109278 127030 109284 127062
rect 109208 126686 109284 127030
rect 108190 126622 108191 126654
rect 108125 126621 108191 126622
rect 109208 126622 109214 126686
rect 109278 126622 109284 126686
rect 110296 127030 110302 127094
rect 110366 127030 110372 127094
rect 110845 127094 110911 127095
rect 110845 127062 110846 127094
rect 110296 126686 110372 127030
rect 110296 126654 110302 126686
rect 109208 126616 109284 126622
rect 110301 126622 110302 126654
rect 110366 126654 110372 126686
rect 110840 127030 110846 127062
rect 110910 127062 110911 127094
rect 111520 127094 111596 127100
rect 110910 127030 110916 127062
rect 110840 126686 110916 127030
rect 110366 126622 110367 126654
rect 110301 126621 110367 126622
rect 110840 126622 110846 126686
rect 110910 126622 110916 126686
rect 111520 127030 111526 127094
rect 111590 127030 111596 127094
rect 112069 127094 112135 127095
rect 112069 127062 112070 127094
rect 111520 126686 111596 127030
rect 111520 126654 111526 126686
rect 110840 126616 110916 126622
rect 111525 126622 111526 126654
rect 111590 126654 111596 126686
rect 112064 127030 112070 127062
rect 112134 127062 112135 127094
rect 112744 127094 112820 127100
rect 112134 127030 112140 127062
rect 112064 126686 112140 127030
rect 111590 126622 111591 126654
rect 111525 126621 111591 126622
rect 112064 126622 112070 126686
rect 112134 126622 112140 126686
rect 112744 127030 112750 127094
rect 112814 127030 112820 127094
rect 113293 127094 113359 127095
rect 113293 127062 113294 127094
rect 112744 126686 112820 127030
rect 112744 126654 112750 126686
rect 112064 126616 112140 126622
rect 112749 126622 112750 126654
rect 112814 126654 112820 126686
rect 113288 127030 113294 127062
rect 113358 127062 113359 127094
rect 114517 127094 114583 127095
rect 114517 127062 114518 127094
rect 113358 127030 113364 127062
rect 113288 126686 113364 127030
rect 112814 126622 112815 126654
rect 112749 126621 112815 126622
rect 113288 126622 113294 126686
rect 113358 126622 113364 126686
rect 113288 126616 113364 126622
rect 114512 127030 114518 127062
rect 114582 127062 114583 127094
rect 115741 127094 115807 127095
rect 115741 127062 115742 127094
rect 114582 127030 114588 127062
rect 114512 126686 114588 127030
rect 114512 126622 114518 126686
rect 114582 126622 114588 126686
rect 114512 126616 114588 126622
rect 115736 127030 115742 127062
rect 115806 127062 115807 127094
rect 116552 127094 116628 127100
rect 115806 127030 115812 127062
rect 115736 126686 115812 127030
rect 115736 126622 115742 126686
rect 115806 126622 115812 126686
rect 116552 127030 116558 127094
rect 116622 127030 116628 127094
rect 117645 127094 117711 127095
rect 117645 127062 117646 127094
rect 116552 126686 116628 127030
rect 116552 126654 116558 126686
rect 115736 126616 115812 126622
rect 116557 126622 116558 126654
rect 116622 126654 116628 126686
rect 117640 127030 117646 127062
rect 117710 127062 117711 127094
rect 117776 127094 117852 127100
rect 117710 127030 117716 127062
rect 117640 126686 117716 127030
rect 116622 126622 116623 126654
rect 116557 126621 116623 126622
rect 117640 126622 117646 126686
rect 117710 126622 117716 126686
rect 117776 127030 117782 127094
rect 117846 127030 117852 127094
rect 118325 127094 118391 127095
rect 118325 127062 118326 127094
rect 117776 126686 117852 127030
rect 117776 126654 117782 126686
rect 117640 126616 117716 126622
rect 117781 126622 117782 126654
rect 117846 126654 117852 126686
rect 118320 127030 118326 127062
rect 118390 127062 118391 127094
rect 119000 127094 119076 127100
rect 118390 127030 118396 127062
rect 118320 126686 118396 127030
rect 117846 126622 117847 126654
rect 117781 126621 117847 126622
rect 118320 126622 118326 126686
rect 118390 126622 118396 126686
rect 119000 127030 119006 127094
rect 119070 127030 119076 127094
rect 119549 127094 119615 127095
rect 119549 127062 119550 127094
rect 119000 126686 119076 127030
rect 119000 126654 119006 126686
rect 118320 126616 118396 126622
rect 119005 126622 119006 126654
rect 119070 126654 119076 126686
rect 119544 127030 119550 127062
rect 119614 127062 119615 127094
rect 120773 127094 120839 127095
rect 120773 127062 120774 127094
rect 119614 127030 119620 127062
rect 119544 126686 119620 127030
rect 119070 126622 119071 126654
rect 119005 126621 119071 126622
rect 119544 126622 119550 126686
rect 119614 126622 119620 126686
rect 119544 126616 119620 126622
rect 120768 127030 120774 127062
rect 120838 127062 120839 127094
rect 121448 127094 121524 127100
rect 120838 127030 120844 127062
rect 120768 126686 120844 127030
rect 120768 126622 120774 126686
rect 120838 126622 120844 126686
rect 121448 127030 121454 127094
rect 121518 127030 121524 127094
rect 121997 127094 122063 127095
rect 121997 127062 121998 127094
rect 121448 126686 121524 127030
rect 121448 126654 121454 126686
rect 120768 126616 120844 126622
rect 121453 126622 121454 126654
rect 121518 126654 121524 126686
rect 121992 127030 121998 127062
rect 122062 127062 122063 127094
rect 122949 127094 123015 127095
rect 122949 127062 122950 127094
rect 122062 127030 122068 127062
rect 121992 126686 122068 127030
rect 121518 126622 121519 126654
rect 121453 126621 121519 126622
rect 121992 126622 121998 126686
rect 122062 126622 122068 126686
rect 121992 126616 122068 126622
rect 122944 127030 122950 127062
rect 123014 127062 123015 127094
rect 123901 127094 123967 127095
rect 123901 127062 123902 127094
rect 123014 127030 123020 127062
rect 122944 126686 123020 127030
rect 122944 126622 122950 126686
rect 123014 126622 123020 126686
rect 122944 126616 123020 126622
rect 123896 127030 123902 127062
rect 123966 127062 123967 127094
rect 124309 127094 124375 127095
rect 124309 127062 124310 127094
rect 123966 127030 123972 127062
rect 123896 126686 123972 127030
rect 123896 126622 123902 126686
rect 123966 126622 123972 126686
rect 123896 126616 123972 126622
rect 124304 127030 124310 127062
rect 124374 127062 124375 127094
rect 125256 127094 125332 127100
rect 124374 127030 124380 127062
rect 124304 126692 124380 127030
rect 125256 127030 125262 127094
rect 125326 127030 125332 127094
rect 125805 127094 125871 127095
rect 125805 127062 125806 127094
rect 124304 126686 124516 126692
rect 124304 126622 124446 126686
rect 124510 126622 124516 126686
rect 125256 126686 125332 127030
rect 125256 126654 125262 126686
rect 124304 126616 124516 126622
rect 125261 126622 125262 126654
rect 125326 126654 125332 126686
rect 125800 127030 125806 127062
rect 125870 127062 125871 127094
rect 126480 127094 126556 127100
rect 125870 127030 125876 127062
rect 125800 126686 125876 127030
rect 125326 126622 125327 126654
rect 125261 126621 125327 126622
rect 125800 126622 125806 126686
rect 125870 126622 125876 126686
rect 126480 127030 126486 127094
rect 126550 127030 126556 127094
rect 127029 127094 127095 127095
rect 127029 127062 127030 127094
rect 126480 126686 126556 127030
rect 126480 126654 126486 126686
rect 125800 126616 125876 126622
rect 126485 126622 126486 126654
rect 126550 126654 126556 126686
rect 127024 127030 127030 127062
rect 127094 127062 127095 127094
rect 128253 127094 128319 127095
rect 128253 127062 128254 127094
rect 127094 127030 127100 127062
rect 127024 126686 127100 127030
rect 126550 126622 126551 126654
rect 126485 126621 126551 126622
rect 127024 126622 127030 126686
rect 127094 126622 127100 126686
rect 127024 126616 127100 126622
rect 128248 127030 128254 127062
rect 128318 127062 128319 127094
rect 128928 127094 129004 127100
rect 128318 127030 128324 127062
rect 128248 126686 128324 127030
rect 128248 126622 128254 126686
rect 128318 126622 128324 126686
rect 128928 127030 128934 127094
rect 128998 127030 129004 127094
rect 129477 127094 129543 127095
rect 129477 127062 129478 127094
rect 128928 126686 129004 127030
rect 128928 126654 128934 126686
rect 128248 126616 128324 126622
rect 128933 126622 128934 126654
rect 128998 126654 129004 126686
rect 129472 127030 129478 127062
rect 129542 127062 129543 127094
rect 130288 127094 130364 127100
rect 129542 127030 129548 127062
rect 129472 126686 129548 127030
rect 128998 126622 128999 126654
rect 128933 126621 128999 126622
rect 129472 126622 129478 126686
rect 129542 126622 129548 126686
rect 130288 127030 130294 127094
rect 130358 127030 130364 127094
rect 130837 127094 130903 127095
rect 130837 127062 130838 127094
rect 130288 126686 130364 127030
rect 130288 126654 130294 126686
rect 129472 126616 129548 126622
rect 130293 126622 130294 126654
rect 130358 126654 130364 126686
rect 130832 127030 130838 127062
rect 130902 127062 130903 127094
rect 132061 127094 132127 127095
rect 132061 127062 132062 127094
rect 130902 127030 130908 127062
rect 130832 126686 130908 127030
rect 130358 126622 130359 126654
rect 130293 126621 130359 126622
rect 130832 126622 130838 126686
rect 130902 126622 130908 126686
rect 130832 126616 130908 126622
rect 132056 127030 132062 127062
rect 132126 127062 132127 127094
rect 133285 127094 133351 127095
rect 133285 127062 133286 127094
rect 132126 127030 132132 127062
rect 132056 126686 132132 127030
rect 132056 126622 132062 126686
rect 132126 126622 132132 126686
rect 132056 126616 132132 126622
rect 133280 127030 133286 127062
rect 133350 127062 133351 127094
rect 133960 127094 134036 127100
rect 133350 127030 133356 127062
rect 133280 126686 133356 127030
rect 133280 126622 133286 126686
rect 133350 126622 133356 126686
rect 133960 127030 133966 127094
rect 134030 127030 134036 127094
rect 134509 127094 134575 127095
rect 134509 127062 134510 127094
rect 133960 126686 134036 127030
rect 133960 126654 133966 126686
rect 133280 126616 133356 126622
rect 133965 126622 133966 126654
rect 134030 126654 134036 126686
rect 134504 127030 134510 127062
rect 134574 127062 134575 127094
rect 135184 127094 135260 127100
rect 134574 127030 134580 127062
rect 134504 126686 134580 127030
rect 134030 126622 134031 126654
rect 133965 126621 134031 126622
rect 134504 126622 134510 126686
rect 134574 126622 134580 126686
rect 135184 127030 135190 127094
rect 135254 127030 135260 127094
rect 135461 127094 135527 127095
rect 135461 127062 135462 127094
rect 135184 126686 135260 127030
rect 135184 126654 135190 126686
rect 134504 126616 134580 126622
rect 135189 126622 135190 126654
rect 135254 126654 135260 126686
rect 135456 127030 135462 127062
rect 135526 127062 135527 127094
rect 137093 127094 137159 127095
rect 137093 127062 137094 127094
rect 135526 127030 135532 127062
rect 135456 126686 135532 127030
rect 135254 126622 135255 126654
rect 135189 126621 135255 126622
rect 135456 126622 135462 126686
rect 135526 126622 135532 126686
rect 135456 126616 135532 126622
rect 137088 127030 137094 127062
rect 137158 127062 137159 127094
rect 138181 127094 138247 127095
rect 138181 127062 138182 127094
rect 137158 127030 137164 127062
rect 137088 126686 137164 127030
rect 137088 126622 137094 126686
rect 137158 126622 137164 126686
rect 137088 126616 137164 126622
rect 138176 127030 138182 127062
rect 138246 127062 138247 127094
rect 139541 127094 139607 127095
rect 139541 127062 139542 127094
rect 138246 127030 138252 127062
rect 138176 126686 138252 127030
rect 138176 126622 138182 126686
rect 138246 126622 138252 126686
rect 138176 126616 138252 126622
rect 139536 127030 139542 127062
rect 139606 127062 139607 127094
rect 140357 127094 140423 127095
rect 140357 127062 140358 127094
rect 139606 127030 139612 127062
rect 139536 126686 139612 127030
rect 139536 126622 139542 126686
rect 139606 126622 139612 126686
rect 139536 126616 139612 126622
rect 140352 127030 140358 127062
rect 140422 127062 140423 127094
rect 141440 127094 141516 127100
rect 140422 127030 140428 127062
rect 140352 126686 140428 127030
rect 140352 126622 140358 126686
rect 140422 126622 140428 126686
rect 141440 127030 141446 127094
rect 141510 127030 141516 127094
rect 141989 127094 142055 127095
rect 141989 127062 141990 127094
rect 141440 126686 141516 127030
rect 141440 126654 141446 126686
rect 140352 126616 140428 126622
rect 141445 126622 141446 126654
rect 141510 126654 141516 126686
rect 141984 127030 141990 127062
rect 142054 127062 142055 127094
rect 142664 127094 142740 127100
rect 142054 127030 142060 127062
rect 141984 126686 142060 127030
rect 141510 126622 141511 126654
rect 141445 126621 141511 126622
rect 141984 126622 141990 126686
rect 142054 126622 142060 126686
rect 142664 127030 142670 127094
rect 142734 127030 142740 127094
rect 144437 127094 144503 127095
rect 144437 127062 144438 127094
rect 142664 126686 142740 127030
rect 142664 126654 142670 126686
rect 141984 126616 142060 126622
rect 142669 126622 142670 126654
rect 142734 126654 142740 126686
rect 144432 127030 144438 127062
rect 144502 127062 144503 127094
rect 145248 127094 145324 127100
rect 144502 127030 144508 127062
rect 144432 126686 144508 127030
rect 142734 126622 142735 126654
rect 142669 126621 142735 126622
rect 144432 126622 144438 126686
rect 144502 126622 144508 126686
rect 145248 127030 145254 127094
rect 145318 127030 145324 127094
rect 145248 126686 145324 127030
rect 145248 126654 145254 126686
rect 144432 126616 144508 126622
rect 145253 126622 145254 126654
rect 145318 126654 145324 126686
rect 146472 127094 146548 127100
rect 146472 127030 146478 127094
rect 146542 127030 146548 127094
rect 147021 127094 147087 127095
rect 147021 127062 147022 127094
rect 146472 126686 146548 127030
rect 146472 126654 146478 126686
rect 145318 126622 145319 126654
rect 145253 126621 145319 126622
rect 146477 126622 146478 126654
rect 146542 126654 146548 126686
rect 147016 127030 147022 127062
rect 147086 127062 147087 127094
rect 147696 127094 147772 127100
rect 147086 127030 147092 127062
rect 147016 126686 147092 127030
rect 146542 126622 146543 126654
rect 146477 126621 146543 126622
rect 147016 126622 147022 126686
rect 147086 126622 147092 126686
rect 147696 127030 147702 127094
rect 147766 127030 147772 127094
rect 148245 127094 148311 127095
rect 148245 127062 148246 127094
rect 147696 126686 147772 127030
rect 147696 126654 147702 126686
rect 147016 126616 147092 126622
rect 147701 126622 147702 126654
rect 147766 126654 147772 126686
rect 148240 127030 148246 127062
rect 148310 127062 148311 127094
rect 150144 127094 150220 127100
rect 148310 127030 148316 127062
rect 148240 126686 148316 127030
rect 150144 127030 150150 127094
rect 150214 127030 150220 127094
rect 149469 126958 149535 126959
rect 149469 126926 149470 126958
rect 147766 126622 147767 126654
rect 147701 126621 147767 126622
rect 148240 126622 148246 126686
rect 148310 126622 148316 126686
rect 148240 126616 148316 126622
rect 149464 126894 149470 126926
rect 149534 126926 149535 126958
rect 149534 126894 149540 126926
rect 149464 126686 149540 126894
rect 149464 126622 149470 126686
rect 149534 126622 149540 126686
rect 150144 126686 150220 127030
rect 150144 126654 150150 126686
rect 149464 126616 149540 126622
rect 150149 126622 150150 126654
rect 150214 126654 150220 126686
rect 151504 127094 151580 127100
rect 151504 127030 151510 127094
rect 151574 127030 151580 127094
rect 151917 127094 151983 127095
rect 151917 127062 151918 127094
rect 151504 126686 151580 127030
rect 151504 126654 151510 126686
rect 150214 126622 150215 126654
rect 150149 126621 150215 126622
rect 151509 126622 151510 126654
rect 151574 126654 151580 126686
rect 151912 127030 151918 127062
rect 151982 127062 151983 127094
rect 153277 127094 153343 127095
rect 153277 127062 153278 127094
rect 151982 127030 151988 127062
rect 151912 126686 151988 127030
rect 151574 126622 151575 126654
rect 151509 126621 151575 126622
rect 151912 126622 151918 126686
rect 151982 126622 151988 126686
rect 151912 126616 151988 126622
rect 153272 127030 153278 127062
rect 153342 127062 153343 127094
rect 153952 127094 154028 127100
rect 153342 127030 153348 127062
rect 153272 126686 153348 127030
rect 153272 126622 153278 126686
rect 153342 126622 153348 126686
rect 153952 127030 153958 127094
rect 154022 127030 154028 127094
rect 154501 127094 154567 127095
rect 154501 127062 154502 127094
rect 153952 126686 154028 127030
rect 153952 126654 153958 126686
rect 153272 126616 153348 126622
rect 153957 126622 153958 126654
rect 154022 126654 154028 126686
rect 154496 127030 154502 127062
rect 154566 127062 154567 127094
rect 155176 127094 155252 127100
rect 154566 127030 154572 127062
rect 154496 126686 154572 127030
rect 154022 126622 154023 126654
rect 153957 126621 154023 126622
rect 154496 126622 154502 126686
rect 154566 126622 154572 126686
rect 155176 127030 155182 127094
rect 155246 127030 155252 127094
rect 155725 127094 155791 127095
rect 155725 127062 155726 127094
rect 155176 126686 155252 127030
rect 155176 126654 155182 126686
rect 154496 126616 154572 126622
rect 155181 126622 155182 126654
rect 155246 126654 155252 126686
rect 155720 127030 155726 127062
rect 155790 127062 155791 127094
rect 156677 127094 156743 127095
rect 156677 127062 156678 127094
rect 155790 127030 155796 127062
rect 155720 126686 155796 127030
rect 155246 126622 155247 126654
rect 155181 126621 155247 126622
rect 155720 126622 155726 126686
rect 155790 126622 155796 126686
rect 155720 126616 155796 126622
rect 156672 127030 156678 127062
rect 156742 127062 156743 127094
rect 157901 127094 157967 127095
rect 157901 127062 157902 127094
rect 156742 127030 156748 127062
rect 156672 126686 156748 127030
rect 156672 126622 156678 126686
rect 156742 126622 156748 126686
rect 156672 126616 156748 126622
rect 157896 127030 157902 127062
rect 157966 127062 157967 127094
rect 158984 127094 159060 127100
rect 157966 127030 157972 127062
rect 97920 126486 97926 126550
rect 97990 126486 97996 126550
rect 97920 126480 97996 126486
rect 157896 126550 157972 127030
rect 158984 127030 158990 127094
rect 159054 127030 159060 127094
rect 158984 126686 159060 127030
rect 158984 126654 158990 126686
rect 158989 126622 158990 126654
rect 159054 126654 159060 126686
rect 160208 127094 160284 127100
rect 160208 127030 160214 127094
rect 160278 127030 160284 127094
rect 160757 127094 160823 127095
rect 160757 127062 160758 127094
rect 160208 126686 160284 127030
rect 160208 126654 160214 126686
rect 159054 126622 159055 126654
rect 158989 126621 159055 126622
rect 160213 126622 160214 126654
rect 160278 126654 160284 126686
rect 160752 127030 160758 127062
rect 160822 127062 160823 127094
rect 161981 127094 162047 127095
rect 161981 127062 161982 127094
rect 160822 127030 160828 127062
rect 160752 126686 160828 127030
rect 160278 126622 160279 126654
rect 160213 126621 160279 126622
rect 160752 126622 160758 126686
rect 160822 126622 160828 126686
rect 160752 126616 160828 126622
rect 161976 127030 161982 127062
rect 162046 127062 162047 127094
rect 163205 127094 163271 127095
rect 163205 127062 163206 127094
rect 162046 127030 162052 127062
rect 161976 126686 162052 127030
rect 161976 126622 161982 126686
rect 162046 126622 162052 126686
rect 161976 126616 162052 126622
rect 163200 127030 163206 127062
rect 163270 127062 163271 127094
rect 163880 127094 163956 127100
rect 163270 127030 163276 127062
rect 163200 126686 163276 127030
rect 163200 126622 163206 126686
rect 163270 126622 163276 126686
rect 163880 127030 163886 127094
rect 163950 127030 163956 127094
rect 164429 127094 164495 127095
rect 164429 127062 164430 127094
rect 163880 126686 163956 127030
rect 163880 126654 163886 126686
rect 163200 126616 163276 126622
rect 163885 126622 163886 126654
rect 163950 126654 163956 126686
rect 164424 127030 164430 127062
rect 164494 127062 164495 127094
rect 165381 127094 165447 127095
rect 165381 127062 165382 127094
rect 164494 127030 164500 127062
rect 164424 126686 164500 127030
rect 163950 126622 163951 126654
rect 163885 126621 163951 126622
rect 164424 126622 164430 126686
rect 164494 126622 164500 126686
rect 164424 126616 164500 126622
rect 165376 127030 165382 127062
rect 165446 127062 165447 127094
rect 166333 127094 166399 127095
rect 166333 127062 166334 127094
rect 165446 127030 165452 127062
rect 165376 126686 165452 127030
rect 165376 126622 165382 126686
rect 165446 126622 165452 126686
rect 165376 126616 165452 126622
rect 166328 127030 166334 127062
rect 166398 127062 166399 127094
rect 166464 127094 166540 127100
rect 166398 127030 166404 127062
rect 166328 126686 166404 127030
rect 166328 126622 166334 126686
rect 166398 126622 166404 126686
rect 166464 127030 166470 127094
rect 166534 127030 166540 127094
rect 168237 127094 168303 127095
rect 168237 127062 168238 127094
rect 166464 126686 166540 127030
rect 166464 126654 166470 126686
rect 166328 126616 166404 126622
rect 166469 126622 166470 126654
rect 166534 126654 166540 126686
rect 168232 127030 168238 127062
rect 168302 127062 168303 127094
rect 168912 127094 168988 127100
rect 168302 127030 168308 127062
rect 168232 126686 168308 127030
rect 166534 126622 166535 126654
rect 166469 126621 166535 126622
rect 168232 126622 168238 126686
rect 168302 126622 168308 126686
rect 168912 127030 168918 127094
rect 168982 127030 168988 127094
rect 169461 127094 169527 127095
rect 169461 127062 169462 127094
rect 168912 126686 168988 127030
rect 168912 126654 168918 126686
rect 168232 126616 168308 126622
rect 168917 126622 168918 126654
rect 168982 126654 168988 126686
rect 169456 127030 169462 127062
rect 169526 127062 169527 127094
rect 170685 127094 170751 127095
rect 170685 127062 170686 127094
rect 169526 127030 169532 127062
rect 169456 126686 169532 127030
rect 168982 126622 168983 126654
rect 168917 126621 168983 126622
rect 169456 126622 169462 126686
rect 169526 126622 169532 126686
rect 169456 126616 169532 126622
rect 170680 127030 170686 127062
rect 170750 127062 170751 127094
rect 171360 127094 171436 127100
rect 170750 127030 170756 127062
rect 170680 126686 170756 127030
rect 170680 126622 170686 126686
rect 170750 126622 170756 126686
rect 171360 127030 171366 127094
rect 171430 127030 171436 127094
rect 171909 127094 171975 127095
rect 171909 127062 171910 127094
rect 171360 126686 171436 127030
rect 171360 126654 171366 126686
rect 170680 126616 170756 126622
rect 171365 126622 171366 126654
rect 171430 126654 171436 126686
rect 171904 127030 171910 127062
rect 171974 127062 171975 127094
rect 173133 127094 173199 127095
rect 173133 127062 173134 127094
rect 171974 127030 171980 127062
rect 171904 126686 171980 127030
rect 171430 126622 171431 126654
rect 171365 126621 171431 126622
rect 171904 126622 171910 126686
rect 171974 126622 171980 126686
rect 171904 126616 171980 126622
rect 173128 127030 173134 127062
rect 173198 127062 173199 127094
rect 174493 127094 174559 127095
rect 174493 127062 174494 127094
rect 173198 127030 173204 127062
rect 173128 126686 173204 127030
rect 173128 126622 173134 126686
rect 173198 126622 173204 126686
rect 173128 126616 173204 126622
rect 174488 127030 174494 127062
rect 174558 127062 174559 127094
rect 175168 127094 175244 127100
rect 174558 127030 174564 127062
rect 174488 126686 174564 127030
rect 174488 126622 174494 126686
rect 174558 126622 174564 126686
rect 175168 127030 175174 127094
rect 175238 127030 175244 127094
rect 175717 127094 175783 127095
rect 175717 127062 175718 127094
rect 175168 126686 175244 127030
rect 175168 126654 175174 126686
rect 174488 126616 174564 126622
rect 175173 126622 175174 126654
rect 175238 126654 175244 126686
rect 175712 127030 175718 127062
rect 175782 127062 175783 127094
rect 176941 127094 177007 127095
rect 176941 127062 176942 127094
rect 175782 127030 175788 127062
rect 175712 126686 175788 127030
rect 175238 126622 175239 126654
rect 175173 126621 175239 126622
rect 175712 126622 175718 126686
rect 175782 126622 175788 126686
rect 175712 126616 175788 126622
rect 176936 127030 176942 127062
rect 177006 127062 177007 127094
rect 178165 127094 178231 127095
rect 178165 127062 178166 127094
rect 177006 127030 177012 127062
rect 176936 126686 177012 127030
rect 176936 126622 176942 126686
rect 177006 126622 177012 126686
rect 176936 126616 177012 126622
rect 178160 127030 178166 127062
rect 178230 127062 178231 127094
rect 178976 127094 179052 127100
rect 178230 127030 178236 127062
rect 178160 126686 178236 127030
rect 178160 126622 178166 126686
rect 178230 126622 178236 126686
rect 178976 127030 178982 127094
rect 179046 127030 179052 127094
rect 178976 126686 179052 127030
rect 178976 126654 178982 126686
rect 178160 126616 178236 126622
rect 178981 126622 178982 126654
rect 179046 126654 179052 126686
rect 180200 127094 180276 127100
rect 180200 127030 180206 127094
rect 180270 127030 180276 127094
rect 180613 127094 180679 127095
rect 180613 127062 180614 127094
rect 180200 126686 180276 127030
rect 180200 126654 180206 126686
rect 179046 126622 179047 126654
rect 178981 126621 179047 126622
rect 180205 126622 180206 126654
rect 180270 126654 180276 126686
rect 180608 127030 180614 127062
rect 180678 127062 180679 127094
rect 181424 127094 181500 127100
rect 180678 127030 180684 127062
rect 180608 126686 180684 127030
rect 180270 126622 180271 126654
rect 180205 126621 180271 126622
rect 180608 126622 180614 126686
rect 180678 126622 180684 126686
rect 181424 127030 181430 127094
rect 181494 127030 181500 127094
rect 181973 127094 182039 127095
rect 181973 127062 181974 127094
rect 181424 126686 181500 127030
rect 181424 126654 181430 126686
rect 180608 126616 180684 126622
rect 181429 126622 181430 126654
rect 181494 126654 181500 126686
rect 181968 127030 181974 127062
rect 182038 127062 182039 127094
rect 183197 127094 183263 127095
rect 183197 127062 183198 127094
rect 182038 127030 182044 127062
rect 181968 126686 182044 127030
rect 181494 126622 181495 126654
rect 181429 126621 181495 126622
rect 181968 126622 181974 126686
rect 182038 126622 182044 126686
rect 181968 126616 182044 126622
rect 183192 127030 183198 127062
rect 183262 127062 183263 127094
rect 184008 127094 184084 127100
rect 183262 127030 183268 127062
rect 183192 126686 183268 127030
rect 183192 126622 183198 126686
rect 183262 126622 183268 126686
rect 184008 127030 184014 127094
rect 184078 127030 184084 127094
rect 184008 126686 184084 127030
rect 184008 126654 184014 126686
rect 183192 126616 183268 126622
rect 184013 126622 184014 126654
rect 184078 126654 184084 126686
rect 184280 127094 184356 127100
rect 184280 127030 184286 127094
rect 184350 127030 184356 127094
rect 184280 126686 184356 127030
rect 184280 126654 184286 126686
rect 184078 126622 184079 126654
rect 184013 126621 184079 126622
rect 184285 126622 184286 126654
rect 184350 126654 184356 126686
rect 184960 127094 185036 127100
rect 184960 127030 184966 127094
rect 185030 127030 185036 127094
rect 184960 126686 185036 127030
rect 184960 126654 184966 126686
rect 184350 126622 184351 126654
rect 184285 126621 184351 126622
rect 184965 126622 184966 126654
rect 185030 126654 185036 126686
rect 185232 127094 185308 127100
rect 185232 127030 185238 127094
rect 185302 127030 185308 127094
rect 185373 127094 185439 127095
rect 185373 127062 185374 127094
rect 185232 126686 185308 127030
rect 185232 126654 185238 126686
rect 185030 126622 185031 126654
rect 184965 126621 185031 126622
rect 185237 126622 185238 126654
rect 185302 126654 185308 126686
rect 185368 127030 185374 127062
rect 185438 127062 185439 127094
rect 187005 127094 187071 127095
rect 187005 127062 187006 127094
rect 185438 127030 185444 127062
rect 185368 126686 185444 127030
rect 185302 126622 185303 126654
rect 185237 126621 185303 126622
rect 185368 126622 185374 126686
rect 185438 126622 185444 126686
rect 185368 126616 185444 126622
rect 187000 127030 187006 127062
rect 187070 127062 187071 127094
rect 188229 127094 188295 127095
rect 188229 127062 188230 127094
rect 187070 127030 187076 127062
rect 187000 126686 187076 127030
rect 187000 126622 187006 126686
rect 187070 126622 187076 126686
rect 187000 126616 187076 126622
rect 188224 127030 188230 127062
rect 188294 127062 188295 127094
rect 188904 127094 188980 127100
rect 188294 127030 188300 127062
rect 188224 126686 188300 127030
rect 188224 126622 188230 126686
rect 188294 126622 188300 126686
rect 188904 127030 188910 127094
rect 188974 127030 188980 127094
rect 189453 127094 189519 127095
rect 189453 127062 189454 127094
rect 188904 126686 188980 127030
rect 188904 126654 188910 126686
rect 188224 126616 188300 126622
rect 188909 126622 188910 126654
rect 188974 126654 188980 126686
rect 189448 127030 189454 127062
rect 189518 127062 189519 127094
rect 189518 127030 189524 127062
rect 189448 126686 189524 127030
rect 188974 126622 188975 126654
rect 188909 126621 188975 126622
rect 189448 126622 189454 126686
rect 189518 126622 189524 126686
rect 189448 126616 189524 126622
rect 157896 126486 157902 126550
rect 157966 126486 157972 126550
rect 157896 126480 157972 126486
rect 28832 126382 28838 126414
rect 28837 126350 28838 126382
rect 28902 126382 28908 126414
rect 190400 126414 190476 128526
rect 191493 126550 191559 126551
rect 191493 126518 191494 126550
rect 28902 126350 28903 126382
rect 28837 126349 28903 126350
rect 190400 126350 190406 126414
rect 190470 126350 190476 126414
rect 190400 126344 190476 126350
rect 191488 126486 191494 126518
rect 191558 126518 191559 126550
rect 191558 126486 191564 126518
rect 28293 126278 28359 126279
rect 28293 126246 28294 126278
rect 28288 126214 28294 126246
rect 28358 126246 28359 126278
rect 190400 126278 190476 126284
rect 28358 126214 28364 126246
rect 28288 126006 28364 126214
rect 28288 125942 28294 126006
rect 28358 125942 28364 126006
rect 190400 126214 190406 126278
rect 190470 126214 190476 126278
rect 190400 126006 190476 126214
rect 191488 126278 191564 126486
rect 191488 126214 191494 126278
rect 191558 126214 191564 126278
rect 196520 126278 196596 129750
rect 197880 128590 197956 131246
rect 203320 129814 203396 132470
rect 203456 132470 203462 132534
rect 203526 132470 203532 132534
rect 203456 131446 203532 132470
rect 203456 131414 203462 131446
rect 203461 131382 203462 131414
rect 203526 131414 203532 131446
rect 203526 131382 203527 131414
rect 203461 131381 203527 131382
rect 203592 131174 203668 133830
rect 203592 131110 203598 131174
rect 203662 131110 203668 131174
rect 203592 131104 203668 131110
rect 217464 133350 217812 134782
rect 217464 133286 217470 133350
rect 217534 133286 217812 133350
rect 217464 131582 217812 133286
rect 217464 131518 217470 131582
rect 217534 131518 217812 131582
rect 203597 131038 203663 131039
rect 203597 131006 203598 131038
rect 203320 129750 203326 129814
rect 203390 129750 203396 129814
rect 203320 129744 203396 129750
rect 203592 130974 203598 131006
rect 203662 131006 203663 131038
rect 203662 130974 203668 131006
rect 203461 129678 203527 129679
rect 203461 129646 203462 129678
rect 197880 128558 197886 128590
rect 197885 128526 197886 128558
rect 197950 128558 197956 128590
rect 203456 129614 203462 129646
rect 203526 129646 203527 129678
rect 203526 129614 203532 129646
rect 197950 128526 197951 128558
rect 197885 128525 197951 128526
rect 196661 128454 196727 128455
rect 196661 128422 196662 128454
rect 196520 126246 196526 126278
rect 191488 126208 191564 126214
rect 196525 126214 196526 126246
rect 196590 126246 196596 126278
rect 196656 128390 196662 128422
rect 196726 128422 196727 128454
rect 196726 128390 196732 128422
rect 196590 126214 196591 126246
rect 196525 126213 196591 126214
rect 194893 126142 194959 126143
rect 194893 126110 194894 126142
rect 190400 125974 190406 126006
rect 28288 125936 28364 125942
rect 190405 125942 190406 125974
rect 190470 125974 190476 126006
rect 194888 126078 194894 126110
rect 194958 126110 194959 126142
rect 195165 126142 195231 126143
rect 195165 126110 195166 126142
rect 194958 126078 194964 126110
rect 190470 125942 190471 125974
rect 190405 125941 190471 125942
rect 28293 125870 28359 125871
rect 28293 125838 28294 125870
rect 28288 125806 28294 125838
rect 28358 125838 28359 125870
rect 28358 125806 28364 125838
rect 21901 125598 21967 125599
rect 21901 125566 21902 125598
rect 21896 125534 21902 125566
rect 21966 125566 21967 125598
rect 22304 125598 22380 125604
rect 21966 125534 21972 125566
rect 21896 125326 21972 125534
rect 21896 125262 21902 125326
rect 21966 125262 21972 125326
rect 22304 125534 22310 125598
rect 22374 125534 22380 125598
rect 22304 125326 22380 125534
rect 22304 125294 22310 125326
rect 21896 125256 21972 125262
rect 22309 125262 22310 125294
rect 22374 125294 22380 125326
rect 22440 125598 22516 125604
rect 22440 125534 22446 125598
rect 22510 125534 22516 125598
rect 22440 125326 22516 125534
rect 28288 125462 28364 125806
rect 28565 125734 28631 125735
rect 28565 125702 28566 125734
rect 28288 125398 28294 125462
rect 28358 125398 28364 125462
rect 28288 125392 28364 125398
rect 28560 125670 28566 125702
rect 28630 125702 28631 125734
rect 190128 125734 190204 125740
rect 28630 125670 28636 125702
rect 28560 125462 28636 125670
rect 28560 125398 28566 125462
rect 28630 125398 28636 125462
rect 28560 125392 28636 125398
rect 190128 125670 190134 125734
rect 190198 125670 190204 125734
rect 22440 125294 22446 125326
rect 22374 125262 22375 125294
rect 22309 125261 22375 125262
rect 22445 125262 22446 125294
rect 22510 125294 22516 125326
rect 28424 125326 28500 125332
rect 22510 125262 22511 125294
rect 22445 125261 22511 125262
rect 28424 125262 28430 125326
rect 28494 125262 28500 125326
rect 190128 125326 190204 125670
rect 194888 125734 194964 126078
rect 194888 125670 194894 125734
rect 194958 125670 194964 125734
rect 194888 125664 194964 125670
rect 195160 126078 195166 126110
rect 195230 126110 195231 126142
rect 195230 126078 195236 126110
rect 195160 125734 195236 126078
rect 195160 125670 195166 125734
rect 195230 125670 195236 125734
rect 195160 125664 195236 125670
rect 196656 125734 196732 128390
rect 203456 126958 203532 129614
rect 203592 128454 203668 130974
rect 203592 128390 203598 128454
rect 203662 128390 203668 128454
rect 203592 128384 203668 128390
rect 217464 129950 217812 131518
rect 217464 129886 217470 129950
rect 217534 129886 217812 129950
rect 217464 128318 217812 129886
rect 217464 128254 217470 128318
rect 217534 128254 217812 128318
rect 216492 127909 216558 127910
rect 216492 127845 216493 127909
rect 216557 127845 216558 127909
rect 216492 127844 216558 127845
rect 203456 126894 203462 126958
rect 203526 126894 203532 126958
rect 203456 126888 203532 126894
rect 196656 125670 196662 125734
rect 196726 125670 196732 125734
rect 196656 125664 196732 125670
rect 196792 125598 196868 125604
rect 196792 125534 196798 125598
rect 196862 125534 196868 125598
rect 190128 125294 190134 125326
rect 952 124854 1230 124918
rect 1294 124854 1300 124918
rect 21760 125190 21836 125196
rect 21760 125126 21766 125190
rect 21830 125126 21836 125190
rect 21760 124918 21836 125126
rect 28424 125054 28500 125262
rect 190133 125262 190134 125294
rect 190198 125294 190204 125326
rect 190269 125326 190335 125327
rect 190269 125294 190270 125326
rect 190198 125262 190199 125294
rect 190133 125261 190199 125262
rect 190264 125262 190270 125294
rect 190334 125294 190335 125326
rect 196792 125326 196868 125534
rect 196792 125294 196798 125326
rect 190334 125262 190340 125294
rect 28424 125022 28430 125054
rect 28429 124990 28430 125022
rect 28494 125022 28500 125054
rect 190264 125054 190340 125262
rect 196797 125262 196798 125294
rect 196862 125294 196868 125326
rect 196862 125262 196863 125294
rect 196797 125261 196863 125262
rect 28494 124990 28495 125022
rect 28429 124989 28495 124990
rect 190264 124990 190270 125054
rect 190334 124990 190340 125054
rect 190264 124984 190340 124990
rect 196656 125190 196732 125196
rect 196656 125126 196662 125190
rect 196726 125126 196732 125190
rect 21760 124886 21766 124918
rect 952 123286 1300 124854
rect 21765 124854 21766 124886
rect 21830 124886 21836 124918
rect 196656 124918 196732 125126
rect 196656 124886 196662 124918
rect 21830 124854 21831 124886
rect 21765 124853 21831 124854
rect 196661 124854 196662 124886
rect 196726 124886 196732 124918
rect 196726 124854 196727 124886
rect 196661 124853 196727 124854
rect 21765 124782 21831 124783
rect 21765 124750 21766 124782
rect 21760 124718 21766 124750
rect 21830 124750 21831 124782
rect 22712 124782 22788 124788
rect 21830 124718 21836 124750
rect 21760 124510 21836 124718
rect 21760 124446 21766 124510
rect 21830 124446 21836 124510
rect 22712 124718 22718 124782
rect 22782 124718 22788 124782
rect 22712 124510 22788 124718
rect 22712 124478 22718 124510
rect 21760 124440 21836 124446
rect 22717 124446 22718 124478
rect 22782 124478 22788 124510
rect 22984 124782 23060 124788
rect 22984 124718 22990 124782
rect 23054 124718 23060 124782
rect 22984 124510 23060 124718
rect 22984 124478 22990 124510
rect 22782 124446 22783 124478
rect 22717 124445 22783 124446
rect 22989 124446 22990 124478
rect 23054 124478 23060 124510
rect 23392 124782 23468 124788
rect 23392 124718 23398 124782
rect 23462 124718 23468 124782
rect 195165 124782 195231 124783
rect 195165 124750 195166 124782
rect 23392 124510 23468 124718
rect 23392 124478 23398 124510
rect 23054 124446 23055 124478
rect 22989 124445 23055 124446
rect 23397 124446 23398 124478
rect 23462 124478 23468 124510
rect 195160 124718 195166 124750
rect 195230 124750 195231 124782
rect 195432 124782 195508 124788
rect 195230 124718 195236 124750
rect 195160 124510 195236 124718
rect 23462 124446 23463 124478
rect 23397 124445 23463 124446
rect 195160 124446 195166 124510
rect 195230 124446 195236 124510
rect 195432 124718 195438 124782
rect 195502 124718 195508 124782
rect 195432 124510 195508 124718
rect 195432 124478 195438 124510
rect 195160 124440 195236 124446
rect 195437 124446 195438 124478
rect 195502 124478 195508 124510
rect 195976 124782 196052 124788
rect 195976 124718 195982 124782
rect 196046 124718 196052 124782
rect 195976 124510 196052 124718
rect 195976 124478 195982 124510
rect 195502 124446 195503 124478
rect 195437 124445 195503 124446
rect 195981 124446 195982 124478
rect 196046 124478 196052 124510
rect 196112 124782 196188 124788
rect 196112 124718 196118 124782
rect 196182 124718 196188 124782
rect 196661 124782 196727 124783
rect 196661 124750 196662 124782
rect 196112 124510 196188 124718
rect 196112 124478 196118 124510
rect 196046 124446 196047 124478
rect 195981 124445 196047 124446
rect 196117 124446 196118 124478
rect 196182 124478 196188 124510
rect 196656 124718 196662 124750
rect 196726 124750 196727 124782
rect 196726 124718 196732 124750
rect 196656 124510 196732 124718
rect 196182 124446 196183 124478
rect 196117 124445 196183 124446
rect 196656 124446 196662 124510
rect 196726 124446 196732 124510
rect 196656 124440 196732 124446
rect 21896 124374 21972 124380
rect 21896 124310 21902 124374
rect 21966 124310 21972 124374
rect 22445 124374 22511 124375
rect 22445 124342 22446 124374
rect 21896 124102 21972 124310
rect 21896 124070 21902 124102
rect 21901 124038 21902 124070
rect 21966 124070 21972 124102
rect 22440 124310 22446 124342
rect 22510 124342 22511 124374
rect 23120 124374 23196 124380
rect 22510 124310 22516 124342
rect 22440 124102 22516 124310
rect 21966 124038 21967 124070
rect 21901 124037 21967 124038
rect 22440 124038 22446 124102
rect 22510 124038 22516 124102
rect 23120 124310 23126 124374
rect 23190 124310 23196 124374
rect 23397 124374 23463 124375
rect 23397 124342 23398 124374
rect 23120 124102 23196 124310
rect 23120 124070 23126 124102
rect 22440 124032 22516 124038
rect 23125 124038 23126 124070
rect 23190 124070 23196 124102
rect 23392 124310 23398 124342
rect 23462 124342 23463 124374
rect 195024 124374 195100 124380
rect 23462 124310 23468 124342
rect 23392 124102 23468 124310
rect 23190 124038 23191 124070
rect 23125 124037 23191 124038
rect 23392 124038 23398 124102
rect 23462 124038 23468 124102
rect 195024 124310 195030 124374
rect 195094 124310 195100 124374
rect 195024 124102 195100 124310
rect 195024 124070 195030 124102
rect 23392 124032 23468 124038
rect 195029 124038 195030 124070
rect 195094 124070 195100 124102
rect 195568 124374 195644 124380
rect 195568 124310 195574 124374
rect 195638 124310 195644 124374
rect 195981 124374 196047 124375
rect 195981 124342 195982 124374
rect 195568 124102 195644 124310
rect 195568 124070 195574 124102
rect 195094 124038 195095 124070
rect 195029 124037 195095 124038
rect 195573 124038 195574 124070
rect 195638 124070 195644 124102
rect 195976 124310 195982 124342
rect 196046 124342 196047 124374
rect 196117 124374 196183 124375
rect 196117 124342 196118 124374
rect 196046 124310 196052 124342
rect 195976 124102 196052 124310
rect 195638 124038 195639 124070
rect 195573 124037 195639 124038
rect 195976 124038 195982 124102
rect 196046 124038 196052 124102
rect 195976 124032 196052 124038
rect 196112 124310 196118 124342
rect 196182 124342 196183 124374
rect 196792 124374 196868 124380
rect 196182 124310 196188 124342
rect 196112 124102 196188 124310
rect 196112 124038 196118 124102
rect 196182 124038 196188 124102
rect 196792 124310 196798 124374
rect 196862 124310 196868 124374
rect 196792 124102 196868 124310
rect 196792 124070 196798 124102
rect 196112 124032 196188 124038
rect 196797 124038 196798 124070
rect 196862 124070 196868 124102
rect 196862 124038 196863 124070
rect 196797 124037 196863 124038
rect 21765 123966 21831 123967
rect 21765 123934 21766 123966
rect 21760 123902 21766 123934
rect 21830 123934 21831 123966
rect 22168 123966 22244 123972
rect 21830 123902 21836 123934
rect 21760 123694 21836 123902
rect 21760 123630 21766 123694
rect 21830 123630 21836 123694
rect 22168 123902 22174 123966
rect 22238 123902 22244 123966
rect 22168 123694 22244 123902
rect 22168 123662 22174 123694
rect 21760 123624 21836 123630
rect 22173 123630 22174 123662
rect 22238 123662 22244 123694
rect 22576 123966 22652 123972
rect 22576 123902 22582 123966
rect 22646 123902 22652 123966
rect 22989 123966 23055 123967
rect 22989 123934 22990 123966
rect 22576 123694 22652 123902
rect 22576 123662 22582 123694
rect 22238 123630 22239 123662
rect 22173 123629 22239 123630
rect 22581 123630 22582 123662
rect 22646 123662 22652 123694
rect 22984 123902 22990 123934
rect 23054 123934 23055 123966
rect 23533 123966 23599 123967
rect 23533 123934 23534 123966
rect 23054 123902 23060 123934
rect 22984 123694 23060 123902
rect 22646 123630 22647 123662
rect 22581 123629 22647 123630
rect 22984 123630 22990 123694
rect 23054 123630 23060 123694
rect 22984 123624 23060 123630
rect 23528 123902 23534 123934
rect 23598 123934 23599 123966
rect 195165 123966 195231 123967
rect 195165 123934 195166 123966
rect 23598 123902 23604 123934
rect 23528 123694 23604 123902
rect 23528 123630 23534 123694
rect 23598 123630 23604 123694
rect 23528 123624 23604 123630
rect 195160 123902 195166 123934
rect 195230 123934 195231 123966
rect 195437 123966 195503 123967
rect 195437 123934 195438 123966
rect 195230 123902 195236 123934
rect 195160 123694 195236 123902
rect 195160 123630 195166 123694
rect 195230 123630 195236 123694
rect 195160 123624 195236 123630
rect 195432 123902 195438 123934
rect 195502 123934 195503 123966
rect 196248 123966 196324 123972
rect 195502 123902 195508 123934
rect 195432 123694 195508 123902
rect 195432 123630 195438 123694
rect 195502 123630 195508 123694
rect 196248 123902 196254 123966
rect 196318 123902 196324 123966
rect 196661 123966 196727 123967
rect 196661 123934 196662 123966
rect 196248 123694 196324 123902
rect 196248 123662 196254 123694
rect 195432 123624 195508 123630
rect 196253 123630 196254 123662
rect 196318 123662 196324 123694
rect 196656 123902 196662 123934
rect 196726 123934 196727 123966
rect 196726 123902 196732 123934
rect 196656 123694 196732 123902
rect 196318 123630 196319 123662
rect 196253 123629 196319 123630
rect 196656 123630 196662 123694
rect 196726 123630 196732 123694
rect 196656 123624 196732 123630
rect 21765 123558 21831 123559
rect 21765 123526 21766 123558
rect 952 123222 1230 123286
rect 1294 123222 1300 123286
rect 952 121382 1300 123222
rect 21760 123494 21766 123526
rect 21830 123526 21831 123558
rect 22440 123558 22516 123564
rect 21830 123494 21836 123526
rect 21760 123286 21836 123494
rect 21760 123222 21766 123286
rect 21830 123222 21836 123286
rect 22440 123494 22446 123558
rect 22510 123494 22516 123558
rect 22581 123558 22647 123559
rect 22581 123526 22582 123558
rect 22440 123286 22516 123494
rect 22440 123254 22446 123286
rect 21760 123216 21836 123222
rect 22445 123222 22446 123254
rect 22510 123254 22516 123286
rect 22576 123494 22582 123526
rect 22646 123526 22647 123558
rect 23125 123558 23191 123559
rect 23125 123526 23126 123558
rect 22646 123494 22652 123526
rect 22576 123286 22652 123494
rect 22510 123222 22511 123254
rect 22445 123221 22511 123222
rect 22576 123222 22582 123286
rect 22646 123222 22652 123286
rect 22576 123216 22652 123222
rect 23120 123494 23126 123526
rect 23190 123526 23191 123558
rect 23533 123558 23599 123559
rect 23533 123526 23534 123558
rect 23190 123494 23196 123526
rect 23120 123286 23196 123494
rect 23120 123222 23126 123286
rect 23190 123222 23196 123286
rect 23120 123216 23196 123222
rect 23528 123494 23534 123526
rect 23598 123526 23599 123558
rect 195165 123558 195231 123559
rect 195165 123526 195166 123558
rect 23598 123494 23604 123526
rect 23528 123286 23604 123494
rect 23528 123222 23534 123286
rect 23598 123222 23604 123286
rect 23528 123216 23604 123222
rect 195160 123494 195166 123526
rect 195230 123526 195231 123558
rect 195573 123558 195639 123559
rect 195573 123526 195574 123558
rect 195230 123494 195236 123526
rect 195160 123286 195236 123494
rect 195160 123222 195166 123286
rect 195230 123222 195236 123286
rect 195160 123216 195236 123222
rect 195568 123494 195574 123526
rect 195638 123526 195639 123558
rect 195976 123558 196052 123564
rect 195638 123494 195644 123526
rect 195568 123286 195644 123494
rect 195568 123222 195574 123286
rect 195638 123222 195644 123286
rect 195976 123494 195982 123558
rect 196046 123494 196052 123558
rect 195976 123286 196052 123494
rect 195976 123254 195982 123286
rect 195568 123216 195644 123222
rect 195981 123222 195982 123254
rect 196046 123254 196052 123286
rect 196112 123558 196188 123564
rect 196112 123494 196118 123558
rect 196182 123494 196188 123558
rect 196112 123286 196188 123494
rect 196112 123254 196118 123286
rect 196046 123222 196047 123254
rect 195981 123221 196047 123222
rect 196117 123222 196118 123254
rect 196182 123254 196188 123286
rect 196792 123558 196868 123564
rect 196792 123494 196798 123558
rect 196862 123494 196868 123558
rect 196792 123286 196868 123494
rect 196792 123254 196798 123286
rect 196182 123222 196183 123254
rect 196117 123221 196183 123222
rect 196797 123222 196798 123254
rect 196862 123254 196868 123286
rect 196862 123222 196863 123254
rect 196797 123221 196863 123222
rect 22309 123150 22375 123151
rect 22309 123118 22310 123150
rect 22304 123086 22310 123118
rect 22374 123118 22375 123150
rect 22445 123150 22511 123151
rect 22445 123118 22446 123150
rect 22374 123086 22380 123118
rect 22304 122878 22380 123086
rect 22304 122814 22310 122878
rect 22374 122814 22380 122878
rect 22304 122808 22380 122814
rect 22440 123086 22446 123118
rect 22510 123118 22511 123150
rect 22984 123150 23060 123156
rect 22510 123086 22516 123118
rect 22440 122878 22516 123086
rect 22440 122814 22446 122878
rect 22510 122814 22516 122878
rect 22984 123086 22990 123150
rect 23054 123086 23060 123150
rect 23397 123150 23463 123151
rect 23397 123118 23398 123150
rect 22984 122878 23060 123086
rect 22984 122846 22990 122878
rect 22440 122808 22516 122814
rect 22989 122814 22990 122846
rect 23054 122846 23060 122878
rect 23392 123086 23398 123118
rect 23462 123118 23463 123150
rect 195160 123150 195236 123156
rect 23462 123086 23468 123118
rect 23392 122878 23468 123086
rect 23054 122814 23055 122846
rect 22989 122813 23055 122814
rect 23392 122814 23398 122878
rect 23462 122814 23468 122878
rect 195160 123086 195166 123150
rect 195230 123086 195236 123150
rect 195160 122878 195236 123086
rect 195160 122846 195166 122878
rect 23392 122808 23468 122814
rect 195165 122814 195166 122846
rect 195230 122846 195236 122878
rect 195432 123150 195508 123156
rect 195432 123086 195438 123150
rect 195502 123086 195508 123150
rect 195432 122878 195508 123086
rect 195432 122846 195438 122878
rect 195230 122814 195231 122846
rect 195165 122813 195231 122814
rect 195437 122814 195438 122846
rect 195502 122846 195508 122878
rect 196248 123150 196324 123156
rect 196248 123086 196254 123150
rect 196318 123086 196324 123150
rect 196248 122878 196324 123086
rect 196248 122846 196254 122878
rect 195502 122814 195503 122846
rect 195437 122813 195503 122814
rect 196253 122814 196254 122846
rect 196318 122846 196324 122878
rect 196318 122814 196319 122846
rect 196253 122813 196319 122814
rect 21760 122742 21836 122748
rect 21760 122678 21766 122742
rect 21830 122678 21836 122742
rect 21760 122470 21836 122678
rect 21760 122438 21766 122470
rect 21765 122406 21766 122438
rect 21830 122438 21836 122470
rect 22304 122742 22380 122748
rect 22304 122678 22310 122742
rect 22374 122678 22380 122742
rect 22304 122470 22380 122678
rect 22304 122438 22310 122470
rect 21830 122406 21831 122438
rect 21765 122405 21831 122406
rect 22309 122406 22310 122438
rect 22374 122438 22380 122470
rect 22576 122742 22652 122748
rect 22576 122678 22582 122742
rect 22646 122678 22652 122742
rect 22989 122742 23055 122743
rect 22989 122710 22990 122742
rect 22576 122470 22652 122678
rect 22576 122438 22582 122470
rect 22374 122406 22375 122438
rect 22309 122405 22375 122406
rect 22581 122406 22582 122438
rect 22646 122438 22652 122470
rect 22984 122678 22990 122710
rect 23054 122710 23055 122742
rect 23528 122742 23604 122748
rect 23054 122678 23060 122710
rect 22984 122470 23060 122678
rect 22646 122406 22647 122438
rect 22581 122405 22647 122406
rect 22984 122406 22990 122470
rect 23054 122406 23060 122470
rect 23528 122678 23534 122742
rect 23598 122678 23604 122742
rect 23528 122470 23604 122678
rect 23528 122438 23534 122470
rect 22984 122400 23060 122406
rect 23533 122406 23534 122438
rect 23598 122438 23604 122470
rect 195160 122742 195236 122748
rect 195160 122678 195166 122742
rect 195230 122678 195236 122742
rect 195160 122470 195236 122678
rect 195160 122438 195166 122470
rect 23598 122406 23599 122438
rect 23533 122405 23599 122406
rect 195165 122406 195166 122438
rect 195230 122438 195236 122470
rect 195568 122742 195644 122748
rect 195568 122678 195574 122742
rect 195638 122678 195644 122742
rect 195845 122742 195911 122743
rect 195845 122710 195846 122742
rect 195568 122470 195644 122678
rect 195568 122438 195574 122470
rect 195230 122406 195231 122438
rect 195165 122405 195231 122406
rect 195573 122406 195574 122438
rect 195638 122438 195644 122470
rect 195840 122678 195846 122710
rect 195910 122710 195911 122742
rect 196656 122742 196732 122748
rect 195910 122678 195916 122710
rect 195840 122470 195916 122678
rect 195638 122406 195639 122438
rect 195573 122405 195639 122406
rect 195840 122406 195846 122470
rect 195910 122406 195916 122470
rect 196656 122678 196662 122742
rect 196726 122678 196732 122742
rect 196656 122470 196732 122678
rect 196656 122438 196662 122470
rect 195840 122400 195916 122406
rect 196661 122406 196662 122438
rect 196726 122438 196732 122470
rect 196726 122406 196727 122438
rect 196661 122405 196727 122406
rect 22717 122334 22783 122335
rect 22717 122302 22718 122334
rect 22712 122270 22718 122302
rect 22782 122302 22783 122334
rect 23120 122334 23196 122340
rect 22782 122270 22788 122302
rect 21760 122062 21836 122068
rect 21760 121998 21766 122062
rect 21830 121998 21836 122062
rect 22445 122062 22511 122063
rect 22445 122030 22446 122062
rect 21760 121790 21836 121998
rect 21760 121758 21766 121790
rect 21765 121726 21766 121758
rect 21830 121758 21836 121790
rect 22440 121998 22446 122030
rect 22510 122030 22511 122062
rect 22712 122062 22788 122270
rect 22510 121998 22516 122030
rect 22440 121790 22516 121998
rect 22712 121998 22718 122062
rect 22782 121998 22788 122062
rect 23120 122270 23126 122334
rect 23190 122270 23196 122334
rect 23397 122334 23463 122335
rect 23397 122302 23398 122334
rect 23120 122062 23196 122270
rect 23120 122030 23126 122062
rect 22712 121992 22788 121998
rect 23125 121998 23126 122030
rect 23190 122030 23196 122062
rect 23392 122270 23398 122302
rect 23462 122302 23463 122334
rect 195029 122334 195095 122335
rect 195029 122302 195030 122334
rect 23462 122270 23468 122302
rect 23392 122062 23468 122270
rect 23190 121998 23191 122030
rect 23125 121997 23191 121998
rect 23392 121998 23398 122062
rect 23462 121998 23468 122062
rect 23392 121992 23468 121998
rect 195024 122270 195030 122302
rect 195094 122302 195095 122334
rect 195437 122334 195503 122335
rect 195437 122302 195438 122334
rect 195094 122270 195100 122302
rect 195024 122062 195100 122270
rect 195024 121998 195030 122062
rect 195094 121998 195100 122062
rect 195024 121992 195100 121998
rect 195432 122270 195438 122302
rect 195502 122302 195503 122334
rect 196112 122334 196188 122340
rect 195502 122270 195508 122302
rect 195432 122062 195508 122270
rect 195432 121998 195438 122062
rect 195502 121998 195508 122062
rect 196112 122270 196118 122334
rect 196182 122270 196188 122334
rect 196112 122062 196188 122270
rect 196112 122030 196118 122062
rect 195432 121992 195508 121998
rect 196117 121998 196118 122030
rect 196182 122030 196188 122062
rect 196797 122062 196863 122063
rect 196797 122030 196798 122062
rect 196182 121998 196183 122030
rect 196117 121997 196183 121998
rect 196792 121998 196798 122030
rect 196862 122030 196863 122062
rect 196862 121998 196868 122030
rect 21830 121726 21831 121758
rect 21765 121725 21831 121726
rect 22440 121726 22446 121790
rect 22510 121726 22516 121790
rect 22440 121720 22516 121726
rect 28288 121790 28364 121796
rect 28288 121726 28294 121790
rect 28358 121726 28364 121790
rect 190133 121790 190199 121791
rect 190133 121758 190134 121790
rect 952 121318 1230 121382
rect 1294 121318 1300 121382
rect 21760 121654 21836 121660
rect 21760 121590 21766 121654
rect 21830 121590 21836 121654
rect 22173 121654 22239 121655
rect 22173 121622 22174 121654
rect 21760 121382 21836 121590
rect 21760 121350 21766 121382
rect 952 119750 1300 121318
rect 21765 121318 21766 121350
rect 21830 121350 21836 121382
rect 22168 121590 22174 121622
rect 22238 121622 22239 121654
rect 22238 121590 22244 121622
rect 22168 121382 22244 121590
rect 28288 121518 28364 121726
rect 28288 121486 28294 121518
rect 28293 121454 28294 121486
rect 28358 121486 28364 121518
rect 190128 121726 190134 121758
rect 190198 121758 190199 121790
rect 196792 121790 196868 121998
rect 190198 121726 190204 121758
rect 190128 121518 190204 121726
rect 196792 121726 196798 121790
rect 196862 121726 196868 121790
rect 196792 121720 196868 121726
rect 196117 121654 196183 121655
rect 196117 121622 196118 121654
rect 28358 121454 28359 121486
rect 28293 121453 28359 121454
rect 190128 121454 190134 121518
rect 190198 121454 190204 121518
rect 190128 121448 190204 121454
rect 196112 121590 196118 121622
rect 196182 121622 196183 121654
rect 196656 121654 196732 121660
rect 196182 121590 196188 121622
rect 21830 121318 21831 121350
rect 21765 121317 21831 121318
rect 22168 121318 22174 121382
rect 22238 121318 22244 121382
rect 28293 121382 28359 121383
rect 28293 121350 28294 121382
rect 22168 121312 22244 121318
rect 28288 121318 28294 121350
rect 28358 121350 28359 121382
rect 190264 121382 190340 121388
rect 28358 121318 28364 121350
rect 21901 121246 21967 121247
rect 21901 121214 21902 121246
rect 21896 121182 21902 121214
rect 21966 121214 21967 121246
rect 21966 121182 21972 121214
rect 21896 120974 21972 121182
rect 28288 121110 28364 121318
rect 28288 121046 28294 121110
rect 28358 121046 28364 121110
rect 190264 121318 190270 121382
rect 190334 121318 190340 121382
rect 190264 121110 190340 121318
rect 196112 121382 196188 121590
rect 196112 121318 196118 121382
rect 196182 121318 196188 121382
rect 196656 121590 196662 121654
rect 196726 121590 196732 121654
rect 196656 121382 196732 121590
rect 196656 121350 196662 121382
rect 196112 121312 196188 121318
rect 196661 121318 196662 121350
rect 196726 121350 196732 121382
rect 196726 121318 196727 121350
rect 196661 121317 196727 121318
rect 196797 121246 196863 121247
rect 196797 121214 196798 121246
rect 190264 121078 190270 121110
rect 28288 121040 28364 121046
rect 190269 121046 190270 121078
rect 190334 121078 190340 121110
rect 196792 121182 196798 121214
rect 196862 121214 196863 121246
rect 196862 121182 196868 121214
rect 190334 121046 190335 121078
rect 190269 121045 190335 121046
rect 21896 120910 21902 120974
rect 21966 120910 21972 120974
rect 28429 120974 28495 120975
rect 28429 120942 28430 120974
rect 21896 120904 21972 120910
rect 28424 120910 28430 120942
rect 28494 120942 28495 120974
rect 190269 120974 190335 120975
rect 190269 120942 190270 120974
rect 28494 120910 28500 120942
rect 21760 120838 21836 120844
rect 21760 120774 21766 120838
rect 21830 120774 21836 120838
rect 22445 120838 22511 120839
rect 22445 120806 22446 120838
rect 21760 120566 21836 120774
rect 21760 120534 21766 120566
rect 21765 120502 21766 120534
rect 21830 120534 21836 120566
rect 22440 120774 22446 120806
rect 22510 120806 22511 120838
rect 23125 120838 23191 120839
rect 23125 120806 23126 120838
rect 22510 120774 22516 120806
rect 22440 120566 22516 120774
rect 21830 120502 21831 120534
rect 21765 120501 21831 120502
rect 22440 120502 22446 120566
rect 22510 120502 22516 120566
rect 22440 120496 22516 120502
rect 23120 120774 23126 120806
rect 23190 120806 23191 120838
rect 23397 120838 23463 120839
rect 23397 120806 23398 120838
rect 23190 120774 23196 120806
rect 23120 120566 23196 120774
rect 23120 120502 23126 120566
rect 23190 120502 23196 120566
rect 23120 120496 23196 120502
rect 23392 120774 23398 120806
rect 23462 120806 23463 120838
rect 23462 120774 23468 120806
rect 23392 120566 23468 120774
rect 23392 120502 23398 120566
rect 23462 120502 23468 120566
rect 28293 120566 28359 120567
rect 28293 120534 28294 120566
rect 23392 120496 23468 120502
rect 28288 120502 28294 120534
rect 28358 120534 28359 120566
rect 28424 120566 28500 120910
rect 190264 120910 190270 120942
rect 190334 120942 190335 120974
rect 196792 120974 196868 121182
rect 190334 120910 190340 120942
rect 28358 120502 28364 120534
rect 21765 120430 21831 120431
rect 21765 120398 21766 120430
rect 21760 120366 21766 120398
rect 21830 120398 21831 120430
rect 22173 120430 22239 120431
rect 22173 120398 22174 120430
rect 21830 120366 21836 120398
rect 21760 120158 21836 120366
rect 21760 120094 21766 120158
rect 21830 120094 21836 120158
rect 21760 120088 21836 120094
rect 22168 120366 22174 120398
rect 22238 120398 22239 120430
rect 22712 120430 22788 120436
rect 22238 120366 22244 120398
rect 22168 120158 22244 120366
rect 22168 120094 22174 120158
rect 22238 120094 22244 120158
rect 22712 120366 22718 120430
rect 22782 120366 22788 120430
rect 23125 120430 23191 120431
rect 23125 120398 23126 120430
rect 22712 120158 22788 120366
rect 22712 120126 22718 120158
rect 22168 120088 22244 120094
rect 22717 120094 22718 120126
rect 22782 120126 22788 120158
rect 23120 120366 23126 120398
rect 23190 120398 23191 120430
rect 23392 120430 23468 120436
rect 23190 120366 23196 120398
rect 23120 120158 23196 120366
rect 22782 120094 22783 120126
rect 22717 120093 22783 120094
rect 23120 120094 23126 120158
rect 23190 120094 23196 120158
rect 23392 120366 23398 120430
rect 23462 120366 23468 120430
rect 23392 120158 23468 120366
rect 28288 120294 28364 120502
rect 28424 120502 28430 120566
rect 28494 120502 28500 120566
rect 190133 120566 190199 120567
rect 190133 120534 190134 120566
rect 28424 120496 28500 120502
rect 190128 120502 190134 120534
rect 190198 120534 190199 120566
rect 190264 120566 190340 120910
rect 196792 120910 196798 120974
rect 196862 120910 196868 120974
rect 196792 120904 196868 120910
rect 190198 120502 190204 120534
rect 28288 120230 28294 120294
rect 28358 120230 28364 120294
rect 28288 120224 28364 120230
rect 190128 120294 190204 120502
rect 190264 120502 190270 120566
rect 190334 120502 190340 120566
rect 195160 120838 195236 120844
rect 195160 120774 195166 120838
rect 195230 120774 195236 120838
rect 195160 120566 195236 120774
rect 195160 120534 195166 120566
rect 190264 120496 190340 120502
rect 195165 120502 195166 120534
rect 195230 120534 195236 120566
rect 195432 120838 195508 120844
rect 195432 120774 195438 120838
rect 195502 120774 195508 120838
rect 195432 120566 195508 120774
rect 195432 120534 195438 120566
rect 195230 120502 195231 120534
rect 195165 120501 195231 120502
rect 195437 120502 195438 120534
rect 195502 120534 195508 120566
rect 195840 120838 195916 120844
rect 195840 120774 195846 120838
rect 195910 120774 195916 120838
rect 195840 120566 195916 120774
rect 195840 120534 195846 120566
rect 195502 120502 195503 120534
rect 195437 120501 195503 120502
rect 195845 120502 195846 120534
rect 195910 120534 195916 120566
rect 196656 120838 196732 120844
rect 196656 120774 196662 120838
rect 196726 120774 196732 120838
rect 196656 120566 196732 120774
rect 196656 120534 196662 120566
rect 195910 120502 195911 120534
rect 195845 120501 195911 120502
rect 196661 120502 196662 120534
rect 196726 120534 196732 120566
rect 196726 120502 196727 120534
rect 196661 120501 196727 120502
rect 195165 120430 195231 120431
rect 195165 120398 195166 120430
rect 190128 120230 190134 120294
rect 190198 120230 190204 120294
rect 190128 120224 190204 120230
rect 195160 120366 195166 120398
rect 195230 120398 195231 120430
rect 195573 120430 195639 120431
rect 195573 120398 195574 120430
rect 195230 120366 195236 120398
rect 23392 120126 23398 120158
rect 23120 120088 23196 120094
rect 23397 120094 23398 120126
rect 23462 120126 23468 120158
rect 195160 120158 195236 120366
rect 23462 120094 23463 120126
rect 23397 120093 23463 120094
rect 195160 120094 195166 120158
rect 195230 120094 195236 120158
rect 195160 120088 195236 120094
rect 195568 120366 195574 120398
rect 195638 120398 195639 120430
rect 195976 120430 196052 120436
rect 195638 120366 195644 120398
rect 195568 120158 195644 120366
rect 195568 120094 195574 120158
rect 195638 120094 195644 120158
rect 195976 120366 195982 120430
rect 196046 120366 196052 120430
rect 195976 120158 196052 120366
rect 195976 120126 195982 120158
rect 195568 120088 195644 120094
rect 195981 120094 195982 120126
rect 196046 120126 196052 120158
rect 196792 120430 196868 120436
rect 196792 120366 196798 120430
rect 196862 120366 196868 120430
rect 196792 120158 196868 120366
rect 196792 120126 196798 120158
rect 196046 120094 196047 120126
rect 195981 120093 196047 120094
rect 196797 120094 196798 120126
rect 196862 120126 196868 120158
rect 196862 120094 196863 120126
rect 196797 120093 196863 120094
rect 21901 120022 21967 120023
rect 21901 119990 21902 120022
rect 952 119686 1230 119750
rect 1294 119686 1300 119750
rect 952 118118 1300 119686
rect 21896 119958 21902 119990
rect 21966 119990 21967 120022
rect 22309 120022 22375 120023
rect 22309 119990 22310 120022
rect 21966 119958 21972 119990
rect 21896 119750 21972 119958
rect 21896 119686 21902 119750
rect 21966 119686 21972 119750
rect 21896 119680 21972 119686
rect 22304 119958 22310 119990
rect 22374 119990 22375 120022
rect 23120 120022 23196 120028
rect 22374 119958 22380 119990
rect 22304 119750 22380 119958
rect 22304 119686 22310 119750
rect 22374 119686 22380 119750
rect 23120 119958 23126 120022
rect 23190 119958 23196 120022
rect 23397 120022 23463 120023
rect 23397 119990 23398 120022
rect 23120 119750 23196 119958
rect 23120 119718 23126 119750
rect 22304 119680 22380 119686
rect 23125 119686 23126 119718
rect 23190 119718 23196 119750
rect 23392 119958 23398 119990
rect 23462 119990 23463 120022
rect 195029 120022 195095 120023
rect 195029 119990 195030 120022
rect 23462 119958 23468 119990
rect 23392 119750 23468 119958
rect 23190 119686 23191 119718
rect 23125 119685 23191 119686
rect 23392 119686 23398 119750
rect 23462 119686 23468 119750
rect 23392 119680 23468 119686
rect 195024 119958 195030 119990
rect 195094 119990 195095 120022
rect 195568 120022 195644 120028
rect 195094 119958 195100 119990
rect 195024 119750 195100 119958
rect 195024 119686 195030 119750
rect 195094 119686 195100 119750
rect 195568 119958 195574 120022
rect 195638 119958 195644 120022
rect 195568 119750 195644 119958
rect 195568 119718 195574 119750
rect 195024 119680 195100 119686
rect 195573 119686 195574 119718
rect 195638 119718 195644 119750
rect 195976 120022 196052 120028
rect 195976 119958 195982 120022
rect 196046 119958 196052 120022
rect 196797 120022 196863 120023
rect 196797 119990 196798 120022
rect 195976 119750 196052 119958
rect 195976 119718 195982 119750
rect 195638 119686 195639 119718
rect 195573 119685 195639 119686
rect 195981 119686 195982 119718
rect 196046 119718 196052 119750
rect 196792 119958 196798 119990
rect 196862 119990 196863 120022
rect 196862 119958 196868 119990
rect 196792 119750 196868 119958
rect 196046 119686 196047 119718
rect 195981 119685 196047 119686
rect 196792 119686 196798 119750
rect 196862 119686 196868 119750
rect 196792 119680 196868 119686
rect 21760 119614 21836 119620
rect 21760 119550 21766 119614
rect 21830 119550 21836 119614
rect 22445 119614 22511 119615
rect 22445 119582 22446 119614
rect 21760 119342 21836 119550
rect 21760 119310 21766 119342
rect 21765 119278 21766 119310
rect 21830 119310 21836 119342
rect 22440 119550 22446 119582
rect 22510 119582 22511 119614
rect 23120 119614 23196 119620
rect 22510 119550 22516 119582
rect 22440 119342 22516 119550
rect 21830 119278 21831 119310
rect 21765 119277 21831 119278
rect 22440 119278 22446 119342
rect 22510 119278 22516 119342
rect 23120 119550 23126 119614
rect 23190 119550 23196 119614
rect 23120 119342 23196 119550
rect 23120 119310 23126 119342
rect 22440 119272 22516 119278
rect 23125 119278 23126 119310
rect 23190 119310 23196 119342
rect 23528 119614 23604 119620
rect 23528 119550 23534 119614
rect 23598 119550 23604 119614
rect 23528 119342 23604 119550
rect 23528 119310 23534 119342
rect 23190 119278 23191 119310
rect 23125 119277 23191 119278
rect 23533 119278 23534 119310
rect 23598 119310 23604 119342
rect 195160 119614 195236 119620
rect 195160 119550 195166 119614
rect 195230 119550 195236 119614
rect 195437 119614 195503 119615
rect 195437 119582 195438 119614
rect 195160 119342 195236 119550
rect 195160 119310 195166 119342
rect 23598 119278 23599 119310
rect 23533 119277 23599 119278
rect 195165 119278 195166 119310
rect 195230 119310 195236 119342
rect 195432 119550 195438 119582
rect 195502 119582 195503 119614
rect 195845 119614 195911 119615
rect 195845 119582 195846 119614
rect 195502 119550 195508 119582
rect 195432 119342 195508 119550
rect 195230 119278 195231 119310
rect 195165 119277 195231 119278
rect 195432 119278 195438 119342
rect 195502 119278 195508 119342
rect 195432 119272 195508 119278
rect 195840 119550 195846 119582
rect 195910 119582 195911 119614
rect 196248 119614 196324 119620
rect 195910 119550 195916 119582
rect 195840 119342 195916 119550
rect 195840 119278 195846 119342
rect 195910 119278 195916 119342
rect 196248 119550 196254 119614
rect 196318 119550 196324 119614
rect 196248 119342 196324 119550
rect 196248 119310 196254 119342
rect 195840 119272 195916 119278
rect 196253 119278 196254 119310
rect 196318 119310 196324 119342
rect 196656 119614 196732 119620
rect 196656 119550 196662 119614
rect 196726 119550 196732 119614
rect 196656 119342 196732 119550
rect 196656 119310 196662 119342
rect 196318 119278 196319 119310
rect 196253 119277 196319 119278
rect 196661 119278 196662 119310
rect 196726 119310 196732 119342
rect 196726 119278 196727 119310
rect 196661 119277 196727 119278
rect 22304 119206 22380 119212
rect 22304 119142 22310 119206
rect 22374 119142 22380 119206
rect 23125 119206 23191 119207
rect 23125 119174 23126 119206
rect 22304 118934 22380 119142
rect 22304 118902 22310 118934
rect 22309 118870 22310 118902
rect 22374 118902 22380 118934
rect 23120 119142 23126 119174
rect 23190 119174 23191 119206
rect 23533 119206 23599 119207
rect 23533 119174 23534 119206
rect 23190 119142 23196 119174
rect 23120 118934 23196 119142
rect 22374 118870 22375 118902
rect 22309 118869 22375 118870
rect 23120 118870 23126 118934
rect 23190 118870 23196 118934
rect 23120 118864 23196 118870
rect 23528 119142 23534 119174
rect 23598 119174 23599 119206
rect 195024 119206 195100 119212
rect 23598 119142 23604 119174
rect 23528 118934 23604 119142
rect 23528 118870 23534 118934
rect 23598 118870 23604 118934
rect 195024 119142 195030 119206
rect 195094 119142 195100 119206
rect 195024 118934 195100 119142
rect 195024 118902 195030 118934
rect 23528 118864 23604 118870
rect 195029 118870 195030 118902
rect 195094 118902 195100 118934
rect 195432 119206 195508 119212
rect 195432 119142 195438 119206
rect 195502 119142 195508 119206
rect 195845 119206 195911 119207
rect 195845 119174 195846 119206
rect 195432 118934 195508 119142
rect 195432 118902 195438 118934
rect 195094 118870 195095 118902
rect 195029 118869 195095 118870
rect 195437 118870 195438 118902
rect 195502 118902 195508 118934
rect 195840 119142 195846 119174
rect 195910 119174 195911 119206
rect 196112 119206 196188 119212
rect 195910 119142 195916 119174
rect 195840 118934 195916 119142
rect 195502 118870 195503 118902
rect 195437 118869 195503 118870
rect 195840 118870 195846 118934
rect 195910 118870 195916 118934
rect 196112 119142 196118 119206
rect 196182 119142 196188 119206
rect 196112 118934 196188 119142
rect 196112 118902 196118 118934
rect 195840 118864 195916 118870
rect 196117 118870 196118 118902
rect 196182 118902 196188 118934
rect 196182 118870 196183 118902
rect 196117 118869 196183 118870
rect 21901 118798 21967 118799
rect 21901 118766 21902 118798
rect 21896 118734 21902 118766
rect 21966 118766 21967 118798
rect 22717 118798 22783 118799
rect 22717 118766 22718 118798
rect 21966 118734 21972 118766
rect 21896 118526 21972 118734
rect 21896 118462 21902 118526
rect 21966 118462 21972 118526
rect 21896 118456 21972 118462
rect 22712 118734 22718 118766
rect 22782 118766 22783 118798
rect 22984 118798 23060 118804
rect 22782 118734 22788 118766
rect 22712 118526 22788 118734
rect 22712 118462 22718 118526
rect 22782 118462 22788 118526
rect 22984 118734 22990 118798
rect 23054 118734 23060 118798
rect 23397 118798 23463 118799
rect 23397 118766 23398 118798
rect 22984 118526 23060 118734
rect 22984 118494 22990 118526
rect 22712 118456 22788 118462
rect 22989 118462 22990 118494
rect 23054 118494 23060 118526
rect 23392 118734 23398 118766
rect 23462 118766 23463 118798
rect 195029 118798 195095 118799
rect 195029 118766 195030 118798
rect 23462 118734 23468 118766
rect 23392 118526 23468 118734
rect 23054 118462 23055 118494
rect 22989 118461 23055 118462
rect 23392 118462 23398 118526
rect 23462 118462 23468 118526
rect 23392 118456 23468 118462
rect 195024 118734 195030 118766
rect 195094 118766 195095 118798
rect 195432 118798 195508 118804
rect 195094 118734 195100 118766
rect 195024 118526 195100 118734
rect 195024 118462 195030 118526
rect 195094 118462 195100 118526
rect 195432 118734 195438 118798
rect 195502 118734 195508 118798
rect 195432 118526 195508 118734
rect 195432 118494 195438 118526
rect 195024 118456 195100 118462
rect 195437 118462 195438 118494
rect 195502 118494 195508 118526
rect 195840 118798 195916 118804
rect 195840 118734 195846 118798
rect 195910 118734 195916 118798
rect 196797 118798 196863 118799
rect 196797 118766 196798 118798
rect 195840 118526 195916 118734
rect 195840 118494 195846 118526
rect 195502 118462 195503 118494
rect 195437 118461 195503 118462
rect 195845 118462 195846 118494
rect 195910 118494 195916 118526
rect 196792 118734 196798 118766
rect 196862 118766 196863 118798
rect 196862 118734 196868 118766
rect 196792 118526 196868 118734
rect 195910 118462 195911 118494
rect 195845 118461 195911 118462
rect 196792 118462 196798 118526
rect 196862 118462 196868 118526
rect 196792 118456 196868 118462
rect 22168 118390 22244 118396
rect 22168 118326 22174 118390
rect 22238 118326 22244 118390
rect 22581 118390 22647 118391
rect 22581 118358 22582 118390
rect 952 118054 1230 118118
rect 1294 118054 1300 118118
rect 21765 118118 21831 118119
rect 21765 118086 21766 118118
rect 952 116486 1300 118054
rect 21760 118054 21766 118086
rect 21830 118086 21831 118118
rect 22168 118118 22244 118326
rect 22168 118086 22174 118118
rect 21830 118054 21836 118086
rect 21760 117846 21836 118054
rect 22173 118054 22174 118086
rect 22238 118086 22244 118118
rect 22576 118326 22582 118358
rect 22646 118358 22647 118390
rect 23120 118390 23196 118396
rect 22646 118326 22652 118358
rect 22576 118118 22652 118326
rect 22238 118054 22239 118086
rect 22173 118053 22239 118054
rect 22576 118054 22582 118118
rect 22646 118054 22652 118118
rect 23120 118326 23126 118390
rect 23190 118326 23196 118390
rect 23533 118390 23599 118391
rect 23533 118358 23534 118390
rect 23120 118118 23196 118326
rect 23120 118086 23126 118118
rect 22576 118048 22652 118054
rect 23125 118054 23126 118086
rect 23190 118086 23196 118118
rect 23528 118326 23534 118358
rect 23598 118358 23599 118390
rect 195160 118390 195236 118396
rect 23598 118326 23604 118358
rect 23528 118118 23604 118326
rect 23190 118054 23191 118086
rect 23125 118053 23191 118054
rect 23528 118054 23534 118118
rect 23598 118054 23604 118118
rect 195160 118326 195166 118390
rect 195230 118326 195236 118390
rect 195437 118390 195503 118391
rect 195437 118358 195438 118390
rect 195160 118118 195236 118326
rect 195160 118086 195166 118118
rect 23528 118048 23604 118054
rect 195165 118054 195166 118086
rect 195230 118086 195236 118118
rect 195432 118326 195438 118358
rect 195502 118358 195503 118390
rect 195845 118390 195911 118391
rect 195845 118358 195846 118390
rect 195502 118326 195508 118358
rect 195432 118118 195508 118326
rect 195230 118054 195231 118086
rect 195165 118053 195231 118054
rect 195432 118054 195438 118118
rect 195502 118054 195508 118118
rect 195432 118048 195508 118054
rect 195840 118326 195846 118358
rect 195910 118358 195911 118390
rect 196112 118390 196188 118396
rect 195910 118326 195916 118358
rect 195840 118118 195916 118326
rect 195840 118054 195846 118118
rect 195910 118054 195916 118118
rect 196112 118326 196118 118390
rect 196182 118326 196188 118390
rect 196112 118118 196188 118326
rect 196112 118086 196118 118118
rect 195840 118048 195916 118054
rect 196117 118054 196118 118086
rect 196182 118086 196188 118118
rect 196661 118118 196727 118119
rect 196661 118086 196662 118118
rect 196182 118054 196183 118086
rect 196117 118053 196183 118054
rect 196656 118054 196662 118086
rect 196726 118086 196727 118118
rect 196726 118054 196732 118086
rect 21760 117782 21766 117846
rect 21830 117782 21836 117846
rect 21760 117776 21836 117782
rect 22440 117982 22516 117988
rect 22440 117918 22446 117982
rect 22510 117918 22516 117982
rect 22440 117710 22516 117918
rect 22440 117678 22446 117710
rect 22445 117646 22446 117678
rect 22510 117678 22516 117710
rect 23120 117982 23196 117988
rect 23120 117918 23126 117982
rect 23190 117918 23196 117982
rect 23397 117982 23463 117983
rect 23397 117950 23398 117982
rect 23120 117710 23196 117918
rect 23120 117678 23126 117710
rect 22510 117646 22511 117678
rect 22445 117645 22511 117646
rect 23125 117646 23126 117678
rect 23190 117678 23196 117710
rect 23392 117918 23398 117950
rect 23462 117950 23463 117982
rect 195029 117982 195095 117983
rect 195029 117950 195030 117982
rect 23462 117918 23468 117950
rect 23392 117710 23468 117918
rect 195024 117918 195030 117950
rect 195094 117950 195095 117982
rect 195437 117982 195503 117983
rect 195437 117950 195438 117982
rect 195094 117918 195100 117950
rect 23190 117646 23191 117678
rect 23125 117645 23191 117646
rect 23392 117646 23398 117710
rect 23462 117646 23468 117710
rect 23392 117640 23468 117646
rect 28288 117710 28364 117716
rect 28288 117646 28294 117710
rect 28358 117646 28364 117710
rect 22576 117574 22652 117580
rect 22576 117510 22582 117574
rect 22646 117510 22652 117574
rect 21765 117302 21831 117303
rect 21765 117270 21766 117302
rect 21760 117238 21766 117270
rect 21830 117270 21831 117302
rect 22576 117302 22652 117510
rect 28288 117438 28364 117646
rect 195024 117710 195100 117918
rect 195024 117646 195030 117710
rect 195094 117646 195100 117710
rect 195024 117640 195100 117646
rect 195432 117918 195438 117950
rect 195502 117950 195503 117982
rect 195502 117918 195508 117950
rect 195432 117710 195508 117918
rect 196656 117846 196732 118054
rect 196656 117782 196662 117846
rect 196726 117782 196732 117846
rect 196656 117776 196732 117782
rect 195432 117646 195438 117710
rect 195502 117646 195508 117710
rect 216495 117675 216555 127844
rect 217464 126414 217812 128254
rect 217464 126350 217470 126414
rect 217534 126350 217812 126414
rect 216789 125462 216855 125463
rect 216789 125430 216790 125462
rect 216784 125398 216790 125430
rect 216854 125430 216855 125462
rect 216854 125398 216860 125430
rect 216784 124918 216860 125398
rect 216784 124854 216790 124918
rect 216854 124854 216860 124918
rect 216784 124848 216860 124854
rect 217464 124782 217812 126350
rect 217464 124718 217470 124782
rect 217534 124718 217812 124782
rect 216784 123150 216860 123156
rect 216784 123086 216790 123150
rect 216854 123086 216860 123150
rect 216784 122742 216860 123086
rect 216784 122710 216790 122742
rect 216789 122678 216790 122710
rect 216854 122710 216860 122742
rect 217464 123150 217812 124718
rect 217464 123086 217470 123150
rect 217534 123086 217812 123150
rect 216854 122678 216855 122710
rect 216789 122677 216855 122678
rect 217464 121518 217812 123086
rect 217464 121454 217470 121518
rect 217534 121454 217812 121518
rect 217464 119886 217812 121454
rect 217464 119822 217470 119886
rect 217534 119822 217812 119886
rect 217464 118254 217812 119822
rect 217464 118190 217470 118254
rect 217534 118190 217812 118254
rect 195432 117640 195508 117646
rect 216492 117674 216558 117675
rect 216492 117610 216493 117674
rect 216557 117610 216558 117674
rect 216492 117609 216558 117610
rect 195840 117574 195916 117580
rect 195840 117510 195846 117574
rect 195910 117510 195916 117574
rect 28288 117406 28294 117438
rect 28293 117374 28294 117406
rect 28358 117406 28364 117438
rect 28429 117438 28495 117439
rect 28429 117406 28430 117438
rect 28358 117374 28359 117406
rect 28293 117373 28359 117374
rect 28424 117374 28430 117406
rect 28494 117406 28495 117438
rect 190128 117438 190204 117444
rect 28494 117374 28500 117406
rect 22576 117270 22582 117302
rect 21830 117238 21836 117270
rect 21760 117030 21836 117238
rect 22581 117238 22582 117270
rect 22646 117270 22652 117302
rect 22646 117238 22647 117270
rect 22581 117237 22647 117238
rect 28424 117166 28500 117374
rect 28424 117102 28430 117166
rect 28494 117102 28500 117166
rect 190128 117374 190134 117438
rect 190198 117374 190204 117438
rect 190128 117166 190204 117374
rect 195840 117302 195916 117510
rect 195840 117270 195846 117302
rect 195845 117238 195846 117270
rect 195910 117270 195916 117302
rect 196661 117302 196727 117303
rect 196661 117270 196662 117302
rect 195910 117238 195911 117270
rect 195845 117237 195911 117238
rect 196656 117238 196662 117270
rect 196726 117270 196727 117302
rect 196726 117238 196732 117270
rect 190128 117134 190134 117166
rect 28424 117096 28500 117102
rect 190133 117102 190134 117134
rect 190198 117134 190204 117166
rect 190198 117102 190199 117134
rect 190133 117101 190199 117102
rect 21760 116966 21766 117030
rect 21830 116966 21836 117030
rect 21760 116960 21836 116966
rect 28560 117030 28636 117036
rect 28560 116966 28566 117030
rect 28630 116966 28636 117030
rect 21901 116894 21967 116895
rect 21901 116862 21902 116894
rect 21896 116830 21902 116862
rect 21966 116862 21967 116894
rect 22304 116894 22380 116900
rect 21966 116830 21972 116862
rect 21896 116622 21972 116830
rect 21896 116558 21902 116622
rect 21966 116558 21972 116622
rect 22304 116830 22310 116894
rect 22374 116830 22380 116894
rect 22304 116622 22380 116830
rect 22304 116590 22310 116622
rect 21896 116552 21972 116558
rect 22309 116558 22310 116590
rect 22374 116590 22380 116622
rect 22440 116894 22516 116900
rect 22440 116830 22446 116894
rect 22510 116830 22516 116894
rect 22440 116622 22516 116830
rect 28560 116758 28636 116966
rect 28560 116726 28566 116758
rect 28565 116694 28566 116726
rect 28630 116726 28636 116758
rect 190264 117030 190340 117036
rect 190264 116966 190270 117030
rect 190334 116966 190340 117030
rect 190264 116758 190340 116966
rect 196656 117030 196732 117238
rect 196656 116966 196662 117030
rect 196726 116966 196732 117030
rect 196656 116960 196732 116966
rect 190264 116726 190270 116758
rect 28630 116694 28631 116726
rect 28565 116693 28631 116694
rect 190269 116694 190270 116726
rect 190334 116726 190340 116758
rect 195840 116894 195916 116900
rect 195840 116830 195846 116894
rect 195910 116830 195916 116894
rect 190334 116694 190335 116726
rect 190269 116693 190335 116694
rect 22440 116590 22446 116622
rect 22374 116558 22375 116590
rect 22309 116557 22375 116558
rect 22445 116558 22446 116590
rect 22510 116590 22516 116622
rect 28429 116622 28495 116623
rect 28429 116590 28430 116622
rect 22510 116558 22511 116590
rect 22445 116557 22511 116558
rect 28424 116558 28430 116590
rect 28494 116590 28495 116622
rect 190269 116622 190335 116623
rect 190269 116590 190270 116622
rect 28494 116558 28500 116590
rect 952 116422 1230 116486
rect 1294 116422 1300 116486
rect 21901 116486 21967 116487
rect 21901 116454 21902 116486
rect 952 114718 1300 116422
rect 21896 116422 21902 116454
rect 21966 116454 21967 116486
rect 23125 116486 23191 116487
rect 23125 116454 23126 116486
rect 21966 116422 21972 116454
rect 21896 116214 21972 116422
rect 21896 116150 21902 116214
rect 21966 116150 21972 116214
rect 21896 116144 21972 116150
rect 23120 116422 23126 116454
rect 23190 116454 23191 116486
rect 23528 116486 23604 116492
rect 23190 116422 23196 116454
rect 23120 116214 23196 116422
rect 23120 116150 23126 116214
rect 23190 116150 23196 116214
rect 23528 116422 23534 116486
rect 23598 116422 23604 116486
rect 23528 116214 23604 116422
rect 28424 116350 28500 116558
rect 28424 116286 28430 116350
rect 28494 116286 28500 116350
rect 28424 116280 28500 116286
rect 190264 116558 190270 116590
rect 190334 116590 190335 116622
rect 195840 116622 195916 116830
rect 195840 116590 195846 116622
rect 190334 116558 190340 116590
rect 190264 116350 190340 116558
rect 195845 116558 195846 116590
rect 195910 116590 195916 116622
rect 196112 116894 196188 116900
rect 196112 116830 196118 116894
rect 196182 116830 196188 116894
rect 196112 116622 196188 116830
rect 196112 116590 196118 116622
rect 195910 116558 195911 116590
rect 195845 116557 195911 116558
rect 196117 116558 196118 116590
rect 196182 116590 196188 116622
rect 196792 116894 196868 116900
rect 196792 116830 196798 116894
rect 196862 116830 196868 116894
rect 216789 116894 216855 116895
rect 216789 116862 216790 116894
rect 196792 116622 196868 116830
rect 196792 116590 196798 116622
rect 196182 116558 196183 116590
rect 196117 116557 196183 116558
rect 196797 116558 196798 116590
rect 196862 116590 196868 116622
rect 216784 116830 216790 116862
rect 216854 116862 216855 116894
rect 216854 116830 216860 116862
rect 196862 116558 196863 116590
rect 196797 116557 196863 116558
rect 190264 116286 190270 116350
rect 190334 116286 190340 116350
rect 190264 116280 190340 116286
rect 195160 116486 195236 116492
rect 195160 116422 195166 116486
rect 195230 116422 195236 116486
rect 23528 116182 23534 116214
rect 23120 116144 23196 116150
rect 23533 116150 23534 116182
rect 23598 116182 23604 116214
rect 195160 116214 195236 116422
rect 195160 116182 195166 116214
rect 23598 116150 23599 116182
rect 23533 116149 23599 116150
rect 195165 116150 195166 116182
rect 195230 116182 195236 116214
rect 195432 116486 195508 116492
rect 195432 116422 195438 116486
rect 195502 116422 195508 116486
rect 196797 116486 196863 116487
rect 196797 116454 196798 116486
rect 195432 116214 195508 116422
rect 195432 116182 195438 116214
rect 195230 116150 195231 116182
rect 195165 116149 195231 116150
rect 195437 116150 195438 116182
rect 195502 116182 195508 116214
rect 196792 116422 196798 116454
rect 196862 116454 196863 116486
rect 216784 116486 216860 116830
rect 196862 116422 196868 116454
rect 196792 116214 196868 116422
rect 216784 116422 216790 116486
rect 216854 116422 216860 116486
rect 216784 116416 216860 116422
rect 195502 116150 195503 116182
rect 195437 116149 195503 116150
rect 196792 116150 196798 116214
rect 196862 116150 196868 116214
rect 196792 116144 196868 116150
rect 217464 116350 217812 118190
rect 217464 116286 217470 116350
rect 217534 116286 217812 116350
rect 21896 116078 21972 116084
rect 21896 116014 21902 116078
rect 21966 116014 21972 116078
rect 22173 116078 22239 116079
rect 22173 116046 22174 116078
rect 21896 115806 21972 116014
rect 21896 115774 21902 115806
rect 21901 115742 21902 115774
rect 21966 115774 21972 115806
rect 22168 116014 22174 116046
rect 22238 116046 22239 116078
rect 22581 116078 22647 116079
rect 22581 116046 22582 116078
rect 22238 116014 22244 116046
rect 22168 115806 22244 116014
rect 21966 115742 21967 115774
rect 21901 115741 21967 115742
rect 22168 115742 22174 115806
rect 22238 115742 22244 115806
rect 22168 115736 22244 115742
rect 22576 116014 22582 116046
rect 22646 116046 22647 116078
rect 22984 116078 23060 116084
rect 22646 116014 22652 116046
rect 22576 115806 22652 116014
rect 22576 115742 22582 115806
rect 22646 115742 22652 115806
rect 22984 116014 22990 116078
rect 23054 116014 23060 116078
rect 22984 115806 23060 116014
rect 22984 115774 22990 115806
rect 22576 115736 22652 115742
rect 22989 115742 22990 115774
rect 23054 115774 23060 115806
rect 23392 116078 23468 116084
rect 23392 116014 23398 116078
rect 23462 116014 23468 116078
rect 195165 116078 195231 116079
rect 195165 116046 195166 116078
rect 23392 115806 23468 116014
rect 23392 115774 23398 115806
rect 23054 115742 23055 115774
rect 22989 115741 23055 115742
rect 23397 115742 23398 115774
rect 23462 115774 23468 115806
rect 195160 116014 195166 116046
rect 195230 116046 195231 116078
rect 195437 116078 195503 116079
rect 195437 116046 195438 116078
rect 195230 116014 195236 116046
rect 195160 115806 195236 116014
rect 23462 115742 23463 115774
rect 23397 115741 23463 115742
rect 195160 115742 195166 115806
rect 195230 115742 195236 115806
rect 195160 115736 195236 115742
rect 195432 116014 195438 116046
rect 195502 116046 195503 116078
rect 195976 116078 196052 116084
rect 195502 116014 195508 116046
rect 195432 115806 195508 116014
rect 195432 115742 195438 115806
rect 195502 115742 195508 115806
rect 195976 116014 195982 116078
rect 196046 116014 196052 116078
rect 195976 115806 196052 116014
rect 195976 115774 195982 115806
rect 195432 115736 195508 115742
rect 195981 115742 195982 115774
rect 196046 115774 196052 115806
rect 196112 116078 196188 116084
rect 196112 116014 196118 116078
rect 196182 116014 196188 116078
rect 196112 115806 196188 116014
rect 196112 115774 196118 115806
rect 196046 115742 196047 115774
rect 195981 115741 196047 115742
rect 196117 115742 196118 115774
rect 196182 115774 196188 115806
rect 196792 116078 196868 116084
rect 196792 116014 196798 116078
rect 196862 116014 196868 116078
rect 196792 115806 196868 116014
rect 196792 115774 196798 115806
rect 196182 115742 196183 115774
rect 196117 115741 196183 115742
rect 196797 115742 196798 115774
rect 196862 115774 196868 115806
rect 196862 115742 196863 115774
rect 196797 115741 196863 115742
rect 21896 115670 21972 115676
rect 21896 115606 21902 115670
rect 21966 115606 21972 115670
rect 22309 115670 22375 115671
rect 22309 115638 22310 115670
rect 21896 115398 21972 115606
rect 21896 115366 21902 115398
rect 21901 115334 21902 115366
rect 21966 115366 21972 115398
rect 22304 115606 22310 115638
rect 22374 115638 22375 115670
rect 22445 115670 22511 115671
rect 22445 115638 22446 115670
rect 22374 115606 22380 115638
rect 22304 115398 22380 115606
rect 21966 115334 21967 115366
rect 21901 115333 21967 115334
rect 22304 115334 22310 115398
rect 22374 115334 22380 115398
rect 22304 115328 22380 115334
rect 22440 115606 22446 115638
rect 22510 115638 22511 115670
rect 22989 115670 23055 115671
rect 22989 115638 22990 115670
rect 22510 115606 22516 115638
rect 22440 115398 22516 115606
rect 22440 115334 22446 115398
rect 22510 115334 22516 115398
rect 22440 115328 22516 115334
rect 22984 115606 22990 115638
rect 23054 115638 23055 115670
rect 23397 115670 23463 115671
rect 23397 115638 23398 115670
rect 23054 115606 23060 115638
rect 22984 115398 23060 115606
rect 22984 115334 22990 115398
rect 23054 115334 23060 115398
rect 22984 115328 23060 115334
rect 23392 115606 23398 115638
rect 23462 115638 23463 115670
rect 195029 115670 195095 115671
rect 195029 115638 195030 115670
rect 23462 115606 23468 115638
rect 23392 115398 23468 115606
rect 23392 115334 23398 115398
rect 23462 115334 23468 115398
rect 23392 115328 23468 115334
rect 195024 115606 195030 115638
rect 195094 115638 195095 115670
rect 195437 115670 195503 115671
rect 195437 115638 195438 115670
rect 195094 115606 195100 115638
rect 195024 115398 195100 115606
rect 195024 115334 195030 115398
rect 195094 115334 195100 115398
rect 195024 115328 195100 115334
rect 195432 115606 195438 115638
rect 195502 115638 195503 115670
rect 196384 115670 196460 115676
rect 195502 115606 195508 115638
rect 195432 115398 195508 115606
rect 195432 115334 195438 115398
rect 195502 115334 195508 115398
rect 196384 115606 196390 115670
rect 196454 115606 196460 115670
rect 196384 115398 196460 115606
rect 196384 115366 196390 115398
rect 195432 115328 195508 115334
rect 196389 115334 196390 115366
rect 196454 115366 196460 115398
rect 196792 115670 196868 115676
rect 196792 115606 196798 115670
rect 196862 115606 196868 115670
rect 196792 115398 196868 115606
rect 196792 115366 196798 115398
rect 196454 115334 196455 115366
rect 196389 115333 196455 115334
rect 196797 115334 196798 115366
rect 196862 115366 196868 115398
rect 196862 115334 196863 115366
rect 196797 115333 196863 115334
rect 21760 115262 21836 115268
rect 21760 115198 21766 115262
rect 21830 115198 21836 115262
rect 21760 114990 21836 115198
rect 21760 114958 21766 114990
rect 21765 114926 21766 114958
rect 21830 114958 21836 114990
rect 22168 115262 22244 115268
rect 22168 115198 22174 115262
rect 22238 115198 22244 115262
rect 22445 115262 22511 115263
rect 22445 115230 22446 115262
rect 22168 114990 22244 115198
rect 22168 114958 22174 114990
rect 21830 114926 21831 114958
rect 21765 114925 21831 114926
rect 22173 114926 22174 114958
rect 22238 114958 22244 114990
rect 22440 115198 22446 115230
rect 22510 115230 22511 115262
rect 23120 115262 23196 115268
rect 22510 115198 22516 115230
rect 22440 114990 22516 115198
rect 22238 114926 22239 114958
rect 22173 114925 22239 114926
rect 22440 114926 22446 114990
rect 22510 114926 22516 114990
rect 23120 115198 23126 115262
rect 23190 115198 23196 115262
rect 23533 115262 23599 115263
rect 23533 115230 23534 115262
rect 23120 114990 23196 115198
rect 23120 114958 23126 114990
rect 22440 114920 22516 114926
rect 23125 114926 23126 114958
rect 23190 114958 23196 114990
rect 23528 115198 23534 115230
rect 23598 115230 23599 115262
rect 195160 115262 195236 115268
rect 23598 115198 23604 115230
rect 23528 114990 23604 115198
rect 23190 114926 23191 114958
rect 23125 114925 23191 114926
rect 23528 114926 23534 114990
rect 23598 114926 23604 114990
rect 195160 115198 195166 115262
rect 195230 115198 195236 115262
rect 195437 115262 195503 115263
rect 195437 115230 195438 115262
rect 195160 114990 195236 115198
rect 195160 114958 195166 114990
rect 23528 114920 23604 114926
rect 195165 114926 195166 114958
rect 195230 114958 195236 114990
rect 195432 115198 195438 115230
rect 195502 115230 195503 115262
rect 195845 115262 195911 115263
rect 195845 115230 195846 115262
rect 195502 115198 195508 115230
rect 195432 114990 195508 115198
rect 195230 114926 195231 114958
rect 195165 114925 195231 114926
rect 195432 114926 195438 114990
rect 195502 114926 195508 114990
rect 195432 114920 195508 114926
rect 195840 115198 195846 115230
rect 195910 115230 195911 115262
rect 196253 115262 196319 115263
rect 196253 115230 196254 115262
rect 195910 115198 195916 115230
rect 195840 114990 195916 115198
rect 195840 114926 195846 114990
rect 195910 114926 195916 114990
rect 195840 114920 195916 114926
rect 196248 115198 196254 115230
rect 196318 115230 196319 115262
rect 196661 115262 196727 115263
rect 196661 115230 196662 115262
rect 196318 115198 196324 115230
rect 196248 114990 196324 115198
rect 196248 114926 196254 114990
rect 196318 114926 196324 114990
rect 196248 114920 196324 114926
rect 196656 115198 196662 115230
rect 196726 115230 196727 115262
rect 196726 115198 196732 115230
rect 196656 114990 196732 115198
rect 196656 114926 196662 114990
rect 196726 114926 196732 114990
rect 196656 114920 196732 114926
rect 21765 114854 21831 114855
rect 21765 114822 21766 114854
rect 952 114654 1230 114718
rect 1294 114654 1300 114718
rect 952 113086 1300 114654
rect 21760 114790 21766 114822
rect 21830 114822 21831 114854
rect 22440 114854 22516 114860
rect 21830 114790 21836 114822
rect 21760 114582 21836 114790
rect 21760 114518 21766 114582
rect 21830 114518 21836 114582
rect 22440 114790 22446 114854
rect 22510 114790 22516 114854
rect 23125 114854 23191 114855
rect 23125 114822 23126 114854
rect 22440 114582 22516 114790
rect 22440 114550 22446 114582
rect 21760 114512 21836 114518
rect 22445 114518 22446 114550
rect 22510 114550 22516 114582
rect 23120 114790 23126 114822
rect 23190 114822 23191 114854
rect 23392 114854 23468 114860
rect 23190 114790 23196 114822
rect 23120 114582 23196 114790
rect 22510 114518 22511 114550
rect 22445 114517 22511 114518
rect 23120 114518 23126 114582
rect 23190 114518 23196 114582
rect 23392 114790 23398 114854
rect 23462 114790 23468 114854
rect 23392 114582 23468 114790
rect 23392 114550 23398 114582
rect 23120 114512 23196 114518
rect 23397 114518 23398 114550
rect 23462 114550 23468 114582
rect 195024 114854 195100 114860
rect 195024 114790 195030 114854
rect 195094 114790 195100 114854
rect 195573 114854 195639 114855
rect 195573 114822 195574 114854
rect 195024 114582 195100 114790
rect 195024 114550 195030 114582
rect 23462 114518 23463 114550
rect 23397 114517 23463 114518
rect 195029 114518 195030 114550
rect 195094 114550 195100 114582
rect 195568 114790 195574 114822
rect 195638 114822 195639 114854
rect 195976 114854 196052 114860
rect 195638 114790 195644 114822
rect 195568 114582 195644 114790
rect 195094 114518 195095 114550
rect 195029 114517 195095 114518
rect 195568 114518 195574 114582
rect 195638 114518 195644 114582
rect 195976 114790 195982 114854
rect 196046 114790 196052 114854
rect 195976 114582 196052 114790
rect 195976 114550 195982 114582
rect 195568 114512 195644 114518
rect 195981 114518 195982 114550
rect 196046 114550 196052 114582
rect 196792 114854 196868 114860
rect 196792 114790 196798 114854
rect 196862 114790 196868 114854
rect 196792 114582 196868 114790
rect 196792 114550 196798 114582
rect 196046 114518 196047 114550
rect 195981 114517 196047 114518
rect 196797 114518 196798 114550
rect 196862 114550 196868 114582
rect 217464 114854 217812 116286
rect 217464 114790 217470 114854
rect 217534 114790 217812 114854
rect 196862 114518 196863 114550
rect 196797 114517 196863 114518
rect 22168 114446 22244 114452
rect 22168 114382 22174 114446
rect 22238 114382 22244 114446
rect 22989 114446 23055 114447
rect 22989 114414 22990 114446
rect 22168 114174 22244 114382
rect 22168 114142 22174 114174
rect 22173 114110 22174 114142
rect 22238 114142 22244 114174
rect 22984 114382 22990 114414
rect 23054 114414 23055 114446
rect 23528 114446 23604 114452
rect 23054 114382 23060 114414
rect 22984 114174 23060 114382
rect 22238 114110 22239 114142
rect 22173 114109 22239 114110
rect 22984 114110 22990 114174
rect 23054 114110 23060 114174
rect 23528 114382 23534 114446
rect 23598 114382 23604 114446
rect 195029 114446 195095 114447
rect 195029 114414 195030 114446
rect 23528 114174 23604 114382
rect 195024 114382 195030 114414
rect 195094 114414 195095 114446
rect 195432 114446 195508 114452
rect 195094 114382 195100 114414
rect 28565 114310 28631 114311
rect 28565 114278 28566 114310
rect 23528 114142 23534 114174
rect 22984 114104 23060 114110
rect 23533 114110 23534 114142
rect 23598 114142 23604 114174
rect 28560 114246 28566 114278
rect 28630 114278 28631 114310
rect 190269 114310 190335 114311
rect 190269 114278 190270 114310
rect 28630 114246 28636 114278
rect 23598 114110 23599 114142
rect 23533 114109 23599 114110
rect 23120 114038 23196 114044
rect 23120 113974 23126 114038
rect 23190 113974 23196 114038
rect 23533 114038 23599 114039
rect 23533 114006 23534 114038
rect 23120 113766 23196 113974
rect 23120 113734 23126 113766
rect 23125 113702 23126 113734
rect 23190 113734 23196 113766
rect 23528 113974 23534 114006
rect 23598 114006 23599 114038
rect 28560 114038 28636 114246
rect 23598 113974 23604 114006
rect 23528 113766 23604 113974
rect 28560 113974 28566 114038
rect 28630 113974 28636 114038
rect 28560 113968 28636 113974
rect 190264 114246 190270 114278
rect 190334 114278 190335 114310
rect 190334 114246 190340 114278
rect 190264 114038 190340 114246
rect 195024 114174 195100 114382
rect 195024 114110 195030 114174
rect 195094 114110 195100 114174
rect 195432 114382 195438 114446
rect 195502 114382 195508 114446
rect 196389 114446 196455 114447
rect 196389 114414 196390 114446
rect 195432 114174 195508 114382
rect 195432 114142 195438 114174
rect 195024 114104 195100 114110
rect 195437 114110 195438 114142
rect 195502 114142 195508 114174
rect 196384 114382 196390 114414
rect 196454 114414 196455 114446
rect 196454 114382 196460 114414
rect 196384 114174 196460 114382
rect 195502 114110 195503 114142
rect 195437 114109 195503 114110
rect 196384 114110 196390 114174
rect 196454 114110 196460 114174
rect 196384 114104 196460 114110
rect 190264 113974 190270 114038
rect 190334 113974 190340 114038
rect 195165 114038 195231 114039
rect 195165 114006 195166 114038
rect 190264 113968 190340 113974
rect 195160 113974 195166 114006
rect 195230 114006 195231 114038
rect 195568 114038 195644 114044
rect 195230 113974 195236 114006
rect 23190 113702 23191 113734
rect 23125 113701 23191 113702
rect 23528 113702 23534 113766
rect 23598 113702 23604 113766
rect 28293 113766 28359 113767
rect 28293 113734 28294 113766
rect 23528 113696 23604 113702
rect 28288 113702 28294 113734
rect 28358 113734 28359 113766
rect 195160 113766 195236 113974
rect 28358 113702 28364 113734
rect 22173 113630 22239 113631
rect 22173 113598 22174 113630
rect 22168 113566 22174 113598
rect 22238 113598 22239 113630
rect 22238 113566 22244 113598
rect 952 113022 1230 113086
rect 1294 113022 1300 113086
rect 21760 113358 21836 113364
rect 21760 113294 21766 113358
rect 21830 113294 21836 113358
rect 21760 113086 21836 113294
rect 22168 113358 22244 113566
rect 28288 113494 28364 113702
rect 195160 113702 195166 113766
rect 195230 113702 195236 113766
rect 195568 113974 195574 114038
rect 195638 113974 195644 114038
rect 195568 113766 195644 113974
rect 195568 113734 195574 113766
rect 195160 113696 195236 113702
rect 195573 113702 195574 113734
rect 195638 113734 195644 113766
rect 195638 113702 195639 113734
rect 195573 113701 195639 113702
rect 195976 113630 196052 113636
rect 195976 113566 195982 113630
rect 196046 113566 196052 113630
rect 28288 113430 28294 113494
rect 28358 113430 28364 113494
rect 190133 113494 190199 113495
rect 190133 113462 190134 113494
rect 28288 113424 28364 113430
rect 190128 113430 190134 113462
rect 190198 113462 190199 113494
rect 190198 113430 190204 113462
rect 22168 113294 22174 113358
rect 22238 113294 22244 113358
rect 22168 113288 22244 113294
rect 190128 113222 190204 113430
rect 195976 113358 196052 113566
rect 195976 113326 195982 113358
rect 195981 113294 195982 113326
rect 196046 113326 196052 113358
rect 196112 113630 196188 113636
rect 196112 113566 196118 113630
rect 196182 113566 196188 113630
rect 196112 113358 196188 113566
rect 196112 113326 196118 113358
rect 196046 113294 196047 113326
rect 195981 113293 196047 113294
rect 196117 113294 196118 113326
rect 196182 113326 196188 113358
rect 196656 113358 196732 113364
rect 196182 113294 196183 113326
rect 196117 113293 196183 113294
rect 196656 113294 196662 113358
rect 196726 113294 196732 113358
rect 190128 113158 190134 113222
rect 190198 113158 190204 113222
rect 190269 113222 190335 113223
rect 190269 113190 190270 113222
rect 190128 113152 190204 113158
rect 190264 113158 190270 113190
rect 190334 113190 190335 113222
rect 190334 113158 190340 113190
rect 21760 113054 21766 113086
rect 952 111318 1300 113022
rect 21765 113022 21766 113054
rect 21830 113054 21836 113086
rect 28429 113086 28495 113087
rect 28429 113054 28430 113086
rect 21830 113022 21831 113054
rect 21765 113021 21831 113022
rect 28424 113022 28430 113054
rect 28494 113054 28495 113086
rect 190128 113086 190204 113092
rect 28494 113022 28500 113054
rect 21760 112950 21836 112956
rect 21760 112886 21766 112950
rect 21830 112886 21836 112950
rect 22581 112950 22647 112951
rect 22581 112918 22582 112950
rect 21760 112678 21836 112886
rect 21760 112646 21766 112678
rect 21765 112614 21766 112646
rect 21830 112646 21836 112678
rect 22576 112886 22582 112918
rect 22646 112918 22647 112950
rect 22646 112886 22652 112918
rect 22576 112678 22652 112886
rect 28424 112814 28500 113022
rect 28424 112750 28430 112814
rect 28494 112750 28500 112814
rect 28424 112744 28500 112750
rect 190128 113022 190134 113086
rect 190198 113022 190204 113086
rect 21830 112614 21831 112646
rect 21765 112613 21831 112614
rect 22576 112614 22582 112678
rect 22646 112614 22652 112678
rect 190128 112678 190204 113022
rect 190264 112814 190340 113158
rect 196656 113086 196732 113294
rect 196656 113054 196662 113086
rect 196661 113022 196662 113054
rect 196726 113054 196732 113086
rect 196726 113022 196727 113054
rect 196661 113021 196727 113022
rect 190264 112750 190270 112814
rect 190334 112750 190340 112814
rect 190264 112744 190340 112750
rect 195976 112950 196052 112956
rect 195976 112886 195982 112950
rect 196046 112886 196052 112950
rect 196661 112950 196727 112951
rect 196661 112918 196662 112950
rect 190128 112646 190134 112678
rect 22576 112608 22652 112614
rect 190133 112614 190134 112646
rect 190198 112646 190204 112678
rect 195976 112678 196052 112886
rect 195976 112646 195982 112678
rect 190198 112614 190199 112646
rect 190133 112613 190199 112614
rect 195981 112614 195982 112646
rect 196046 112646 196052 112678
rect 196656 112886 196662 112918
rect 196726 112918 196727 112950
rect 217464 112950 217812 114790
rect 196726 112886 196732 112918
rect 196656 112678 196732 112886
rect 196046 112614 196047 112646
rect 195981 112613 196047 112614
rect 196656 112614 196662 112678
rect 196726 112614 196732 112678
rect 196656 112608 196732 112614
rect 217464 112886 217470 112950
rect 217534 112886 217812 112950
rect 21901 112542 21967 112543
rect 21901 112510 21902 112542
rect 21896 112478 21902 112510
rect 21966 112510 21967 112542
rect 23120 112542 23196 112548
rect 21966 112478 21972 112510
rect 21896 112270 21972 112478
rect 21896 112206 21902 112270
rect 21966 112206 21972 112270
rect 23120 112478 23126 112542
rect 23190 112478 23196 112542
rect 23120 112270 23196 112478
rect 23120 112238 23126 112270
rect 21896 112200 21972 112206
rect 23125 112206 23126 112238
rect 23190 112238 23196 112270
rect 23392 112542 23468 112548
rect 23392 112478 23398 112542
rect 23462 112478 23468 112542
rect 195029 112542 195095 112543
rect 195029 112510 195030 112542
rect 23392 112270 23468 112478
rect 23392 112238 23398 112270
rect 23190 112206 23191 112238
rect 23125 112205 23191 112206
rect 23397 112206 23398 112238
rect 23462 112238 23468 112270
rect 195024 112478 195030 112510
rect 195094 112510 195095 112542
rect 195568 112542 195644 112548
rect 195094 112478 195100 112510
rect 195024 112270 195100 112478
rect 23462 112206 23463 112238
rect 23397 112205 23463 112206
rect 195024 112206 195030 112270
rect 195094 112206 195100 112270
rect 195568 112478 195574 112542
rect 195638 112478 195644 112542
rect 196797 112542 196863 112543
rect 196797 112510 196798 112542
rect 195568 112270 195644 112478
rect 195568 112238 195574 112270
rect 195024 112200 195100 112206
rect 195573 112206 195574 112238
rect 195638 112238 195644 112270
rect 196792 112478 196798 112510
rect 196862 112510 196863 112542
rect 196862 112478 196868 112510
rect 196792 112270 196868 112478
rect 195638 112206 195639 112238
rect 195573 112205 195639 112206
rect 196792 112206 196798 112270
rect 196862 112206 196868 112270
rect 196792 112200 196868 112206
rect 21901 112134 21967 112135
rect 21901 112102 21902 112134
rect 21896 112070 21902 112102
rect 21966 112102 21967 112134
rect 22309 112134 22375 112135
rect 22309 112102 22310 112134
rect 21966 112070 21972 112102
rect 21896 111862 21972 112070
rect 21896 111798 21902 111862
rect 21966 111798 21972 111862
rect 21896 111792 21972 111798
rect 22304 112070 22310 112102
rect 22374 112102 22375 112134
rect 22445 112134 22511 112135
rect 22445 112102 22446 112134
rect 22374 112070 22380 112102
rect 22304 111862 22380 112070
rect 22304 111798 22310 111862
rect 22374 111798 22380 111862
rect 22304 111792 22380 111798
rect 22440 112070 22446 112102
rect 22510 112102 22511 112134
rect 22984 112134 23060 112140
rect 22510 112070 22516 112102
rect 22440 111862 22516 112070
rect 22440 111798 22446 111862
rect 22510 111798 22516 111862
rect 22984 112070 22990 112134
rect 23054 112070 23060 112134
rect 23397 112134 23463 112135
rect 23397 112102 23398 112134
rect 22984 111862 23060 112070
rect 22984 111830 22990 111862
rect 22440 111792 22516 111798
rect 22989 111798 22990 111830
rect 23054 111830 23060 111862
rect 23392 112070 23398 112102
rect 23462 112102 23463 112134
rect 195029 112134 195095 112135
rect 195029 112102 195030 112134
rect 23462 112070 23468 112102
rect 23392 111862 23468 112070
rect 195024 112070 195030 112102
rect 195094 112102 195095 112134
rect 195432 112134 195508 112140
rect 195094 112070 195100 112102
rect 23054 111798 23055 111830
rect 22989 111797 23055 111798
rect 23392 111798 23398 111862
rect 23462 111798 23468 111862
rect 28293 111862 28359 111863
rect 28293 111830 28294 111862
rect 23392 111792 23468 111798
rect 28288 111798 28294 111830
rect 28358 111830 28359 111862
rect 195024 111862 195100 112070
rect 28358 111798 28364 111830
rect 21896 111726 21972 111732
rect 21896 111662 21902 111726
rect 21966 111662 21972 111726
rect 22173 111726 22239 111727
rect 22173 111694 22174 111726
rect 21896 111454 21972 111662
rect 21896 111422 21902 111454
rect 21901 111390 21902 111422
rect 21966 111422 21972 111454
rect 22168 111662 22174 111694
rect 22238 111694 22239 111726
rect 22581 111726 22647 111727
rect 22581 111694 22582 111726
rect 22238 111662 22244 111694
rect 22168 111454 22244 111662
rect 21966 111390 21967 111422
rect 21901 111389 21967 111390
rect 22168 111390 22174 111454
rect 22238 111390 22244 111454
rect 22168 111384 22244 111390
rect 22576 111662 22582 111694
rect 22646 111694 22647 111726
rect 23125 111726 23191 111727
rect 23125 111694 23126 111726
rect 22646 111662 22652 111694
rect 22576 111454 22652 111662
rect 22576 111390 22582 111454
rect 22646 111390 22652 111454
rect 22576 111384 22652 111390
rect 23120 111662 23126 111694
rect 23190 111694 23191 111726
rect 23533 111726 23599 111727
rect 23533 111694 23534 111726
rect 23190 111662 23196 111694
rect 23120 111454 23196 111662
rect 23120 111390 23126 111454
rect 23190 111390 23196 111454
rect 23120 111384 23196 111390
rect 23528 111662 23534 111694
rect 23598 111694 23599 111726
rect 23598 111662 23604 111694
rect 23528 111454 23604 111662
rect 28288 111590 28364 111798
rect 195024 111798 195030 111862
rect 195094 111798 195100 111862
rect 195432 112070 195438 112134
rect 195502 112070 195508 112134
rect 195432 111862 195508 112070
rect 195432 111830 195438 111862
rect 195024 111792 195100 111798
rect 195437 111798 195438 111830
rect 195502 111830 195508 111862
rect 196656 112134 196732 112140
rect 196656 112070 196662 112134
rect 196726 112070 196732 112134
rect 196656 111862 196732 112070
rect 196656 111830 196662 111862
rect 195502 111798 195503 111830
rect 195437 111797 195503 111798
rect 196661 111798 196662 111830
rect 196726 111830 196732 111862
rect 196726 111798 196727 111830
rect 196661 111797 196727 111798
rect 28288 111526 28294 111590
rect 28358 111526 28364 111590
rect 28288 111520 28364 111526
rect 195024 111726 195100 111732
rect 195024 111662 195030 111726
rect 195094 111662 195100 111726
rect 195573 111726 195639 111727
rect 195573 111694 195574 111726
rect 23528 111390 23534 111454
rect 23598 111390 23604 111454
rect 195024 111454 195100 111662
rect 195024 111422 195030 111454
rect 23528 111384 23604 111390
rect 195029 111390 195030 111422
rect 195094 111422 195100 111454
rect 195568 111662 195574 111694
rect 195638 111694 195639 111726
rect 195976 111726 196052 111732
rect 195638 111662 195644 111694
rect 195568 111454 195644 111662
rect 195094 111390 195095 111422
rect 195029 111389 195095 111390
rect 195568 111390 195574 111454
rect 195638 111390 195644 111454
rect 195976 111662 195982 111726
rect 196046 111662 196052 111726
rect 196661 111726 196727 111727
rect 196661 111694 196662 111726
rect 195976 111454 196052 111662
rect 195976 111422 195982 111454
rect 195568 111384 195644 111390
rect 195981 111390 195982 111422
rect 196046 111422 196052 111454
rect 196656 111662 196662 111694
rect 196726 111694 196727 111726
rect 196726 111662 196732 111694
rect 196656 111454 196732 111662
rect 196046 111390 196047 111422
rect 195981 111389 196047 111390
rect 196656 111390 196662 111454
rect 196726 111390 196732 111454
rect 196656 111384 196732 111390
rect 217464 111454 217812 112886
rect 217464 111390 217470 111454
rect 217534 111390 217812 111454
rect 952 111254 1230 111318
rect 1294 111254 1300 111318
rect 21901 111318 21967 111319
rect 21901 111286 21902 111318
rect 952 109686 1300 111254
rect 21896 111254 21902 111286
rect 21966 111286 21967 111318
rect 22445 111318 22511 111319
rect 22445 111286 22446 111318
rect 21966 111254 21972 111286
rect 21896 111046 21972 111254
rect 21896 110982 21902 111046
rect 21966 110982 21972 111046
rect 21896 110976 21972 110982
rect 22440 111254 22446 111286
rect 22510 111286 22511 111318
rect 23120 111318 23196 111324
rect 22510 111254 22516 111286
rect 22440 111046 22516 111254
rect 22440 110982 22446 111046
rect 22510 110982 22516 111046
rect 23120 111254 23126 111318
rect 23190 111254 23196 111318
rect 23120 111046 23196 111254
rect 23120 111014 23126 111046
rect 22440 110976 22516 110982
rect 23125 110982 23126 111014
rect 23190 111014 23196 111046
rect 23392 111318 23468 111324
rect 23392 111254 23398 111318
rect 23462 111254 23468 111318
rect 23392 111046 23468 111254
rect 23392 111014 23398 111046
rect 23190 110982 23191 111014
rect 23125 110981 23191 110982
rect 23397 110982 23398 111014
rect 23462 111014 23468 111046
rect 195024 111318 195100 111324
rect 195024 111254 195030 111318
rect 195094 111254 195100 111318
rect 195437 111318 195503 111319
rect 195437 111286 195438 111318
rect 195024 111046 195100 111254
rect 195024 111014 195030 111046
rect 23462 110982 23463 111014
rect 23397 110981 23463 110982
rect 195029 110982 195030 111014
rect 195094 111014 195100 111046
rect 195432 111254 195438 111286
rect 195502 111286 195503 111318
rect 196389 111318 196455 111319
rect 196389 111286 196390 111318
rect 195502 111254 195508 111286
rect 195432 111046 195508 111254
rect 195094 110982 195095 111014
rect 195029 110981 195095 110982
rect 195432 110982 195438 111046
rect 195502 110982 195508 111046
rect 195432 110976 195508 110982
rect 196384 111254 196390 111286
rect 196454 111286 196455 111318
rect 196792 111318 196868 111324
rect 196454 111254 196460 111286
rect 196384 111046 196460 111254
rect 196384 110982 196390 111046
rect 196454 110982 196460 111046
rect 196792 111254 196798 111318
rect 196862 111254 196868 111318
rect 196792 111046 196868 111254
rect 196792 111014 196798 111046
rect 196384 110976 196460 110982
rect 196797 110982 196798 111014
rect 196862 111014 196868 111046
rect 196862 110982 196863 111014
rect 196797 110981 196863 110982
rect 21760 110910 21836 110916
rect 21760 110846 21766 110910
rect 21830 110846 21836 110910
rect 22173 110910 22239 110911
rect 22173 110878 22174 110910
rect 21760 110638 21836 110846
rect 21760 110606 21766 110638
rect 21765 110574 21766 110606
rect 21830 110606 21836 110638
rect 22168 110846 22174 110878
rect 22238 110878 22239 110910
rect 22581 110910 22647 110911
rect 22581 110878 22582 110910
rect 22238 110846 22244 110878
rect 22168 110638 22244 110846
rect 21830 110574 21831 110606
rect 21765 110573 21831 110574
rect 22168 110574 22174 110638
rect 22238 110574 22244 110638
rect 22168 110568 22244 110574
rect 22576 110846 22582 110878
rect 22646 110878 22647 110910
rect 23120 110910 23196 110916
rect 22646 110846 22652 110878
rect 22576 110638 22652 110846
rect 22576 110574 22582 110638
rect 22646 110574 22652 110638
rect 23120 110846 23126 110910
rect 23190 110846 23196 110910
rect 23120 110638 23196 110846
rect 23120 110606 23126 110638
rect 22576 110568 22652 110574
rect 23125 110574 23126 110606
rect 23190 110606 23196 110638
rect 23528 110910 23604 110916
rect 23528 110846 23534 110910
rect 23598 110846 23604 110910
rect 195165 110910 195231 110911
rect 195165 110878 195166 110910
rect 23528 110638 23604 110846
rect 23528 110606 23534 110638
rect 23190 110574 23191 110606
rect 23125 110573 23191 110574
rect 23533 110574 23534 110606
rect 23598 110606 23604 110638
rect 195160 110846 195166 110878
rect 195230 110878 195231 110910
rect 195568 110910 195644 110916
rect 195230 110846 195236 110878
rect 195160 110638 195236 110846
rect 23598 110574 23599 110606
rect 23533 110573 23599 110574
rect 195160 110574 195166 110638
rect 195230 110574 195236 110638
rect 195568 110846 195574 110910
rect 195638 110846 195644 110910
rect 195568 110638 195644 110846
rect 195568 110606 195574 110638
rect 195160 110568 195236 110574
rect 195573 110574 195574 110606
rect 195638 110606 195644 110638
rect 196248 110910 196324 110916
rect 196248 110846 196254 110910
rect 196318 110846 196324 110910
rect 196661 110910 196727 110911
rect 196661 110878 196662 110910
rect 196248 110638 196324 110846
rect 196248 110606 196254 110638
rect 195638 110574 195639 110606
rect 195573 110573 195639 110574
rect 196253 110574 196254 110606
rect 196318 110606 196324 110638
rect 196656 110846 196662 110878
rect 196726 110878 196727 110910
rect 196726 110846 196732 110878
rect 196656 110638 196732 110846
rect 196318 110574 196319 110606
rect 196253 110573 196319 110574
rect 196656 110574 196662 110638
rect 196726 110574 196732 110638
rect 196656 110568 196732 110574
rect 22173 110502 22239 110503
rect 22173 110470 22174 110502
rect 22168 110438 22174 110470
rect 22238 110470 22239 110502
rect 22440 110502 22516 110508
rect 22238 110438 22244 110470
rect 22168 110230 22244 110438
rect 22168 110166 22174 110230
rect 22238 110166 22244 110230
rect 22440 110438 22446 110502
rect 22510 110438 22516 110502
rect 23125 110502 23191 110503
rect 23125 110470 23126 110502
rect 22440 110230 22516 110438
rect 22440 110198 22446 110230
rect 22168 110160 22244 110166
rect 22445 110166 22446 110198
rect 22510 110198 22516 110230
rect 23120 110438 23126 110470
rect 23190 110470 23191 110502
rect 23533 110502 23599 110503
rect 23533 110470 23534 110502
rect 23190 110438 23196 110470
rect 23120 110230 23196 110438
rect 22510 110166 22511 110198
rect 22445 110165 22511 110166
rect 23120 110166 23126 110230
rect 23190 110166 23196 110230
rect 23120 110160 23196 110166
rect 23528 110438 23534 110470
rect 23598 110470 23599 110502
rect 195165 110502 195231 110503
rect 195165 110470 195166 110502
rect 23598 110438 23604 110470
rect 23528 110230 23604 110438
rect 195160 110438 195166 110470
rect 195230 110470 195231 110502
rect 195432 110502 195508 110508
rect 195230 110438 195236 110470
rect 23528 110166 23534 110230
rect 23598 110166 23604 110230
rect 23528 110160 23604 110166
rect 190264 110366 190340 110372
rect 190264 110302 190270 110366
rect 190334 110302 190340 110366
rect 22440 110094 22516 110100
rect 22440 110030 22446 110094
rect 22510 110030 22516 110094
rect 22440 109822 22516 110030
rect 22440 109790 22446 109822
rect 22445 109758 22446 109790
rect 22510 109790 22516 109822
rect 22984 110094 23060 110100
rect 22984 110030 22990 110094
rect 23054 110030 23060 110094
rect 23397 110094 23463 110095
rect 23397 110062 23398 110094
rect 22984 109822 23060 110030
rect 22984 109790 22990 109822
rect 22510 109758 22511 109790
rect 22445 109757 22511 109758
rect 22989 109758 22990 109790
rect 23054 109790 23060 109822
rect 23392 110030 23398 110062
rect 23462 110062 23463 110094
rect 190133 110094 190199 110095
rect 190133 110062 190134 110094
rect 23462 110030 23468 110062
rect 23392 109822 23468 110030
rect 23054 109758 23055 109790
rect 22989 109757 23055 109758
rect 23392 109758 23398 109822
rect 23462 109758 23468 109822
rect 23392 109752 23468 109758
rect 190128 110030 190134 110062
rect 190198 110062 190199 110094
rect 190264 110094 190340 110302
rect 195160 110230 195236 110438
rect 195160 110166 195166 110230
rect 195230 110166 195236 110230
rect 195432 110438 195438 110502
rect 195502 110438 195508 110502
rect 195845 110502 195911 110503
rect 195845 110470 195846 110502
rect 195432 110230 195508 110438
rect 195432 110198 195438 110230
rect 195160 110160 195236 110166
rect 195437 110166 195438 110198
rect 195502 110198 195508 110230
rect 195840 110438 195846 110470
rect 195910 110470 195911 110502
rect 195910 110438 195916 110470
rect 195840 110230 195916 110438
rect 195502 110166 195503 110198
rect 195437 110165 195503 110166
rect 195840 110166 195846 110230
rect 195910 110166 195916 110230
rect 195840 110160 195916 110166
rect 190264 110062 190270 110094
rect 190198 110030 190204 110062
rect 952 109622 1230 109686
rect 1294 109622 1300 109686
rect 22581 109686 22647 109687
rect 22581 109654 22582 109686
rect 952 108190 1300 109622
rect 22576 109622 22582 109654
rect 22646 109654 22647 109686
rect 22989 109686 23055 109687
rect 22989 109654 22990 109686
rect 22646 109622 22652 109654
rect 21765 109414 21831 109415
rect 21765 109382 21766 109414
rect 21760 109350 21766 109382
rect 21830 109382 21831 109414
rect 22576 109414 22652 109622
rect 21830 109350 21836 109382
rect 21760 109142 21836 109350
rect 22576 109350 22582 109414
rect 22646 109350 22652 109414
rect 22576 109344 22652 109350
rect 22984 109622 22990 109654
rect 23054 109654 23055 109686
rect 23528 109686 23604 109692
rect 23054 109622 23060 109654
rect 22984 109414 23060 109622
rect 22984 109350 22990 109414
rect 23054 109350 23060 109414
rect 23528 109622 23534 109686
rect 23598 109622 23604 109686
rect 23528 109414 23604 109622
rect 190128 109686 190204 110030
rect 190269 110030 190270 110062
rect 190334 110062 190340 110094
rect 195029 110094 195095 110095
rect 195029 110062 195030 110094
rect 190334 110030 190335 110062
rect 190269 110029 190335 110030
rect 195024 110030 195030 110062
rect 195094 110062 195095 110094
rect 195573 110094 195639 110095
rect 195573 110062 195574 110094
rect 195094 110030 195100 110062
rect 195024 109822 195100 110030
rect 195024 109758 195030 109822
rect 195094 109758 195100 109822
rect 195024 109752 195100 109758
rect 195568 110030 195574 110062
rect 195638 110062 195639 110094
rect 195638 110030 195644 110062
rect 195568 109822 195644 110030
rect 195568 109758 195574 109822
rect 195638 109758 195644 109822
rect 195568 109752 195644 109758
rect 217464 109822 217812 111390
rect 217464 109758 217470 109822
rect 217534 109758 217812 109822
rect 190128 109622 190134 109686
rect 190198 109622 190204 109686
rect 190128 109616 190204 109622
rect 195160 109686 195236 109692
rect 195160 109622 195166 109686
rect 195230 109622 195236 109686
rect 23528 109382 23534 109414
rect 22984 109344 23060 109350
rect 23533 109350 23534 109382
rect 23598 109382 23604 109414
rect 190264 109550 190340 109556
rect 190264 109486 190270 109550
rect 190334 109486 190340 109550
rect 23598 109350 23599 109382
rect 23533 109349 23599 109350
rect 190264 109278 190340 109486
rect 195160 109414 195236 109622
rect 195160 109382 195166 109414
rect 195165 109350 195166 109382
rect 195230 109382 195236 109414
rect 195568 109686 195644 109692
rect 195568 109622 195574 109686
rect 195638 109622 195644 109686
rect 196117 109686 196183 109687
rect 196117 109654 196118 109686
rect 195568 109414 195644 109622
rect 195568 109382 195574 109414
rect 195230 109350 195231 109382
rect 195165 109349 195231 109350
rect 195573 109350 195574 109382
rect 195638 109382 195644 109414
rect 196112 109622 196118 109654
rect 196182 109654 196183 109686
rect 196182 109622 196188 109654
rect 196112 109414 196188 109622
rect 195638 109350 195639 109382
rect 195573 109349 195639 109350
rect 196112 109350 196118 109414
rect 196182 109350 196188 109414
rect 196112 109344 196188 109350
rect 196792 109414 196868 109420
rect 196792 109350 196798 109414
rect 196862 109350 196868 109414
rect 190264 109246 190270 109278
rect 190269 109214 190270 109246
rect 190334 109246 190340 109278
rect 190334 109214 190335 109246
rect 190269 109213 190335 109214
rect 21760 109078 21766 109142
rect 21830 109078 21836 109142
rect 21760 109072 21836 109078
rect 28424 109142 28500 109148
rect 28424 109078 28430 109142
rect 28494 109078 28500 109142
rect 190269 109142 190335 109143
rect 190269 109110 190270 109142
rect 21760 109006 21836 109012
rect 21760 108942 21766 109006
rect 21830 108942 21836 109006
rect 22445 109006 22511 109007
rect 22445 108974 22446 109006
rect 21760 108734 21836 108942
rect 21760 108702 21766 108734
rect 21765 108670 21766 108702
rect 21830 108702 21836 108734
rect 22440 108942 22446 108974
rect 22510 108974 22511 109006
rect 22510 108942 22516 108974
rect 22440 108734 22516 108942
rect 28424 108870 28500 109078
rect 28424 108838 28430 108870
rect 28429 108806 28430 108838
rect 28494 108838 28500 108870
rect 190264 109078 190270 109110
rect 190334 109110 190335 109142
rect 196792 109142 196868 109350
rect 196792 109110 196798 109142
rect 190334 109078 190340 109110
rect 190264 108870 190340 109078
rect 196797 109078 196798 109110
rect 196862 109110 196868 109142
rect 196862 109078 196863 109110
rect 196797 109077 196863 109078
rect 28494 108806 28495 108838
rect 28429 108805 28495 108806
rect 190264 108806 190270 108870
rect 190334 108806 190340 108870
rect 190264 108800 190340 108806
rect 196112 109006 196188 109012
rect 196112 108942 196118 109006
rect 196182 108942 196188 109006
rect 196797 109006 196863 109007
rect 196797 108974 196798 109006
rect 21830 108670 21831 108702
rect 21765 108669 21831 108670
rect 22440 108670 22446 108734
rect 22510 108670 22516 108734
rect 22440 108664 22516 108670
rect 28288 108734 28364 108740
rect 28288 108670 28294 108734
rect 28358 108670 28364 108734
rect 21760 108598 21836 108604
rect 21760 108534 21766 108598
rect 21830 108534 21836 108598
rect 21760 108326 21836 108534
rect 28288 108462 28364 108670
rect 28288 108430 28294 108462
rect 28293 108398 28294 108430
rect 28358 108430 28364 108462
rect 190128 108734 190204 108740
rect 190128 108670 190134 108734
rect 190198 108670 190204 108734
rect 196112 108734 196188 108942
rect 196112 108702 196118 108734
rect 190128 108462 190204 108670
rect 196117 108670 196118 108702
rect 196182 108702 196188 108734
rect 196792 108942 196798 108974
rect 196862 108974 196863 109006
rect 196862 108942 196868 108974
rect 196792 108734 196868 108942
rect 196182 108670 196183 108702
rect 196117 108669 196183 108670
rect 196792 108670 196798 108734
rect 196862 108670 196868 108734
rect 196792 108664 196868 108670
rect 196656 108598 196732 108604
rect 196656 108534 196662 108598
rect 196726 108534 196732 108598
rect 190128 108430 190134 108462
rect 28358 108398 28359 108430
rect 28293 108397 28359 108398
rect 190133 108398 190134 108430
rect 190198 108430 190204 108462
rect 196112 108462 196324 108468
rect 190198 108398 190199 108430
rect 190133 108397 190199 108398
rect 196112 108398 196254 108462
rect 196318 108398 196324 108462
rect 196112 108392 196324 108398
rect 21760 108294 21766 108326
rect 21765 108262 21766 108294
rect 21830 108294 21836 108326
rect 190128 108326 190204 108332
rect 21830 108262 21831 108294
rect 21765 108261 21831 108262
rect 190128 108262 190134 108326
rect 190198 108262 190204 108326
rect 196112 108326 196188 108392
rect 196112 108294 196118 108326
rect 952 108126 1230 108190
rect 1294 108126 1300 108190
rect 952 106422 1300 108126
rect 21896 108190 21972 108196
rect 21896 108126 21902 108190
rect 21966 108126 21972 108190
rect 22717 108190 22783 108191
rect 22717 108158 22718 108190
rect 21896 107918 21972 108126
rect 21896 107886 21902 107918
rect 21901 107854 21902 107886
rect 21966 107886 21972 107918
rect 22712 108126 22718 108158
rect 22782 108158 22783 108190
rect 23120 108190 23196 108196
rect 22782 108126 22788 108158
rect 22712 107918 22788 108126
rect 21966 107854 21967 107886
rect 21901 107853 21967 107854
rect 22712 107854 22718 107918
rect 22782 107854 22788 107918
rect 23120 108126 23126 108190
rect 23190 108126 23196 108190
rect 23120 107918 23196 108126
rect 23120 107886 23126 107918
rect 22712 107848 22788 107854
rect 23125 107854 23126 107886
rect 23190 107886 23196 107918
rect 23392 108190 23468 108196
rect 23392 108126 23398 108190
rect 23462 108126 23468 108190
rect 23392 107918 23468 108126
rect 23392 107886 23398 107918
rect 23190 107854 23191 107886
rect 23125 107853 23191 107854
rect 23397 107854 23398 107886
rect 23462 107886 23468 107918
rect 28424 107918 28500 107924
rect 23462 107854 23463 107886
rect 23397 107853 23463 107854
rect 28424 107854 28430 107918
rect 28494 107854 28500 107918
rect 190128 107918 190204 108262
rect 196117 108262 196118 108294
rect 196182 108294 196188 108326
rect 196656 108326 196732 108534
rect 196656 108294 196662 108326
rect 196182 108262 196183 108294
rect 196117 108261 196183 108262
rect 196661 108262 196662 108294
rect 196726 108294 196732 108326
rect 196726 108262 196727 108294
rect 196661 108261 196727 108262
rect 195029 108190 195095 108191
rect 195029 108158 195030 108190
rect 195024 108126 195030 108158
rect 195094 108158 195095 108190
rect 195437 108190 195503 108191
rect 195437 108158 195438 108190
rect 195094 108126 195100 108158
rect 190128 107886 190134 107918
rect 21901 107782 21967 107783
rect 21901 107750 21902 107782
rect 21896 107718 21902 107750
rect 21966 107750 21967 107782
rect 22445 107782 22511 107783
rect 22445 107750 22446 107782
rect 21966 107718 21972 107750
rect 21896 107510 21972 107718
rect 21896 107446 21902 107510
rect 21966 107446 21972 107510
rect 21896 107440 21972 107446
rect 22440 107718 22446 107750
rect 22510 107750 22511 107782
rect 22984 107782 23060 107788
rect 22510 107718 22516 107750
rect 22440 107510 22516 107718
rect 22440 107446 22446 107510
rect 22510 107446 22516 107510
rect 22984 107718 22990 107782
rect 23054 107718 23060 107782
rect 23397 107782 23463 107783
rect 23397 107750 23398 107782
rect 22984 107510 23060 107718
rect 22984 107478 22990 107510
rect 22440 107440 22516 107446
rect 22989 107446 22990 107478
rect 23054 107478 23060 107510
rect 23392 107718 23398 107750
rect 23462 107750 23463 107782
rect 23462 107718 23468 107750
rect 23392 107510 23468 107718
rect 28424 107646 28500 107854
rect 190133 107854 190134 107886
rect 190198 107886 190204 107918
rect 190269 107918 190335 107919
rect 190269 107886 190270 107918
rect 190198 107854 190199 107886
rect 190133 107853 190199 107854
rect 190264 107854 190270 107886
rect 190334 107886 190335 107918
rect 195024 107918 195100 108126
rect 190334 107854 190340 107886
rect 28424 107614 28430 107646
rect 28429 107582 28430 107614
rect 28494 107614 28500 107646
rect 190264 107646 190340 107854
rect 195024 107854 195030 107918
rect 195094 107854 195100 107918
rect 195024 107848 195100 107854
rect 195432 108126 195438 108158
rect 195502 108158 195503 108190
rect 196112 108190 196188 108196
rect 195502 108126 195508 108158
rect 195432 107918 195508 108126
rect 195432 107854 195438 107918
rect 195502 107854 195508 107918
rect 196112 108126 196118 108190
rect 196182 108126 196188 108190
rect 196112 107918 196188 108126
rect 196112 107886 196118 107918
rect 195432 107848 195508 107854
rect 196117 107854 196118 107886
rect 196182 107886 196188 107918
rect 196792 108190 196868 108196
rect 196792 108126 196798 108190
rect 196862 108126 196868 108190
rect 196792 107918 196868 108126
rect 196792 107886 196798 107918
rect 196182 107854 196183 107886
rect 196117 107853 196183 107854
rect 196797 107854 196798 107886
rect 196862 107886 196868 107918
rect 217464 108190 217812 109758
rect 217464 108126 217470 108190
rect 217534 108126 217812 108190
rect 196862 107854 196863 107886
rect 196797 107853 196863 107854
rect 28494 107582 28495 107614
rect 28429 107581 28495 107582
rect 190264 107582 190270 107646
rect 190334 107582 190340 107646
rect 190264 107576 190340 107582
rect 195160 107782 195236 107788
rect 195160 107718 195166 107782
rect 195230 107718 195236 107782
rect 195573 107782 195639 107783
rect 195573 107750 195574 107782
rect 23054 107446 23055 107478
rect 22989 107445 23055 107446
rect 23392 107446 23398 107510
rect 23462 107446 23468 107510
rect 195160 107510 195236 107718
rect 195160 107478 195166 107510
rect 23392 107440 23468 107446
rect 195165 107446 195166 107478
rect 195230 107478 195236 107510
rect 195568 107718 195574 107750
rect 195638 107750 195639 107782
rect 196389 107782 196455 107783
rect 196389 107750 196390 107782
rect 195638 107718 195644 107750
rect 195568 107510 195644 107718
rect 195230 107446 195231 107478
rect 195165 107445 195231 107446
rect 195568 107446 195574 107510
rect 195638 107446 195644 107510
rect 195568 107440 195644 107446
rect 196384 107718 196390 107750
rect 196454 107750 196455 107782
rect 196797 107782 196863 107783
rect 196797 107750 196798 107782
rect 196454 107718 196460 107750
rect 196384 107510 196460 107718
rect 196384 107446 196390 107510
rect 196454 107446 196460 107510
rect 196384 107440 196460 107446
rect 196792 107718 196798 107750
rect 196862 107750 196863 107782
rect 196862 107718 196868 107750
rect 196792 107510 196868 107718
rect 196792 107446 196798 107510
rect 196862 107446 196868 107510
rect 196792 107440 196868 107446
rect 21896 107374 21972 107380
rect 21896 107310 21902 107374
rect 21966 107310 21972 107374
rect 22173 107374 22239 107375
rect 22173 107342 22174 107374
rect 21896 107102 21972 107310
rect 21896 107070 21902 107102
rect 21901 107038 21902 107070
rect 21966 107070 21972 107102
rect 22168 107310 22174 107342
rect 22238 107342 22239 107374
rect 22581 107374 22647 107375
rect 22581 107342 22582 107374
rect 22238 107310 22244 107342
rect 22168 107102 22244 107310
rect 21966 107038 21967 107070
rect 21901 107037 21967 107038
rect 22168 107038 22174 107102
rect 22238 107038 22244 107102
rect 22168 107032 22244 107038
rect 22576 107310 22582 107342
rect 22646 107342 22647 107374
rect 22989 107374 23055 107375
rect 22989 107342 22990 107374
rect 22646 107310 22652 107342
rect 22576 107102 22652 107310
rect 22576 107038 22582 107102
rect 22646 107038 22652 107102
rect 22576 107032 22652 107038
rect 22984 107310 22990 107342
rect 23054 107342 23055 107374
rect 23392 107374 23468 107380
rect 23054 107310 23060 107342
rect 22984 107102 23060 107310
rect 22984 107038 22990 107102
rect 23054 107038 23060 107102
rect 23392 107310 23398 107374
rect 23462 107310 23468 107374
rect 23392 107102 23468 107310
rect 23392 107070 23398 107102
rect 22984 107032 23060 107038
rect 23397 107038 23398 107070
rect 23462 107070 23468 107102
rect 195024 107374 195100 107380
rect 195024 107310 195030 107374
rect 195094 107310 195100 107374
rect 195024 107102 195100 107310
rect 195024 107070 195030 107102
rect 23462 107038 23463 107070
rect 23397 107037 23463 107038
rect 195029 107038 195030 107070
rect 195094 107070 195100 107102
rect 195432 107374 195508 107380
rect 195432 107310 195438 107374
rect 195502 107310 195508 107374
rect 195432 107102 195508 107310
rect 195432 107070 195438 107102
rect 195094 107038 195095 107070
rect 195029 107037 195095 107038
rect 195437 107038 195438 107070
rect 195502 107070 195508 107102
rect 195976 107374 196052 107380
rect 195976 107310 195982 107374
rect 196046 107310 196052 107374
rect 196253 107374 196319 107375
rect 196253 107342 196254 107374
rect 195976 107102 196052 107310
rect 195976 107070 195982 107102
rect 195502 107038 195503 107070
rect 195437 107037 195503 107038
rect 195981 107038 195982 107070
rect 196046 107070 196052 107102
rect 196248 107310 196254 107342
rect 196318 107342 196319 107374
rect 196792 107374 196868 107380
rect 196318 107310 196324 107342
rect 196248 107102 196324 107310
rect 196046 107038 196047 107070
rect 195981 107037 196047 107038
rect 196248 107038 196254 107102
rect 196318 107038 196324 107102
rect 196792 107310 196798 107374
rect 196862 107310 196868 107374
rect 196792 107102 196868 107310
rect 196792 107070 196798 107102
rect 196248 107032 196324 107038
rect 196797 107038 196798 107070
rect 196862 107070 196868 107102
rect 196862 107038 196863 107070
rect 196797 107037 196863 107038
rect 21896 106966 21972 106972
rect 21896 106902 21902 106966
rect 21966 106902 21972 106966
rect 22309 106966 22375 106967
rect 22309 106934 22310 106966
rect 21896 106694 21972 106902
rect 21896 106662 21902 106694
rect 21901 106630 21902 106662
rect 21966 106662 21972 106694
rect 22304 106902 22310 106934
rect 22374 106934 22375 106966
rect 23120 106966 23196 106972
rect 22374 106902 22380 106934
rect 22304 106694 22380 106902
rect 21966 106630 21967 106662
rect 21901 106629 21967 106630
rect 22304 106630 22310 106694
rect 22374 106630 22380 106694
rect 23120 106902 23126 106966
rect 23190 106902 23196 106966
rect 23397 106966 23463 106967
rect 23397 106934 23398 106966
rect 23120 106694 23196 106902
rect 23120 106662 23126 106694
rect 22304 106624 22380 106630
rect 23125 106630 23126 106662
rect 23190 106662 23196 106694
rect 23392 106902 23398 106934
rect 23462 106934 23463 106966
rect 195029 106966 195095 106967
rect 195029 106934 195030 106966
rect 23462 106902 23468 106934
rect 23392 106694 23468 106902
rect 23190 106630 23191 106662
rect 23125 106629 23191 106630
rect 23392 106630 23398 106694
rect 23462 106630 23468 106694
rect 23392 106624 23468 106630
rect 195024 106902 195030 106934
rect 195094 106934 195095 106966
rect 195437 106966 195503 106967
rect 195437 106934 195438 106966
rect 195094 106902 195100 106934
rect 195024 106694 195100 106902
rect 195024 106630 195030 106694
rect 195094 106630 195100 106694
rect 195024 106624 195100 106630
rect 195432 106902 195438 106934
rect 195502 106934 195503 106966
rect 196117 106966 196183 106967
rect 196117 106934 196118 106966
rect 195502 106902 195508 106934
rect 195432 106694 195508 106902
rect 195432 106630 195438 106694
rect 195502 106630 195508 106694
rect 195432 106624 195508 106630
rect 196112 106902 196118 106934
rect 196182 106934 196183 106966
rect 196797 106966 196863 106967
rect 196797 106934 196798 106966
rect 196182 106902 196188 106934
rect 196112 106694 196188 106902
rect 196112 106630 196118 106694
rect 196182 106630 196188 106694
rect 196112 106624 196188 106630
rect 196792 106902 196798 106934
rect 196862 106934 196863 106966
rect 196862 106902 196868 106934
rect 196792 106694 196868 106902
rect 196792 106630 196798 106694
rect 196862 106630 196868 106694
rect 196792 106624 196868 106630
rect 952 106358 1230 106422
rect 1294 106358 1300 106422
rect 952 104790 1300 106358
rect 22168 106558 22244 106564
rect 22168 106494 22174 106558
rect 22238 106494 22244 106558
rect 22168 106286 22244 106494
rect 22168 106254 22174 106286
rect 22173 106222 22174 106254
rect 22238 106254 22244 106286
rect 23120 106558 23196 106564
rect 23120 106494 23126 106558
rect 23190 106494 23196 106558
rect 23533 106558 23599 106559
rect 23533 106526 23534 106558
rect 23120 106286 23196 106494
rect 23120 106254 23126 106286
rect 22238 106222 22239 106254
rect 22173 106221 22239 106222
rect 23125 106222 23126 106254
rect 23190 106254 23196 106286
rect 23528 106494 23534 106526
rect 23598 106526 23599 106558
rect 195160 106558 195236 106564
rect 23598 106494 23604 106526
rect 23528 106286 23604 106494
rect 23190 106222 23191 106254
rect 23125 106221 23191 106222
rect 23528 106222 23534 106286
rect 23598 106222 23604 106286
rect 195160 106494 195166 106558
rect 195230 106494 195236 106558
rect 195160 106286 195236 106494
rect 195160 106254 195166 106286
rect 23528 106216 23604 106222
rect 195165 106222 195166 106254
rect 195230 106254 195236 106286
rect 195568 106558 195644 106564
rect 195568 106494 195574 106558
rect 195638 106494 195644 106558
rect 195568 106286 195644 106494
rect 195568 106254 195574 106286
rect 195230 106222 195231 106254
rect 195165 106221 195231 106222
rect 195573 106222 195574 106254
rect 195638 106254 195644 106286
rect 195840 106558 195916 106564
rect 195840 106494 195846 106558
rect 195910 106494 195916 106558
rect 195840 106286 195916 106494
rect 195840 106254 195846 106286
rect 195638 106222 195639 106254
rect 195573 106221 195639 106222
rect 195845 106222 195846 106254
rect 195910 106254 195916 106286
rect 196248 106558 196324 106564
rect 196248 106494 196254 106558
rect 196318 106494 196324 106558
rect 196248 106286 196324 106494
rect 196248 106254 196254 106286
rect 195910 106222 195911 106254
rect 195845 106221 195911 106222
rect 196253 106222 196254 106254
rect 196318 106254 196324 106286
rect 217464 106286 217812 108126
rect 196318 106222 196319 106254
rect 196253 106221 196319 106222
rect 217464 106222 217470 106286
rect 217534 106222 217812 106286
rect 23120 106150 23196 106156
rect 23120 106086 23126 106150
rect 23190 106086 23196 106150
rect 23533 106150 23599 106151
rect 23533 106118 23534 106150
rect 23120 105878 23196 106086
rect 23120 105846 23126 105878
rect 23125 105814 23126 105846
rect 23190 105846 23196 105878
rect 23528 106086 23534 106118
rect 23598 106118 23599 106150
rect 195165 106150 195231 106151
rect 195165 106118 195166 106150
rect 23598 106086 23604 106118
rect 23528 105878 23604 106086
rect 23190 105814 23191 105846
rect 23125 105813 23191 105814
rect 23528 105814 23534 105878
rect 23598 105814 23604 105878
rect 23528 105808 23604 105814
rect 195160 106086 195166 106118
rect 195230 106118 195231 106150
rect 195568 106150 195644 106156
rect 195230 106086 195236 106118
rect 195160 105878 195236 106086
rect 195160 105814 195166 105878
rect 195230 105814 195236 105878
rect 195568 106086 195574 106150
rect 195638 106086 195644 106150
rect 195568 105878 195644 106086
rect 195568 105846 195574 105878
rect 195160 105808 195236 105814
rect 195573 105814 195574 105846
rect 195638 105846 195644 105878
rect 195638 105814 195639 105846
rect 195573 105813 195639 105814
rect 22168 105742 22244 105748
rect 22168 105678 22174 105742
rect 22238 105678 22244 105742
rect 21760 105470 21836 105476
rect 21760 105406 21766 105470
rect 21830 105406 21836 105470
rect 22168 105470 22244 105678
rect 22168 105438 22174 105470
rect 21760 105198 21836 105406
rect 22173 105406 22174 105438
rect 22238 105438 22244 105470
rect 22576 105742 22652 105748
rect 22576 105678 22582 105742
rect 22646 105678 22652 105742
rect 23125 105742 23191 105743
rect 23125 105710 23126 105742
rect 22576 105470 22652 105678
rect 22576 105438 22582 105470
rect 22238 105406 22239 105438
rect 22173 105405 22239 105406
rect 22581 105406 22582 105438
rect 22646 105438 22652 105470
rect 23120 105678 23126 105710
rect 23190 105710 23191 105742
rect 23528 105742 23604 105748
rect 23190 105678 23196 105710
rect 23120 105470 23196 105678
rect 22646 105406 22647 105438
rect 22581 105405 22647 105406
rect 23120 105406 23126 105470
rect 23190 105406 23196 105470
rect 23528 105678 23534 105742
rect 23598 105678 23604 105742
rect 23528 105470 23604 105678
rect 195160 105742 195236 105748
rect 195160 105678 195166 105742
rect 195230 105678 195236 105742
rect 28565 105606 28631 105607
rect 28565 105574 28566 105606
rect 23528 105438 23534 105470
rect 23120 105400 23196 105406
rect 23533 105406 23534 105438
rect 23598 105438 23604 105470
rect 28560 105542 28566 105574
rect 28630 105574 28631 105606
rect 190269 105606 190335 105607
rect 190269 105574 190270 105606
rect 28630 105542 28636 105574
rect 23598 105406 23599 105438
rect 23533 105405 23599 105406
rect 28560 105334 28636 105542
rect 28560 105270 28566 105334
rect 28630 105270 28636 105334
rect 28560 105264 28636 105270
rect 190264 105542 190270 105574
rect 190334 105574 190335 105606
rect 190334 105542 190340 105574
rect 190264 105334 190340 105542
rect 195160 105470 195236 105678
rect 195160 105438 195166 105470
rect 195165 105406 195166 105438
rect 195230 105438 195236 105470
rect 195432 105742 195508 105748
rect 195432 105678 195438 105742
rect 195502 105678 195508 105742
rect 195432 105470 195508 105678
rect 195432 105438 195438 105470
rect 195230 105406 195231 105438
rect 195165 105405 195231 105406
rect 195437 105406 195438 105438
rect 195502 105438 195508 105470
rect 196248 105742 196324 105748
rect 196248 105678 196254 105742
rect 196318 105678 196324 105742
rect 196248 105470 196324 105678
rect 196248 105438 196254 105470
rect 195502 105406 195503 105438
rect 195437 105405 195503 105406
rect 196253 105406 196254 105438
rect 196318 105438 196324 105470
rect 196656 105470 196732 105476
rect 196318 105406 196319 105438
rect 196253 105405 196319 105406
rect 196656 105406 196662 105470
rect 196726 105406 196732 105470
rect 190264 105270 190270 105334
rect 190334 105270 190340 105334
rect 190264 105264 190340 105270
rect 21760 105166 21766 105198
rect 21765 105134 21766 105166
rect 21830 105166 21836 105198
rect 28429 105198 28495 105199
rect 28429 105166 28430 105198
rect 21830 105134 21831 105166
rect 21765 105133 21831 105134
rect 28424 105134 28430 105166
rect 28494 105166 28495 105198
rect 190264 105198 190340 105204
rect 28494 105134 28500 105166
rect 21765 105062 21831 105063
rect 21765 105030 21766 105062
rect 952 104726 1230 104790
rect 1294 104726 1300 104790
rect 952 103158 1300 104726
rect 21760 104998 21766 105030
rect 21830 105030 21831 105062
rect 22440 105062 22516 105068
rect 21830 104998 21836 105030
rect 21760 104790 21836 104998
rect 21760 104726 21766 104790
rect 21830 104726 21836 104790
rect 22440 104998 22446 105062
rect 22510 104998 22516 105062
rect 22581 105062 22647 105063
rect 22581 105030 22582 105062
rect 22440 104790 22516 104998
rect 22440 104758 22446 104790
rect 21760 104720 21836 104726
rect 22445 104726 22446 104758
rect 22510 104758 22516 104790
rect 22576 104998 22582 105030
rect 22646 105030 22647 105062
rect 22646 104998 22652 105030
rect 22576 104790 22652 104998
rect 28424 104926 28500 105134
rect 28424 104862 28430 104926
rect 28494 104862 28500 104926
rect 190264 105134 190270 105198
rect 190334 105134 190340 105198
rect 196656 105198 196732 105406
rect 196656 105166 196662 105198
rect 190264 104926 190340 105134
rect 196661 105134 196662 105166
rect 196726 105166 196732 105198
rect 196726 105134 196727 105166
rect 196661 105133 196727 105134
rect 195845 105062 195911 105063
rect 195845 105030 195846 105062
rect 190264 104894 190270 104926
rect 28424 104856 28500 104862
rect 190269 104862 190270 104894
rect 190334 104894 190340 104926
rect 195840 104998 195846 105030
rect 195910 105030 195911 105062
rect 196112 105062 196188 105068
rect 195910 104998 195916 105030
rect 190334 104862 190335 104894
rect 190269 104861 190335 104862
rect 22510 104726 22511 104758
rect 22445 104725 22511 104726
rect 22576 104726 22582 104790
rect 22646 104726 22652 104790
rect 22576 104720 22652 104726
rect 195840 104790 195916 104998
rect 195840 104726 195846 104790
rect 195910 104726 195916 104790
rect 196112 104998 196118 105062
rect 196182 104998 196188 105062
rect 196112 104790 196188 104998
rect 196112 104758 196118 104790
rect 195840 104720 195916 104726
rect 196117 104726 196118 104758
rect 196182 104758 196188 104790
rect 196792 105062 196868 105068
rect 196792 104998 196798 105062
rect 196862 104998 196868 105062
rect 196792 104790 196868 104998
rect 196792 104758 196798 104790
rect 196182 104726 196183 104758
rect 196117 104725 196183 104726
rect 196797 104726 196798 104758
rect 196862 104758 196868 104790
rect 196862 104726 196863 104758
rect 196797 104725 196863 104726
rect 21760 104654 21836 104660
rect 21760 104590 21766 104654
rect 21830 104590 21836 104654
rect 21760 104382 21836 104590
rect 196656 104654 196732 104660
rect 196656 104590 196662 104654
rect 196726 104590 196732 104654
rect 190269 104518 190335 104519
rect 190269 104486 190270 104518
rect 21760 104350 21766 104382
rect 21765 104318 21766 104350
rect 21830 104350 21836 104382
rect 190264 104454 190270 104486
rect 190334 104486 190335 104518
rect 190334 104454 190340 104486
rect 21830 104318 21831 104350
rect 21765 104317 21831 104318
rect 21760 104246 21836 104252
rect 21760 104182 21766 104246
rect 21830 104182 21836 104246
rect 21760 103974 21836 104182
rect 21760 103942 21766 103974
rect 21765 103910 21766 103942
rect 21830 103942 21836 103974
rect 22576 104246 22652 104252
rect 22576 104182 22582 104246
rect 22646 104182 22652 104246
rect 22989 104246 23055 104247
rect 22989 104214 22990 104246
rect 22576 103974 22652 104182
rect 22576 103942 22582 103974
rect 21830 103910 21831 103942
rect 21765 103909 21831 103910
rect 22581 103910 22582 103942
rect 22646 103942 22652 103974
rect 22984 104182 22990 104214
rect 23054 104214 23055 104246
rect 23528 104246 23604 104252
rect 23054 104182 23060 104214
rect 22984 103974 23060 104182
rect 22646 103910 22647 103942
rect 22581 103909 22647 103910
rect 22984 103910 22990 103974
rect 23054 103910 23060 103974
rect 23528 104182 23534 104246
rect 23598 104182 23604 104246
rect 23528 103974 23604 104182
rect 190264 104246 190340 104454
rect 196656 104382 196732 104590
rect 196656 104350 196662 104382
rect 196661 104318 196662 104350
rect 196726 104350 196732 104382
rect 217464 104654 217812 106222
rect 217464 104590 217470 104654
rect 217534 104590 217812 104654
rect 196726 104318 196727 104350
rect 196661 104317 196727 104318
rect 190264 104182 190270 104246
rect 190334 104182 190340 104246
rect 195165 104246 195231 104247
rect 195165 104214 195166 104246
rect 190264 104176 190340 104182
rect 195160 104182 195166 104214
rect 195230 104214 195231 104246
rect 195568 104246 195644 104252
rect 195230 104182 195236 104214
rect 23528 103942 23534 103974
rect 22984 103904 23060 103910
rect 23533 103910 23534 103942
rect 23598 103942 23604 103974
rect 195160 103974 195236 104182
rect 23598 103910 23599 103942
rect 23533 103909 23599 103910
rect 195160 103910 195166 103974
rect 195230 103910 195236 103974
rect 195568 104182 195574 104246
rect 195638 104182 195644 104246
rect 195845 104246 195911 104247
rect 195845 104214 195846 104246
rect 195568 103974 195644 104182
rect 195568 103942 195574 103974
rect 195160 103904 195236 103910
rect 195573 103910 195574 103942
rect 195638 103942 195644 103974
rect 195840 104182 195846 104214
rect 195910 104214 195911 104246
rect 196661 104246 196727 104247
rect 196661 104214 196662 104246
rect 195910 104182 195916 104214
rect 195840 103974 195916 104182
rect 195638 103910 195639 103942
rect 195573 103909 195639 103910
rect 195840 103910 195846 103974
rect 195910 103910 195916 103974
rect 195840 103904 195916 103910
rect 196656 104182 196662 104214
rect 196726 104214 196727 104246
rect 196726 104182 196732 104214
rect 196656 103974 196732 104182
rect 196656 103910 196662 103974
rect 196726 103910 196732 103974
rect 196656 103904 196732 103910
rect 21901 103838 21967 103839
rect 21901 103806 21902 103838
rect 21896 103774 21902 103806
rect 21966 103806 21967 103838
rect 22989 103838 23055 103839
rect 22989 103806 22990 103838
rect 21966 103774 21972 103806
rect 21896 103566 21972 103774
rect 21896 103502 21902 103566
rect 21966 103502 21972 103566
rect 21896 103496 21972 103502
rect 22984 103774 22990 103806
rect 23054 103806 23055 103838
rect 23392 103838 23468 103844
rect 23054 103774 23060 103806
rect 22984 103566 23060 103774
rect 22984 103502 22990 103566
rect 23054 103502 23060 103566
rect 23392 103774 23398 103838
rect 23462 103774 23468 103838
rect 23392 103566 23468 103774
rect 23392 103534 23398 103566
rect 22984 103496 23060 103502
rect 23397 103502 23398 103534
rect 23462 103534 23468 103566
rect 195024 103838 195100 103844
rect 195024 103774 195030 103838
rect 195094 103774 195100 103838
rect 195437 103838 195503 103839
rect 195437 103806 195438 103838
rect 195024 103566 195100 103774
rect 195024 103534 195030 103566
rect 23462 103502 23463 103534
rect 23397 103501 23463 103502
rect 195029 103502 195030 103534
rect 195094 103534 195100 103566
rect 195432 103774 195438 103806
rect 195502 103806 195503 103838
rect 196792 103838 196868 103844
rect 195502 103774 195508 103806
rect 195432 103566 195508 103774
rect 195094 103502 195095 103534
rect 195029 103501 195095 103502
rect 195432 103502 195438 103566
rect 195502 103502 195508 103566
rect 196792 103774 196798 103838
rect 196862 103774 196868 103838
rect 196792 103566 196868 103774
rect 196792 103534 196798 103566
rect 195432 103496 195508 103502
rect 196797 103502 196798 103534
rect 196862 103534 196868 103566
rect 196862 103502 196863 103534
rect 196797 103501 196863 103502
rect 952 103094 1230 103158
rect 1294 103094 1300 103158
rect 21760 103430 21836 103436
rect 21760 103366 21766 103430
rect 21830 103366 21836 103430
rect 22445 103430 22511 103431
rect 22445 103398 22446 103430
rect 21760 103158 21836 103366
rect 21760 103126 21766 103158
rect 952 101254 1300 103094
rect 21765 103094 21766 103126
rect 21830 103126 21836 103158
rect 22440 103366 22446 103398
rect 22510 103398 22511 103430
rect 23120 103430 23196 103436
rect 22510 103366 22516 103398
rect 22440 103158 22516 103366
rect 21830 103094 21831 103126
rect 21765 103093 21831 103094
rect 22440 103094 22446 103158
rect 22510 103094 22516 103158
rect 23120 103366 23126 103430
rect 23190 103366 23196 103430
rect 23397 103430 23463 103431
rect 23397 103398 23398 103430
rect 23120 103158 23196 103366
rect 23120 103126 23126 103158
rect 22440 103088 22516 103094
rect 23125 103094 23126 103126
rect 23190 103126 23196 103158
rect 23392 103366 23398 103398
rect 23462 103398 23463 103430
rect 195160 103430 195236 103436
rect 23462 103366 23468 103398
rect 23392 103158 23468 103366
rect 23190 103094 23191 103126
rect 23125 103093 23191 103094
rect 23392 103094 23398 103158
rect 23462 103094 23468 103158
rect 195160 103366 195166 103430
rect 195230 103366 195236 103430
rect 195573 103430 195639 103431
rect 195573 103398 195574 103430
rect 195160 103158 195236 103366
rect 195160 103126 195166 103158
rect 23392 103088 23468 103094
rect 195165 103094 195166 103126
rect 195230 103126 195236 103158
rect 195568 103366 195574 103398
rect 195638 103398 195639 103430
rect 195840 103430 195916 103436
rect 195638 103366 195644 103398
rect 195568 103158 195644 103366
rect 195230 103094 195231 103126
rect 195165 103093 195231 103094
rect 195568 103094 195574 103158
rect 195638 103094 195644 103158
rect 195840 103366 195846 103430
rect 195910 103366 195916 103430
rect 196797 103430 196863 103431
rect 196797 103398 196798 103430
rect 195840 103158 195916 103366
rect 195840 103126 195846 103158
rect 195568 103088 195644 103094
rect 195845 103094 195846 103126
rect 195910 103126 195916 103158
rect 196792 103366 196798 103398
rect 196862 103398 196863 103430
rect 196862 103366 196868 103398
rect 196792 103158 196868 103366
rect 195910 103094 195911 103126
rect 195845 103093 195911 103094
rect 196792 103094 196798 103158
rect 196862 103094 196868 103158
rect 196792 103088 196868 103094
rect 21896 103022 21972 103028
rect 21896 102958 21902 103022
rect 21966 102958 21972 103022
rect 21896 102750 21972 102958
rect 21896 102718 21902 102750
rect 21901 102686 21902 102718
rect 21966 102718 21972 102750
rect 22304 103022 22380 103028
rect 22304 102958 22310 103022
rect 22374 102958 22380 103022
rect 22304 102750 22380 102958
rect 22304 102718 22310 102750
rect 21966 102686 21967 102718
rect 21901 102685 21967 102686
rect 22309 102686 22310 102718
rect 22374 102718 22380 102750
rect 22712 103022 22788 103028
rect 22712 102958 22718 103022
rect 22782 102958 22788 103022
rect 22712 102750 22788 102958
rect 22712 102718 22718 102750
rect 22374 102686 22375 102718
rect 22309 102685 22375 102686
rect 22717 102686 22718 102718
rect 22782 102718 22788 102750
rect 22984 103022 23060 103028
rect 22984 102958 22990 103022
rect 23054 102958 23060 103022
rect 22984 102750 23060 102958
rect 22984 102718 22990 102750
rect 22782 102686 22783 102718
rect 22717 102685 22783 102686
rect 22989 102686 22990 102718
rect 23054 102718 23060 102750
rect 23392 103022 23468 103028
rect 23392 102958 23398 103022
rect 23462 102958 23468 103022
rect 195165 103022 195231 103023
rect 195165 102990 195166 103022
rect 23392 102750 23468 102958
rect 23392 102718 23398 102750
rect 23054 102686 23055 102718
rect 22989 102685 23055 102686
rect 23397 102686 23398 102718
rect 23462 102718 23468 102750
rect 195160 102958 195166 102990
rect 195230 102990 195231 103022
rect 195432 103022 195508 103028
rect 195230 102958 195236 102990
rect 195160 102750 195236 102958
rect 23462 102686 23463 102718
rect 23397 102685 23463 102686
rect 195160 102686 195166 102750
rect 195230 102686 195236 102750
rect 195432 102958 195438 103022
rect 195502 102958 195508 103022
rect 195432 102750 195508 102958
rect 195432 102718 195438 102750
rect 195160 102680 195236 102686
rect 195437 102686 195438 102718
rect 195502 102718 195508 102750
rect 196792 103022 196868 103028
rect 196792 102958 196798 103022
rect 196862 102958 196868 103022
rect 196792 102750 196868 102958
rect 196792 102718 196798 102750
rect 195502 102686 195503 102718
rect 195437 102685 195503 102686
rect 196797 102686 196798 102718
rect 196862 102718 196868 102750
rect 217464 103022 217812 104590
rect 217464 102958 217470 103022
rect 217534 102958 217812 103022
rect 196862 102686 196863 102718
rect 196797 102685 196863 102686
rect 22445 102614 22511 102615
rect 22445 102582 22446 102614
rect 22440 102550 22446 102582
rect 22510 102582 22511 102614
rect 22989 102614 23055 102615
rect 22989 102582 22990 102614
rect 22510 102550 22516 102582
rect 22440 102342 22516 102550
rect 22440 102278 22446 102342
rect 22510 102278 22516 102342
rect 22440 102272 22516 102278
rect 22984 102550 22990 102582
rect 23054 102582 23055 102614
rect 23397 102614 23463 102615
rect 23397 102582 23398 102614
rect 23054 102550 23060 102582
rect 22984 102342 23060 102550
rect 22984 102278 22990 102342
rect 23054 102278 23060 102342
rect 22984 102272 23060 102278
rect 23392 102550 23398 102582
rect 23462 102582 23463 102614
rect 195024 102614 195100 102620
rect 23462 102550 23468 102582
rect 23392 102342 23468 102550
rect 23392 102278 23398 102342
rect 23462 102278 23468 102342
rect 195024 102550 195030 102614
rect 195094 102550 195100 102614
rect 195024 102342 195100 102550
rect 195024 102310 195030 102342
rect 23392 102272 23468 102278
rect 195029 102278 195030 102310
rect 195094 102310 195100 102342
rect 195568 102614 195644 102620
rect 195568 102550 195574 102614
rect 195638 102550 195644 102614
rect 195981 102614 196047 102615
rect 195981 102582 195982 102614
rect 195568 102342 195644 102550
rect 195568 102310 195574 102342
rect 195094 102278 195095 102310
rect 195029 102277 195095 102278
rect 195573 102278 195574 102310
rect 195638 102310 195644 102342
rect 195976 102550 195982 102582
rect 196046 102582 196047 102614
rect 196389 102614 196455 102615
rect 196389 102582 196390 102614
rect 196046 102550 196052 102582
rect 195976 102342 196052 102550
rect 195638 102278 195639 102310
rect 195573 102277 195639 102278
rect 195976 102278 195982 102342
rect 196046 102278 196052 102342
rect 195976 102272 196052 102278
rect 196384 102550 196390 102582
rect 196454 102582 196455 102614
rect 196454 102550 196460 102582
rect 196384 102342 196460 102550
rect 196384 102278 196390 102342
rect 196454 102278 196460 102342
rect 196384 102272 196460 102278
rect 21901 102206 21967 102207
rect 21901 102174 21902 102206
rect 21896 102142 21902 102174
rect 21966 102174 21967 102206
rect 23120 102206 23196 102212
rect 21966 102142 21972 102174
rect 21896 101934 21972 102142
rect 21896 101870 21902 101934
rect 21966 101870 21972 101934
rect 23120 102142 23126 102206
rect 23190 102142 23196 102206
rect 23120 101934 23196 102142
rect 23120 101902 23126 101934
rect 21896 101864 21972 101870
rect 23125 101870 23126 101902
rect 23190 101902 23196 101934
rect 23528 102206 23604 102212
rect 23528 102142 23534 102206
rect 23598 102142 23604 102206
rect 195165 102206 195231 102207
rect 195165 102174 195166 102206
rect 23528 101934 23604 102142
rect 23528 101902 23534 101934
rect 23190 101870 23191 101902
rect 23125 101869 23191 101870
rect 23533 101870 23534 101902
rect 23598 101902 23604 101934
rect 195160 102142 195166 102174
rect 195230 102174 195231 102206
rect 195437 102206 195503 102207
rect 195437 102174 195438 102206
rect 195230 102142 195236 102174
rect 195160 101934 195236 102142
rect 23598 101870 23599 101902
rect 23533 101869 23599 101870
rect 195160 101870 195166 101934
rect 195230 101870 195236 101934
rect 195160 101864 195236 101870
rect 195432 102142 195438 102174
rect 195502 102174 195503 102206
rect 196117 102206 196183 102207
rect 196117 102174 196118 102206
rect 195502 102142 195508 102174
rect 195432 101934 195508 102142
rect 195432 101870 195438 101934
rect 195502 101870 195508 101934
rect 195432 101864 195508 101870
rect 196112 102142 196118 102174
rect 196182 102174 196183 102206
rect 196656 102206 196732 102212
rect 196182 102142 196188 102174
rect 196112 101934 196188 102142
rect 196112 101870 196118 101934
rect 196182 101870 196188 101934
rect 196656 102142 196662 102206
rect 196726 102142 196732 102206
rect 196656 101934 196732 102142
rect 196656 101902 196662 101934
rect 196112 101864 196188 101870
rect 196661 101870 196662 101902
rect 196726 101902 196732 101934
rect 196726 101870 196727 101902
rect 196661 101869 196727 101870
rect 22304 101798 22380 101804
rect 22304 101734 22310 101798
rect 22374 101734 22380 101798
rect 21901 101526 21967 101527
rect 21901 101494 21902 101526
rect 952 101190 1230 101254
rect 1294 101190 1300 101254
rect 952 99622 1300 101190
rect 21896 101462 21902 101494
rect 21966 101494 21967 101526
rect 22304 101526 22380 101734
rect 22304 101494 22310 101526
rect 21966 101462 21972 101494
rect 21896 101254 21972 101462
rect 22309 101462 22310 101494
rect 22374 101494 22380 101526
rect 22440 101798 22516 101804
rect 22440 101734 22446 101798
rect 22510 101734 22516 101798
rect 23125 101798 23191 101799
rect 23125 101766 23126 101798
rect 22440 101526 22516 101734
rect 22440 101494 22446 101526
rect 22374 101462 22375 101494
rect 22309 101461 22375 101462
rect 22445 101462 22446 101494
rect 22510 101494 22516 101526
rect 23120 101734 23126 101766
rect 23190 101766 23191 101798
rect 23533 101798 23599 101799
rect 23533 101766 23534 101798
rect 23190 101734 23196 101766
rect 23120 101526 23196 101734
rect 22510 101462 22511 101494
rect 22445 101461 22511 101462
rect 23120 101462 23126 101526
rect 23190 101462 23196 101526
rect 23120 101456 23196 101462
rect 23528 101734 23534 101766
rect 23598 101766 23599 101798
rect 195024 101798 195100 101804
rect 23598 101734 23604 101766
rect 23528 101526 23604 101734
rect 195024 101734 195030 101798
rect 195094 101734 195100 101798
rect 28429 101662 28495 101663
rect 28429 101630 28430 101662
rect 23528 101462 23534 101526
rect 23598 101462 23604 101526
rect 23528 101456 23604 101462
rect 28424 101598 28430 101630
rect 28494 101630 28495 101662
rect 28494 101598 28500 101630
rect 21896 101190 21902 101254
rect 21966 101190 21972 101254
rect 21896 101184 21972 101190
rect 22984 101390 23060 101396
rect 22984 101326 22990 101390
rect 23054 101326 23060 101390
rect 22984 101118 23060 101326
rect 22984 101086 22990 101118
rect 22989 101054 22990 101086
rect 23054 101086 23060 101118
rect 23528 101390 23604 101396
rect 23528 101326 23534 101390
rect 23598 101326 23604 101390
rect 23528 101118 23604 101326
rect 28424 101390 28500 101598
rect 195024 101526 195100 101734
rect 195024 101494 195030 101526
rect 195029 101462 195030 101494
rect 195094 101494 195100 101526
rect 195432 101798 195508 101804
rect 195432 101734 195438 101798
rect 195502 101734 195508 101798
rect 195845 101798 195911 101799
rect 195845 101766 195846 101798
rect 195432 101526 195508 101734
rect 195432 101494 195438 101526
rect 195094 101462 195095 101494
rect 195029 101461 195095 101462
rect 195437 101462 195438 101494
rect 195502 101494 195508 101526
rect 195840 101734 195846 101766
rect 195910 101766 195911 101798
rect 195910 101734 195916 101766
rect 195840 101526 195916 101734
rect 195502 101462 195503 101494
rect 195437 101461 195503 101462
rect 195840 101462 195846 101526
rect 195910 101462 195916 101526
rect 196797 101526 196863 101527
rect 196797 101494 196798 101526
rect 195840 101456 195916 101462
rect 196792 101462 196798 101494
rect 196862 101494 196863 101526
rect 196862 101462 196868 101494
rect 28424 101326 28430 101390
rect 28494 101326 28500 101390
rect 190269 101390 190335 101391
rect 190269 101358 190270 101390
rect 28424 101320 28500 101326
rect 190264 101326 190270 101358
rect 190334 101358 190335 101390
rect 195029 101390 195095 101391
rect 195029 101358 195030 101390
rect 190334 101326 190340 101358
rect 23528 101086 23534 101118
rect 23054 101054 23055 101086
rect 22989 101053 23055 101054
rect 23533 101054 23534 101086
rect 23598 101086 23604 101118
rect 23598 101054 23599 101086
rect 23533 101053 23599 101054
rect 22173 100982 22239 100983
rect 22173 100950 22174 100982
rect 22168 100918 22174 100950
rect 22238 100950 22239 100982
rect 22576 100982 22652 100988
rect 22238 100918 22244 100950
rect 21765 100710 21831 100711
rect 21765 100678 21766 100710
rect 21760 100646 21766 100678
rect 21830 100678 21831 100710
rect 22168 100710 22244 100918
rect 21830 100646 21836 100678
rect 21760 100438 21836 100646
rect 22168 100646 22174 100710
rect 22238 100646 22244 100710
rect 22576 100918 22582 100982
rect 22646 100918 22652 100982
rect 22576 100710 22652 100918
rect 190264 100982 190340 101326
rect 195024 101326 195030 101358
rect 195094 101358 195095 101390
rect 195437 101390 195503 101391
rect 195437 101358 195438 101390
rect 195094 101326 195100 101358
rect 195024 101118 195100 101326
rect 195024 101054 195030 101118
rect 195094 101054 195100 101118
rect 195024 101048 195100 101054
rect 195432 101326 195438 101358
rect 195502 101358 195503 101390
rect 195502 101326 195508 101358
rect 195432 101118 195508 101326
rect 196792 101254 196868 101462
rect 196792 101190 196798 101254
rect 196862 101190 196868 101254
rect 196792 101184 196868 101190
rect 217464 101390 217812 102958
rect 217464 101326 217470 101390
rect 217534 101326 217812 101390
rect 195432 101054 195438 101118
rect 195502 101054 195508 101118
rect 195432 101048 195508 101054
rect 190264 100918 190270 100982
rect 190334 100918 190340 100982
rect 195845 100982 195911 100983
rect 195845 100950 195846 100982
rect 190264 100912 190340 100918
rect 195840 100918 195846 100950
rect 195910 100950 195911 100982
rect 196248 100982 196324 100988
rect 195910 100918 195916 100950
rect 22576 100678 22582 100710
rect 22168 100640 22244 100646
rect 22581 100646 22582 100678
rect 22646 100678 22652 100710
rect 195840 100710 195916 100918
rect 22646 100646 22647 100678
rect 22581 100645 22647 100646
rect 195840 100646 195846 100710
rect 195910 100646 195916 100710
rect 196248 100918 196254 100982
rect 196318 100918 196324 100982
rect 196248 100710 196324 100918
rect 196248 100678 196254 100710
rect 195840 100640 195916 100646
rect 196253 100646 196254 100678
rect 196318 100678 196324 100710
rect 196661 100710 196727 100711
rect 196661 100678 196662 100710
rect 196318 100646 196319 100678
rect 196253 100645 196319 100646
rect 196656 100646 196662 100678
rect 196726 100678 196727 100710
rect 196726 100646 196732 100678
rect 21760 100374 21766 100438
rect 21830 100374 21836 100438
rect 21760 100368 21836 100374
rect 196656 100438 196732 100646
rect 196656 100374 196662 100438
rect 196726 100374 196732 100438
rect 196656 100368 196732 100374
rect 21760 100302 21836 100308
rect 21760 100238 21766 100302
rect 21830 100238 21836 100302
rect 22445 100302 22511 100303
rect 22445 100270 22446 100302
rect 21760 100030 21836 100238
rect 21760 99998 21766 100030
rect 21765 99966 21766 99998
rect 21830 99998 21836 100030
rect 22440 100238 22446 100270
rect 22510 100270 22511 100302
rect 23125 100302 23191 100303
rect 23125 100270 23126 100302
rect 22510 100238 22516 100270
rect 22440 100030 22516 100238
rect 21830 99966 21831 99998
rect 21765 99965 21831 99966
rect 22440 99966 22446 100030
rect 22510 99966 22516 100030
rect 22440 99960 22516 99966
rect 23120 100238 23126 100270
rect 23190 100270 23191 100302
rect 23397 100302 23463 100303
rect 23397 100270 23398 100302
rect 23190 100238 23196 100270
rect 23120 100030 23196 100238
rect 23120 99966 23126 100030
rect 23190 99966 23196 100030
rect 23120 99960 23196 99966
rect 23392 100238 23398 100270
rect 23462 100270 23463 100302
rect 195029 100302 195095 100303
rect 195029 100270 195030 100302
rect 23462 100238 23468 100270
rect 23392 100030 23468 100238
rect 23392 99966 23398 100030
rect 23462 99966 23468 100030
rect 23392 99960 23468 99966
rect 195024 100238 195030 100270
rect 195094 100270 195095 100302
rect 195573 100302 195639 100303
rect 195573 100270 195574 100302
rect 195094 100238 195100 100270
rect 195024 100030 195100 100238
rect 195024 99966 195030 100030
rect 195094 99966 195100 100030
rect 195024 99960 195100 99966
rect 195568 100238 195574 100270
rect 195638 100270 195639 100302
rect 195840 100302 195916 100308
rect 195638 100238 195644 100270
rect 195568 100030 195644 100238
rect 195568 99966 195574 100030
rect 195638 99966 195644 100030
rect 195840 100238 195846 100302
rect 195910 100238 195916 100302
rect 196797 100302 196863 100303
rect 196797 100270 196798 100302
rect 195840 100030 195916 100238
rect 195840 99998 195846 100030
rect 195568 99960 195644 99966
rect 195845 99966 195846 99998
rect 195910 99998 195916 100030
rect 196792 100238 196798 100270
rect 196862 100270 196863 100302
rect 196862 100238 196868 100270
rect 196792 100030 196868 100238
rect 195910 99966 195911 99998
rect 195845 99965 195911 99966
rect 196792 99966 196798 100030
rect 196862 99966 196868 100030
rect 196792 99960 196868 99966
rect 21765 99894 21831 99895
rect 21765 99862 21766 99894
rect 952 99558 1230 99622
rect 1294 99558 1300 99622
rect 952 97990 1300 99558
rect 21760 99830 21766 99862
rect 21830 99862 21831 99894
rect 23120 99894 23196 99900
rect 21830 99830 21836 99862
rect 21760 99622 21836 99830
rect 21760 99558 21766 99622
rect 21830 99558 21836 99622
rect 23120 99830 23126 99894
rect 23190 99830 23196 99894
rect 23120 99622 23196 99830
rect 23120 99590 23126 99622
rect 21760 99552 21836 99558
rect 23125 99558 23126 99590
rect 23190 99590 23196 99622
rect 23528 99894 23604 99900
rect 23528 99830 23534 99894
rect 23598 99830 23604 99894
rect 23528 99622 23604 99830
rect 23528 99590 23534 99622
rect 23190 99558 23191 99590
rect 23125 99557 23191 99558
rect 23533 99558 23534 99590
rect 23598 99590 23604 99622
rect 195160 99894 195236 99900
rect 195160 99830 195166 99894
rect 195230 99830 195236 99894
rect 195160 99622 195236 99830
rect 195160 99590 195166 99622
rect 23598 99558 23599 99590
rect 23533 99557 23599 99558
rect 195165 99558 195166 99590
rect 195230 99590 195236 99622
rect 195568 99894 195644 99900
rect 195568 99830 195574 99894
rect 195638 99830 195644 99894
rect 195568 99622 195644 99830
rect 195568 99590 195574 99622
rect 195230 99558 195231 99590
rect 195165 99557 195231 99558
rect 195573 99558 195574 99590
rect 195638 99590 195644 99622
rect 196656 99894 196732 99900
rect 196656 99830 196662 99894
rect 196726 99830 196732 99894
rect 196656 99622 196732 99830
rect 196656 99590 196662 99622
rect 195638 99558 195639 99590
rect 195573 99557 195639 99558
rect 196661 99558 196662 99590
rect 196726 99590 196732 99622
rect 217464 99758 217812 101326
rect 217464 99694 217470 99758
rect 217534 99694 217812 99758
rect 196726 99558 196727 99590
rect 196661 99557 196727 99558
rect 21896 99486 21972 99492
rect 21896 99422 21902 99486
rect 21966 99422 21972 99486
rect 21896 99214 21972 99422
rect 21896 99182 21902 99214
rect 21901 99150 21902 99182
rect 21966 99182 21972 99214
rect 22712 99486 22788 99492
rect 22712 99422 22718 99486
rect 22782 99422 22788 99486
rect 22712 99214 22788 99422
rect 22712 99182 22718 99214
rect 21966 99150 21967 99182
rect 21901 99149 21967 99150
rect 22717 99150 22718 99182
rect 22782 99182 22788 99214
rect 23120 99486 23196 99492
rect 23120 99422 23126 99486
rect 23190 99422 23196 99486
rect 23397 99486 23463 99487
rect 23397 99454 23398 99486
rect 23120 99214 23196 99422
rect 23120 99182 23126 99214
rect 22782 99150 22783 99182
rect 22717 99149 22783 99150
rect 23125 99150 23126 99182
rect 23190 99182 23196 99214
rect 23392 99422 23398 99454
rect 23462 99454 23463 99486
rect 195029 99486 195095 99487
rect 195029 99454 195030 99486
rect 23462 99422 23468 99454
rect 23392 99214 23468 99422
rect 23190 99150 23191 99182
rect 23125 99149 23191 99150
rect 23392 99150 23398 99214
rect 23462 99150 23468 99214
rect 23392 99144 23468 99150
rect 195024 99422 195030 99454
rect 195094 99454 195095 99486
rect 195568 99486 195644 99492
rect 195094 99422 195100 99454
rect 195024 99214 195100 99422
rect 195024 99150 195030 99214
rect 195094 99150 195100 99214
rect 195568 99422 195574 99486
rect 195638 99422 195644 99486
rect 196797 99486 196863 99487
rect 196797 99454 196798 99486
rect 195568 99214 195644 99422
rect 195568 99182 195574 99214
rect 195024 99144 195100 99150
rect 195573 99150 195574 99182
rect 195638 99182 195644 99214
rect 196792 99422 196798 99454
rect 196862 99454 196863 99486
rect 196862 99422 196868 99454
rect 196792 99214 196868 99422
rect 195638 99150 195639 99182
rect 195573 99149 195639 99150
rect 196792 99150 196798 99214
rect 196862 99150 196868 99214
rect 196792 99144 196868 99150
rect 21760 99078 21836 99084
rect 21760 99014 21766 99078
rect 21830 99014 21836 99078
rect 23125 99078 23191 99079
rect 23125 99046 23126 99078
rect 21760 98806 21836 99014
rect 21760 98774 21766 98806
rect 21765 98742 21766 98774
rect 21830 98774 21836 98806
rect 23120 99014 23126 99046
rect 23190 99046 23191 99078
rect 23528 99078 23604 99084
rect 23190 99014 23196 99046
rect 23120 98806 23196 99014
rect 21830 98742 21831 98774
rect 21765 98741 21831 98742
rect 23120 98742 23126 98806
rect 23190 98742 23196 98806
rect 23528 99014 23534 99078
rect 23598 99014 23604 99078
rect 195029 99078 195095 99079
rect 195029 99046 195030 99078
rect 23528 98806 23604 99014
rect 23528 98774 23534 98806
rect 23120 98736 23196 98742
rect 23533 98742 23534 98774
rect 23598 98774 23604 98806
rect 195024 99014 195030 99046
rect 195094 99046 195095 99078
rect 195573 99078 195639 99079
rect 195573 99046 195574 99078
rect 195094 99014 195100 99046
rect 195024 98806 195100 99014
rect 23598 98742 23599 98774
rect 23533 98741 23599 98742
rect 195024 98742 195030 98806
rect 195094 98742 195100 98806
rect 195024 98736 195100 98742
rect 195568 99014 195574 99046
rect 195638 99046 195639 99078
rect 196117 99078 196183 99079
rect 196117 99046 196118 99078
rect 195638 99014 195644 99046
rect 195568 98806 195644 99014
rect 195568 98742 195574 98806
rect 195638 98742 195644 98806
rect 195568 98736 195644 98742
rect 196112 99014 196118 99046
rect 196182 99046 196183 99078
rect 196797 99078 196863 99079
rect 196797 99046 196798 99078
rect 196182 99014 196188 99046
rect 196112 98806 196188 99014
rect 196112 98742 196118 98806
rect 196182 98742 196188 98806
rect 196112 98736 196188 98742
rect 196792 99014 196798 99046
rect 196862 99046 196863 99078
rect 196862 99014 196868 99046
rect 196792 98806 196868 99014
rect 196792 98742 196798 98806
rect 196862 98742 196868 98806
rect 196792 98736 196868 98742
rect 21765 98670 21831 98671
rect 21765 98638 21766 98670
rect 21760 98606 21766 98638
rect 21830 98638 21831 98670
rect 22173 98670 22239 98671
rect 22173 98638 22174 98670
rect 21830 98606 21836 98638
rect 21760 98398 21836 98606
rect 21760 98334 21766 98398
rect 21830 98334 21836 98398
rect 21760 98328 21836 98334
rect 22168 98606 22174 98638
rect 22238 98638 22239 98670
rect 22712 98670 22788 98676
rect 22238 98606 22244 98638
rect 22168 98398 22244 98606
rect 22168 98334 22174 98398
rect 22238 98334 22244 98398
rect 22712 98606 22718 98670
rect 22782 98606 22788 98670
rect 22989 98670 23055 98671
rect 22989 98638 22990 98670
rect 22712 98398 22788 98606
rect 22712 98366 22718 98398
rect 22168 98328 22244 98334
rect 22717 98334 22718 98366
rect 22782 98366 22788 98398
rect 22984 98606 22990 98638
rect 23054 98638 23055 98670
rect 23533 98670 23599 98671
rect 23533 98638 23534 98670
rect 23054 98606 23060 98638
rect 22984 98398 23060 98606
rect 22782 98334 22783 98366
rect 22717 98333 22783 98334
rect 22984 98334 22990 98398
rect 23054 98334 23060 98398
rect 22984 98328 23060 98334
rect 23528 98606 23534 98638
rect 23598 98638 23599 98670
rect 195024 98670 195100 98676
rect 23598 98606 23604 98638
rect 23528 98398 23604 98606
rect 23528 98334 23534 98398
rect 23598 98334 23604 98398
rect 195024 98606 195030 98670
rect 195094 98606 195100 98670
rect 195573 98670 195639 98671
rect 195573 98638 195574 98670
rect 195024 98398 195100 98606
rect 195024 98366 195030 98398
rect 23528 98328 23604 98334
rect 195029 98334 195030 98366
rect 195094 98366 195100 98398
rect 195568 98606 195574 98638
rect 195638 98638 195639 98670
rect 195976 98670 196052 98676
rect 195638 98606 195644 98638
rect 195568 98398 195644 98606
rect 195094 98334 195095 98366
rect 195029 98333 195095 98334
rect 195568 98334 195574 98398
rect 195638 98334 195644 98398
rect 195976 98606 195982 98670
rect 196046 98606 196052 98670
rect 196661 98670 196727 98671
rect 196661 98638 196662 98670
rect 195976 98398 196052 98606
rect 195976 98366 195982 98398
rect 195568 98328 195644 98334
rect 195981 98334 195982 98366
rect 196046 98366 196052 98398
rect 196656 98606 196662 98638
rect 196726 98638 196727 98670
rect 196726 98606 196732 98638
rect 196656 98398 196732 98606
rect 196046 98334 196047 98366
rect 195981 98333 196047 98334
rect 196656 98334 196662 98398
rect 196726 98334 196732 98398
rect 196656 98328 196732 98334
rect 21901 98262 21967 98263
rect 21901 98230 21902 98262
rect 952 97926 1230 97990
rect 1294 97926 1300 97990
rect 952 96222 1300 97926
rect 21896 98198 21902 98230
rect 21966 98230 21967 98262
rect 22309 98262 22375 98263
rect 22309 98230 22310 98262
rect 21966 98198 21972 98230
rect 21896 97990 21972 98198
rect 21896 97926 21902 97990
rect 21966 97926 21972 97990
rect 21896 97920 21972 97926
rect 22304 98198 22310 98230
rect 22374 98230 22375 98262
rect 22445 98262 22511 98263
rect 22445 98230 22446 98262
rect 22374 98198 22380 98230
rect 22304 97990 22380 98198
rect 22304 97926 22310 97990
rect 22374 97926 22380 97990
rect 22304 97920 22380 97926
rect 22440 98198 22446 98230
rect 22510 98230 22511 98262
rect 23120 98262 23196 98268
rect 22510 98198 22516 98230
rect 22440 97990 22516 98198
rect 22440 97926 22446 97990
rect 22510 97926 22516 97990
rect 23120 98198 23126 98262
rect 23190 98198 23196 98262
rect 23120 97990 23196 98198
rect 23120 97958 23126 97990
rect 22440 97920 22516 97926
rect 23125 97926 23126 97958
rect 23190 97958 23196 97990
rect 23392 98262 23468 98268
rect 23392 98198 23398 98262
rect 23462 98198 23468 98262
rect 23392 97990 23468 98198
rect 23392 97958 23398 97990
rect 23190 97926 23191 97958
rect 23125 97925 23191 97926
rect 23397 97926 23398 97958
rect 23462 97958 23468 97990
rect 195024 98262 195100 98268
rect 195024 98198 195030 98262
rect 195094 98198 195100 98262
rect 195024 97990 195100 98198
rect 195024 97958 195030 97990
rect 23462 97926 23463 97958
rect 23397 97925 23463 97926
rect 195029 97926 195030 97958
rect 195094 97958 195100 97990
rect 195568 98262 195644 98268
rect 195568 98198 195574 98262
rect 195638 98198 195644 98262
rect 196389 98262 196455 98263
rect 196389 98230 196390 98262
rect 195568 97990 195644 98198
rect 195568 97958 195574 97990
rect 195094 97926 195095 97958
rect 195029 97925 195095 97926
rect 195573 97926 195574 97958
rect 195638 97958 195644 97990
rect 196384 98198 196390 98230
rect 196454 98230 196455 98262
rect 196792 98262 196868 98268
rect 196454 98198 196460 98230
rect 196384 97990 196460 98198
rect 195638 97926 195639 97958
rect 195573 97925 195639 97926
rect 196384 97926 196390 97990
rect 196454 97926 196460 97990
rect 196792 98198 196798 98262
rect 196862 98198 196868 98262
rect 196792 97990 196868 98198
rect 196792 97958 196798 97990
rect 196384 97920 196460 97926
rect 196797 97926 196798 97958
rect 196862 97958 196868 97990
rect 196862 97926 196863 97958
rect 196797 97925 196863 97926
rect 22168 97854 22244 97860
rect 22168 97790 22174 97854
rect 22238 97790 22244 97854
rect 22989 97854 23055 97855
rect 22989 97822 22990 97854
rect 22168 97582 22244 97790
rect 22168 97550 22174 97582
rect 22173 97518 22174 97550
rect 22238 97550 22244 97582
rect 22984 97790 22990 97822
rect 23054 97822 23055 97854
rect 23528 97854 23604 97860
rect 23054 97790 23060 97822
rect 22984 97582 23060 97790
rect 22238 97518 22239 97550
rect 22173 97517 22239 97518
rect 22984 97518 22990 97582
rect 23054 97518 23060 97582
rect 23528 97790 23534 97854
rect 23598 97790 23604 97854
rect 195165 97854 195231 97855
rect 195165 97822 195166 97854
rect 23528 97582 23604 97790
rect 23528 97550 23534 97582
rect 22984 97512 23060 97518
rect 23533 97518 23534 97550
rect 23598 97550 23604 97582
rect 195160 97790 195166 97822
rect 195230 97822 195231 97854
rect 195437 97854 195503 97855
rect 195437 97822 195438 97854
rect 195230 97790 195236 97822
rect 195160 97582 195236 97790
rect 23598 97518 23599 97550
rect 23533 97517 23599 97518
rect 195160 97518 195166 97582
rect 195230 97518 195236 97582
rect 195160 97512 195236 97518
rect 195432 97790 195438 97822
rect 195502 97822 195503 97854
rect 195845 97854 195911 97855
rect 195845 97822 195846 97854
rect 195502 97790 195508 97822
rect 195432 97582 195508 97790
rect 195432 97518 195438 97582
rect 195502 97518 195508 97582
rect 195432 97512 195508 97518
rect 195840 97790 195846 97822
rect 195910 97822 195911 97854
rect 196248 97854 196324 97860
rect 195910 97790 195916 97822
rect 195840 97582 195916 97790
rect 195840 97518 195846 97582
rect 195910 97518 195916 97582
rect 196248 97790 196254 97854
rect 196318 97790 196324 97854
rect 196248 97582 196324 97790
rect 196248 97550 196254 97582
rect 195840 97512 195916 97518
rect 196253 97518 196254 97550
rect 196318 97550 196324 97582
rect 217464 97854 217812 99694
rect 217464 97790 217470 97854
rect 217534 97790 217812 97854
rect 196318 97518 196319 97550
rect 196253 97517 196319 97518
rect 22984 97446 23060 97452
rect 22984 97382 22990 97446
rect 23054 97382 23060 97446
rect 23533 97446 23599 97447
rect 23533 97414 23534 97446
rect 22984 97174 23060 97382
rect 22984 97142 22990 97174
rect 22989 97110 22990 97142
rect 23054 97142 23060 97174
rect 23528 97382 23534 97414
rect 23598 97414 23599 97446
rect 195024 97446 195100 97452
rect 23598 97382 23604 97414
rect 23528 97174 23604 97382
rect 23054 97110 23055 97142
rect 22989 97109 23055 97110
rect 23528 97110 23534 97174
rect 23598 97110 23604 97174
rect 195024 97382 195030 97446
rect 195094 97382 195100 97446
rect 195573 97446 195639 97447
rect 195573 97414 195574 97446
rect 195024 97174 195100 97382
rect 195024 97142 195030 97174
rect 23528 97104 23604 97110
rect 195029 97110 195030 97142
rect 195094 97142 195100 97174
rect 195568 97382 195574 97414
rect 195638 97414 195639 97446
rect 195638 97382 195644 97414
rect 195568 97174 195644 97382
rect 195094 97110 195095 97142
rect 195029 97109 195095 97110
rect 195568 97110 195574 97174
rect 195638 97110 195644 97174
rect 195568 97104 195644 97110
rect 22717 97038 22783 97039
rect 22717 97006 22718 97038
rect 22712 96974 22718 97006
rect 22782 97006 22783 97038
rect 196248 97038 196324 97044
rect 22782 96974 22788 97006
rect 21760 96766 21836 96772
rect 21760 96702 21766 96766
rect 21830 96702 21836 96766
rect 21760 96494 21836 96702
rect 22712 96766 22788 96974
rect 196248 96974 196254 97038
rect 196318 96974 196324 97038
rect 28565 96902 28631 96903
rect 28565 96870 28566 96902
rect 22712 96702 22718 96766
rect 22782 96702 22788 96766
rect 22712 96696 22788 96702
rect 28560 96838 28566 96870
rect 28630 96870 28631 96902
rect 28630 96838 28636 96870
rect 28560 96630 28636 96838
rect 196248 96766 196324 96974
rect 196248 96734 196254 96766
rect 196253 96702 196254 96734
rect 196318 96734 196324 96766
rect 196656 96766 196732 96772
rect 196318 96702 196319 96734
rect 196253 96701 196319 96702
rect 196656 96702 196662 96766
rect 196726 96702 196732 96766
rect 28560 96566 28566 96630
rect 28630 96566 28636 96630
rect 28560 96560 28636 96566
rect 21760 96462 21766 96494
rect 21765 96430 21766 96462
rect 21830 96462 21836 96494
rect 28429 96494 28495 96495
rect 28429 96462 28430 96494
rect 21830 96430 21831 96462
rect 21765 96429 21831 96430
rect 28424 96430 28430 96462
rect 28494 96462 28495 96494
rect 190133 96494 190199 96495
rect 190133 96462 190134 96494
rect 28494 96430 28500 96462
rect 21765 96358 21831 96359
rect 21765 96326 21766 96358
rect 952 96158 1230 96222
rect 1294 96158 1300 96222
rect 952 94726 1300 96158
rect 21760 96294 21766 96326
rect 21830 96326 21831 96358
rect 22304 96358 22380 96364
rect 21830 96294 21836 96326
rect 21760 96086 21836 96294
rect 21760 96022 21766 96086
rect 21830 96022 21836 96086
rect 22304 96294 22310 96358
rect 22374 96294 22380 96358
rect 22304 96086 22380 96294
rect 28424 96222 28500 96430
rect 28424 96158 28430 96222
rect 28494 96158 28500 96222
rect 28424 96152 28500 96158
rect 190128 96430 190134 96462
rect 190198 96462 190199 96494
rect 196656 96494 196732 96702
rect 196656 96462 196662 96494
rect 190198 96430 190204 96462
rect 190128 96222 190204 96430
rect 196661 96430 196662 96462
rect 196726 96462 196732 96494
rect 196726 96430 196727 96462
rect 196661 96429 196727 96430
rect 190128 96158 190134 96222
rect 190198 96158 190204 96222
rect 190128 96152 190204 96158
rect 195976 96358 196052 96364
rect 195976 96294 195982 96358
rect 196046 96294 196052 96358
rect 22304 96054 22310 96086
rect 21760 96016 21836 96022
rect 22309 96022 22310 96054
rect 22374 96054 22380 96086
rect 28424 96086 28500 96092
rect 22374 96022 22375 96054
rect 22309 96021 22375 96022
rect 28424 96022 28430 96086
rect 28494 96022 28500 96086
rect 195976 96086 196052 96294
rect 195976 96054 195982 96086
rect 21760 95950 21836 95956
rect 21760 95886 21766 95950
rect 21830 95886 21836 95950
rect 21760 95678 21836 95886
rect 21760 95646 21766 95678
rect 21765 95614 21766 95646
rect 21830 95646 21836 95678
rect 22984 95950 23060 95956
rect 22984 95886 22990 95950
rect 23054 95886 23060 95950
rect 23397 95950 23463 95951
rect 23397 95918 23398 95950
rect 22984 95678 23060 95886
rect 22984 95646 22990 95678
rect 21830 95614 21831 95646
rect 21765 95613 21831 95614
rect 22989 95614 22990 95646
rect 23054 95646 23060 95678
rect 23392 95886 23398 95918
rect 23462 95918 23463 95950
rect 23462 95886 23468 95918
rect 23392 95678 23468 95886
rect 28424 95814 28500 96022
rect 195981 96022 195982 96054
rect 196046 96054 196052 96086
rect 196112 96358 196188 96364
rect 196112 96294 196118 96358
rect 196182 96294 196188 96358
rect 196661 96358 196727 96359
rect 196661 96326 196662 96358
rect 196112 96086 196188 96294
rect 196112 96054 196118 96086
rect 196046 96022 196047 96054
rect 195981 96021 196047 96022
rect 196117 96022 196118 96054
rect 196182 96054 196188 96086
rect 196656 96294 196662 96326
rect 196726 96326 196727 96358
rect 217464 96358 217812 97790
rect 196726 96294 196732 96326
rect 196656 96086 196732 96294
rect 196182 96022 196183 96054
rect 196117 96021 196183 96022
rect 196656 96022 196662 96086
rect 196726 96022 196732 96086
rect 196656 96016 196732 96022
rect 217464 96294 217470 96358
rect 217534 96294 217812 96358
rect 195029 95950 195095 95951
rect 195029 95918 195030 95950
rect 28424 95782 28430 95814
rect 28429 95750 28430 95782
rect 28494 95782 28500 95814
rect 195024 95886 195030 95918
rect 195094 95918 195095 95950
rect 195573 95950 195639 95951
rect 195573 95918 195574 95950
rect 195094 95886 195100 95918
rect 28494 95750 28495 95782
rect 28429 95749 28495 95750
rect 23054 95614 23055 95646
rect 22989 95613 23055 95614
rect 23392 95614 23398 95678
rect 23462 95614 23468 95678
rect 23392 95608 23468 95614
rect 195024 95678 195100 95886
rect 195024 95614 195030 95678
rect 195094 95614 195100 95678
rect 195024 95608 195100 95614
rect 195568 95886 195574 95918
rect 195638 95918 195639 95950
rect 196797 95950 196863 95951
rect 196797 95918 196798 95950
rect 195638 95886 195644 95918
rect 195568 95678 195644 95886
rect 196792 95886 196798 95918
rect 196862 95918 196863 95950
rect 196862 95886 196868 95918
rect 195568 95614 195574 95678
rect 195638 95614 195644 95678
rect 196112 95814 196324 95820
rect 196112 95750 196254 95814
rect 196318 95750 196324 95814
rect 196112 95744 196324 95750
rect 196112 95678 196188 95744
rect 196112 95646 196118 95678
rect 195568 95608 195644 95614
rect 196117 95614 196118 95646
rect 196182 95646 196188 95678
rect 196792 95678 196868 95886
rect 196182 95614 196183 95646
rect 196117 95613 196183 95614
rect 196792 95614 196798 95678
rect 196862 95614 196868 95678
rect 196792 95608 196868 95614
rect 21765 95542 21831 95543
rect 21765 95510 21766 95542
rect 21760 95478 21766 95510
rect 21830 95510 21831 95542
rect 22576 95542 22652 95548
rect 21830 95478 21836 95510
rect 21760 95270 21836 95478
rect 21760 95206 21766 95270
rect 21830 95206 21836 95270
rect 22576 95478 22582 95542
rect 22646 95478 22652 95542
rect 22989 95542 23055 95543
rect 22989 95510 22990 95542
rect 22576 95270 22652 95478
rect 22576 95238 22582 95270
rect 21760 95200 21836 95206
rect 22581 95206 22582 95238
rect 22646 95238 22652 95270
rect 22984 95478 22990 95510
rect 23054 95510 23055 95542
rect 23528 95542 23604 95548
rect 23054 95478 23060 95510
rect 22984 95270 23060 95478
rect 22646 95206 22647 95238
rect 22581 95205 22647 95206
rect 22984 95206 22990 95270
rect 23054 95206 23060 95270
rect 23528 95478 23534 95542
rect 23598 95478 23604 95542
rect 195165 95542 195231 95543
rect 195165 95510 195166 95542
rect 23528 95270 23604 95478
rect 195160 95478 195166 95510
rect 195230 95510 195231 95542
rect 195568 95542 195644 95548
rect 195230 95478 195236 95510
rect 23528 95238 23534 95270
rect 22984 95200 23060 95206
rect 23533 95206 23534 95238
rect 23598 95238 23604 95270
rect 190269 95270 190335 95271
rect 190269 95238 190270 95270
rect 23598 95206 23599 95238
rect 23533 95205 23599 95206
rect 190264 95206 190270 95238
rect 190334 95238 190335 95270
rect 195160 95270 195236 95478
rect 190334 95206 190340 95238
rect 21901 95134 21967 95135
rect 21901 95102 21902 95134
rect 21896 95070 21902 95102
rect 21966 95102 21967 95134
rect 22717 95134 22783 95135
rect 22717 95102 22718 95134
rect 21966 95070 21972 95102
rect 21896 94862 21972 95070
rect 21896 94798 21902 94862
rect 21966 94798 21972 94862
rect 21896 94792 21972 94798
rect 22712 95070 22718 95102
rect 22782 95102 22783 95134
rect 23120 95134 23196 95140
rect 22782 95070 22788 95102
rect 22712 94862 22788 95070
rect 22712 94798 22718 94862
rect 22782 94798 22788 94862
rect 23120 95070 23126 95134
rect 23190 95070 23196 95134
rect 23397 95134 23463 95135
rect 23397 95102 23398 95134
rect 23120 94862 23196 95070
rect 23120 94830 23126 94862
rect 22712 94792 22788 94798
rect 23125 94798 23126 94830
rect 23190 94830 23196 94862
rect 23392 95070 23398 95102
rect 23462 95102 23463 95134
rect 23462 95070 23468 95102
rect 23392 94862 23468 95070
rect 190264 94998 190340 95206
rect 195160 95206 195166 95270
rect 195230 95206 195236 95270
rect 195568 95478 195574 95542
rect 195638 95478 195644 95542
rect 196117 95542 196183 95543
rect 196117 95510 196118 95542
rect 195568 95270 195644 95478
rect 195568 95238 195574 95270
rect 195160 95200 195236 95206
rect 195573 95206 195574 95238
rect 195638 95238 195644 95270
rect 196112 95478 196118 95510
rect 196182 95510 196183 95542
rect 196656 95542 196732 95548
rect 196182 95478 196188 95510
rect 196112 95270 196188 95478
rect 195638 95206 195639 95238
rect 195573 95205 195639 95206
rect 196112 95206 196118 95270
rect 196182 95206 196188 95270
rect 196656 95478 196662 95542
rect 196726 95478 196732 95542
rect 196656 95270 196732 95478
rect 196656 95238 196662 95270
rect 196112 95200 196188 95206
rect 196661 95206 196662 95238
rect 196726 95238 196732 95270
rect 196726 95206 196727 95238
rect 196661 95205 196727 95206
rect 190264 94934 190270 94998
rect 190334 94934 190340 94998
rect 190264 94928 190340 94934
rect 195024 95134 195100 95140
rect 195024 95070 195030 95134
rect 195094 95070 195100 95134
rect 23190 94798 23191 94830
rect 23125 94797 23191 94798
rect 23392 94798 23398 94862
rect 23462 94798 23468 94862
rect 195024 94862 195100 95070
rect 195024 94830 195030 94862
rect 23392 94792 23468 94798
rect 195029 94798 195030 94830
rect 195094 94830 195100 94862
rect 195568 95134 195644 95140
rect 195568 95070 195574 95134
rect 195638 95070 195644 95134
rect 195568 94862 195644 95070
rect 195568 94830 195574 94862
rect 195094 94798 195095 94830
rect 195029 94797 195095 94798
rect 195573 94798 195574 94830
rect 195638 94830 195644 94862
rect 195976 95134 196052 95140
rect 195976 95070 195982 95134
rect 196046 95070 196052 95134
rect 196797 95134 196863 95135
rect 196797 95102 196798 95134
rect 195976 94862 196052 95070
rect 195976 94830 195982 94862
rect 195638 94798 195639 94830
rect 195573 94797 195639 94798
rect 195981 94798 195982 94830
rect 196046 94830 196052 94862
rect 196792 95070 196798 95102
rect 196862 95102 196863 95134
rect 196862 95070 196868 95102
rect 196792 94862 196868 95070
rect 196046 94798 196047 94830
rect 195981 94797 196047 94798
rect 196792 94798 196798 94862
rect 196862 94798 196868 94862
rect 196792 94792 196868 94798
rect 952 94662 1230 94726
rect 1294 94662 1300 94726
rect 952 92822 1300 94662
rect 21760 94726 21836 94732
rect 21760 94662 21766 94726
rect 21830 94662 21836 94726
rect 22309 94726 22375 94727
rect 22309 94694 22310 94726
rect 21760 94454 21836 94662
rect 21760 94422 21766 94454
rect 21765 94390 21766 94422
rect 21830 94422 21836 94454
rect 22304 94662 22310 94694
rect 22374 94694 22375 94726
rect 22445 94726 22511 94727
rect 22445 94694 22446 94726
rect 22374 94662 22380 94694
rect 22304 94454 22380 94662
rect 21830 94390 21831 94422
rect 21765 94389 21831 94390
rect 22304 94390 22310 94454
rect 22374 94390 22380 94454
rect 22304 94384 22380 94390
rect 22440 94662 22446 94694
rect 22510 94694 22511 94726
rect 22984 94726 23060 94732
rect 22510 94662 22516 94694
rect 22440 94454 22516 94662
rect 22440 94390 22446 94454
rect 22510 94390 22516 94454
rect 22984 94662 22990 94726
rect 23054 94662 23060 94726
rect 22984 94454 23060 94662
rect 22984 94422 22990 94454
rect 22440 94384 22516 94390
rect 22989 94390 22990 94422
rect 23054 94422 23060 94454
rect 23528 94726 23604 94732
rect 23528 94662 23534 94726
rect 23598 94662 23604 94726
rect 195029 94726 195095 94727
rect 195029 94694 195030 94726
rect 23528 94454 23604 94662
rect 23528 94422 23534 94454
rect 23054 94390 23055 94422
rect 22989 94389 23055 94390
rect 23533 94390 23534 94422
rect 23598 94422 23604 94454
rect 195024 94662 195030 94694
rect 195094 94694 195095 94726
rect 195573 94726 195639 94727
rect 195573 94694 195574 94726
rect 195094 94662 195100 94694
rect 195024 94454 195100 94662
rect 23598 94390 23599 94422
rect 23533 94389 23599 94390
rect 195024 94390 195030 94454
rect 195094 94390 195100 94454
rect 195024 94384 195100 94390
rect 195568 94662 195574 94694
rect 195638 94694 195639 94726
rect 196117 94726 196183 94727
rect 196117 94694 196118 94726
rect 195638 94662 195644 94694
rect 195568 94454 195644 94662
rect 195568 94390 195574 94454
rect 195638 94390 195644 94454
rect 195568 94384 195644 94390
rect 196112 94662 196118 94694
rect 196182 94694 196183 94726
rect 196656 94726 196732 94732
rect 196182 94662 196188 94694
rect 196112 94454 196188 94662
rect 196112 94390 196118 94454
rect 196182 94390 196188 94454
rect 196656 94662 196662 94726
rect 196726 94662 196732 94726
rect 196656 94454 196732 94662
rect 196656 94422 196662 94454
rect 196112 94384 196188 94390
rect 196661 94390 196662 94422
rect 196726 94422 196732 94454
rect 217464 94590 217812 96294
rect 217464 94526 217470 94590
rect 217534 94526 217812 94590
rect 196726 94390 196727 94422
rect 196661 94389 196727 94390
rect 21765 94318 21831 94319
rect 21765 94286 21766 94318
rect 21760 94254 21766 94286
rect 21830 94286 21831 94318
rect 22712 94318 22788 94324
rect 21830 94254 21836 94286
rect 21760 94046 21836 94254
rect 21760 93982 21766 94046
rect 21830 93982 21836 94046
rect 22712 94254 22718 94318
rect 22782 94254 22788 94318
rect 22712 94046 22788 94254
rect 22712 94014 22718 94046
rect 21760 93976 21836 93982
rect 22717 93982 22718 94014
rect 22782 94014 22788 94046
rect 22984 94318 23060 94324
rect 22984 94254 22990 94318
rect 23054 94254 23060 94318
rect 23533 94318 23599 94319
rect 23533 94286 23534 94318
rect 22984 94046 23060 94254
rect 22984 94014 22990 94046
rect 22782 93982 22783 94014
rect 22717 93981 22783 93982
rect 22989 93982 22990 94014
rect 23054 94014 23060 94046
rect 23528 94254 23534 94286
rect 23598 94286 23599 94318
rect 195024 94318 195100 94324
rect 23598 94254 23604 94286
rect 23528 94046 23604 94254
rect 23054 93982 23055 94014
rect 22989 93981 23055 93982
rect 23528 93982 23534 94046
rect 23598 93982 23604 94046
rect 195024 94254 195030 94318
rect 195094 94254 195100 94318
rect 195024 94046 195100 94254
rect 195024 94014 195030 94046
rect 23528 93976 23604 93982
rect 195029 93982 195030 94014
rect 195094 94014 195100 94046
rect 195432 94318 195508 94324
rect 195432 94254 195438 94318
rect 195502 94254 195508 94318
rect 195432 94046 195508 94254
rect 195432 94014 195438 94046
rect 195094 93982 195095 94014
rect 195029 93981 195095 93982
rect 195437 93982 195438 94014
rect 195502 94014 195508 94046
rect 195976 94318 196052 94324
rect 195976 94254 195982 94318
rect 196046 94254 196052 94318
rect 195976 94046 196052 94254
rect 195976 94014 195982 94046
rect 195502 93982 195503 94014
rect 195437 93981 195503 93982
rect 195981 93982 195982 94014
rect 196046 94014 196052 94046
rect 196112 94318 196188 94324
rect 196112 94254 196118 94318
rect 196182 94254 196188 94318
rect 196253 94318 196319 94319
rect 196253 94286 196254 94318
rect 196112 94046 196188 94254
rect 196112 94014 196118 94046
rect 196046 93982 196047 94014
rect 195981 93981 196047 93982
rect 196117 93982 196118 94014
rect 196182 94014 196188 94046
rect 196248 94254 196254 94286
rect 196318 94286 196319 94318
rect 196661 94318 196727 94319
rect 196661 94286 196662 94318
rect 196318 94254 196324 94286
rect 196248 94046 196324 94254
rect 196182 93982 196183 94014
rect 196117 93981 196183 93982
rect 196248 93982 196254 94046
rect 196318 93982 196324 94046
rect 196248 93976 196324 93982
rect 196656 94254 196662 94286
rect 196726 94286 196727 94318
rect 196726 94254 196732 94286
rect 196656 94046 196732 94254
rect 196656 93982 196662 94046
rect 196726 93982 196732 94046
rect 196656 93976 196732 93982
rect 22309 93910 22375 93911
rect 22309 93878 22310 93910
rect 22304 93846 22310 93878
rect 22374 93878 22375 93910
rect 22989 93910 23055 93911
rect 22989 93878 22990 93910
rect 22374 93846 22380 93878
rect 22304 93638 22380 93846
rect 22304 93574 22310 93638
rect 22374 93574 22380 93638
rect 22304 93568 22380 93574
rect 22984 93846 22990 93878
rect 23054 93878 23055 93910
rect 23397 93910 23463 93911
rect 23397 93878 23398 93910
rect 23054 93846 23060 93878
rect 22984 93638 23060 93846
rect 22984 93574 22990 93638
rect 23054 93574 23060 93638
rect 22984 93568 23060 93574
rect 23392 93846 23398 93878
rect 23462 93878 23463 93910
rect 195029 93910 195095 93911
rect 195029 93878 195030 93910
rect 23462 93846 23468 93878
rect 23392 93638 23468 93846
rect 195024 93846 195030 93878
rect 195094 93878 195095 93910
rect 195437 93910 195503 93911
rect 195437 93878 195438 93910
rect 195094 93846 195100 93878
rect 23392 93574 23398 93638
rect 23462 93574 23468 93638
rect 23392 93568 23468 93574
rect 28288 93774 28364 93780
rect 28288 93710 28294 93774
rect 28358 93710 28364 93774
rect 22989 93502 23055 93503
rect 22989 93470 22990 93502
rect 22984 93438 22990 93470
rect 23054 93470 23055 93502
rect 23528 93502 23604 93508
rect 23054 93438 23060 93470
rect 22984 93230 23060 93438
rect 22984 93166 22990 93230
rect 23054 93166 23060 93230
rect 23528 93438 23534 93502
rect 23598 93438 23604 93502
rect 28288 93502 28364 93710
rect 195024 93638 195100 93846
rect 195024 93574 195030 93638
rect 195094 93574 195100 93638
rect 195024 93568 195100 93574
rect 195432 93846 195438 93878
rect 195502 93878 195503 93910
rect 195981 93910 196047 93911
rect 195981 93878 195982 93910
rect 195502 93846 195508 93878
rect 195432 93638 195508 93846
rect 195432 93574 195438 93638
rect 195502 93574 195508 93638
rect 195432 93568 195508 93574
rect 195976 93846 195982 93878
rect 196046 93878 196047 93910
rect 196046 93846 196052 93878
rect 195976 93638 196052 93846
rect 195976 93574 195982 93638
rect 196046 93574 196052 93638
rect 195976 93568 196052 93574
rect 28288 93470 28294 93502
rect 23528 93230 23604 93438
rect 28293 93438 28294 93470
rect 28358 93470 28364 93502
rect 195165 93502 195231 93503
rect 195165 93470 195166 93502
rect 28358 93438 28359 93470
rect 28293 93437 28359 93438
rect 195160 93438 195166 93470
rect 195230 93470 195231 93502
rect 195568 93502 195644 93508
rect 195230 93438 195236 93470
rect 23528 93198 23534 93230
rect 22984 93160 23060 93166
rect 23533 93166 23534 93198
rect 23598 93198 23604 93230
rect 195160 93230 195236 93438
rect 23598 93166 23599 93198
rect 23533 93165 23599 93166
rect 195160 93166 195166 93230
rect 195230 93166 195236 93230
rect 195568 93438 195574 93502
rect 195638 93438 195644 93502
rect 195568 93230 195644 93438
rect 195568 93198 195574 93230
rect 195160 93160 195236 93166
rect 195573 93166 195574 93198
rect 195638 93198 195644 93230
rect 195638 93166 195639 93198
rect 195573 93165 195639 93166
rect 23125 93094 23191 93095
rect 23125 93062 23126 93094
rect 23120 93030 23126 93062
rect 23190 93062 23191 93094
rect 23392 93094 23468 93100
rect 23190 93030 23196 93062
rect 952 92758 1230 92822
rect 1294 92758 1300 92822
rect 21901 92822 21967 92823
rect 21901 92790 21902 92822
rect 952 91190 1300 92758
rect 21896 92758 21902 92790
rect 21966 92790 21967 92822
rect 23120 92822 23196 93030
rect 21966 92758 21972 92790
rect 21896 92550 21972 92758
rect 23120 92758 23126 92822
rect 23190 92758 23196 92822
rect 23392 93030 23398 93094
rect 23462 93030 23468 93094
rect 23392 92822 23468 93030
rect 195024 93094 195100 93100
rect 195024 93030 195030 93094
rect 195094 93030 195100 93094
rect 195573 93094 195639 93095
rect 195573 93062 195574 93094
rect 190269 92958 190335 92959
rect 190269 92926 190270 92958
rect 23392 92790 23398 92822
rect 23120 92752 23196 92758
rect 23397 92758 23398 92790
rect 23462 92790 23468 92822
rect 190264 92894 190270 92926
rect 190334 92926 190335 92958
rect 190334 92894 190340 92926
rect 23462 92758 23463 92790
rect 23397 92757 23463 92758
rect 190264 92686 190340 92894
rect 195024 92822 195100 93030
rect 195024 92790 195030 92822
rect 195029 92758 195030 92790
rect 195094 92790 195100 92822
rect 195568 93030 195574 93062
rect 195638 93062 195639 93094
rect 195638 93030 195644 93062
rect 195568 92822 195644 93030
rect 217464 92958 217812 94526
rect 217464 92894 217470 92958
rect 217534 92894 217812 92958
rect 195094 92758 195095 92790
rect 195029 92757 195095 92758
rect 195568 92758 195574 92822
rect 195638 92758 195644 92822
rect 196797 92822 196863 92823
rect 196797 92790 196798 92822
rect 195568 92752 195644 92758
rect 196792 92758 196798 92790
rect 196862 92790 196863 92822
rect 196862 92758 196868 92790
rect 190264 92622 190270 92686
rect 190334 92622 190340 92686
rect 190264 92616 190340 92622
rect 21896 92486 21902 92550
rect 21966 92486 21972 92550
rect 28565 92550 28631 92551
rect 28565 92518 28566 92550
rect 21896 92480 21972 92486
rect 28560 92486 28566 92518
rect 28630 92518 28631 92550
rect 190128 92550 190204 92556
rect 28630 92486 28636 92518
rect 21760 92414 21836 92420
rect 21760 92350 21766 92414
rect 21830 92350 21836 92414
rect 22445 92414 22511 92415
rect 22445 92382 22446 92414
rect 21760 92142 21836 92350
rect 21760 92110 21766 92142
rect 21765 92078 21766 92110
rect 21830 92110 21836 92142
rect 22440 92350 22446 92382
rect 22510 92382 22511 92414
rect 22510 92350 22516 92382
rect 22440 92142 22516 92350
rect 28560 92278 28636 92486
rect 28560 92214 28566 92278
rect 28630 92214 28636 92278
rect 190128 92486 190134 92550
rect 190198 92486 190204 92550
rect 190128 92278 190204 92486
rect 196792 92550 196868 92758
rect 196792 92486 196798 92550
rect 196862 92486 196868 92550
rect 196792 92480 196868 92486
rect 196117 92414 196183 92415
rect 196117 92382 196118 92414
rect 190128 92246 190134 92278
rect 28560 92208 28636 92214
rect 190133 92214 190134 92246
rect 190198 92246 190204 92278
rect 196112 92350 196118 92382
rect 196182 92382 196183 92414
rect 196661 92414 196727 92415
rect 196661 92382 196662 92414
rect 196182 92350 196188 92382
rect 190198 92214 190199 92246
rect 190133 92213 190199 92214
rect 21830 92078 21831 92110
rect 21765 92077 21831 92078
rect 22440 92078 22446 92142
rect 22510 92078 22516 92142
rect 22440 92072 22516 92078
rect 196112 92142 196188 92350
rect 196112 92078 196118 92142
rect 196182 92078 196188 92142
rect 196112 92072 196188 92078
rect 196656 92350 196662 92382
rect 196726 92382 196727 92414
rect 196726 92350 196732 92382
rect 196656 92142 196732 92350
rect 196656 92078 196662 92142
rect 196726 92078 196732 92142
rect 196656 92072 196732 92078
rect 21765 92006 21831 92007
rect 21765 91974 21766 92006
rect 21760 91942 21766 91974
rect 21830 91974 21831 92006
rect 22984 92006 23060 92012
rect 21830 91942 21836 91974
rect 21760 91734 21836 91942
rect 22984 91942 22990 92006
rect 23054 91942 23060 92006
rect 23533 92006 23599 92007
rect 23533 91974 23534 92006
rect 21760 91670 21766 91734
rect 21830 91670 21836 91734
rect 21760 91664 21836 91670
rect 22440 91870 22516 91876
rect 22440 91806 22446 91870
rect 22510 91806 22516 91870
rect 21901 91598 21967 91599
rect 21901 91566 21902 91598
rect 21896 91534 21902 91566
rect 21966 91566 21967 91598
rect 22440 91598 22516 91806
rect 22984 91734 23060 91942
rect 22984 91702 22990 91734
rect 22989 91670 22990 91702
rect 23054 91702 23060 91734
rect 23528 91942 23534 91974
rect 23598 91974 23599 92006
rect 195165 92006 195231 92007
rect 195165 91974 195166 92006
rect 23598 91942 23604 91974
rect 23528 91734 23604 91942
rect 23054 91670 23055 91702
rect 22989 91669 23055 91670
rect 23528 91670 23534 91734
rect 23598 91670 23604 91734
rect 23528 91664 23604 91670
rect 195160 91942 195166 91974
rect 195230 91974 195231 92006
rect 195432 92006 195508 92012
rect 195230 91942 195236 91974
rect 195160 91734 195236 91942
rect 195160 91670 195166 91734
rect 195230 91670 195236 91734
rect 195432 91942 195438 92006
rect 195502 91942 195508 92006
rect 195432 91734 195508 91942
rect 195432 91702 195438 91734
rect 195160 91664 195236 91670
rect 195437 91670 195438 91702
rect 195502 91702 195508 91734
rect 196792 92006 196868 92012
rect 196792 91942 196798 92006
rect 196862 91942 196868 92006
rect 196792 91734 196868 91942
rect 196792 91702 196798 91734
rect 195502 91670 195503 91702
rect 195437 91669 195503 91670
rect 196797 91670 196798 91702
rect 196862 91702 196868 91734
rect 196862 91670 196863 91702
rect 196797 91669 196863 91670
rect 22440 91566 22446 91598
rect 21966 91534 21972 91566
rect 21896 91326 21972 91534
rect 22445 91534 22446 91566
rect 22510 91566 22516 91598
rect 22717 91598 22783 91599
rect 22717 91566 22718 91598
rect 22510 91534 22511 91566
rect 22445 91533 22511 91534
rect 22712 91534 22718 91566
rect 22782 91566 22783 91598
rect 23125 91598 23191 91599
rect 23125 91566 23126 91598
rect 22782 91534 22788 91566
rect 21896 91262 21902 91326
rect 21966 91262 21972 91326
rect 21896 91256 21972 91262
rect 22712 91326 22788 91534
rect 22712 91262 22718 91326
rect 22782 91262 22788 91326
rect 22712 91256 22788 91262
rect 23120 91534 23126 91566
rect 23190 91566 23191 91598
rect 23528 91598 23604 91604
rect 23190 91534 23196 91566
rect 23120 91326 23196 91534
rect 23120 91262 23126 91326
rect 23190 91262 23196 91326
rect 23528 91534 23534 91598
rect 23598 91534 23604 91598
rect 195029 91598 195095 91599
rect 195029 91566 195030 91598
rect 23528 91326 23604 91534
rect 23528 91294 23534 91326
rect 23120 91256 23196 91262
rect 23533 91262 23534 91294
rect 23598 91294 23604 91326
rect 195024 91534 195030 91566
rect 195094 91566 195095 91598
rect 195437 91598 195503 91599
rect 195437 91566 195438 91598
rect 195094 91534 195100 91566
rect 195024 91326 195100 91534
rect 23598 91262 23599 91294
rect 23533 91261 23599 91262
rect 195024 91262 195030 91326
rect 195094 91262 195100 91326
rect 195024 91256 195100 91262
rect 195432 91534 195438 91566
rect 195502 91566 195503 91598
rect 196248 91598 196324 91604
rect 195502 91534 195508 91566
rect 195432 91326 195508 91534
rect 195432 91262 195438 91326
rect 195502 91262 195508 91326
rect 196248 91534 196254 91598
rect 196318 91534 196324 91598
rect 196248 91326 196324 91534
rect 196248 91294 196254 91326
rect 195432 91256 195508 91262
rect 196253 91262 196254 91294
rect 196318 91294 196324 91326
rect 196656 91598 196732 91604
rect 196656 91534 196662 91598
rect 196726 91534 196732 91598
rect 196656 91326 196732 91534
rect 196656 91294 196662 91326
rect 196318 91262 196319 91294
rect 196253 91261 196319 91262
rect 196661 91262 196662 91294
rect 196726 91294 196732 91326
rect 217464 91326 217812 92894
rect 196726 91262 196727 91294
rect 196661 91261 196727 91262
rect 217464 91262 217470 91326
rect 217534 91262 217812 91326
rect 952 91126 1230 91190
rect 1294 91126 1300 91190
rect 952 89558 1300 91126
rect 21760 91190 21836 91196
rect 21760 91126 21766 91190
rect 21830 91126 21836 91190
rect 21760 90918 21836 91126
rect 21760 90886 21766 90918
rect 21765 90854 21766 90886
rect 21830 90886 21836 90918
rect 22168 91190 22244 91196
rect 22168 91126 22174 91190
rect 22238 91126 22244 91190
rect 22168 90918 22244 91126
rect 22168 90886 22174 90918
rect 21830 90854 21831 90886
rect 21765 90853 21831 90854
rect 22173 90854 22174 90886
rect 22238 90886 22244 90918
rect 22576 91190 22652 91196
rect 22576 91126 22582 91190
rect 22646 91126 22652 91190
rect 22989 91190 23055 91191
rect 22989 91158 22990 91190
rect 22576 90918 22652 91126
rect 22576 90886 22582 90918
rect 22238 90854 22239 90886
rect 22173 90853 22239 90854
rect 22581 90854 22582 90886
rect 22646 90886 22652 90918
rect 22984 91126 22990 91158
rect 23054 91158 23055 91190
rect 23528 91190 23604 91196
rect 23054 91126 23060 91158
rect 22984 90918 23060 91126
rect 22646 90854 22647 90886
rect 22581 90853 22647 90854
rect 22984 90854 22990 90918
rect 23054 90854 23060 90918
rect 23528 91126 23534 91190
rect 23598 91126 23604 91190
rect 23528 90918 23604 91126
rect 23528 90886 23534 90918
rect 22984 90848 23060 90854
rect 23533 90854 23534 90886
rect 23598 90886 23604 90918
rect 195160 91190 195236 91196
rect 195160 91126 195166 91190
rect 195230 91126 195236 91190
rect 195160 90918 195236 91126
rect 195160 90886 195166 90918
rect 23598 90854 23599 90886
rect 23533 90853 23599 90854
rect 195165 90854 195166 90886
rect 195230 90886 195236 90918
rect 195568 91190 195644 91196
rect 195568 91126 195574 91190
rect 195638 91126 195644 91190
rect 195845 91190 195911 91191
rect 195845 91158 195846 91190
rect 195568 90918 195644 91126
rect 195568 90886 195574 90918
rect 195230 90854 195231 90886
rect 195165 90853 195231 90854
rect 195573 90854 195574 90886
rect 195638 90886 195644 90918
rect 195840 91126 195846 91158
rect 195910 91158 195911 91190
rect 196661 91190 196727 91191
rect 196661 91158 196662 91190
rect 195910 91126 195916 91158
rect 195840 90918 195916 91126
rect 195638 90854 195639 90886
rect 195573 90853 195639 90854
rect 195840 90854 195846 90918
rect 195910 90854 195916 90918
rect 195840 90848 195916 90854
rect 196656 91126 196662 91158
rect 196726 91158 196727 91190
rect 196726 91126 196732 91158
rect 196656 90918 196732 91126
rect 196656 90854 196662 90918
rect 196726 90854 196732 90918
rect 196656 90848 196732 90854
rect 21896 90782 21972 90788
rect 21896 90718 21902 90782
rect 21966 90718 21972 90782
rect 22717 90782 22783 90783
rect 22717 90750 22718 90782
rect 21896 90510 21972 90718
rect 21896 90478 21902 90510
rect 21901 90446 21902 90478
rect 21966 90478 21972 90510
rect 22712 90718 22718 90750
rect 22782 90750 22783 90782
rect 23120 90782 23196 90788
rect 22782 90718 22788 90750
rect 22712 90510 22788 90718
rect 21966 90446 21967 90478
rect 21901 90445 21967 90446
rect 22712 90446 22718 90510
rect 22782 90446 22788 90510
rect 23120 90718 23126 90782
rect 23190 90718 23196 90782
rect 23397 90782 23463 90783
rect 23397 90750 23398 90782
rect 23120 90510 23196 90718
rect 23120 90478 23126 90510
rect 22712 90440 22788 90446
rect 23125 90446 23126 90478
rect 23190 90478 23196 90510
rect 23392 90718 23398 90750
rect 23462 90750 23463 90782
rect 195029 90782 195095 90783
rect 195029 90750 195030 90782
rect 23462 90718 23468 90750
rect 23392 90510 23468 90718
rect 23190 90446 23191 90478
rect 23125 90445 23191 90446
rect 23392 90446 23398 90510
rect 23462 90446 23468 90510
rect 23392 90440 23468 90446
rect 195024 90718 195030 90750
rect 195094 90750 195095 90782
rect 195568 90782 195644 90788
rect 195094 90718 195100 90750
rect 195024 90510 195100 90718
rect 195024 90446 195030 90510
rect 195094 90446 195100 90510
rect 195568 90718 195574 90782
rect 195638 90718 195644 90782
rect 195568 90510 195644 90718
rect 195568 90478 195574 90510
rect 195024 90440 195100 90446
rect 195573 90446 195574 90478
rect 195638 90478 195644 90510
rect 196112 90782 196188 90788
rect 196112 90718 196118 90782
rect 196182 90718 196188 90782
rect 196112 90510 196188 90718
rect 196112 90478 196118 90510
rect 195638 90446 195639 90478
rect 195573 90445 195639 90446
rect 196117 90446 196118 90478
rect 196182 90478 196188 90510
rect 196792 90782 196868 90788
rect 196792 90718 196798 90782
rect 196862 90718 196868 90782
rect 196792 90510 196868 90718
rect 196792 90478 196798 90510
rect 196182 90446 196183 90478
rect 196117 90445 196183 90446
rect 196797 90446 196798 90478
rect 196862 90478 196868 90510
rect 196862 90446 196863 90478
rect 196797 90445 196863 90446
rect 21901 90374 21967 90375
rect 21901 90342 21902 90374
rect 21896 90310 21902 90342
rect 21966 90342 21967 90374
rect 22309 90374 22375 90375
rect 22309 90342 22310 90374
rect 21966 90310 21972 90342
rect 21896 90102 21972 90310
rect 21896 90038 21902 90102
rect 21966 90038 21972 90102
rect 21896 90032 21972 90038
rect 22304 90310 22310 90342
rect 22374 90342 22375 90374
rect 22984 90374 23060 90380
rect 22374 90310 22380 90342
rect 22304 90102 22380 90310
rect 22304 90038 22310 90102
rect 22374 90038 22380 90102
rect 22984 90310 22990 90374
rect 23054 90310 23060 90374
rect 22984 90102 23060 90310
rect 22984 90070 22990 90102
rect 22304 90032 22380 90038
rect 22989 90038 22990 90070
rect 23054 90070 23060 90102
rect 23528 90374 23604 90380
rect 23528 90310 23534 90374
rect 23598 90310 23604 90374
rect 195029 90374 195095 90375
rect 195029 90342 195030 90374
rect 23528 90102 23604 90310
rect 23528 90070 23534 90102
rect 23054 90038 23055 90070
rect 22989 90037 23055 90038
rect 23533 90038 23534 90070
rect 23598 90070 23604 90102
rect 195024 90310 195030 90342
rect 195094 90342 195095 90374
rect 195573 90374 195639 90375
rect 195573 90342 195574 90374
rect 195094 90310 195100 90342
rect 195024 90102 195100 90310
rect 23598 90038 23599 90070
rect 23533 90037 23599 90038
rect 195024 90038 195030 90102
rect 195094 90038 195100 90102
rect 195024 90032 195100 90038
rect 195568 90310 195574 90342
rect 195638 90342 195639 90374
rect 195840 90374 195916 90380
rect 195638 90310 195644 90342
rect 195568 90102 195644 90310
rect 195568 90038 195574 90102
rect 195638 90038 195644 90102
rect 195840 90310 195846 90374
rect 195910 90310 195916 90374
rect 196797 90374 196863 90375
rect 196797 90342 196798 90374
rect 195840 90102 195916 90310
rect 195840 90070 195846 90102
rect 195568 90032 195644 90038
rect 195845 90038 195846 90070
rect 195910 90070 195916 90102
rect 196792 90310 196798 90342
rect 196862 90342 196863 90374
rect 196862 90310 196868 90342
rect 196792 90102 196868 90310
rect 195910 90038 195911 90070
rect 195845 90037 195911 90038
rect 196792 90038 196798 90102
rect 196862 90038 196868 90102
rect 196792 90032 196868 90038
rect 22173 89966 22239 89967
rect 22173 89934 22174 89966
rect 22168 89902 22174 89934
rect 22238 89934 22239 89966
rect 22712 89966 22788 89972
rect 22238 89902 22244 89934
rect 22168 89694 22244 89902
rect 22168 89630 22174 89694
rect 22238 89630 22244 89694
rect 22712 89902 22718 89966
rect 22782 89902 22788 89966
rect 22989 89966 23055 89967
rect 22989 89934 22990 89966
rect 22712 89694 22788 89902
rect 22712 89662 22718 89694
rect 22168 89624 22244 89630
rect 22717 89630 22718 89662
rect 22782 89662 22788 89694
rect 22984 89902 22990 89934
rect 23054 89934 23055 89966
rect 23533 89966 23599 89967
rect 23533 89934 23534 89966
rect 23054 89902 23060 89934
rect 22984 89694 23060 89902
rect 22782 89630 22783 89662
rect 22717 89629 22783 89630
rect 22984 89630 22990 89694
rect 23054 89630 23060 89694
rect 22984 89624 23060 89630
rect 23528 89902 23534 89934
rect 23598 89934 23599 89966
rect 195024 89966 195100 89972
rect 23598 89902 23604 89934
rect 23528 89694 23604 89902
rect 195024 89902 195030 89966
rect 195094 89902 195100 89966
rect 28565 89830 28631 89831
rect 28565 89798 28566 89830
rect 23528 89630 23534 89694
rect 23598 89630 23604 89694
rect 23528 89624 23604 89630
rect 28560 89766 28566 89798
rect 28630 89798 28631 89830
rect 28630 89766 28636 89798
rect 952 89494 1230 89558
rect 1294 89494 1300 89558
rect 952 87926 1300 89494
rect 23120 89558 23196 89564
rect 23120 89494 23126 89558
rect 23190 89494 23196 89558
rect 23120 89286 23196 89494
rect 23120 89254 23126 89286
rect 23125 89222 23126 89254
rect 23190 89254 23196 89286
rect 23392 89558 23468 89564
rect 23392 89494 23398 89558
rect 23462 89494 23468 89558
rect 23392 89286 23468 89494
rect 28560 89558 28636 89766
rect 195024 89694 195100 89902
rect 195024 89662 195030 89694
rect 195029 89630 195030 89662
rect 195094 89662 195100 89694
rect 195432 89966 195508 89972
rect 195432 89902 195438 89966
rect 195502 89902 195508 89966
rect 195432 89694 195508 89902
rect 195432 89662 195438 89694
rect 195094 89630 195095 89662
rect 195029 89629 195095 89630
rect 195437 89630 195438 89662
rect 195502 89662 195508 89694
rect 195976 89966 196052 89972
rect 195976 89902 195982 89966
rect 196046 89902 196052 89966
rect 195976 89694 196052 89902
rect 195976 89662 195982 89694
rect 195502 89630 195503 89662
rect 195437 89629 195503 89630
rect 195981 89630 195982 89662
rect 196046 89662 196052 89694
rect 196112 89966 196188 89972
rect 196112 89902 196118 89966
rect 196182 89902 196188 89966
rect 196112 89694 196188 89902
rect 196112 89662 196118 89694
rect 196046 89630 196047 89662
rect 195981 89629 196047 89630
rect 196117 89630 196118 89662
rect 196182 89662 196188 89694
rect 217464 89694 217812 91262
rect 196182 89630 196183 89662
rect 196117 89629 196183 89630
rect 217464 89630 217470 89694
rect 217534 89630 217812 89694
rect 28560 89494 28566 89558
rect 28630 89494 28636 89558
rect 28560 89488 28636 89494
rect 195024 89558 195100 89564
rect 195024 89494 195030 89558
rect 195094 89494 195100 89558
rect 195437 89558 195503 89559
rect 195437 89526 195438 89558
rect 23392 89254 23398 89286
rect 23190 89222 23191 89254
rect 23125 89221 23191 89222
rect 23397 89222 23398 89254
rect 23462 89254 23468 89286
rect 195024 89286 195100 89494
rect 195024 89254 195030 89286
rect 23462 89222 23463 89254
rect 23397 89221 23463 89222
rect 195029 89222 195030 89254
rect 195094 89254 195100 89286
rect 195432 89494 195438 89526
rect 195502 89526 195503 89558
rect 195502 89494 195508 89526
rect 195432 89286 195508 89494
rect 195094 89222 195095 89254
rect 195029 89221 195095 89222
rect 195432 89222 195438 89286
rect 195502 89222 195508 89286
rect 195432 89216 195508 89222
rect 22173 89150 22239 89151
rect 22173 89118 22174 89150
rect 22168 89086 22174 89118
rect 22238 89118 22239 89150
rect 23120 89150 23196 89156
rect 22238 89086 22244 89118
rect 21896 88878 21972 88884
rect 21896 88814 21902 88878
rect 21966 88814 21972 88878
rect 21896 88606 21972 88814
rect 22168 88878 22244 89086
rect 22168 88814 22174 88878
rect 22238 88814 22244 88878
rect 23120 89086 23126 89150
rect 23190 89086 23196 89150
rect 23120 88878 23196 89086
rect 23120 88846 23126 88878
rect 22168 88808 22244 88814
rect 23125 88814 23126 88846
rect 23190 88846 23196 88878
rect 23528 89150 23604 89156
rect 23528 89086 23534 89150
rect 23598 89086 23604 89150
rect 195165 89150 195231 89151
rect 195165 89118 195166 89150
rect 23528 88878 23604 89086
rect 195160 89086 195166 89118
rect 195230 89118 195231 89150
rect 195437 89150 195503 89151
rect 195437 89118 195438 89150
rect 195230 89086 195236 89118
rect 23528 88846 23534 88878
rect 23190 88814 23191 88846
rect 23125 88813 23191 88814
rect 23533 88814 23534 88846
rect 23598 88846 23604 88878
rect 190128 89014 190204 89020
rect 190128 88950 190134 89014
rect 190198 88950 190204 89014
rect 23598 88814 23599 88846
rect 23533 88813 23599 88814
rect 190128 88742 190204 88950
rect 195160 88878 195236 89086
rect 195160 88814 195166 88878
rect 195230 88814 195236 88878
rect 195160 88808 195236 88814
rect 195432 89086 195438 89118
rect 195502 89118 195503 89150
rect 195981 89150 196047 89151
rect 195981 89118 195982 89150
rect 195502 89086 195508 89118
rect 195432 88878 195508 89086
rect 195432 88814 195438 88878
rect 195502 88814 195508 88878
rect 195432 88808 195508 88814
rect 195976 89086 195982 89118
rect 196046 89118 196047 89150
rect 196248 89150 196324 89156
rect 196046 89086 196052 89118
rect 195976 88878 196052 89086
rect 195976 88814 195982 88878
rect 196046 88814 196052 88878
rect 196248 89086 196254 89150
rect 196318 89086 196324 89150
rect 196248 88878 196324 89086
rect 196248 88846 196254 88878
rect 195976 88808 196052 88814
rect 196253 88814 196254 88846
rect 196318 88846 196324 88878
rect 196661 88878 196727 88879
rect 196661 88846 196662 88878
rect 196318 88814 196319 88846
rect 196253 88813 196319 88814
rect 196656 88814 196662 88846
rect 196726 88846 196727 88878
rect 196726 88814 196732 88846
rect 190128 88710 190134 88742
rect 190133 88678 190134 88710
rect 190198 88710 190204 88742
rect 190269 88742 190335 88743
rect 190269 88710 190270 88742
rect 190198 88678 190199 88710
rect 190133 88677 190199 88678
rect 190264 88678 190270 88710
rect 190334 88710 190335 88742
rect 190334 88678 190340 88710
rect 21896 88574 21902 88606
rect 21901 88542 21902 88574
rect 21966 88574 21972 88606
rect 28429 88606 28495 88607
rect 28429 88574 28430 88606
rect 21966 88542 21967 88574
rect 21901 88541 21967 88542
rect 28424 88542 28430 88574
rect 28494 88574 28495 88606
rect 28494 88542 28500 88574
rect 21901 88470 21967 88471
rect 21901 88438 21902 88470
rect 21896 88406 21902 88438
rect 21966 88438 21967 88470
rect 22168 88470 22244 88476
rect 21966 88406 21972 88438
rect 21896 88198 21972 88406
rect 21896 88134 21902 88198
rect 21966 88134 21972 88198
rect 22168 88406 22174 88470
rect 22238 88406 22244 88470
rect 22168 88198 22244 88406
rect 22168 88166 22174 88198
rect 21896 88128 21972 88134
rect 22173 88134 22174 88166
rect 22238 88166 22244 88198
rect 22440 88470 22516 88476
rect 22440 88406 22446 88470
rect 22510 88406 22516 88470
rect 22440 88198 22516 88406
rect 28424 88334 28500 88542
rect 28424 88270 28430 88334
rect 28494 88270 28500 88334
rect 28424 88264 28500 88270
rect 190264 88334 190340 88678
rect 196656 88606 196732 88814
rect 196656 88542 196662 88606
rect 196726 88542 196732 88606
rect 196656 88536 196732 88542
rect 196117 88470 196183 88471
rect 196117 88438 196118 88470
rect 190264 88270 190270 88334
rect 190334 88270 190340 88334
rect 190264 88264 190340 88270
rect 196112 88406 196118 88438
rect 196182 88438 196183 88470
rect 196792 88470 196868 88476
rect 196182 88406 196188 88438
rect 22440 88166 22446 88198
rect 22238 88134 22239 88166
rect 22173 88133 22239 88134
rect 22445 88134 22446 88166
rect 22510 88166 22516 88198
rect 28565 88198 28631 88199
rect 28565 88166 28566 88198
rect 22510 88134 22511 88166
rect 22445 88133 22511 88134
rect 28560 88134 28566 88166
rect 28630 88166 28631 88198
rect 196112 88198 196188 88406
rect 28630 88134 28636 88166
rect 952 87862 1230 87926
rect 1294 87862 1300 87926
rect 952 86294 1300 87862
rect 21760 88062 21836 88068
rect 21760 87998 21766 88062
rect 21830 87998 21836 88062
rect 21760 87790 21836 87998
rect 28560 87926 28636 88134
rect 196112 88134 196118 88198
rect 196182 88134 196188 88198
rect 196792 88406 196798 88470
rect 196862 88406 196868 88470
rect 196792 88198 196868 88406
rect 196792 88166 196798 88198
rect 196112 88128 196188 88134
rect 196797 88134 196798 88166
rect 196862 88166 196868 88198
rect 196862 88134 196863 88166
rect 196797 88133 196863 88134
rect 196656 88062 196732 88068
rect 196656 87998 196662 88062
rect 196726 87998 196732 88062
rect 28560 87862 28566 87926
rect 28630 87862 28636 87926
rect 28560 87856 28636 87862
rect 190128 87926 190204 87932
rect 190128 87862 190134 87926
rect 190198 87862 190204 87926
rect 21760 87758 21766 87790
rect 21765 87726 21766 87758
rect 21830 87758 21836 87790
rect 21830 87726 21831 87758
rect 21765 87725 21831 87726
rect 21765 87654 21831 87655
rect 21765 87622 21766 87654
rect 21760 87590 21766 87622
rect 21830 87622 21831 87654
rect 22304 87654 22380 87660
rect 21830 87590 21836 87622
rect 21760 87382 21836 87590
rect 21760 87318 21766 87382
rect 21830 87318 21836 87382
rect 22304 87590 22310 87654
rect 22374 87590 22380 87654
rect 22304 87382 22380 87590
rect 22304 87350 22310 87382
rect 21760 87312 21836 87318
rect 22309 87318 22310 87350
rect 22374 87350 22380 87382
rect 22440 87654 22516 87660
rect 22440 87590 22446 87654
rect 22510 87590 22516 87654
rect 22581 87654 22647 87655
rect 22581 87622 22582 87654
rect 22440 87382 22516 87590
rect 22440 87350 22446 87382
rect 22374 87318 22375 87350
rect 22309 87317 22375 87318
rect 22445 87318 22446 87350
rect 22510 87350 22516 87382
rect 22576 87590 22582 87622
rect 22646 87622 22647 87654
rect 23125 87654 23191 87655
rect 23125 87622 23126 87654
rect 22646 87590 22652 87622
rect 22576 87382 22652 87590
rect 22510 87318 22511 87350
rect 22445 87317 22511 87318
rect 22576 87318 22582 87382
rect 22646 87318 22652 87382
rect 22576 87312 22652 87318
rect 23120 87590 23126 87622
rect 23190 87622 23191 87654
rect 23533 87654 23599 87655
rect 23533 87622 23534 87654
rect 23190 87590 23196 87622
rect 23120 87382 23196 87590
rect 23120 87318 23126 87382
rect 23190 87318 23196 87382
rect 23120 87312 23196 87318
rect 23528 87590 23534 87622
rect 23598 87622 23599 87654
rect 190128 87654 190204 87862
rect 196656 87790 196732 87998
rect 196656 87758 196662 87790
rect 196661 87726 196662 87758
rect 196726 87758 196732 87790
rect 217464 87790 217812 89630
rect 196726 87726 196727 87758
rect 196661 87725 196727 87726
rect 217464 87726 217470 87790
rect 217534 87726 217812 87790
rect 190128 87622 190134 87654
rect 23598 87590 23604 87622
rect 23528 87382 23604 87590
rect 190133 87590 190134 87622
rect 190198 87622 190204 87654
rect 195024 87654 195100 87660
rect 190198 87590 190199 87622
rect 190133 87589 190199 87590
rect 195024 87590 195030 87654
rect 195094 87590 195100 87654
rect 195573 87654 195639 87655
rect 195573 87622 195574 87654
rect 23528 87318 23534 87382
rect 23598 87318 23604 87382
rect 23528 87312 23604 87318
rect 28424 87382 28500 87388
rect 28424 87318 28430 87382
rect 28494 87318 28500 87382
rect 21760 87246 21836 87252
rect 21760 87182 21766 87246
rect 21830 87182 21836 87246
rect 21760 86974 21836 87182
rect 21760 86942 21766 86974
rect 21765 86910 21766 86942
rect 21830 86942 21836 86974
rect 22168 87246 22244 87252
rect 22168 87182 22174 87246
rect 22238 87182 22244 87246
rect 22445 87246 22511 87247
rect 22445 87214 22446 87246
rect 22168 86974 22244 87182
rect 22168 86942 22174 86974
rect 21830 86910 21831 86942
rect 21765 86909 21831 86910
rect 22173 86910 22174 86942
rect 22238 86942 22244 86974
rect 22440 87182 22446 87214
rect 22510 87214 22511 87246
rect 22984 87246 23060 87252
rect 22510 87182 22516 87214
rect 22440 86974 22516 87182
rect 22238 86910 22239 86942
rect 22173 86909 22239 86910
rect 22440 86910 22446 86974
rect 22510 86910 22516 86974
rect 22984 87182 22990 87246
rect 23054 87182 23060 87246
rect 23397 87246 23463 87247
rect 23397 87214 23398 87246
rect 22984 86974 23060 87182
rect 22984 86942 22990 86974
rect 22440 86904 22516 86910
rect 22989 86910 22990 86942
rect 23054 86942 23060 86974
rect 23392 87182 23398 87214
rect 23462 87214 23463 87246
rect 23462 87182 23468 87214
rect 23392 86974 23468 87182
rect 28424 87110 28500 87318
rect 28424 87078 28430 87110
rect 28429 87046 28430 87078
rect 28494 87078 28500 87110
rect 190264 87382 190340 87388
rect 190264 87318 190270 87382
rect 190334 87318 190340 87382
rect 195024 87382 195100 87590
rect 195024 87350 195030 87382
rect 190264 87110 190340 87318
rect 195029 87318 195030 87350
rect 195094 87350 195100 87382
rect 195568 87590 195574 87622
rect 195638 87622 195639 87654
rect 195976 87654 196052 87660
rect 195638 87590 195644 87622
rect 195568 87382 195644 87590
rect 195094 87318 195095 87350
rect 195029 87317 195095 87318
rect 195568 87318 195574 87382
rect 195638 87318 195644 87382
rect 195976 87590 195982 87654
rect 196046 87590 196052 87654
rect 195976 87382 196052 87590
rect 195976 87350 195982 87382
rect 195568 87312 195644 87318
rect 195981 87318 195982 87350
rect 196046 87350 196052 87382
rect 196384 87654 196460 87660
rect 196384 87590 196390 87654
rect 196454 87590 196460 87654
rect 196661 87654 196727 87655
rect 196661 87622 196662 87654
rect 196384 87382 196460 87590
rect 196384 87350 196390 87382
rect 196046 87318 196047 87350
rect 195981 87317 196047 87318
rect 196389 87318 196390 87350
rect 196454 87350 196460 87382
rect 196656 87590 196662 87622
rect 196726 87622 196727 87654
rect 196726 87590 196732 87622
rect 196656 87382 196732 87590
rect 196454 87318 196455 87350
rect 196389 87317 196455 87318
rect 196656 87318 196662 87382
rect 196726 87318 196732 87382
rect 196656 87312 196732 87318
rect 195029 87246 195095 87247
rect 195029 87214 195030 87246
rect 190264 87078 190270 87110
rect 28494 87046 28495 87078
rect 28429 87045 28495 87046
rect 190269 87046 190270 87078
rect 190334 87078 190340 87110
rect 195024 87182 195030 87214
rect 195094 87214 195095 87246
rect 195437 87246 195503 87247
rect 195437 87214 195438 87246
rect 195094 87182 195100 87214
rect 190334 87046 190335 87078
rect 190269 87045 190335 87046
rect 23054 86910 23055 86942
rect 22989 86909 23055 86910
rect 23392 86910 23398 86974
rect 23462 86910 23468 86974
rect 23392 86904 23468 86910
rect 195024 86974 195100 87182
rect 195024 86910 195030 86974
rect 195094 86910 195100 86974
rect 195024 86904 195100 86910
rect 195432 87182 195438 87214
rect 195502 87214 195503 87246
rect 196248 87246 196324 87252
rect 195502 87182 195508 87214
rect 195432 86974 195508 87182
rect 195432 86910 195438 86974
rect 195502 86910 195508 86974
rect 196248 87182 196254 87246
rect 196318 87182 196324 87246
rect 196248 86974 196324 87182
rect 196248 86942 196254 86974
rect 195432 86904 195508 86910
rect 196253 86910 196254 86942
rect 196318 86942 196324 86974
rect 196656 87246 196732 87252
rect 196656 87182 196662 87246
rect 196726 87182 196732 87246
rect 196656 86974 196732 87182
rect 196656 86942 196662 86974
rect 196318 86910 196319 86942
rect 196253 86909 196319 86910
rect 196661 86910 196662 86942
rect 196726 86942 196732 86974
rect 196726 86910 196727 86942
rect 196661 86909 196727 86910
rect 21760 86838 21836 86844
rect 21760 86774 21766 86838
rect 21830 86774 21836 86838
rect 21760 86566 21836 86774
rect 21760 86534 21766 86566
rect 21765 86502 21766 86534
rect 21830 86534 21836 86566
rect 22576 86838 22652 86844
rect 22576 86774 22582 86838
rect 22646 86774 22652 86838
rect 22576 86566 22652 86774
rect 22576 86534 22582 86566
rect 21830 86502 21831 86534
rect 21765 86501 21831 86502
rect 22581 86502 22582 86534
rect 22646 86534 22652 86566
rect 23120 86838 23196 86844
rect 23120 86774 23126 86838
rect 23190 86774 23196 86838
rect 23120 86566 23196 86774
rect 23120 86534 23126 86566
rect 22646 86502 22647 86534
rect 22581 86501 22647 86502
rect 23125 86502 23126 86534
rect 23190 86534 23196 86566
rect 23528 86838 23604 86844
rect 23528 86774 23534 86838
rect 23598 86774 23604 86838
rect 23528 86566 23604 86774
rect 23528 86534 23534 86566
rect 23190 86502 23191 86534
rect 23125 86501 23191 86502
rect 23533 86502 23534 86534
rect 23598 86534 23604 86566
rect 195160 86838 195236 86844
rect 195160 86774 195166 86838
rect 195230 86774 195236 86838
rect 195160 86566 195236 86774
rect 195160 86534 195166 86566
rect 23598 86502 23599 86534
rect 23533 86501 23599 86502
rect 195165 86502 195166 86534
rect 195230 86534 195236 86566
rect 195568 86838 195644 86844
rect 195568 86774 195574 86838
rect 195638 86774 195644 86838
rect 195845 86838 195911 86839
rect 195845 86806 195846 86838
rect 195568 86566 195644 86774
rect 195568 86534 195574 86566
rect 195230 86502 195231 86534
rect 195165 86501 195231 86502
rect 195573 86502 195574 86534
rect 195638 86534 195644 86566
rect 195840 86774 195846 86806
rect 195910 86806 195911 86838
rect 196112 86838 196188 86844
rect 195910 86774 195916 86806
rect 195840 86566 195916 86774
rect 195638 86502 195639 86534
rect 195573 86501 195639 86502
rect 195840 86502 195846 86566
rect 195910 86502 195916 86566
rect 196112 86774 196118 86838
rect 196182 86774 196188 86838
rect 196661 86838 196727 86839
rect 196661 86806 196662 86838
rect 196112 86566 196188 86774
rect 196112 86534 196118 86566
rect 195840 86496 195916 86502
rect 196117 86502 196118 86534
rect 196182 86534 196188 86566
rect 196656 86774 196662 86806
rect 196726 86806 196727 86838
rect 196726 86774 196732 86806
rect 196656 86566 196732 86774
rect 196182 86502 196183 86534
rect 196117 86501 196183 86502
rect 196656 86502 196662 86566
rect 196726 86502 196732 86566
rect 196656 86496 196732 86502
rect 952 86230 1230 86294
rect 1294 86230 1300 86294
rect 952 84526 1300 86230
rect 21896 86430 21972 86436
rect 21896 86366 21902 86430
rect 21966 86366 21972 86430
rect 22309 86430 22375 86431
rect 22309 86398 22310 86430
rect 21896 86158 21972 86366
rect 21896 86126 21902 86158
rect 21901 86094 21902 86126
rect 21966 86126 21972 86158
rect 22304 86366 22310 86398
rect 22374 86398 22375 86430
rect 23120 86430 23196 86436
rect 22374 86366 22380 86398
rect 22304 86158 22380 86366
rect 21966 86094 21967 86126
rect 21901 86093 21967 86094
rect 22304 86094 22310 86158
rect 22374 86094 22380 86158
rect 23120 86366 23126 86430
rect 23190 86366 23196 86430
rect 23120 86158 23196 86366
rect 23120 86126 23126 86158
rect 22304 86088 22380 86094
rect 23125 86094 23126 86126
rect 23190 86126 23196 86158
rect 23392 86430 23468 86436
rect 23392 86366 23398 86430
rect 23462 86366 23468 86430
rect 23392 86158 23468 86366
rect 23392 86126 23398 86158
rect 23190 86094 23191 86126
rect 23125 86093 23191 86094
rect 23397 86094 23398 86126
rect 23462 86126 23468 86158
rect 195024 86430 195100 86436
rect 195024 86366 195030 86430
rect 195094 86366 195100 86430
rect 195437 86430 195503 86431
rect 195437 86398 195438 86430
rect 195024 86158 195100 86366
rect 195024 86126 195030 86158
rect 23462 86094 23463 86126
rect 23397 86093 23463 86094
rect 195029 86094 195030 86126
rect 195094 86126 195100 86158
rect 195432 86366 195438 86398
rect 195502 86398 195503 86430
rect 195981 86430 196047 86431
rect 195981 86398 195982 86430
rect 195502 86366 195508 86398
rect 195432 86158 195508 86366
rect 195094 86094 195095 86126
rect 195029 86093 195095 86094
rect 195432 86094 195438 86158
rect 195502 86094 195508 86158
rect 195432 86088 195508 86094
rect 195976 86366 195982 86398
rect 196046 86398 196047 86430
rect 196117 86430 196183 86431
rect 196117 86398 196118 86430
rect 196046 86366 196052 86398
rect 195976 86158 196052 86366
rect 195976 86094 195982 86158
rect 196046 86094 196052 86158
rect 195976 86088 196052 86094
rect 196112 86366 196118 86398
rect 196182 86398 196183 86430
rect 196792 86430 196868 86436
rect 196182 86366 196188 86398
rect 196112 86158 196188 86366
rect 196112 86094 196118 86158
rect 196182 86094 196188 86158
rect 196792 86366 196798 86430
rect 196862 86366 196868 86430
rect 196792 86158 196868 86366
rect 196792 86126 196798 86158
rect 196112 86088 196188 86094
rect 196797 86094 196798 86126
rect 196862 86126 196868 86158
rect 217464 86158 217812 87726
rect 196862 86094 196863 86126
rect 196797 86093 196863 86094
rect 217464 86094 217470 86158
rect 217534 86094 217812 86158
rect 23125 86022 23191 86023
rect 23125 85990 23126 86022
rect 23120 85958 23126 85990
rect 23190 85990 23191 86022
rect 23397 86022 23463 86023
rect 23397 85990 23398 86022
rect 23190 85958 23196 85990
rect 23120 85750 23196 85958
rect 23120 85686 23126 85750
rect 23190 85686 23196 85750
rect 23120 85680 23196 85686
rect 23392 85958 23398 85990
rect 23462 85990 23463 86022
rect 195029 86022 195095 86023
rect 195029 85990 195030 86022
rect 23462 85958 23468 85990
rect 23392 85750 23468 85958
rect 23392 85686 23398 85750
rect 23462 85686 23468 85750
rect 23392 85680 23468 85686
rect 195024 85958 195030 85990
rect 195094 85990 195095 86022
rect 195573 86022 195639 86023
rect 195573 85990 195574 86022
rect 195094 85958 195100 85990
rect 195024 85750 195100 85958
rect 195024 85686 195030 85750
rect 195094 85686 195100 85750
rect 195024 85680 195100 85686
rect 195568 85958 195574 85990
rect 195638 85990 195639 86022
rect 195840 86022 195916 86028
rect 195638 85958 195644 85990
rect 195568 85750 195644 85958
rect 195568 85686 195574 85750
rect 195638 85686 195644 85750
rect 195840 85958 195846 86022
rect 195910 85958 195916 86022
rect 195840 85750 195916 85958
rect 195840 85718 195846 85750
rect 195568 85680 195644 85686
rect 195845 85686 195846 85718
rect 195910 85718 195916 85750
rect 195910 85686 195911 85718
rect 195845 85685 195911 85686
rect 21896 85614 21972 85620
rect 21896 85550 21902 85614
rect 21966 85550 21972 85614
rect 22173 85614 22239 85615
rect 22173 85582 22174 85614
rect 21896 85342 21972 85550
rect 21896 85310 21902 85342
rect 21901 85278 21902 85310
rect 21966 85310 21972 85342
rect 22168 85550 22174 85582
rect 22238 85582 22239 85614
rect 22581 85614 22647 85615
rect 22581 85582 22582 85614
rect 22238 85550 22244 85582
rect 22168 85342 22244 85550
rect 21966 85278 21967 85310
rect 21901 85277 21967 85278
rect 22168 85278 22174 85342
rect 22238 85278 22244 85342
rect 22168 85272 22244 85278
rect 22576 85550 22582 85582
rect 22646 85582 22647 85614
rect 23125 85614 23191 85615
rect 23125 85582 23126 85614
rect 22646 85550 22652 85582
rect 22576 85342 22652 85550
rect 22576 85278 22582 85342
rect 22646 85278 22652 85342
rect 22576 85272 22652 85278
rect 23120 85550 23126 85582
rect 23190 85582 23191 85614
rect 23392 85614 23468 85620
rect 23190 85550 23196 85582
rect 23120 85342 23196 85550
rect 23120 85278 23126 85342
rect 23190 85278 23196 85342
rect 23392 85550 23398 85614
rect 23462 85550 23468 85614
rect 23392 85342 23468 85550
rect 23392 85310 23398 85342
rect 23120 85272 23196 85278
rect 23397 85278 23398 85310
rect 23462 85310 23468 85342
rect 195024 85614 195100 85620
rect 195024 85550 195030 85614
rect 195094 85550 195100 85614
rect 195024 85342 195100 85550
rect 195024 85310 195030 85342
rect 23462 85278 23463 85310
rect 23397 85277 23463 85278
rect 195029 85278 195030 85310
rect 195094 85310 195100 85342
rect 195432 85614 195508 85620
rect 195432 85550 195438 85614
rect 195502 85550 195508 85614
rect 195432 85342 195508 85550
rect 195432 85310 195438 85342
rect 195094 85278 195095 85310
rect 195029 85277 195095 85278
rect 195437 85278 195438 85310
rect 195502 85310 195508 85342
rect 195976 85614 196052 85620
rect 195976 85550 195982 85614
rect 196046 85550 196052 85614
rect 195976 85342 196052 85550
rect 195976 85310 195982 85342
rect 195502 85278 195503 85310
rect 195437 85277 195503 85278
rect 195981 85278 195982 85310
rect 196046 85310 196052 85342
rect 196792 85614 196868 85620
rect 196792 85550 196798 85614
rect 196862 85550 196868 85614
rect 196792 85342 196868 85550
rect 196792 85310 196798 85342
rect 196046 85278 196047 85310
rect 195981 85277 196047 85278
rect 196797 85278 196798 85310
rect 196862 85310 196868 85342
rect 196862 85278 196863 85310
rect 196797 85277 196863 85278
rect 22309 85206 22375 85207
rect 22309 85174 22310 85206
rect 22304 85142 22310 85174
rect 22374 85174 22375 85206
rect 23120 85206 23196 85212
rect 22374 85142 22380 85174
rect 21901 84934 21967 84935
rect 21901 84902 21902 84934
rect 21896 84870 21902 84902
rect 21966 84902 21967 84934
rect 22304 84934 22380 85142
rect 21966 84870 21972 84902
rect 21896 84662 21972 84870
rect 22304 84870 22310 84934
rect 22374 84870 22380 84934
rect 23120 85142 23126 85206
rect 23190 85142 23196 85206
rect 23120 84934 23196 85142
rect 23120 84902 23126 84934
rect 22304 84864 22380 84870
rect 23125 84870 23126 84902
rect 23190 84902 23196 84934
rect 23392 85206 23468 85212
rect 23392 85142 23398 85206
rect 23462 85142 23468 85206
rect 195029 85206 195095 85207
rect 195029 85174 195030 85206
rect 23392 84934 23468 85142
rect 195024 85142 195030 85174
rect 195094 85174 195095 85206
rect 195568 85206 195644 85212
rect 195094 85142 195100 85174
rect 23392 84902 23398 84934
rect 23190 84870 23191 84902
rect 23125 84869 23191 84870
rect 23397 84870 23398 84902
rect 23462 84902 23468 84934
rect 28288 85070 28364 85076
rect 28288 85006 28294 85070
rect 28358 85006 28364 85070
rect 23462 84870 23463 84902
rect 23397 84869 23463 84870
rect 21896 84598 21902 84662
rect 21966 84598 21972 84662
rect 21896 84592 21972 84598
rect 23120 84798 23196 84804
rect 23120 84734 23126 84798
rect 23190 84734 23196 84798
rect 23533 84798 23599 84799
rect 23533 84766 23534 84798
rect 952 84462 1230 84526
rect 1294 84462 1300 84526
rect 23120 84526 23196 84734
rect 23120 84494 23126 84526
rect 952 82758 1300 84462
rect 23125 84462 23126 84494
rect 23190 84494 23196 84526
rect 23528 84734 23534 84766
rect 23598 84766 23599 84798
rect 28288 84798 28364 85006
rect 195024 84934 195100 85142
rect 195024 84870 195030 84934
rect 195094 84870 195100 84934
rect 195568 85142 195574 85206
rect 195638 85142 195644 85206
rect 196389 85206 196455 85207
rect 196389 85174 196390 85206
rect 195568 84934 195644 85142
rect 195568 84902 195574 84934
rect 195024 84864 195100 84870
rect 195573 84870 195574 84902
rect 195638 84902 195644 84934
rect 196384 85142 196390 85174
rect 196454 85174 196455 85206
rect 196454 85142 196460 85174
rect 196384 84934 196460 85142
rect 195638 84870 195639 84902
rect 195573 84869 195639 84870
rect 196384 84870 196390 84934
rect 196454 84870 196460 84934
rect 196797 84934 196863 84935
rect 196797 84902 196798 84934
rect 196384 84864 196460 84870
rect 196792 84870 196798 84902
rect 196862 84902 196863 84934
rect 196862 84870 196868 84902
rect 28288 84766 28294 84798
rect 23598 84734 23604 84766
rect 23528 84526 23604 84734
rect 28293 84734 28294 84766
rect 28358 84766 28364 84798
rect 195165 84798 195231 84799
rect 195165 84766 195166 84798
rect 28358 84734 28359 84766
rect 28293 84733 28359 84734
rect 195160 84734 195166 84766
rect 195230 84766 195231 84798
rect 195437 84798 195503 84799
rect 195437 84766 195438 84798
rect 195230 84734 195236 84766
rect 23190 84462 23191 84494
rect 23125 84461 23191 84462
rect 23528 84462 23534 84526
rect 23598 84462 23604 84526
rect 23528 84456 23604 84462
rect 28424 84526 28500 84532
rect 28424 84462 28430 84526
rect 28494 84462 28500 84526
rect 22304 84390 22380 84396
rect 22304 84326 22310 84390
rect 22374 84326 22380 84390
rect 21896 84118 21972 84124
rect 21896 84054 21902 84118
rect 21966 84054 21972 84118
rect 22304 84118 22380 84326
rect 22304 84086 22310 84118
rect 21896 83846 21972 84054
rect 22309 84054 22310 84086
rect 22374 84086 22380 84118
rect 22440 84390 22516 84396
rect 22440 84326 22446 84390
rect 22510 84326 22516 84390
rect 22440 84118 22516 84326
rect 28424 84254 28500 84462
rect 195160 84526 195236 84734
rect 195160 84462 195166 84526
rect 195230 84462 195236 84526
rect 195160 84456 195236 84462
rect 195432 84734 195438 84766
rect 195502 84766 195503 84798
rect 195502 84734 195508 84766
rect 195432 84526 195508 84734
rect 196792 84662 196868 84870
rect 196792 84598 196798 84662
rect 196862 84598 196868 84662
rect 196792 84592 196868 84598
rect 195432 84462 195438 84526
rect 195502 84462 195508 84526
rect 195432 84456 195508 84462
rect 195845 84390 195911 84391
rect 195845 84358 195846 84390
rect 195840 84326 195846 84358
rect 195910 84358 195911 84390
rect 196112 84390 196188 84396
rect 195910 84326 195916 84358
rect 28424 84222 28430 84254
rect 28429 84190 28430 84222
rect 28494 84222 28500 84254
rect 28565 84254 28631 84255
rect 28565 84222 28566 84254
rect 28494 84190 28495 84222
rect 28429 84189 28495 84190
rect 28560 84190 28566 84222
rect 28630 84222 28631 84254
rect 190264 84254 190340 84260
rect 28630 84190 28636 84222
rect 22440 84086 22446 84118
rect 22374 84054 22375 84086
rect 22309 84053 22375 84054
rect 22445 84054 22446 84086
rect 22510 84086 22516 84118
rect 22510 84054 22511 84086
rect 22445 84053 22511 84054
rect 28560 83982 28636 84190
rect 28560 83918 28566 83982
rect 28630 83918 28636 83982
rect 190264 84190 190270 84254
rect 190334 84190 190340 84254
rect 190264 83982 190340 84190
rect 195840 84118 195916 84326
rect 195840 84054 195846 84118
rect 195910 84054 195916 84118
rect 196112 84326 196118 84390
rect 196182 84326 196188 84390
rect 196112 84118 196188 84326
rect 217464 84390 217812 86094
rect 217464 84326 217470 84390
rect 217534 84326 217812 84390
rect 196112 84086 196118 84118
rect 195840 84048 195916 84054
rect 196117 84054 196118 84086
rect 196182 84086 196188 84118
rect 196797 84118 196863 84119
rect 196797 84086 196798 84118
rect 196182 84054 196183 84086
rect 196117 84053 196183 84054
rect 196792 84054 196798 84086
rect 196862 84086 196863 84118
rect 196862 84054 196868 84086
rect 190264 83950 190270 83982
rect 28560 83912 28636 83918
rect 190269 83918 190270 83950
rect 190334 83950 190340 83982
rect 190334 83918 190335 83950
rect 190269 83917 190335 83918
rect 21896 83814 21902 83846
rect 21901 83782 21902 83814
rect 21966 83814 21972 83846
rect 28565 83846 28631 83847
rect 28565 83814 28566 83846
rect 21966 83782 21967 83814
rect 21901 83781 21967 83782
rect 28560 83782 28566 83814
rect 28630 83814 28631 83846
rect 196792 83846 196868 84054
rect 28630 83782 28636 83814
rect 21760 83710 21836 83716
rect 21760 83646 21766 83710
rect 21830 83646 21836 83710
rect 22309 83710 22375 83711
rect 22309 83678 22310 83710
rect 21760 83438 21836 83646
rect 21760 83406 21766 83438
rect 21765 83374 21766 83406
rect 21830 83406 21836 83438
rect 22304 83646 22310 83678
rect 22374 83678 22375 83710
rect 22581 83710 22647 83711
rect 22581 83678 22582 83710
rect 22374 83646 22380 83678
rect 22304 83438 22380 83646
rect 21830 83374 21831 83406
rect 21765 83373 21831 83374
rect 22304 83374 22310 83438
rect 22374 83374 22380 83438
rect 22304 83368 22380 83374
rect 22576 83646 22582 83678
rect 22646 83678 22647 83710
rect 23120 83710 23196 83716
rect 22646 83646 22652 83678
rect 22576 83438 22652 83646
rect 22576 83374 22582 83438
rect 22646 83374 22652 83438
rect 23120 83646 23126 83710
rect 23190 83646 23196 83710
rect 23120 83438 23196 83646
rect 23120 83406 23126 83438
rect 22576 83368 22652 83374
rect 23125 83374 23126 83406
rect 23190 83406 23196 83438
rect 23528 83710 23604 83716
rect 23528 83646 23534 83710
rect 23598 83646 23604 83710
rect 23528 83438 23604 83646
rect 23528 83406 23534 83438
rect 23190 83374 23191 83406
rect 23125 83373 23191 83374
rect 23533 83374 23534 83406
rect 23598 83406 23604 83438
rect 28429 83438 28495 83439
rect 28429 83406 28430 83438
rect 23598 83374 23599 83406
rect 23533 83373 23599 83374
rect 28424 83374 28430 83406
rect 28494 83406 28495 83438
rect 28560 83438 28636 83782
rect 196792 83782 196798 83846
rect 196862 83782 196868 83846
rect 196792 83776 196868 83782
rect 28494 83374 28500 83406
rect 21765 83302 21831 83303
rect 21765 83270 21766 83302
rect 21760 83238 21766 83270
rect 21830 83270 21831 83302
rect 23125 83302 23191 83303
rect 23125 83270 23126 83302
rect 21830 83238 21836 83270
rect 21760 83030 21836 83238
rect 21760 82966 21766 83030
rect 21830 82966 21836 83030
rect 21760 82960 21836 82966
rect 23120 83238 23126 83270
rect 23190 83270 23191 83302
rect 23533 83302 23599 83303
rect 23533 83270 23534 83302
rect 23190 83238 23196 83270
rect 23120 83030 23196 83238
rect 23120 82966 23126 83030
rect 23190 82966 23196 83030
rect 23120 82960 23196 82966
rect 23528 83238 23534 83270
rect 23598 83270 23599 83302
rect 23598 83238 23604 83270
rect 23528 83030 23604 83238
rect 28424 83166 28500 83374
rect 28560 83374 28566 83438
rect 28630 83374 28636 83438
rect 195160 83710 195236 83716
rect 195160 83646 195166 83710
rect 195230 83646 195236 83710
rect 195437 83710 195503 83711
rect 195437 83678 195438 83710
rect 195160 83438 195236 83646
rect 195160 83406 195166 83438
rect 28560 83368 28636 83374
rect 195165 83374 195166 83406
rect 195230 83406 195236 83438
rect 195432 83646 195438 83678
rect 195502 83678 195503 83710
rect 195845 83710 195911 83711
rect 195845 83678 195846 83710
rect 195502 83646 195508 83678
rect 195432 83438 195508 83646
rect 195230 83374 195231 83406
rect 195165 83373 195231 83374
rect 195432 83374 195438 83438
rect 195502 83374 195508 83438
rect 195432 83368 195508 83374
rect 195840 83646 195846 83678
rect 195910 83678 195911 83710
rect 196656 83710 196732 83716
rect 195910 83646 195916 83678
rect 195840 83438 195916 83646
rect 195840 83374 195846 83438
rect 195910 83374 195916 83438
rect 196656 83646 196662 83710
rect 196726 83646 196732 83710
rect 196656 83438 196732 83646
rect 196656 83406 196662 83438
rect 195840 83368 195916 83374
rect 196661 83374 196662 83406
rect 196726 83406 196732 83438
rect 196726 83374 196727 83406
rect 196661 83373 196727 83374
rect 195165 83302 195231 83303
rect 195165 83270 195166 83302
rect 28424 83102 28430 83166
rect 28494 83102 28500 83166
rect 28424 83096 28500 83102
rect 195160 83238 195166 83270
rect 195230 83270 195231 83302
rect 195573 83302 195639 83303
rect 195573 83270 195574 83302
rect 195230 83238 195236 83270
rect 23528 82966 23534 83030
rect 23598 82966 23604 83030
rect 23528 82960 23604 82966
rect 195160 83030 195236 83238
rect 195160 82966 195166 83030
rect 195230 82966 195236 83030
rect 195160 82960 195236 82966
rect 195568 83238 195574 83270
rect 195638 83270 195639 83302
rect 195976 83302 196052 83308
rect 195638 83238 195644 83270
rect 195568 83030 195644 83238
rect 195568 82966 195574 83030
rect 195638 82966 195644 83030
rect 195976 83238 195982 83302
rect 196046 83238 196052 83302
rect 195976 83030 196052 83238
rect 195976 82998 195982 83030
rect 195568 82960 195644 82966
rect 195981 82966 195982 82998
rect 196046 82998 196052 83030
rect 196384 83302 196460 83308
rect 196384 83238 196390 83302
rect 196454 83238 196460 83302
rect 196661 83302 196727 83303
rect 196661 83270 196662 83302
rect 196384 83030 196460 83238
rect 196384 82998 196390 83030
rect 196046 82966 196047 82998
rect 195981 82965 196047 82966
rect 196389 82966 196390 82998
rect 196454 82998 196460 83030
rect 196656 83238 196662 83270
rect 196726 83270 196727 83302
rect 196726 83238 196732 83270
rect 196656 83030 196732 83238
rect 196454 82966 196455 82998
rect 196389 82965 196455 82966
rect 196656 82966 196662 83030
rect 196726 82966 196732 83030
rect 196656 82960 196732 82966
rect 952 82694 1230 82758
rect 1294 82694 1300 82758
rect 952 81126 1300 82694
rect 21760 82894 21836 82900
rect 21760 82830 21766 82894
rect 21830 82830 21836 82894
rect 22717 82894 22783 82895
rect 22717 82862 22718 82894
rect 21760 82622 21836 82830
rect 21760 82590 21766 82622
rect 21765 82558 21766 82590
rect 21830 82590 21836 82622
rect 22712 82830 22718 82862
rect 22782 82862 22783 82894
rect 23125 82894 23191 82895
rect 23125 82862 23126 82894
rect 22782 82830 22788 82862
rect 22712 82622 22788 82830
rect 21830 82558 21831 82590
rect 21765 82557 21831 82558
rect 22712 82558 22718 82622
rect 22782 82558 22788 82622
rect 22712 82552 22788 82558
rect 23120 82830 23126 82862
rect 23190 82862 23191 82894
rect 23528 82894 23604 82900
rect 23190 82830 23196 82862
rect 23120 82622 23196 82830
rect 23120 82558 23126 82622
rect 23190 82558 23196 82622
rect 23528 82830 23534 82894
rect 23598 82830 23604 82894
rect 23528 82622 23604 82830
rect 23528 82590 23534 82622
rect 23120 82552 23196 82558
rect 23533 82558 23534 82590
rect 23598 82590 23604 82622
rect 195160 82894 195236 82900
rect 195160 82830 195166 82894
rect 195230 82830 195236 82894
rect 195160 82622 195236 82830
rect 195160 82590 195166 82622
rect 23598 82558 23599 82590
rect 23533 82557 23599 82558
rect 195165 82558 195166 82590
rect 195230 82590 195236 82622
rect 195432 82894 195508 82900
rect 195432 82830 195438 82894
rect 195502 82830 195508 82894
rect 195432 82622 195508 82830
rect 195432 82590 195438 82622
rect 195230 82558 195231 82590
rect 195165 82557 195231 82558
rect 195437 82558 195438 82590
rect 195502 82590 195508 82622
rect 196248 82894 196324 82900
rect 196248 82830 196254 82894
rect 196318 82830 196324 82894
rect 196797 82894 196863 82895
rect 196797 82862 196798 82894
rect 196248 82622 196324 82830
rect 196248 82590 196254 82622
rect 195502 82558 195503 82590
rect 195437 82557 195503 82558
rect 196253 82558 196254 82590
rect 196318 82590 196324 82622
rect 196792 82830 196798 82862
rect 196862 82862 196863 82894
rect 217464 82894 217812 84326
rect 196862 82830 196868 82862
rect 196792 82622 196868 82830
rect 196318 82558 196319 82590
rect 196253 82557 196319 82558
rect 196792 82558 196798 82622
rect 196862 82558 196868 82622
rect 196792 82552 196868 82558
rect 217464 82830 217470 82894
rect 217534 82830 217812 82894
rect 21765 82486 21831 82487
rect 21765 82454 21766 82486
rect 21760 82422 21766 82454
rect 21830 82454 21831 82486
rect 22168 82486 22244 82492
rect 21830 82422 21836 82454
rect 21760 82214 21836 82422
rect 21760 82150 21766 82214
rect 21830 82150 21836 82214
rect 22168 82422 22174 82486
rect 22238 82422 22244 82486
rect 22168 82214 22244 82422
rect 22168 82182 22174 82214
rect 21760 82144 21836 82150
rect 22173 82150 22174 82182
rect 22238 82182 22244 82214
rect 22576 82486 22652 82492
rect 22576 82422 22582 82486
rect 22646 82422 22652 82486
rect 22576 82214 22652 82422
rect 22576 82182 22582 82214
rect 22238 82150 22239 82182
rect 22173 82149 22239 82150
rect 22581 82150 22582 82182
rect 22646 82182 22652 82214
rect 23120 82486 23196 82492
rect 23120 82422 23126 82486
rect 23190 82422 23196 82486
rect 23533 82486 23599 82487
rect 23533 82454 23534 82486
rect 23120 82214 23196 82422
rect 23120 82182 23126 82214
rect 22646 82150 22647 82182
rect 22581 82149 22647 82150
rect 23125 82150 23126 82182
rect 23190 82182 23196 82214
rect 23528 82422 23534 82454
rect 23598 82454 23599 82486
rect 195160 82486 195236 82492
rect 23598 82422 23604 82454
rect 23528 82214 23604 82422
rect 23190 82150 23191 82182
rect 23125 82149 23191 82150
rect 23528 82150 23534 82214
rect 23598 82150 23604 82214
rect 195160 82422 195166 82486
rect 195230 82422 195236 82486
rect 195437 82486 195503 82487
rect 195437 82454 195438 82486
rect 195160 82214 195236 82422
rect 195160 82182 195166 82214
rect 23528 82144 23604 82150
rect 195165 82150 195166 82182
rect 195230 82182 195236 82214
rect 195432 82422 195438 82454
rect 195502 82454 195503 82486
rect 195840 82486 195916 82492
rect 195502 82422 195508 82454
rect 195432 82214 195508 82422
rect 195230 82150 195231 82182
rect 195165 82149 195231 82150
rect 195432 82150 195438 82214
rect 195502 82150 195508 82214
rect 195840 82422 195846 82486
rect 195910 82422 195916 82486
rect 196253 82486 196319 82487
rect 196253 82454 196254 82486
rect 195840 82214 195916 82422
rect 195840 82182 195846 82214
rect 195432 82144 195508 82150
rect 195845 82150 195846 82182
rect 195910 82182 195916 82214
rect 196248 82422 196254 82454
rect 196318 82454 196319 82486
rect 196661 82486 196727 82487
rect 196661 82454 196662 82486
rect 196318 82422 196324 82454
rect 196248 82214 196324 82422
rect 195910 82150 195911 82182
rect 195845 82149 195911 82150
rect 196248 82150 196254 82214
rect 196318 82150 196324 82214
rect 196248 82144 196324 82150
rect 196656 82422 196662 82454
rect 196726 82454 196727 82486
rect 196726 82422 196732 82454
rect 196656 82214 196732 82422
rect 196656 82150 196662 82214
rect 196726 82150 196732 82214
rect 196656 82144 196732 82150
rect 21896 82078 21972 82084
rect 21896 82014 21902 82078
rect 21966 82014 21972 82078
rect 22717 82078 22783 82079
rect 22717 82046 22718 82078
rect 21896 81806 21972 82014
rect 21896 81774 21902 81806
rect 21901 81742 21902 81774
rect 21966 81774 21972 81806
rect 22712 82014 22718 82046
rect 22782 82046 22783 82078
rect 23120 82078 23196 82084
rect 22782 82014 22788 82046
rect 22712 81806 22788 82014
rect 21966 81742 21967 81774
rect 21901 81741 21967 81742
rect 22712 81742 22718 81806
rect 22782 81742 22788 81806
rect 23120 82014 23126 82078
rect 23190 82014 23196 82078
rect 23397 82078 23463 82079
rect 23397 82046 23398 82078
rect 23120 81806 23196 82014
rect 23120 81774 23126 81806
rect 22712 81736 22788 81742
rect 23125 81742 23126 81774
rect 23190 81774 23196 81806
rect 23392 82014 23398 82046
rect 23462 82046 23463 82078
rect 195029 82078 195095 82079
rect 195029 82046 195030 82078
rect 23462 82014 23468 82046
rect 23392 81806 23468 82014
rect 23190 81742 23191 81774
rect 23125 81741 23191 81742
rect 23392 81742 23398 81806
rect 23462 81742 23468 81806
rect 23392 81736 23468 81742
rect 195024 82014 195030 82046
rect 195094 82046 195095 82078
rect 195437 82078 195503 82079
rect 195437 82046 195438 82078
rect 195094 82014 195100 82046
rect 195024 81806 195100 82014
rect 195024 81742 195030 81806
rect 195094 81742 195100 81806
rect 195024 81736 195100 81742
rect 195432 82014 195438 82046
rect 195502 82046 195503 82078
rect 195981 82078 196047 82079
rect 195981 82046 195982 82078
rect 195502 82014 195508 82046
rect 195432 81806 195508 82014
rect 195432 81742 195438 81806
rect 195502 81742 195508 81806
rect 195432 81736 195508 81742
rect 195976 82014 195982 82046
rect 196046 82046 196047 82078
rect 196792 82078 196868 82084
rect 196046 82014 196052 82046
rect 195976 81806 196052 82014
rect 195976 81742 195982 81806
rect 196046 81742 196052 81806
rect 196792 82014 196798 82078
rect 196862 82014 196868 82078
rect 196792 81806 196868 82014
rect 196792 81774 196798 81806
rect 195976 81736 196052 81742
rect 196797 81742 196798 81774
rect 196862 81774 196868 81806
rect 196862 81742 196863 81774
rect 196797 81741 196863 81742
rect 21760 81670 21836 81676
rect 21760 81606 21766 81670
rect 21830 81606 21836 81670
rect 22309 81670 22375 81671
rect 22309 81638 22310 81670
rect 21760 81398 21836 81606
rect 21760 81366 21766 81398
rect 21765 81334 21766 81366
rect 21830 81366 21836 81398
rect 22304 81606 22310 81638
rect 22374 81638 22375 81670
rect 22445 81670 22511 81671
rect 22445 81638 22446 81670
rect 22374 81606 22380 81638
rect 22304 81398 22380 81606
rect 21830 81334 21831 81366
rect 21765 81333 21831 81334
rect 22304 81334 22310 81398
rect 22374 81334 22380 81398
rect 22304 81328 22380 81334
rect 22440 81606 22446 81638
rect 22510 81638 22511 81670
rect 23125 81670 23191 81671
rect 23125 81638 23126 81670
rect 22510 81606 22516 81638
rect 22440 81398 22516 81606
rect 22440 81334 22446 81398
rect 22510 81334 22516 81398
rect 22440 81328 22516 81334
rect 23120 81606 23126 81638
rect 23190 81638 23191 81670
rect 23528 81670 23604 81676
rect 23190 81606 23196 81638
rect 23120 81398 23196 81606
rect 23120 81334 23126 81398
rect 23190 81334 23196 81398
rect 23528 81606 23534 81670
rect 23598 81606 23604 81670
rect 23528 81398 23604 81606
rect 23528 81366 23534 81398
rect 23120 81328 23196 81334
rect 23533 81334 23534 81366
rect 23598 81366 23604 81398
rect 195160 81670 195236 81676
rect 195160 81606 195166 81670
rect 195230 81606 195236 81670
rect 195160 81398 195236 81606
rect 195160 81366 195166 81398
rect 23598 81334 23599 81366
rect 23533 81333 23599 81334
rect 195165 81334 195166 81366
rect 195230 81366 195236 81398
rect 195432 81670 195508 81676
rect 195432 81606 195438 81670
rect 195502 81606 195508 81670
rect 196117 81670 196183 81671
rect 196117 81638 196118 81670
rect 195432 81398 195508 81606
rect 195432 81366 195438 81398
rect 195230 81334 195231 81366
rect 195165 81333 195231 81334
rect 195437 81334 195438 81366
rect 195502 81366 195508 81398
rect 196112 81606 196118 81638
rect 196182 81638 196183 81670
rect 196656 81670 196732 81676
rect 196182 81606 196188 81638
rect 196112 81398 196188 81606
rect 195502 81334 195503 81366
rect 195437 81333 195503 81334
rect 196112 81334 196118 81398
rect 196182 81334 196188 81398
rect 196656 81606 196662 81670
rect 196726 81606 196732 81670
rect 196656 81398 196732 81606
rect 196656 81366 196662 81398
rect 196112 81328 196188 81334
rect 196661 81334 196662 81366
rect 196726 81366 196732 81398
rect 196726 81334 196727 81366
rect 196661 81333 196727 81334
rect 22581 81262 22647 81263
rect 22581 81230 22582 81262
rect 952 81062 1230 81126
rect 1294 81062 1300 81126
rect 952 79630 1300 81062
rect 22576 81198 22582 81230
rect 22646 81230 22647 81262
rect 22984 81262 23060 81268
rect 22646 81198 22652 81230
rect 21901 80990 21967 80991
rect 21901 80958 21902 80990
rect 21896 80926 21902 80958
rect 21966 80958 21967 80990
rect 22445 80990 22511 80991
rect 22445 80958 22446 80990
rect 21966 80926 21972 80958
rect 21896 80718 21972 80926
rect 21896 80654 21902 80718
rect 21966 80654 21972 80718
rect 21896 80648 21972 80654
rect 22440 80926 22446 80958
rect 22510 80958 22511 80990
rect 22576 80990 22652 81198
rect 22510 80926 22516 80958
rect 22440 80718 22516 80926
rect 22576 80926 22582 80990
rect 22646 80926 22652 80990
rect 22984 81198 22990 81262
rect 23054 81198 23060 81262
rect 23533 81262 23599 81263
rect 23533 81230 23534 81262
rect 22984 80990 23060 81198
rect 22984 80958 22990 80990
rect 22576 80920 22652 80926
rect 22989 80926 22990 80958
rect 23054 80958 23060 80990
rect 23528 81198 23534 81230
rect 23598 81230 23599 81262
rect 195165 81262 195231 81263
rect 195165 81230 195166 81262
rect 23598 81198 23604 81230
rect 23528 80990 23604 81198
rect 195160 81198 195166 81230
rect 195230 81230 195231 81262
rect 195437 81262 195503 81263
rect 195437 81230 195438 81262
rect 195230 81198 195236 81230
rect 23054 80926 23055 80958
rect 22989 80925 23055 80926
rect 23528 80926 23534 80990
rect 23598 80926 23604 80990
rect 23528 80920 23604 80926
rect 28560 81126 28636 81132
rect 28560 81062 28566 81126
rect 28630 81062 28636 81126
rect 22989 80854 23055 80855
rect 22989 80822 22990 80854
rect 22440 80654 22446 80718
rect 22510 80654 22516 80718
rect 22440 80648 22516 80654
rect 22984 80790 22990 80822
rect 23054 80822 23055 80854
rect 23397 80854 23463 80855
rect 23397 80822 23398 80854
rect 23054 80790 23060 80822
rect 22984 80582 23060 80790
rect 22984 80518 22990 80582
rect 23054 80518 23060 80582
rect 22984 80512 23060 80518
rect 23392 80790 23398 80822
rect 23462 80822 23463 80854
rect 28429 80854 28495 80855
rect 28429 80822 28430 80854
rect 23462 80790 23468 80822
rect 23392 80582 23468 80790
rect 23392 80518 23398 80582
rect 23462 80518 23468 80582
rect 23392 80512 23468 80518
rect 28424 80790 28430 80822
rect 28494 80822 28495 80854
rect 28560 80854 28636 81062
rect 195160 80990 195236 81198
rect 195160 80926 195166 80990
rect 195230 80926 195236 80990
rect 195160 80920 195236 80926
rect 195432 81198 195438 81230
rect 195502 81230 195503 81262
rect 195976 81262 196052 81268
rect 195502 81198 195508 81230
rect 195432 80990 195508 81198
rect 195432 80926 195438 80990
rect 195502 80926 195508 80990
rect 195976 81198 195982 81262
rect 196046 81198 196052 81262
rect 195976 80990 196052 81198
rect 195976 80958 195982 80990
rect 195432 80920 195508 80926
rect 195981 80926 195982 80958
rect 196046 80958 196052 80990
rect 196112 81262 196188 81268
rect 196112 81198 196118 81262
rect 196182 81198 196188 81262
rect 196112 80990 196188 81198
rect 217464 81262 217812 82830
rect 217464 81198 217470 81262
rect 217534 81198 217812 81262
rect 196112 80958 196118 80990
rect 196046 80926 196047 80958
rect 195981 80925 196047 80926
rect 196117 80926 196118 80958
rect 196182 80958 196188 80990
rect 196656 80990 196732 80996
rect 196182 80926 196183 80958
rect 196117 80925 196183 80926
rect 196656 80926 196662 80990
rect 196726 80926 196732 80990
rect 28560 80822 28566 80854
rect 28494 80790 28500 80822
rect 22440 80446 22516 80452
rect 22440 80382 22446 80446
rect 22510 80382 22516 80446
rect 21765 80174 21831 80175
rect 21765 80142 21766 80174
rect 21760 80110 21766 80142
rect 21830 80142 21831 80174
rect 22440 80174 22516 80382
rect 28424 80446 28500 80790
rect 28565 80790 28566 80822
rect 28630 80822 28636 80854
rect 195029 80854 195095 80855
rect 195029 80822 195030 80854
rect 28630 80790 28631 80822
rect 28565 80789 28631 80790
rect 195024 80790 195030 80822
rect 195094 80822 195095 80854
rect 195568 80854 195644 80860
rect 195094 80790 195100 80822
rect 195024 80582 195100 80790
rect 195024 80518 195030 80582
rect 195094 80518 195100 80582
rect 195568 80790 195574 80854
rect 195638 80790 195644 80854
rect 195568 80582 195644 80790
rect 196656 80718 196732 80926
rect 196656 80686 196662 80718
rect 196661 80654 196662 80686
rect 196726 80686 196732 80718
rect 196726 80654 196727 80686
rect 196661 80653 196727 80654
rect 195568 80550 195574 80582
rect 195024 80512 195100 80518
rect 195573 80518 195574 80550
rect 195638 80550 195644 80582
rect 195638 80518 195639 80550
rect 195573 80517 195639 80518
rect 28424 80382 28430 80446
rect 28494 80382 28500 80446
rect 195981 80446 196047 80447
rect 195981 80414 195982 80446
rect 28424 80376 28500 80382
rect 195976 80382 195982 80414
rect 196046 80414 196047 80446
rect 196046 80382 196052 80414
rect 28293 80310 28359 80311
rect 28293 80278 28294 80310
rect 22440 80142 22446 80174
rect 21830 80110 21836 80142
rect 21760 79902 21836 80110
rect 22445 80110 22446 80142
rect 22510 80142 22516 80174
rect 28288 80246 28294 80278
rect 28358 80278 28359 80310
rect 190128 80310 190204 80316
rect 28358 80246 28364 80278
rect 22510 80110 22511 80142
rect 22445 80109 22511 80110
rect 28288 80038 28364 80246
rect 190128 80246 190134 80310
rect 190198 80246 190204 80310
rect 28288 79974 28294 80038
rect 28358 79974 28364 80038
rect 28429 80038 28495 80039
rect 28429 80006 28430 80038
rect 28288 79968 28364 79974
rect 28424 79974 28430 80006
rect 28494 80006 28495 80038
rect 190128 80038 190204 80246
rect 195976 80174 196052 80382
rect 195976 80110 195982 80174
rect 196046 80110 196052 80174
rect 195976 80104 196052 80110
rect 196792 80174 196868 80180
rect 196792 80110 196798 80174
rect 196862 80110 196868 80174
rect 190128 80006 190134 80038
rect 28494 79974 28500 80006
rect 21760 79838 21766 79902
rect 21830 79838 21836 79902
rect 21760 79832 21836 79838
rect 952 79566 1230 79630
rect 1294 79566 1300 79630
rect 952 77726 1300 79566
rect 21896 79766 21972 79772
rect 21896 79702 21902 79766
rect 21966 79702 21972 79766
rect 22309 79766 22375 79767
rect 22309 79734 22310 79766
rect 21896 79494 21972 79702
rect 21896 79462 21902 79494
rect 21901 79430 21902 79462
rect 21966 79462 21972 79494
rect 22304 79702 22310 79734
rect 22374 79734 22375 79766
rect 22445 79766 22511 79767
rect 22445 79734 22446 79766
rect 22374 79702 22380 79734
rect 22304 79494 22380 79702
rect 21966 79430 21967 79462
rect 21901 79429 21967 79430
rect 22304 79430 22310 79494
rect 22374 79430 22380 79494
rect 22304 79424 22380 79430
rect 22440 79702 22446 79734
rect 22510 79734 22511 79766
rect 22510 79702 22516 79734
rect 22440 79494 22516 79702
rect 28424 79630 28500 79974
rect 190133 79974 190134 80006
rect 190198 80006 190204 80038
rect 190198 79974 190199 80006
rect 190133 79973 190199 79974
rect 190269 79902 190335 79903
rect 190269 79870 190270 79902
rect 28424 79566 28430 79630
rect 28494 79566 28500 79630
rect 28424 79560 28500 79566
rect 190264 79838 190270 79870
rect 190334 79870 190335 79902
rect 196792 79902 196868 80110
rect 196792 79870 196798 79902
rect 190334 79838 190340 79870
rect 190264 79630 190340 79838
rect 196797 79838 196798 79870
rect 196862 79870 196868 79902
rect 196862 79838 196863 79870
rect 196797 79837 196863 79838
rect 196389 79766 196455 79767
rect 196389 79734 196390 79766
rect 190264 79566 190270 79630
rect 190334 79566 190340 79630
rect 190264 79560 190340 79566
rect 196384 79702 196390 79734
rect 196454 79734 196455 79766
rect 196797 79766 196863 79767
rect 196797 79734 196798 79766
rect 196454 79702 196460 79734
rect 22440 79430 22446 79494
rect 22510 79430 22516 79494
rect 22440 79424 22516 79430
rect 28560 79494 28636 79500
rect 28560 79430 28566 79494
rect 28630 79430 28636 79494
rect 190269 79494 190335 79495
rect 190269 79462 190270 79494
rect 21765 79358 21831 79359
rect 21765 79326 21766 79358
rect 21760 79294 21766 79326
rect 21830 79326 21831 79358
rect 23120 79358 23196 79364
rect 21830 79294 21836 79326
rect 21760 79086 21836 79294
rect 21760 79022 21766 79086
rect 21830 79022 21836 79086
rect 23120 79294 23126 79358
rect 23190 79294 23196 79358
rect 23533 79358 23599 79359
rect 23533 79326 23534 79358
rect 23120 79086 23196 79294
rect 23120 79054 23126 79086
rect 21760 79016 21836 79022
rect 23125 79022 23126 79054
rect 23190 79054 23196 79086
rect 23528 79294 23534 79326
rect 23598 79326 23599 79358
rect 23598 79294 23604 79326
rect 23528 79086 23604 79294
rect 28560 79222 28636 79430
rect 28560 79190 28566 79222
rect 28565 79158 28566 79190
rect 28630 79190 28636 79222
rect 190264 79430 190270 79462
rect 190334 79462 190335 79494
rect 196384 79494 196460 79702
rect 190334 79430 190340 79462
rect 190264 79222 190340 79430
rect 196384 79430 196390 79494
rect 196454 79430 196460 79494
rect 196384 79424 196460 79430
rect 196792 79702 196798 79734
rect 196862 79734 196863 79766
rect 196862 79702 196868 79734
rect 196792 79494 196868 79702
rect 196792 79430 196798 79494
rect 196862 79430 196868 79494
rect 196792 79424 196868 79430
rect 28630 79158 28631 79190
rect 28565 79157 28631 79158
rect 190264 79158 190270 79222
rect 190334 79158 190340 79222
rect 190264 79152 190340 79158
rect 195160 79358 195236 79364
rect 195160 79294 195166 79358
rect 195230 79294 195236 79358
rect 23190 79022 23191 79054
rect 23125 79021 23191 79022
rect 23528 79022 23534 79086
rect 23598 79022 23604 79086
rect 195160 79086 195236 79294
rect 195160 79054 195166 79086
rect 23528 79016 23604 79022
rect 195165 79022 195166 79054
rect 195230 79054 195236 79086
rect 195568 79358 195644 79364
rect 195568 79294 195574 79358
rect 195638 79294 195644 79358
rect 196661 79358 196727 79359
rect 196661 79326 196662 79358
rect 195568 79086 195644 79294
rect 195568 79054 195574 79086
rect 195230 79022 195231 79054
rect 195165 79021 195231 79022
rect 195573 79022 195574 79054
rect 195638 79054 195644 79086
rect 196656 79294 196662 79326
rect 196726 79326 196727 79358
rect 217464 79358 217812 81198
rect 196726 79294 196732 79326
rect 196656 79086 196732 79294
rect 195638 79022 195639 79054
rect 195573 79021 195639 79022
rect 196656 79022 196662 79086
rect 196726 79022 196732 79086
rect 196656 79016 196732 79022
rect 217464 79294 217470 79358
rect 217534 79294 217812 79358
rect 21896 78950 21972 78956
rect 21896 78886 21902 78950
rect 21966 78886 21972 78950
rect 22581 78950 22647 78951
rect 22581 78918 22582 78950
rect 21896 78678 21972 78886
rect 21896 78646 21902 78678
rect 21901 78614 21902 78646
rect 21966 78646 21972 78678
rect 22576 78886 22582 78918
rect 22646 78918 22647 78950
rect 22984 78950 23060 78956
rect 22646 78886 22652 78918
rect 22576 78678 22652 78886
rect 21966 78614 21967 78646
rect 21901 78613 21967 78614
rect 22576 78614 22582 78678
rect 22646 78614 22652 78678
rect 22984 78886 22990 78950
rect 23054 78886 23060 78950
rect 22984 78678 23060 78886
rect 22984 78646 22990 78678
rect 22576 78608 22652 78614
rect 22989 78614 22990 78646
rect 23054 78646 23060 78678
rect 23392 78950 23468 78956
rect 23392 78886 23398 78950
rect 23462 78886 23468 78950
rect 195165 78950 195231 78951
rect 195165 78918 195166 78950
rect 23392 78678 23468 78886
rect 23392 78646 23398 78678
rect 23054 78614 23055 78646
rect 22989 78613 23055 78614
rect 23397 78614 23398 78646
rect 23462 78646 23468 78678
rect 195160 78886 195166 78918
rect 195230 78918 195231 78950
rect 195432 78950 195508 78956
rect 195230 78886 195236 78918
rect 195160 78678 195236 78886
rect 23462 78614 23463 78646
rect 23397 78613 23463 78614
rect 195160 78614 195166 78678
rect 195230 78614 195236 78678
rect 195432 78886 195438 78950
rect 195502 78886 195508 78950
rect 195845 78950 195911 78951
rect 195845 78918 195846 78950
rect 195432 78678 195508 78886
rect 195432 78646 195438 78678
rect 195160 78608 195236 78614
rect 195437 78614 195438 78646
rect 195502 78646 195508 78678
rect 195840 78886 195846 78918
rect 195910 78918 195911 78950
rect 196112 78950 196188 78956
rect 195910 78886 195916 78918
rect 195840 78678 195916 78886
rect 195502 78614 195503 78646
rect 195437 78613 195503 78614
rect 195840 78614 195846 78678
rect 195910 78614 195916 78678
rect 196112 78886 196118 78950
rect 196182 78886 196188 78950
rect 196112 78678 196188 78886
rect 196112 78646 196118 78678
rect 195840 78608 195916 78614
rect 196117 78614 196118 78646
rect 196182 78646 196188 78678
rect 196792 78950 196868 78956
rect 196792 78886 196798 78950
rect 196862 78886 196868 78950
rect 196792 78678 196868 78886
rect 196792 78646 196798 78678
rect 196182 78614 196183 78646
rect 196117 78613 196183 78614
rect 196797 78614 196798 78646
rect 196862 78646 196868 78678
rect 196862 78614 196863 78646
rect 196797 78613 196863 78614
rect 21901 78542 21967 78543
rect 21901 78510 21902 78542
rect 21896 78478 21902 78510
rect 21966 78510 21967 78542
rect 22168 78542 22244 78548
rect 21966 78478 21972 78510
rect 21896 78270 21972 78478
rect 21896 78206 21902 78270
rect 21966 78206 21972 78270
rect 22168 78478 22174 78542
rect 22238 78478 22244 78542
rect 22717 78542 22783 78543
rect 22717 78510 22718 78542
rect 22168 78270 22244 78478
rect 22168 78238 22174 78270
rect 21896 78200 21972 78206
rect 22173 78206 22174 78238
rect 22238 78238 22244 78270
rect 22712 78478 22718 78510
rect 22782 78510 22783 78542
rect 22989 78542 23055 78543
rect 22989 78510 22990 78542
rect 22782 78478 22788 78510
rect 22712 78270 22788 78478
rect 22238 78206 22239 78238
rect 22173 78205 22239 78206
rect 22712 78206 22718 78270
rect 22782 78206 22788 78270
rect 22712 78200 22788 78206
rect 22984 78478 22990 78510
rect 23054 78510 23055 78542
rect 23397 78542 23463 78543
rect 23397 78510 23398 78542
rect 23054 78478 23060 78510
rect 22984 78270 23060 78478
rect 22984 78206 22990 78270
rect 23054 78206 23060 78270
rect 22984 78200 23060 78206
rect 23392 78478 23398 78510
rect 23462 78510 23463 78542
rect 195160 78542 195236 78548
rect 23462 78478 23468 78510
rect 23392 78270 23468 78478
rect 23392 78206 23398 78270
rect 23462 78206 23468 78270
rect 195160 78478 195166 78542
rect 195230 78478 195236 78542
rect 195573 78542 195639 78543
rect 195573 78510 195574 78542
rect 195160 78270 195236 78478
rect 195160 78238 195166 78270
rect 23392 78200 23468 78206
rect 195165 78206 195166 78238
rect 195230 78238 195236 78270
rect 195568 78478 195574 78510
rect 195638 78510 195639 78542
rect 195840 78542 195916 78548
rect 195638 78478 195644 78510
rect 195568 78270 195644 78478
rect 195230 78206 195231 78238
rect 195165 78205 195231 78206
rect 195568 78206 195574 78270
rect 195638 78206 195644 78270
rect 195840 78478 195846 78542
rect 195910 78478 195916 78542
rect 196797 78542 196863 78543
rect 196797 78510 196798 78542
rect 195840 78270 195916 78478
rect 195840 78238 195846 78270
rect 195568 78200 195644 78206
rect 195845 78206 195846 78238
rect 195910 78238 195916 78270
rect 196792 78478 196798 78510
rect 196862 78510 196863 78542
rect 196862 78478 196868 78510
rect 196792 78270 196868 78478
rect 195910 78206 195911 78238
rect 195845 78205 195911 78206
rect 196792 78206 196798 78270
rect 196862 78206 196868 78270
rect 196792 78200 196868 78206
rect 21760 78134 21836 78140
rect 21760 78070 21766 78134
rect 21830 78070 21836 78134
rect 21760 77862 21836 78070
rect 21760 77830 21766 77862
rect 21765 77798 21766 77830
rect 21830 77830 21836 77862
rect 22576 78134 22652 78140
rect 22576 78070 22582 78134
rect 22646 78070 22652 78134
rect 22989 78134 23055 78135
rect 22989 78102 22990 78134
rect 22576 77862 22652 78070
rect 22576 77830 22582 77862
rect 21830 77798 21831 77830
rect 21765 77797 21831 77798
rect 22581 77798 22582 77830
rect 22646 77830 22652 77862
rect 22984 78070 22990 78102
rect 23054 78102 23055 78134
rect 23528 78134 23604 78140
rect 23054 78070 23060 78102
rect 22984 77862 23060 78070
rect 22646 77798 22647 77830
rect 22581 77797 22647 77798
rect 22984 77798 22990 77862
rect 23054 77798 23060 77862
rect 23528 78070 23534 78134
rect 23598 78070 23604 78134
rect 195165 78134 195231 78135
rect 195165 78102 195166 78134
rect 23528 77862 23604 78070
rect 23528 77830 23534 77862
rect 22984 77792 23060 77798
rect 23533 77798 23534 77830
rect 23598 77830 23604 77862
rect 195160 78070 195166 78102
rect 195230 78102 195231 78134
rect 195437 78134 195503 78135
rect 195437 78102 195438 78134
rect 195230 78070 195236 78102
rect 195160 77862 195236 78070
rect 23598 77798 23599 77830
rect 23533 77797 23599 77798
rect 195160 77798 195166 77862
rect 195230 77798 195236 77862
rect 195160 77792 195236 77798
rect 195432 78070 195438 78102
rect 195502 78102 195503 78134
rect 195845 78134 195911 78135
rect 195845 78102 195846 78134
rect 195502 78070 195508 78102
rect 195432 77862 195508 78070
rect 195432 77798 195438 77862
rect 195502 77798 195508 77862
rect 195432 77792 195508 77798
rect 195840 78070 195846 78102
rect 195910 78102 195911 78134
rect 196656 78134 196732 78140
rect 195910 78070 195916 78102
rect 195840 77862 195916 78070
rect 195840 77798 195846 77862
rect 195910 77798 195916 77862
rect 196656 78070 196662 78134
rect 196726 78070 196732 78134
rect 196656 77862 196732 78070
rect 196656 77830 196662 77862
rect 195840 77792 195916 77798
rect 196661 77798 196662 77830
rect 196726 77830 196732 77862
rect 217464 77862 217812 79294
rect 196726 77798 196727 77830
rect 196661 77797 196727 77798
rect 217464 77798 217470 77862
rect 217534 77798 217812 77862
rect 952 77662 1230 77726
rect 1294 77662 1300 77726
rect 21901 77726 21967 77727
rect 21901 77694 21902 77726
rect 952 76230 1300 77662
rect 21896 77662 21902 77694
rect 21966 77694 21967 77726
rect 22445 77726 22511 77727
rect 22445 77694 22446 77726
rect 21966 77662 21972 77694
rect 21896 77454 21972 77662
rect 21896 77390 21902 77454
rect 21966 77390 21972 77454
rect 21896 77384 21972 77390
rect 22440 77662 22446 77694
rect 22510 77694 22511 77726
rect 22989 77726 23055 77727
rect 22989 77694 22990 77726
rect 22510 77662 22516 77694
rect 22440 77454 22516 77662
rect 22440 77390 22446 77454
rect 22510 77390 22516 77454
rect 22440 77384 22516 77390
rect 22984 77662 22990 77694
rect 23054 77694 23055 77726
rect 23392 77726 23468 77732
rect 23054 77662 23060 77694
rect 22984 77454 23060 77662
rect 22984 77390 22990 77454
rect 23054 77390 23060 77454
rect 23392 77662 23398 77726
rect 23462 77662 23468 77726
rect 195029 77726 195095 77727
rect 195029 77694 195030 77726
rect 23392 77454 23468 77662
rect 23392 77422 23398 77454
rect 22984 77384 23060 77390
rect 23397 77390 23398 77422
rect 23462 77422 23468 77454
rect 195024 77662 195030 77694
rect 195094 77694 195095 77726
rect 195437 77726 195503 77727
rect 195437 77694 195438 77726
rect 195094 77662 195100 77694
rect 195024 77454 195100 77662
rect 23462 77390 23463 77422
rect 23397 77389 23463 77390
rect 195024 77390 195030 77454
rect 195094 77390 195100 77454
rect 195024 77384 195100 77390
rect 195432 77662 195438 77694
rect 195502 77694 195503 77726
rect 195981 77726 196047 77727
rect 195981 77694 195982 77726
rect 195502 77662 195508 77694
rect 195432 77454 195508 77662
rect 195432 77390 195438 77454
rect 195502 77390 195508 77454
rect 195432 77384 195508 77390
rect 195976 77662 195982 77694
rect 196046 77694 196047 77726
rect 196389 77726 196455 77727
rect 196389 77694 196390 77726
rect 196046 77662 196052 77694
rect 195976 77454 196052 77662
rect 195976 77390 195982 77454
rect 196046 77390 196052 77454
rect 195976 77384 196052 77390
rect 196384 77662 196390 77694
rect 196454 77694 196455 77726
rect 196792 77726 196868 77732
rect 196454 77662 196460 77694
rect 196384 77454 196460 77662
rect 196384 77390 196390 77454
rect 196454 77390 196460 77454
rect 196792 77662 196798 77726
rect 196862 77662 196868 77726
rect 196792 77454 196868 77662
rect 196792 77422 196798 77454
rect 196384 77384 196460 77390
rect 196797 77390 196798 77422
rect 196862 77422 196868 77454
rect 196862 77390 196863 77422
rect 196797 77389 196863 77390
rect 22309 77318 22375 77319
rect 22309 77286 22310 77318
rect 22304 77254 22310 77286
rect 22374 77286 22375 77318
rect 22984 77318 23060 77324
rect 22374 77254 22380 77286
rect 22304 77046 22380 77254
rect 22304 76982 22310 77046
rect 22374 76982 22380 77046
rect 22984 77254 22990 77318
rect 23054 77254 23060 77318
rect 22984 77046 23060 77254
rect 22984 77014 22990 77046
rect 22304 76976 22380 76982
rect 22989 76982 22990 77014
rect 23054 77014 23060 77046
rect 23528 77318 23604 77324
rect 23528 77254 23534 77318
rect 23598 77254 23604 77318
rect 23528 77046 23604 77254
rect 195160 77318 195236 77324
rect 195160 77254 195166 77318
rect 195230 77254 195236 77318
rect 190133 77182 190199 77183
rect 190133 77150 190134 77182
rect 23528 77014 23534 77046
rect 23054 76982 23055 77014
rect 22989 76981 23055 76982
rect 23533 76982 23534 77014
rect 23598 77014 23604 77046
rect 190128 77118 190134 77150
rect 190198 77150 190199 77182
rect 190198 77118 190204 77150
rect 23598 76982 23599 77014
rect 23533 76981 23599 76982
rect 22984 76910 23060 76916
rect 22984 76846 22990 76910
rect 23054 76846 23060 76910
rect 23533 76910 23599 76911
rect 23533 76878 23534 76910
rect 22984 76638 23060 76846
rect 22984 76606 22990 76638
rect 22989 76574 22990 76606
rect 23054 76606 23060 76638
rect 23528 76846 23534 76878
rect 23598 76878 23599 76910
rect 190128 76910 190204 77118
rect 195160 77046 195236 77254
rect 195160 77014 195166 77046
rect 195165 76982 195166 77014
rect 195230 77014 195236 77046
rect 195432 77318 195508 77324
rect 195432 77254 195438 77318
rect 195502 77254 195508 77318
rect 195432 77046 195508 77254
rect 195432 77014 195438 77046
rect 195230 76982 195231 77014
rect 195165 76981 195231 76982
rect 195437 76982 195438 77014
rect 195502 77014 195508 77046
rect 195840 77318 195916 77324
rect 195840 77254 195846 77318
rect 195910 77254 195916 77318
rect 196389 77318 196455 77319
rect 196389 77286 196390 77318
rect 195840 77046 195916 77254
rect 195840 77014 195846 77046
rect 195502 76982 195503 77014
rect 195437 76981 195503 76982
rect 195845 76982 195846 77014
rect 195910 77014 195916 77046
rect 196384 77254 196390 77286
rect 196454 77286 196455 77318
rect 196454 77254 196460 77286
rect 196384 77046 196460 77254
rect 195910 76982 195911 77014
rect 195845 76981 195911 76982
rect 196384 76982 196390 77046
rect 196454 76982 196460 77046
rect 196384 76976 196460 76982
rect 23598 76846 23604 76878
rect 23528 76638 23604 76846
rect 190128 76846 190134 76910
rect 190198 76846 190204 76910
rect 195165 76910 195231 76911
rect 195165 76878 195166 76910
rect 190128 76840 190204 76846
rect 195160 76846 195166 76878
rect 195230 76878 195231 76910
rect 195437 76910 195503 76911
rect 195437 76878 195438 76910
rect 195230 76846 195236 76878
rect 23054 76574 23055 76606
rect 22989 76573 23055 76574
rect 23528 76574 23534 76638
rect 23598 76574 23604 76638
rect 23528 76568 23604 76574
rect 195160 76638 195236 76846
rect 195160 76574 195166 76638
rect 195230 76574 195236 76638
rect 195160 76568 195236 76574
rect 195432 76846 195438 76878
rect 195502 76878 195503 76910
rect 195502 76846 195508 76878
rect 195432 76638 195508 76846
rect 195432 76574 195438 76638
rect 195502 76574 195508 76638
rect 195432 76568 195508 76574
rect 22309 76502 22375 76503
rect 22309 76470 22310 76502
rect 22304 76438 22310 76470
rect 22374 76470 22375 76502
rect 22445 76502 22511 76503
rect 22445 76470 22446 76502
rect 22374 76438 22380 76470
rect 952 76166 1230 76230
rect 1294 76166 1300 76230
rect 952 74598 1300 76166
rect 21760 76230 21836 76236
rect 21760 76166 21766 76230
rect 21830 76166 21836 76230
rect 21760 75958 21836 76166
rect 22304 76230 22380 76438
rect 22304 76166 22310 76230
rect 22374 76166 22380 76230
rect 22304 76160 22380 76166
rect 22440 76438 22446 76470
rect 22510 76470 22511 76502
rect 195845 76502 195911 76503
rect 195845 76470 195846 76502
rect 22510 76438 22516 76470
rect 22440 76230 22516 76438
rect 195840 76438 195846 76470
rect 195910 76470 195911 76502
rect 196117 76502 196183 76503
rect 196117 76470 196118 76502
rect 195910 76438 195916 76470
rect 28565 76366 28631 76367
rect 28565 76334 28566 76366
rect 22440 76166 22446 76230
rect 22510 76166 22516 76230
rect 22440 76160 22516 76166
rect 28560 76302 28566 76334
rect 28630 76334 28631 76366
rect 190269 76366 190335 76367
rect 190269 76334 190270 76366
rect 28630 76302 28636 76334
rect 28560 76094 28636 76302
rect 28560 76030 28566 76094
rect 28630 76030 28636 76094
rect 28560 76024 28636 76030
rect 190264 76302 190270 76334
rect 190334 76334 190335 76366
rect 190334 76302 190340 76334
rect 190264 76094 190340 76302
rect 195840 76230 195916 76438
rect 195840 76166 195846 76230
rect 195910 76166 195916 76230
rect 195840 76160 195916 76166
rect 196112 76438 196118 76470
rect 196182 76470 196183 76502
rect 196182 76438 196188 76470
rect 196112 76230 196188 76438
rect 196112 76166 196118 76230
rect 196182 76166 196188 76230
rect 196797 76230 196863 76231
rect 196797 76198 196798 76230
rect 196112 76160 196188 76166
rect 196792 76166 196798 76198
rect 196862 76198 196863 76230
rect 196862 76166 196868 76198
rect 190264 76030 190270 76094
rect 190334 76030 190340 76094
rect 190264 76024 190340 76030
rect 21760 75926 21766 75958
rect 21765 75894 21766 75926
rect 21830 75926 21836 75958
rect 28424 75958 28500 75964
rect 21830 75894 21831 75926
rect 21765 75893 21831 75894
rect 28424 75894 28430 75958
rect 28494 75894 28500 75958
rect 190133 75958 190199 75959
rect 190133 75926 190134 75958
rect 21765 75822 21831 75823
rect 21765 75790 21766 75822
rect 21760 75758 21766 75790
rect 21830 75790 21831 75822
rect 22173 75822 22239 75823
rect 22173 75790 22174 75822
rect 21830 75758 21836 75790
rect 21760 75550 21836 75758
rect 21760 75486 21766 75550
rect 21830 75486 21836 75550
rect 21760 75480 21836 75486
rect 22168 75758 22174 75790
rect 22238 75790 22239 75822
rect 22440 75822 22516 75828
rect 22238 75758 22244 75790
rect 22168 75550 22244 75758
rect 22168 75486 22174 75550
rect 22238 75486 22244 75550
rect 22440 75758 22446 75822
rect 22510 75758 22516 75822
rect 22440 75550 22516 75758
rect 23261 75686 23327 75687
rect 23261 75654 23262 75686
rect 22440 75518 22446 75550
rect 22168 75480 22244 75486
rect 22445 75486 22446 75518
rect 22510 75518 22516 75550
rect 23256 75622 23262 75654
rect 23326 75654 23327 75686
rect 28424 75686 28500 75894
rect 28424 75654 28430 75686
rect 23326 75622 23332 75654
rect 22510 75486 22511 75518
rect 22445 75485 22511 75486
rect 21901 75414 21967 75415
rect 21901 75382 21902 75414
rect 21896 75350 21902 75382
rect 21966 75382 21967 75414
rect 23120 75414 23196 75420
rect 21966 75350 21972 75382
rect 21896 75142 21972 75350
rect 21896 75078 21902 75142
rect 21966 75078 21972 75142
rect 23120 75350 23126 75414
rect 23190 75350 23196 75414
rect 23120 75142 23196 75350
rect 23256 75278 23332 75622
rect 28429 75622 28430 75654
rect 28494 75654 28500 75686
rect 190128 75894 190134 75926
rect 190198 75926 190199 75958
rect 196792 75958 196868 76166
rect 190198 75894 190204 75926
rect 190128 75686 190204 75894
rect 196792 75894 196798 75958
rect 196862 75894 196868 75958
rect 196792 75888 196868 75894
rect 217464 76094 217812 77798
rect 217464 76030 217470 76094
rect 217534 76030 217812 76094
rect 28494 75622 28495 75654
rect 28429 75621 28495 75622
rect 190128 75622 190134 75686
rect 190198 75622 190204 75686
rect 190128 75616 190204 75622
rect 196112 75822 196188 75828
rect 196112 75758 196118 75822
rect 196182 75758 196188 75822
rect 28429 75550 28495 75551
rect 28429 75518 28430 75550
rect 28424 75486 28430 75518
rect 28494 75518 28495 75550
rect 190264 75550 190340 75556
rect 28494 75486 28500 75518
rect 23256 75214 23262 75278
rect 23326 75214 23332 75278
rect 23256 75208 23332 75214
rect 23392 75414 23468 75420
rect 23392 75350 23398 75414
rect 23462 75350 23468 75414
rect 23120 75110 23126 75142
rect 21896 75072 21972 75078
rect 23125 75078 23126 75110
rect 23190 75110 23196 75142
rect 23392 75142 23468 75350
rect 23392 75110 23398 75142
rect 23190 75078 23191 75110
rect 23125 75077 23191 75078
rect 23397 75078 23398 75110
rect 23462 75110 23468 75142
rect 25296 75414 25372 75420
rect 25296 75350 25302 75414
rect 25366 75350 25372 75414
rect 25296 75142 25372 75350
rect 28424 75278 28500 75486
rect 28424 75214 28430 75278
rect 28494 75214 28500 75278
rect 190264 75486 190270 75550
rect 190334 75486 190340 75550
rect 196112 75550 196188 75758
rect 196112 75518 196118 75550
rect 190264 75278 190340 75486
rect 196117 75486 196118 75518
rect 196182 75518 196188 75550
rect 196384 75822 196460 75828
rect 196384 75758 196390 75822
rect 196454 75758 196460 75822
rect 196661 75822 196727 75823
rect 196661 75790 196662 75822
rect 196384 75550 196460 75758
rect 196384 75518 196390 75550
rect 196182 75486 196183 75518
rect 196117 75485 196183 75486
rect 196389 75486 196390 75518
rect 196454 75518 196460 75550
rect 196656 75758 196662 75790
rect 196726 75790 196727 75822
rect 196726 75758 196732 75790
rect 196656 75550 196732 75758
rect 196454 75486 196455 75518
rect 196389 75485 196455 75486
rect 196656 75486 196662 75550
rect 196726 75486 196732 75550
rect 196656 75480 196732 75486
rect 190264 75246 190270 75278
rect 28424 75208 28500 75214
rect 190269 75214 190270 75246
rect 190334 75246 190340 75278
rect 193120 75414 193196 75420
rect 193120 75350 193126 75414
rect 193190 75350 193196 75414
rect 195029 75414 195095 75415
rect 195029 75382 195030 75414
rect 190334 75214 190335 75246
rect 190269 75213 190335 75214
rect 25296 75110 25302 75142
rect 23462 75078 23463 75110
rect 23397 75077 23463 75078
rect 25301 75078 25302 75110
rect 25366 75110 25372 75142
rect 193120 75142 193196 75350
rect 193120 75110 193126 75142
rect 25366 75078 25367 75110
rect 25301 75077 25367 75078
rect 193125 75078 193126 75110
rect 193190 75110 193196 75142
rect 195024 75350 195030 75382
rect 195094 75382 195095 75414
rect 195437 75414 195503 75415
rect 195437 75382 195438 75414
rect 195094 75350 195100 75382
rect 195024 75142 195100 75350
rect 193190 75078 193191 75110
rect 193125 75077 193191 75078
rect 195024 75078 195030 75142
rect 195094 75078 195100 75142
rect 195024 75072 195100 75078
rect 195432 75350 195438 75382
rect 195502 75382 195503 75414
rect 196792 75414 196868 75420
rect 195502 75350 195508 75382
rect 195432 75142 195508 75350
rect 195432 75078 195438 75142
rect 195502 75078 195508 75142
rect 196792 75350 196798 75414
rect 196862 75350 196868 75414
rect 196792 75142 196868 75350
rect 196792 75110 196798 75142
rect 195432 75072 195508 75078
rect 196797 75078 196798 75110
rect 196862 75110 196868 75142
rect 196862 75078 196863 75110
rect 196797 75077 196863 75078
rect 21760 75006 21836 75012
rect 21760 74942 21766 75006
rect 21830 74942 21836 75006
rect 21760 74734 21836 74942
rect 21760 74702 21766 74734
rect 21765 74670 21766 74702
rect 21830 74702 21836 74734
rect 22168 75006 22244 75012
rect 22168 74942 22174 75006
rect 22238 74942 22244 75006
rect 22989 75006 23055 75007
rect 22989 74974 22990 75006
rect 22168 74734 22244 74942
rect 22168 74702 22174 74734
rect 21830 74670 21831 74702
rect 21765 74669 21831 74670
rect 22173 74670 22174 74702
rect 22238 74702 22244 74734
rect 22984 74942 22990 74974
rect 23054 74974 23055 75006
rect 23533 75006 23599 75007
rect 23533 74974 23534 75006
rect 23054 74942 23060 74974
rect 22984 74734 23060 74942
rect 22238 74670 22239 74702
rect 22173 74669 22239 74670
rect 22984 74670 22990 74734
rect 23054 74670 23060 74734
rect 22984 74664 23060 74670
rect 23528 74942 23534 74974
rect 23598 74974 23599 75006
rect 195160 75006 195236 75012
rect 23598 74942 23604 74974
rect 23528 74734 23604 74942
rect 23528 74670 23534 74734
rect 23598 74670 23604 74734
rect 195160 74942 195166 75006
rect 195230 74942 195236 75006
rect 195437 75006 195503 75007
rect 195437 74974 195438 75006
rect 195160 74734 195236 74942
rect 195160 74702 195166 74734
rect 23528 74664 23604 74670
rect 195165 74670 195166 74702
rect 195230 74702 195236 74734
rect 195432 74942 195438 74974
rect 195502 74974 195503 75006
rect 196248 75006 196324 75012
rect 195502 74942 195508 74974
rect 195432 74734 195508 74942
rect 195230 74670 195231 74702
rect 195165 74669 195231 74670
rect 195432 74670 195438 74734
rect 195502 74670 195508 74734
rect 196248 74942 196254 75006
rect 196318 74942 196324 75006
rect 196661 75006 196727 75007
rect 196661 74974 196662 75006
rect 196248 74734 196324 74942
rect 196248 74702 196254 74734
rect 195432 74664 195508 74670
rect 196253 74670 196254 74702
rect 196318 74702 196324 74734
rect 196656 74942 196662 74974
rect 196726 74974 196727 75006
rect 196726 74942 196732 74974
rect 196656 74734 196732 74942
rect 196318 74670 196319 74702
rect 196253 74669 196319 74670
rect 196656 74670 196662 74734
rect 196726 74670 196732 74734
rect 196656 74664 196732 74670
rect 952 74534 1230 74598
rect 1294 74534 1300 74598
rect 21765 74598 21831 74599
rect 21765 74566 21766 74598
rect 952 72694 1300 74534
rect 21760 74534 21766 74566
rect 21830 74566 21831 74598
rect 22984 74598 23060 74604
rect 21830 74534 21836 74566
rect 21760 74326 21836 74534
rect 21760 74262 21766 74326
rect 21830 74262 21836 74326
rect 22984 74534 22990 74598
rect 23054 74534 23060 74598
rect 23533 74598 23599 74599
rect 23533 74566 23534 74598
rect 22984 74326 23060 74534
rect 22984 74294 22990 74326
rect 21760 74256 21836 74262
rect 22989 74262 22990 74294
rect 23054 74294 23060 74326
rect 23528 74534 23534 74566
rect 23598 74566 23599 74598
rect 195165 74598 195231 74599
rect 195165 74566 195166 74598
rect 23598 74534 23604 74566
rect 23528 74326 23604 74534
rect 23054 74262 23055 74294
rect 22989 74261 23055 74262
rect 23528 74262 23534 74326
rect 23598 74262 23604 74326
rect 23528 74256 23604 74262
rect 195160 74534 195166 74566
rect 195230 74566 195231 74598
rect 195432 74598 195508 74604
rect 195230 74534 195236 74566
rect 195160 74326 195236 74534
rect 195160 74262 195166 74326
rect 195230 74262 195236 74326
rect 195432 74534 195438 74598
rect 195502 74534 195508 74598
rect 195845 74598 195911 74599
rect 195845 74566 195846 74598
rect 195432 74326 195508 74534
rect 195432 74294 195438 74326
rect 195160 74256 195236 74262
rect 195437 74262 195438 74294
rect 195502 74294 195508 74326
rect 195840 74534 195846 74566
rect 195910 74566 195911 74598
rect 196384 74598 196460 74604
rect 195910 74534 195916 74566
rect 195840 74326 195916 74534
rect 195502 74262 195503 74294
rect 195437 74261 195503 74262
rect 195840 74262 195846 74326
rect 195910 74262 195916 74326
rect 196384 74534 196390 74598
rect 196454 74534 196460 74598
rect 196384 74326 196460 74534
rect 196384 74294 196390 74326
rect 195840 74256 195916 74262
rect 196389 74262 196390 74294
rect 196454 74294 196460 74326
rect 196792 74598 196868 74604
rect 196792 74534 196798 74598
rect 196862 74534 196868 74598
rect 196792 74326 196868 74534
rect 196792 74294 196798 74326
rect 196454 74262 196455 74294
rect 196389 74261 196455 74262
rect 196797 74262 196798 74294
rect 196862 74294 196868 74326
rect 217464 74598 217812 76030
rect 217464 74534 217470 74598
rect 217534 74534 217812 74598
rect 196862 74262 196863 74294
rect 196797 74261 196863 74262
rect 21760 74190 21836 74196
rect 21760 74126 21766 74190
rect 21830 74126 21836 74190
rect 21760 73918 21836 74126
rect 21760 73886 21766 73918
rect 21765 73854 21766 73886
rect 21830 73886 21836 73918
rect 22168 74190 22244 74196
rect 22168 74126 22174 74190
rect 22238 74126 22244 74190
rect 22717 74190 22783 74191
rect 22717 74158 22718 74190
rect 22168 73918 22244 74126
rect 22168 73886 22174 73918
rect 21830 73854 21831 73886
rect 21765 73853 21831 73854
rect 22173 73854 22174 73886
rect 22238 73886 22244 73918
rect 22712 74126 22718 74158
rect 22782 74158 22783 74190
rect 22989 74190 23055 74191
rect 22989 74158 22990 74190
rect 22782 74126 22788 74158
rect 22712 73918 22788 74126
rect 22238 73854 22239 73886
rect 22173 73853 22239 73854
rect 22712 73854 22718 73918
rect 22782 73854 22788 73918
rect 22712 73848 22788 73854
rect 22984 74126 22990 74158
rect 23054 74158 23055 74190
rect 23528 74190 23604 74196
rect 23054 74126 23060 74158
rect 22984 73918 23060 74126
rect 22984 73854 22990 73918
rect 23054 73854 23060 73918
rect 23528 74126 23534 74190
rect 23598 74126 23604 74190
rect 23528 73918 23604 74126
rect 23528 73886 23534 73918
rect 22984 73848 23060 73854
rect 23533 73854 23534 73886
rect 23598 73886 23604 73918
rect 195160 74190 195236 74196
rect 195160 74126 195166 74190
rect 195230 74126 195236 74190
rect 195160 73918 195236 74126
rect 195160 73886 195166 73918
rect 23598 73854 23599 73886
rect 23533 73853 23599 73854
rect 195165 73854 195166 73886
rect 195230 73886 195236 73918
rect 195432 74190 195508 74196
rect 195432 74126 195438 74190
rect 195502 74126 195508 74190
rect 196117 74190 196183 74191
rect 196117 74158 196118 74190
rect 195432 73918 195508 74126
rect 195432 73886 195438 73918
rect 195230 73854 195231 73886
rect 195165 73853 195231 73854
rect 195437 73854 195438 73886
rect 195502 73886 195508 73918
rect 196112 74126 196118 74158
rect 196182 74158 196183 74190
rect 196656 74190 196732 74196
rect 196182 74126 196188 74158
rect 196112 73918 196188 74126
rect 195502 73854 195503 73886
rect 195437 73853 195503 73854
rect 196112 73854 196118 73918
rect 196182 73854 196188 73918
rect 196656 74126 196662 74190
rect 196726 74126 196732 74190
rect 196656 73918 196732 74126
rect 196656 73886 196662 73918
rect 196112 73848 196188 73854
rect 196661 73854 196662 73886
rect 196726 73886 196732 73918
rect 196726 73854 196727 73886
rect 196661 73853 196727 73854
rect 21765 73782 21831 73783
rect 21765 73750 21766 73782
rect 21760 73718 21766 73750
rect 21830 73750 21831 73782
rect 22576 73782 22652 73788
rect 21830 73718 21836 73750
rect 21760 73510 21836 73718
rect 21760 73446 21766 73510
rect 21830 73446 21836 73510
rect 22576 73718 22582 73782
rect 22646 73718 22652 73782
rect 22576 73510 22652 73718
rect 22576 73478 22582 73510
rect 21760 73440 21836 73446
rect 22581 73446 22582 73478
rect 22646 73478 22652 73510
rect 23120 73782 23196 73788
rect 23120 73718 23126 73782
rect 23190 73718 23196 73782
rect 23533 73782 23599 73783
rect 23533 73750 23534 73782
rect 23120 73510 23196 73718
rect 23120 73478 23126 73510
rect 22646 73446 22647 73478
rect 22581 73445 22647 73446
rect 23125 73446 23126 73478
rect 23190 73478 23196 73510
rect 23528 73718 23534 73750
rect 23598 73750 23599 73782
rect 195165 73782 195231 73783
rect 195165 73750 195166 73782
rect 23598 73718 23604 73750
rect 23528 73510 23604 73718
rect 23190 73446 23191 73478
rect 23125 73445 23191 73446
rect 23528 73446 23534 73510
rect 23598 73446 23604 73510
rect 23528 73440 23604 73446
rect 195160 73718 195166 73750
rect 195230 73750 195231 73782
rect 195568 73782 195644 73788
rect 195230 73718 195236 73750
rect 195160 73510 195236 73718
rect 195160 73446 195166 73510
rect 195230 73446 195236 73510
rect 195568 73718 195574 73782
rect 195638 73718 195644 73782
rect 195568 73510 195644 73718
rect 195568 73478 195574 73510
rect 195160 73440 195236 73446
rect 195573 73446 195574 73478
rect 195638 73478 195644 73510
rect 195840 73782 195916 73788
rect 195840 73718 195846 73782
rect 195910 73718 195916 73782
rect 195840 73510 195916 73718
rect 195840 73478 195846 73510
rect 195638 73446 195639 73478
rect 195573 73445 195639 73446
rect 195845 73446 195846 73478
rect 195910 73478 195916 73510
rect 196248 73782 196324 73788
rect 196248 73718 196254 73782
rect 196318 73718 196324 73782
rect 196661 73782 196727 73783
rect 196661 73750 196662 73782
rect 196248 73510 196324 73718
rect 196248 73478 196254 73510
rect 195910 73446 195911 73478
rect 195845 73445 195911 73446
rect 196253 73446 196254 73478
rect 196318 73478 196324 73510
rect 196656 73718 196662 73750
rect 196726 73750 196727 73782
rect 196726 73718 196732 73750
rect 196656 73510 196732 73718
rect 196318 73446 196319 73478
rect 196253 73445 196319 73446
rect 196656 73446 196662 73510
rect 196726 73446 196732 73510
rect 196656 73440 196732 73446
rect 22173 73374 22239 73375
rect 22173 73342 22174 73374
rect 22168 73310 22174 73342
rect 22238 73342 22239 73374
rect 22712 73374 22788 73380
rect 22238 73310 22244 73342
rect 22168 73102 22244 73310
rect 22168 73038 22174 73102
rect 22238 73038 22244 73102
rect 22712 73310 22718 73374
rect 22782 73310 22788 73374
rect 22712 73102 22788 73310
rect 22712 73070 22718 73102
rect 22168 73032 22244 73038
rect 22717 73038 22718 73070
rect 22782 73070 22788 73102
rect 23120 73374 23196 73380
rect 23120 73310 23126 73374
rect 23190 73310 23196 73374
rect 23397 73374 23463 73375
rect 23397 73342 23398 73374
rect 23120 73102 23196 73310
rect 23120 73070 23126 73102
rect 22782 73038 22783 73070
rect 22717 73037 22783 73038
rect 23125 73038 23126 73070
rect 23190 73070 23196 73102
rect 23392 73310 23398 73342
rect 23462 73342 23463 73374
rect 195024 73374 195100 73380
rect 23462 73310 23468 73342
rect 23392 73102 23468 73310
rect 23190 73038 23191 73070
rect 23125 73037 23191 73038
rect 23392 73038 23398 73102
rect 23462 73038 23468 73102
rect 195024 73310 195030 73374
rect 195094 73310 195100 73374
rect 195437 73374 195503 73375
rect 195437 73342 195438 73374
rect 195024 73102 195100 73310
rect 195024 73070 195030 73102
rect 23392 73032 23468 73038
rect 195029 73038 195030 73070
rect 195094 73070 195100 73102
rect 195432 73310 195438 73342
rect 195502 73342 195503 73374
rect 195981 73374 196047 73375
rect 195981 73342 195982 73374
rect 195502 73310 195508 73342
rect 195432 73102 195508 73310
rect 195094 73038 195095 73070
rect 195029 73037 195095 73038
rect 195432 73038 195438 73102
rect 195502 73038 195508 73102
rect 195432 73032 195508 73038
rect 195976 73310 195982 73342
rect 196046 73342 196047 73374
rect 196112 73374 196188 73380
rect 196046 73310 196052 73342
rect 195976 73102 196052 73310
rect 195976 73038 195982 73102
rect 196046 73038 196052 73102
rect 196112 73310 196118 73374
rect 196182 73310 196188 73374
rect 196112 73102 196188 73310
rect 196112 73070 196118 73102
rect 195976 73032 196052 73038
rect 196117 73038 196118 73070
rect 196182 73070 196188 73102
rect 196182 73038 196183 73070
rect 196117 73037 196183 73038
rect 23125 72966 23191 72967
rect 23125 72934 23126 72966
rect 952 72630 1230 72694
rect 1294 72630 1300 72694
rect 952 71062 1300 72630
rect 23120 72902 23126 72934
rect 23190 72934 23191 72966
rect 23528 72966 23604 72972
rect 23190 72902 23196 72934
rect 23120 72694 23196 72902
rect 23120 72630 23126 72694
rect 23190 72630 23196 72694
rect 23528 72902 23534 72966
rect 23598 72902 23604 72966
rect 28293 72966 28359 72967
rect 28293 72934 28294 72966
rect 23528 72694 23604 72902
rect 23528 72662 23534 72694
rect 23120 72624 23196 72630
rect 23533 72630 23534 72662
rect 23598 72662 23604 72694
rect 28288 72902 28294 72934
rect 28358 72934 28359 72966
rect 195029 72966 195095 72967
rect 195029 72934 195030 72966
rect 28358 72902 28364 72934
rect 23598 72630 23599 72662
rect 23533 72629 23599 72630
rect 22717 72558 22783 72559
rect 22717 72526 22718 72558
rect 22712 72494 22718 72526
rect 22782 72526 22783 72558
rect 22984 72558 23060 72564
rect 22782 72494 22788 72526
rect 21901 72286 21967 72287
rect 21901 72254 21902 72286
rect 21896 72222 21902 72254
rect 21966 72254 21967 72286
rect 22712 72286 22788 72494
rect 21966 72222 21972 72254
rect 21896 72014 21972 72222
rect 22712 72222 22718 72286
rect 22782 72222 22788 72286
rect 22984 72494 22990 72558
rect 23054 72494 23060 72558
rect 22984 72286 23060 72494
rect 22984 72254 22990 72286
rect 22712 72216 22788 72222
rect 22989 72222 22990 72254
rect 23054 72254 23060 72286
rect 23392 72558 23468 72564
rect 23392 72494 23398 72558
rect 23462 72494 23468 72558
rect 23392 72286 23468 72494
rect 28288 72558 28364 72902
rect 195024 72902 195030 72934
rect 195094 72934 195095 72966
rect 195573 72966 195639 72967
rect 195573 72934 195574 72966
rect 195094 72902 195100 72934
rect 195024 72694 195100 72902
rect 195024 72630 195030 72694
rect 195094 72630 195100 72694
rect 195024 72624 195100 72630
rect 195568 72902 195574 72934
rect 195638 72934 195639 72966
rect 195638 72902 195644 72934
rect 195568 72694 195644 72902
rect 195568 72630 195574 72694
rect 195638 72630 195644 72694
rect 195568 72624 195644 72630
rect 217464 72830 217812 74534
rect 217464 72766 217470 72830
rect 217534 72766 217812 72830
rect 28288 72494 28294 72558
rect 28358 72494 28364 72558
rect 28288 72488 28364 72494
rect 195024 72558 195100 72564
rect 195024 72494 195030 72558
rect 195094 72494 195100 72558
rect 195437 72558 195503 72559
rect 195437 72526 195438 72558
rect 28565 72422 28631 72423
rect 28565 72390 28566 72422
rect 23392 72254 23398 72286
rect 23054 72222 23055 72254
rect 22989 72221 23055 72222
rect 23397 72222 23398 72254
rect 23462 72254 23468 72286
rect 28560 72358 28566 72390
rect 28630 72390 28631 72422
rect 28630 72358 28636 72390
rect 23462 72222 23463 72254
rect 23397 72221 23463 72222
rect 28560 72150 28636 72358
rect 195024 72286 195100 72494
rect 195024 72254 195030 72286
rect 195029 72222 195030 72254
rect 195094 72254 195100 72286
rect 195432 72494 195438 72526
rect 195502 72526 195503 72558
rect 196112 72558 196188 72564
rect 195502 72494 195508 72526
rect 195432 72286 195508 72494
rect 195094 72222 195095 72254
rect 195029 72221 195095 72222
rect 195432 72222 195438 72286
rect 195502 72222 195508 72286
rect 196112 72494 196118 72558
rect 196182 72494 196188 72558
rect 196112 72286 196188 72494
rect 196112 72254 196118 72286
rect 195432 72216 195508 72222
rect 196117 72222 196118 72254
rect 196182 72254 196188 72286
rect 196792 72286 196868 72292
rect 196182 72222 196183 72254
rect 196117 72221 196183 72222
rect 196792 72222 196798 72286
rect 196862 72222 196868 72286
rect 28560 72086 28566 72150
rect 28630 72086 28636 72150
rect 28560 72080 28636 72086
rect 21896 71950 21902 72014
rect 21966 71950 21972 72014
rect 28565 72014 28631 72015
rect 28565 71982 28566 72014
rect 21896 71944 21972 71950
rect 28560 71950 28566 71982
rect 28630 71982 28631 72014
rect 190128 72014 190204 72020
rect 28630 71950 28636 71982
rect 21901 71878 21967 71879
rect 21901 71846 21902 71878
rect 21896 71814 21902 71846
rect 21966 71846 21967 71878
rect 22309 71878 22375 71879
rect 22309 71846 22310 71878
rect 21966 71814 21972 71846
rect 21896 71606 21972 71814
rect 21896 71542 21902 71606
rect 21966 71542 21972 71606
rect 21896 71536 21972 71542
rect 22304 71814 22310 71846
rect 22374 71846 22375 71878
rect 22445 71878 22511 71879
rect 22445 71846 22446 71878
rect 22374 71814 22380 71846
rect 22304 71606 22380 71814
rect 22304 71542 22310 71606
rect 22374 71542 22380 71606
rect 22304 71536 22380 71542
rect 22440 71814 22446 71846
rect 22510 71846 22511 71878
rect 22510 71814 22516 71846
rect 22440 71606 22516 71814
rect 28560 71742 28636 71950
rect 28560 71678 28566 71742
rect 28630 71678 28636 71742
rect 190128 71950 190134 72014
rect 190198 71950 190204 72014
rect 196792 72014 196868 72222
rect 196792 71982 196798 72014
rect 190128 71742 190204 71950
rect 196797 71950 196798 71982
rect 196862 71982 196868 72014
rect 196862 71950 196863 71982
rect 196797 71949 196863 71950
rect 196389 71878 196455 71879
rect 196389 71846 196390 71878
rect 190128 71710 190134 71742
rect 28560 71672 28636 71678
rect 190133 71678 190134 71710
rect 190198 71710 190204 71742
rect 196384 71814 196390 71846
rect 196454 71846 196455 71878
rect 196797 71878 196863 71879
rect 196797 71846 196798 71878
rect 196454 71814 196460 71846
rect 190198 71678 190199 71710
rect 190133 71677 190199 71678
rect 22440 71542 22446 71606
rect 22510 71542 22516 71606
rect 22440 71536 22516 71542
rect 190128 71606 190204 71612
rect 190128 71542 190134 71606
rect 190198 71542 190204 71606
rect 21896 71470 21972 71476
rect 21896 71406 21902 71470
rect 21966 71406 21972 71470
rect 21896 71198 21972 71406
rect 28429 71334 28495 71335
rect 28429 71302 28430 71334
rect 28424 71270 28430 71302
rect 28494 71302 28495 71334
rect 190128 71334 190204 71542
rect 196384 71606 196460 71814
rect 196384 71542 196390 71606
rect 196454 71542 196460 71606
rect 196384 71536 196460 71542
rect 196792 71814 196798 71846
rect 196862 71846 196863 71878
rect 196862 71814 196868 71846
rect 196792 71606 196868 71814
rect 196792 71542 196798 71606
rect 196862 71542 196868 71606
rect 196792 71536 196868 71542
rect 196661 71470 196727 71471
rect 196661 71438 196662 71470
rect 196656 71406 196662 71438
rect 196726 71438 196727 71470
rect 196726 71406 196732 71438
rect 190128 71302 190134 71334
rect 28494 71270 28500 71302
rect 21896 71166 21902 71198
rect 21901 71134 21902 71166
rect 21966 71166 21972 71198
rect 28288 71198 28364 71204
rect 21966 71134 21967 71166
rect 21901 71133 21967 71134
rect 28288 71134 28294 71198
rect 28358 71134 28364 71198
rect 952 70998 1230 71062
rect 1294 70998 1300 71062
rect 21901 71062 21967 71063
rect 21901 71030 21902 71062
rect 952 69430 1300 70998
rect 21896 70998 21902 71030
rect 21966 71030 21967 71062
rect 22989 71062 23055 71063
rect 22989 71030 22990 71062
rect 21966 70998 21972 71030
rect 21896 70790 21972 70998
rect 21896 70726 21902 70790
rect 21966 70726 21972 70790
rect 21896 70720 21972 70726
rect 22984 70998 22990 71030
rect 23054 71030 23055 71062
rect 23392 71062 23468 71068
rect 23054 70998 23060 71030
rect 22984 70790 23060 70998
rect 22984 70726 22990 70790
rect 23054 70726 23060 70790
rect 23392 70998 23398 71062
rect 23462 70998 23468 71062
rect 23392 70790 23468 70998
rect 23392 70758 23398 70790
rect 22984 70720 23060 70726
rect 23397 70726 23398 70758
rect 23462 70758 23468 70790
rect 28288 70790 28364 71134
rect 28424 71062 28500 71270
rect 190133 71270 190134 71302
rect 190198 71302 190204 71334
rect 190264 71334 190340 71340
rect 190198 71270 190199 71302
rect 190133 71269 190199 71270
rect 190264 71270 190270 71334
rect 190334 71270 190340 71334
rect 28424 70998 28430 71062
rect 28494 70998 28500 71062
rect 190264 71062 190340 71270
rect 196656 71198 196732 71406
rect 196656 71134 196662 71198
rect 196726 71134 196732 71198
rect 196656 71128 196732 71134
rect 217464 71198 217812 72766
rect 217464 71134 217470 71198
rect 217534 71134 217812 71198
rect 190264 71030 190270 71062
rect 28424 70992 28500 70998
rect 190269 70998 190270 71030
rect 190334 71030 190340 71062
rect 195029 71062 195095 71063
rect 195029 71030 195030 71062
rect 190334 70998 190335 71030
rect 190269 70997 190335 70998
rect 195024 70998 195030 71030
rect 195094 71030 195095 71062
rect 195568 71062 195644 71068
rect 195094 70998 195100 71030
rect 28288 70758 28294 70790
rect 23462 70726 23463 70758
rect 23397 70725 23463 70726
rect 28293 70726 28294 70758
rect 28358 70758 28364 70790
rect 28565 70790 28631 70791
rect 28565 70758 28566 70790
rect 28358 70726 28359 70758
rect 28293 70725 28359 70726
rect 28560 70726 28566 70758
rect 28630 70758 28631 70790
rect 190128 70790 190204 70796
rect 28630 70726 28636 70758
rect 21765 70654 21831 70655
rect 21765 70622 21766 70654
rect 21760 70590 21766 70622
rect 21830 70622 21831 70654
rect 22440 70654 22516 70660
rect 21830 70590 21836 70622
rect 21760 70382 21836 70590
rect 21760 70318 21766 70382
rect 21830 70318 21836 70382
rect 22440 70590 22446 70654
rect 22510 70590 22516 70654
rect 22989 70654 23055 70655
rect 22989 70622 22990 70654
rect 22440 70382 22516 70590
rect 22440 70350 22446 70382
rect 21760 70312 21836 70318
rect 22445 70318 22446 70350
rect 22510 70350 22516 70382
rect 22984 70590 22990 70622
rect 23054 70622 23055 70654
rect 23533 70654 23599 70655
rect 23533 70622 23534 70654
rect 23054 70590 23060 70622
rect 22984 70382 23060 70590
rect 22510 70318 22511 70350
rect 22445 70317 22511 70318
rect 22984 70318 22990 70382
rect 23054 70318 23060 70382
rect 22984 70312 23060 70318
rect 23528 70590 23534 70622
rect 23598 70622 23599 70654
rect 23598 70590 23604 70622
rect 23528 70382 23604 70590
rect 28560 70518 28636 70726
rect 28560 70454 28566 70518
rect 28630 70454 28636 70518
rect 190128 70726 190134 70790
rect 190198 70726 190204 70790
rect 190128 70518 190204 70726
rect 195024 70790 195100 70998
rect 195024 70726 195030 70790
rect 195094 70726 195100 70790
rect 195568 70998 195574 71062
rect 195638 70998 195644 71062
rect 196389 71062 196455 71063
rect 196389 71030 196390 71062
rect 195568 70790 195644 70998
rect 195568 70758 195574 70790
rect 195024 70720 195100 70726
rect 195573 70726 195574 70758
rect 195638 70758 195644 70790
rect 196384 70998 196390 71030
rect 196454 71030 196455 71062
rect 196792 71062 196868 71068
rect 196454 70998 196460 71030
rect 196384 70790 196460 70998
rect 195638 70726 195639 70758
rect 195573 70725 195639 70726
rect 196384 70726 196390 70790
rect 196454 70726 196460 70790
rect 196792 70998 196798 71062
rect 196862 70998 196868 71062
rect 196792 70790 196868 70998
rect 196792 70758 196798 70790
rect 196384 70720 196460 70726
rect 196797 70726 196798 70758
rect 196862 70758 196868 70790
rect 196862 70726 196863 70758
rect 196797 70725 196863 70726
rect 195165 70654 195231 70655
rect 195165 70622 195166 70654
rect 190128 70486 190134 70518
rect 28560 70448 28636 70454
rect 190133 70454 190134 70486
rect 190198 70486 190204 70518
rect 195160 70590 195166 70622
rect 195230 70622 195231 70654
rect 195437 70654 195503 70655
rect 195437 70622 195438 70654
rect 195230 70590 195236 70622
rect 190198 70454 190199 70486
rect 190133 70453 190199 70454
rect 23528 70318 23534 70382
rect 23598 70318 23604 70382
rect 23528 70312 23604 70318
rect 195160 70382 195236 70590
rect 195160 70318 195166 70382
rect 195230 70318 195236 70382
rect 195160 70312 195236 70318
rect 195432 70590 195438 70622
rect 195502 70622 195503 70654
rect 196117 70654 196183 70655
rect 196117 70622 196118 70654
rect 195502 70590 195508 70622
rect 195432 70382 195508 70590
rect 195432 70318 195438 70382
rect 195502 70318 195508 70382
rect 195432 70312 195508 70318
rect 196112 70590 196118 70622
rect 196182 70622 196183 70654
rect 196248 70654 196324 70660
rect 196182 70590 196188 70622
rect 196112 70382 196188 70590
rect 196112 70318 196118 70382
rect 196182 70318 196188 70382
rect 196248 70590 196254 70654
rect 196318 70590 196324 70654
rect 196248 70382 196324 70590
rect 196248 70350 196254 70382
rect 196112 70312 196188 70318
rect 196253 70318 196254 70350
rect 196318 70350 196324 70382
rect 196656 70654 196732 70660
rect 196656 70590 196662 70654
rect 196726 70590 196732 70654
rect 196656 70382 196732 70590
rect 196656 70350 196662 70382
rect 196318 70318 196319 70350
rect 196253 70317 196319 70318
rect 196661 70318 196662 70350
rect 196726 70350 196732 70382
rect 196726 70318 196727 70350
rect 196661 70317 196727 70318
rect 21896 70246 21972 70252
rect 21896 70182 21902 70246
rect 21966 70182 21972 70246
rect 21896 69974 21972 70182
rect 21896 69942 21902 69974
rect 21901 69910 21902 69942
rect 21966 69942 21972 69974
rect 22304 70246 22380 70252
rect 22304 70182 22310 70246
rect 22374 70182 22380 70246
rect 22581 70246 22647 70247
rect 22581 70214 22582 70246
rect 22304 69974 22380 70182
rect 22304 69942 22310 69974
rect 21966 69910 21967 69942
rect 21901 69909 21967 69910
rect 22309 69910 22310 69942
rect 22374 69942 22380 69974
rect 22576 70182 22582 70214
rect 22646 70214 22647 70246
rect 22984 70246 23060 70252
rect 22646 70182 22652 70214
rect 22576 69974 22652 70182
rect 22374 69910 22375 69942
rect 22309 69909 22375 69910
rect 22576 69910 22582 69974
rect 22646 69910 22652 69974
rect 22984 70182 22990 70246
rect 23054 70182 23060 70246
rect 23533 70246 23599 70247
rect 23533 70214 23534 70246
rect 22984 69974 23060 70182
rect 22984 69942 22990 69974
rect 22576 69904 22652 69910
rect 22989 69910 22990 69942
rect 23054 69942 23060 69974
rect 23528 70182 23534 70214
rect 23598 70214 23599 70246
rect 195024 70246 195100 70252
rect 23598 70182 23604 70214
rect 23528 69974 23604 70182
rect 23054 69910 23055 69942
rect 22989 69909 23055 69910
rect 23528 69910 23534 69974
rect 23598 69910 23604 69974
rect 195024 70182 195030 70246
rect 195094 70182 195100 70246
rect 195024 69974 195100 70182
rect 195024 69942 195030 69974
rect 23528 69904 23604 69910
rect 195029 69910 195030 69942
rect 195094 69942 195100 69974
rect 195432 70246 195508 70252
rect 195432 70182 195438 70246
rect 195502 70182 195508 70246
rect 195432 69974 195508 70182
rect 195432 69942 195438 69974
rect 195094 69910 195095 69942
rect 195029 69909 195095 69910
rect 195437 69910 195438 69942
rect 195502 69942 195508 69974
rect 195976 70246 196052 70252
rect 195976 70182 195982 70246
rect 196046 70182 196052 70246
rect 195976 69974 196052 70182
rect 195976 69942 195982 69974
rect 195502 69910 195503 69942
rect 195437 69909 195503 69910
rect 195981 69910 195982 69942
rect 196046 69942 196052 69974
rect 196112 70246 196188 70252
rect 196112 70182 196118 70246
rect 196182 70182 196188 70246
rect 196661 70246 196727 70247
rect 196661 70214 196662 70246
rect 196112 69974 196188 70182
rect 196112 69942 196118 69974
rect 196046 69910 196047 69942
rect 195981 69909 196047 69910
rect 196117 69910 196118 69942
rect 196182 69942 196188 69974
rect 196656 70182 196662 70214
rect 196726 70214 196727 70246
rect 196726 70182 196732 70214
rect 196656 69974 196732 70182
rect 196182 69910 196183 69942
rect 196117 69909 196183 69910
rect 196656 69910 196662 69974
rect 196726 69910 196732 69974
rect 196656 69904 196732 69910
rect 21760 69838 21836 69844
rect 21760 69774 21766 69838
rect 21830 69774 21836 69838
rect 22309 69838 22375 69839
rect 22309 69806 22310 69838
rect 21760 69566 21836 69774
rect 21760 69534 21766 69566
rect 21765 69502 21766 69534
rect 21830 69534 21836 69566
rect 22304 69774 22310 69806
rect 22374 69806 22375 69838
rect 22576 69838 22652 69844
rect 22374 69774 22380 69806
rect 22304 69566 22380 69774
rect 21830 69502 21831 69534
rect 21765 69501 21831 69502
rect 22304 69502 22310 69566
rect 22374 69502 22380 69566
rect 22576 69774 22582 69838
rect 22646 69774 22652 69838
rect 22989 69838 23055 69839
rect 22989 69806 22990 69838
rect 22576 69566 22652 69774
rect 22576 69534 22582 69566
rect 22304 69496 22380 69502
rect 22581 69502 22582 69534
rect 22646 69534 22652 69566
rect 22984 69774 22990 69806
rect 23054 69806 23055 69838
rect 23528 69838 23604 69844
rect 23054 69774 23060 69806
rect 22984 69566 23060 69774
rect 22646 69502 22647 69534
rect 22581 69501 22647 69502
rect 22984 69502 22990 69566
rect 23054 69502 23060 69566
rect 23528 69774 23534 69838
rect 23598 69774 23604 69838
rect 195029 69838 195095 69839
rect 195029 69806 195030 69838
rect 23528 69566 23604 69774
rect 23528 69534 23534 69566
rect 22984 69496 23060 69502
rect 23533 69502 23534 69534
rect 23598 69534 23604 69566
rect 195024 69774 195030 69806
rect 195094 69806 195095 69838
rect 195437 69838 195503 69839
rect 195437 69806 195438 69838
rect 195094 69774 195100 69806
rect 195024 69566 195100 69774
rect 23598 69502 23599 69534
rect 23533 69501 23599 69502
rect 195024 69502 195030 69566
rect 195094 69502 195100 69566
rect 195024 69496 195100 69502
rect 195432 69774 195438 69806
rect 195502 69806 195503 69838
rect 196248 69838 196324 69844
rect 195502 69774 195508 69806
rect 195432 69566 195508 69774
rect 195432 69502 195438 69566
rect 195502 69502 195508 69566
rect 196248 69774 196254 69838
rect 196318 69774 196324 69838
rect 196797 69838 196863 69839
rect 196797 69806 196798 69838
rect 196248 69566 196324 69774
rect 196248 69534 196254 69566
rect 195432 69496 195508 69502
rect 196253 69502 196254 69534
rect 196318 69534 196324 69566
rect 196792 69774 196798 69806
rect 196862 69806 196863 69838
rect 196862 69774 196868 69806
rect 196792 69566 196868 69774
rect 196318 69502 196319 69534
rect 196253 69501 196319 69502
rect 196792 69502 196798 69566
rect 196862 69502 196868 69566
rect 196792 69496 196868 69502
rect 952 69366 1230 69430
rect 1294 69366 1300 69430
rect 22581 69430 22647 69431
rect 22581 69398 22582 69430
rect 952 67798 1300 69366
rect 22576 69366 22582 69398
rect 22646 69398 22647 69430
rect 22989 69430 23055 69431
rect 22989 69398 22990 69430
rect 22646 69366 22652 69398
rect 22576 69158 22652 69366
rect 22576 69094 22582 69158
rect 22646 69094 22652 69158
rect 22576 69088 22652 69094
rect 22984 69366 22990 69398
rect 23054 69398 23055 69430
rect 23528 69430 23604 69436
rect 23054 69366 23060 69398
rect 22984 69158 23060 69366
rect 22984 69094 22990 69158
rect 23054 69094 23060 69158
rect 23528 69366 23534 69430
rect 23598 69366 23604 69430
rect 23528 69158 23604 69366
rect 23528 69126 23534 69158
rect 22984 69088 23060 69094
rect 23533 69094 23534 69126
rect 23598 69126 23604 69158
rect 195160 69430 195236 69436
rect 195160 69366 195166 69430
rect 195230 69366 195236 69430
rect 195160 69158 195236 69366
rect 195160 69126 195166 69158
rect 23598 69094 23599 69126
rect 23533 69093 23599 69094
rect 195165 69094 195166 69126
rect 195230 69126 195236 69158
rect 195568 69430 195644 69436
rect 195568 69366 195574 69430
rect 195638 69366 195644 69430
rect 195845 69430 195911 69431
rect 195845 69398 195846 69430
rect 195568 69158 195644 69366
rect 195568 69126 195574 69158
rect 195230 69094 195231 69126
rect 195165 69093 195231 69094
rect 195573 69094 195574 69126
rect 195638 69126 195644 69158
rect 195840 69366 195846 69398
rect 195910 69398 195911 69430
rect 196112 69430 196188 69436
rect 195910 69366 195916 69398
rect 195840 69158 195916 69366
rect 195638 69094 195639 69126
rect 195573 69093 195639 69094
rect 195840 69094 195846 69158
rect 195910 69094 195916 69158
rect 196112 69366 196118 69430
rect 196182 69366 196188 69430
rect 196112 69158 196188 69366
rect 196112 69126 196118 69158
rect 195840 69088 195916 69094
rect 196117 69094 196118 69126
rect 196182 69126 196188 69158
rect 217464 69294 217812 71134
rect 217464 69230 217470 69294
rect 217534 69230 217812 69294
rect 196182 69094 196183 69126
rect 196117 69093 196183 69094
rect 21896 69022 21972 69028
rect 21896 68958 21902 69022
rect 21966 68958 21972 69022
rect 21896 68750 21972 68958
rect 21896 68718 21902 68750
rect 21901 68686 21902 68718
rect 21966 68718 21972 68750
rect 22712 69022 22788 69028
rect 22712 68958 22718 69022
rect 22782 68958 22788 69022
rect 22712 68750 22788 68958
rect 22712 68718 22718 68750
rect 21966 68686 21967 68718
rect 21901 68685 21967 68686
rect 22717 68686 22718 68718
rect 22782 68718 22788 68750
rect 23120 69022 23196 69028
rect 23120 68958 23126 69022
rect 23190 68958 23196 69022
rect 23397 69022 23463 69023
rect 23397 68990 23398 69022
rect 23120 68750 23196 68958
rect 23120 68718 23126 68750
rect 22782 68686 22783 68718
rect 22717 68685 22783 68686
rect 23125 68686 23126 68718
rect 23190 68718 23196 68750
rect 23392 68958 23398 68990
rect 23462 68990 23463 69022
rect 195024 69022 195100 69028
rect 23462 68958 23468 68990
rect 23392 68750 23468 68958
rect 23190 68686 23191 68718
rect 23125 68685 23191 68686
rect 23392 68686 23398 68750
rect 23462 68686 23468 68750
rect 195024 68958 195030 69022
rect 195094 68958 195100 69022
rect 195437 69022 195503 69023
rect 195437 68990 195438 69022
rect 195024 68750 195100 68958
rect 195024 68718 195030 68750
rect 23392 68680 23468 68686
rect 195029 68686 195030 68718
rect 195094 68718 195100 68750
rect 195432 68958 195438 68990
rect 195502 68990 195503 69022
rect 196797 69022 196863 69023
rect 196797 68990 196798 69022
rect 195502 68958 195508 68990
rect 195432 68750 195508 68958
rect 195094 68686 195095 68718
rect 195029 68685 195095 68686
rect 195432 68686 195438 68750
rect 195502 68686 195508 68750
rect 195432 68680 195508 68686
rect 196792 68958 196798 68990
rect 196862 68990 196863 69022
rect 196862 68958 196868 68990
rect 196792 68750 196868 68958
rect 196792 68686 196798 68750
rect 196862 68686 196868 68750
rect 196792 68680 196868 68686
rect 22309 68614 22375 68615
rect 22309 68582 22310 68614
rect 22304 68550 22310 68582
rect 22374 68582 22375 68614
rect 22984 68614 23060 68620
rect 22374 68550 22380 68582
rect 21765 68342 21831 68343
rect 21765 68310 21766 68342
rect 21760 68278 21766 68310
rect 21830 68310 21831 68342
rect 22304 68342 22380 68550
rect 21830 68278 21836 68310
rect 21760 68070 21836 68278
rect 22304 68278 22310 68342
rect 22374 68278 22380 68342
rect 22984 68550 22990 68614
rect 23054 68550 23060 68614
rect 22984 68342 23060 68550
rect 22984 68310 22990 68342
rect 22304 68272 22380 68278
rect 22989 68278 22990 68310
rect 23054 68310 23060 68342
rect 23528 68614 23604 68620
rect 23528 68550 23534 68614
rect 23598 68550 23604 68614
rect 195029 68614 195095 68615
rect 195029 68582 195030 68614
rect 23528 68342 23604 68550
rect 195024 68550 195030 68582
rect 195094 68582 195095 68614
rect 195573 68614 195639 68615
rect 195573 68582 195574 68614
rect 195094 68550 195100 68582
rect 190133 68478 190199 68479
rect 190133 68446 190134 68478
rect 23528 68310 23534 68342
rect 23054 68278 23055 68310
rect 22989 68277 23055 68278
rect 23533 68278 23534 68310
rect 23598 68310 23604 68342
rect 190128 68414 190134 68446
rect 190198 68446 190199 68478
rect 190198 68414 190204 68446
rect 23598 68278 23599 68310
rect 23533 68277 23599 68278
rect 190128 68206 190204 68414
rect 195024 68342 195100 68550
rect 195024 68278 195030 68342
rect 195094 68278 195100 68342
rect 195024 68272 195100 68278
rect 195568 68550 195574 68582
rect 195638 68582 195639 68614
rect 195840 68614 195916 68620
rect 195638 68550 195644 68582
rect 195568 68342 195644 68550
rect 195568 68278 195574 68342
rect 195638 68278 195644 68342
rect 195840 68550 195846 68614
rect 195910 68550 195916 68614
rect 195840 68342 195916 68550
rect 195840 68310 195846 68342
rect 195568 68272 195644 68278
rect 195845 68278 195846 68310
rect 195910 68310 195916 68342
rect 196656 68342 196732 68348
rect 195910 68278 195911 68310
rect 195845 68277 195911 68278
rect 196656 68278 196662 68342
rect 196726 68278 196732 68342
rect 190128 68142 190134 68206
rect 190198 68142 190204 68206
rect 190128 68136 190204 68142
rect 21760 68006 21766 68070
rect 21830 68006 21836 68070
rect 21760 68000 21836 68006
rect 28424 68070 28500 68076
rect 28424 68006 28430 68070
rect 28494 68006 28500 68070
rect 190133 68070 190199 68071
rect 190133 68038 190134 68070
rect 21901 67934 21967 67935
rect 21901 67902 21902 67934
rect 952 67734 1230 67798
rect 1294 67734 1300 67798
rect 952 66166 1300 67734
rect 21896 67870 21902 67902
rect 21966 67902 21967 67934
rect 22440 67934 22516 67940
rect 21966 67870 21972 67902
rect 21896 67662 21972 67870
rect 21896 67598 21902 67662
rect 21966 67598 21972 67662
rect 22440 67870 22446 67934
rect 22510 67870 22516 67934
rect 22440 67662 22516 67870
rect 28424 67798 28500 68006
rect 28424 67766 28430 67798
rect 28429 67734 28430 67766
rect 28494 67766 28500 67798
rect 190128 68006 190134 68038
rect 190198 68038 190199 68070
rect 196656 68070 196732 68278
rect 196656 68038 196662 68070
rect 190198 68006 190204 68038
rect 190128 67798 190204 68006
rect 196661 68006 196662 68038
rect 196726 68038 196732 68070
rect 196726 68006 196727 68038
rect 196661 68005 196727 68006
rect 28494 67734 28495 67766
rect 28429 67733 28495 67734
rect 190128 67734 190134 67798
rect 190198 67734 190204 67798
rect 190128 67728 190204 67734
rect 196792 67934 196868 67940
rect 196792 67870 196798 67934
rect 196862 67870 196868 67934
rect 22440 67630 22446 67662
rect 21896 67592 21972 67598
rect 22445 67598 22446 67630
rect 22510 67630 22516 67662
rect 28288 67662 28364 67668
rect 22510 67598 22511 67630
rect 22445 67597 22511 67598
rect 28288 67598 28294 67662
rect 28358 67598 28364 67662
rect 196792 67662 196868 67870
rect 196792 67630 196798 67662
rect 21901 67526 21967 67527
rect 21901 67494 21902 67526
rect 21896 67462 21902 67494
rect 21966 67494 21967 67526
rect 21966 67462 21972 67494
rect 21896 67254 21972 67462
rect 28288 67390 28364 67598
rect 196797 67598 196798 67630
rect 196862 67630 196868 67662
rect 217464 67662 217812 69230
rect 196862 67598 196863 67630
rect 196797 67597 196863 67598
rect 217464 67598 217470 67662
rect 217534 67598 217812 67662
rect 28288 67358 28294 67390
rect 28293 67326 28294 67358
rect 28358 67358 28364 67390
rect 196656 67526 196732 67532
rect 196656 67462 196662 67526
rect 196726 67462 196732 67526
rect 28358 67326 28359 67358
rect 28293 67325 28359 67326
rect 21896 67190 21902 67254
rect 21966 67190 21972 67254
rect 196656 67254 196732 67462
rect 196656 67222 196662 67254
rect 21896 67184 21972 67190
rect 196661 67190 196662 67222
rect 196726 67222 196732 67254
rect 196726 67190 196727 67222
rect 196661 67189 196727 67190
rect 21896 67118 21972 67124
rect 21896 67054 21902 67118
rect 21966 67054 21972 67118
rect 22581 67118 22647 67119
rect 22581 67086 22582 67118
rect 21896 66846 21972 67054
rect 21896 66814 21902 66846
rect 21901 66782 21902 66814
rect 21966 66814 21972 66846
rect 22576 67054 22582 67086
rect 22646 67086 22647 67118
rect 23125 67118 23191 67119
rect 23125 67086 23126 67118
rect 22646 67054 22652 67086
rect 22576 66846 22652 67054
rect 21966 66782 21967 66814
rect 21901 66781 21967 66782
rect 22576 66782 22582 66846
rect 22646 66782 22652 66846
rect 22576 66776 22652 66782
rect 23120 67054 23126 67086
rect 23190 67086 23191 67118
rect 23392 67118 23468 67124
rect 23190 67054 23196 67086
rect 23120 66846 23196 67054
rect 23120 66782 23126 66846
rect 23190 66782 23196 66846
rect 23392 67054 23398 67118
rect 23462 67054 23468 67118
rect 23392 66846 23468 67054
rect 195024 67118 195100 67124
rect 195024 67054 195030 67118
rect 195094 67054 195100 67118
rect 23392 66814 23398 66846
rect 23120 66776 23196 66782
rect 23397 66782 23398 66814
rect 23462 66814 23468 66846
rect 28288 66846 28364 66852
rect 23462 66782 23463 66814
rect 23397 66781 23463 66782
rect 28288 66782 28294 66846
rect 28358 66782 28364 66846
rect 21901 66710 21967 66711
rect 21901 66678 21902 66710
rect 21896 66646 21902 66678
rect 21966 66678 21967 66710
rect 22309 66710 22375 66711
rect 22309 66678 22310 66710
rect 21966 66646 21972 66678
rect 21896 66438 21972 66646
rect 21896 66374 21902 66438
rect 21966 66374 21972 66438
rect 21896 66368 21972 66374
rect 22304 66646 22310 66678
rect 22374 66678 22375 66710
rect 22712 66710 22788 66716
rect 22374 66646 22380 66678
rect 22304 66438 22380 66646
rect 22304 66374 22310 66438
rect 22374 66374 22380 66438
rect 22712 66646 22718 66710
rect 22782 66646 22788 66710
rect 22989 66710 23055 66711
rect 22989 66678 22990 66710
rect 22712 66438 22788 66646
rect 22712 66406 22718 66438
rect 22304 66368 22380 66374
rect 22717 66374 22718 66406
rect 22782 66406 22788 66438
rect 22984 66646 22990 66678
rect 23054 66678 23055 66710
rect 23397 66710 23463 66711
rect 23397 66678 23398 66710
rect 23054 66646 23060 66678
rect 22984 66438 23060 66646
rect 22782 66374 22783 66406
rect 22717 66373 22783 66374
rect 22984 66374 22990 66438
rect 23054 66374 23060 66438
rect 22984 66368 23060 66374
rect 23392 66646 23398 66678
rect 23462 66678 23463 66710
rect 23462 66646 23468 66678
rect 23392 66438 23468 66646
rect 28288 66574 28364 66782
rect 28288 66542 28294 66574
rect 28293 66510 28294 66542
rect 28358 66542 28364 66574
rect 190264 66846 190340 66852
rect 190264 66782 190270 66846
rect 190334 66782 190340 66846
rect 195024 66846 195100 67054
rect 195024 66814 195030 66846
rect 190264 66574 190340 66782
rect 195029 66782 195030 66814
rect 195094 66814 195100 66846
rect 195432 67118 195508 67124
rect 195432 67054 195438 67118
rect 195502 67054 195508 67118
rect 195432 66846 195508 67054
rect 195432 66814 195438 66846
rect 195094 66782 195095 66814
rect 195029 66781 195095 66782
rect 195437 66782 195438 66814
rect 195502 66814 195508 66846
rect 196792 67118 196868 67124
rect 196792 67054 196798 67118
rect 196862 67054 196868 67118
rect 196792 66846 196868 67054
rect 196792 66814 196798 66846
rect 195502 66782 195503 66814
rect 195437 66781 195503 66782
rect 196797 66782 196798 66814
rect 196862 66814 196868 66846
rect 196862 66782 196863 66814
rect 196797 66781 196863 66782
rect 195029 66710 195095 66711
rect 195029 66678 195030 66710
rect 190264 66542 190270 66574
rect 28358 66510 28359 66542
rect 28293 66509 28359 66510
rect 190269 66510 190270 66542
rect 190334 66542 190340 66574
rect 195024 66646 195030 66678
rect 195094 66678 195095 66710
rect 195437 66710 195503 66711
rect 195437 66678 195438 66710
rect 195094 66646 195100 66678
rect 190334 66510 190335 66542
rect 190269 66509 190335 66510
rect 23392 66374 23398 66438
rect 23462 66374 23468 66438
rect 23392 66368 23468 66374
rect 195024 66438 195100 66646
rect 195024 66374 195030 66438
rect 195094 66374 195100 66438
rect 195024 66368 195100 66374
rect 195432 66646 195438 66678
rect 195502 66678 195503 66710
rect 196389 66710 196455 66711
rect 196389 66678 196390 66710
rect 195502 66646 195508 66678
rect 195432 66438 195508 66646
rect 195432 66374 195438 66438
rect 195502 66374 195508 66438
rect 195432 66368 195508 66374
rect 196384 66646 196390 66678
rect 196454 66678 196455 66710
rect 196797 66710 196863 66711
rect 196797 66678 196798 66710
rect 196454 66646 196460 66678
rect 196384 66438 196460 66646
rect 196384 66374 196390 66438
rect 196454 66374 196460 66438
rect 196384 66368 196460 66374
rect 196792 66646 196798 66678
rect 196862 66678 196863 66710
rect 196862 66646 196868 66678
rect 196792 66438 196868 66646
rect 196792 66374 196798 66438
rect 196862 66374 196868 66438
rect 196792 66368 196868 66374
rect 952 66102 1230 66166
rect 1294 66102 1300 66166
rect 952 64262 1300 66102
rect 21760 66302 21836 66308
rect 21760 66238 21766 66302
rect 21830 66238 21836 66302
rect 21760 66030 21836 66238
rect 21760 65998 21766 66030
rect 21765 65966 21766 65998
rect 21830 65998 21836 66030
rect 22168 66302 22244 66308
rect 22168 66238 22174 66302
rect 22238 66238 22244 66302
rect 22445 66302 22511 66303
rect 22445 66270 22446 66302
rect 22168 66030 22244 66238
rect 22168 65998 22174 66030
rect 21830 65966 21831 65998
rect 21765 65965 21831 65966
rect 22173 65966 22174 65998
rect 22238 65998 22244 66030
rect 22440 66238 22446 66270
rect 22510 66270 22511 66302
rect 23120 66302 23196 66308
rect 22510 66238 22516 66270
rect 22440 66030 22516 66238
rect 22238 65966 22239 65998
rect 22173 65965 22239 65966
rect 22440 65966 22446 66030
rect 22510 65966 22516 66030
rect 23120 66238 23126 66302
rect 23190 66238 23196 66302
rect 23120 66030 23196 66238
rect 23120 65998 23126 66030
rect 22440 65960 22516 65966
rect 23125 65966 23126 65998
rect 23190 65998 23196 66030
rect 23528 66302 23604 66308
rect 23528 66238 23534 66302
rect 23598 66238 23604 66302
rect 23528 66030 23604 66238
rect 23528 65998 23534 66030
rect 23190 65966 23191 65998
rect 23125 65965 23191 65966
rect 23533 65966 23534 65998
rect 23598 65998 23604 66030
rect 195160 66302 195236 66308
rect 195160 66238 195166 66302
rect 195230 66238 195236 66302
rect 195437 66302 195503 66303
rect 195437 66270 195438 66302
rect 195160 66030 195236 66238
rect 195160 65998 195166 66030
rect 23598 65966 23599 65998
rect 23533 65965 23599 65966
rect 195165 65966 195166 65998
rect 195230 65998 195236 66030
rect 195432 66238 195438 66270
rect 195502 66270 195503 66302
rect 195845 66302 195911 66303
rect 195845 66270 195846 66302
rect 195502 66238 195508 66270
rect 195432 66030 195508 66238
rect 195230 65966 195231 65998
rect 195165 65965 195231 65966
rect 195432 65966 195438 66030
rect 195502 65966 195508 66030
rect 195432 65960 195508 65966
rect 195840 66238 195846 66270
rect 195910 66270 195911 66302
rect 196248 66302 196324 66308
rect 195910 66238 195916 66270
rect 195840 66030 195916 66238
rect 195840 65966 195846 66030
rect 195910 65966 195916 66030
rect 196248 66238 196254 66302
rect 196318 66238 196324 66302
rect 196248 66030 196324 66238
rect 196248 65998 196254 66030
rect 195840 65960 195916 65966
rect 196253 65966 196254 65998
rect 196318 65998 196324 66030
rect 196656 66302 196732 66308
rect 196656 66238 196662 66302
rect 196726 66238 196732 66302
rect 196656 66030 196732 66238
rect 196656 65998 196662 66030
rect 196318 65966 196319 65998
rect 196253 65965 196319 65966
rect 196661 65966 196662 65998
rect 196726 65998 196732 66030
rect 217464 66030 217812 67598
rect 196726 65966 196727 65998
rect 196661 65965 196727 65966
rect 217464 65966 217470 66030
rect 217534 65966 217812 66030
rect 21765 65894 21831 65895
rect 21765 65862 21766 65894
rect 21760 65830 21766 65862
rect 21830 65862 21831 65894
rect 22581 65894 22647 65895
rect 22581 65862 22582 65894
rect 21830 65830 21836 65862
rect 21760 65622 21836 65830
rect 21760 65558 21766 65622
rect 21830 65558 21836 65622
rect 21760 65552 21836 65558
rect 22576 65830 22582 65862
rect 22646 65862 22647 65894
rect 23125 65894 23191 65895
rect 23125 65862 23126 65894
rect 22646 65830 22652 65862
rect 22576 65622 22652 65830
rect 22576 65558 22582 65622
rect 22646 65558 22652 65622
rect 22576 65552 22652 65558
rect 23120 65830 23126 65862
rect 23190 65862 23191 65894
rect 23392 65894 23468 65900
rect 23190 65830 23196 65862
rect 23120 65622 23196 65830
rect 23120 65558 23126 65622
rect 23190 65558 23196 65622
rect 23392 65830 23398 65894
rect 23462 65830 23468 65894
rect 195165 65894 195231 65895
rect 195165 65862 195166 65894
rect 23392 65622 23468 65830
rect 23392 65590 23398 65622
rect 23120 65552 23196 65558
rect 23397 65558 23398 65590
rect 23462 65590 23468 65622
rect 195160 65830 195166 65862
rect 195230 65862 195231 65894
rect 195568 65894 195644 65900
rect 195230 65830 195236 65862
rect 195160 65622 195236 65830
rect 23462 65558 23463 65590
rect 23397 65557 23463 65558
rect 195160 65558 195166 65622
rect 195230 65558 195236 65622
rect 195568 65830 195574 65894
rect 195638 65830 195644 65894
rect 195568 65622 195644 65830
rect 195568 65590 195574 65622
rect 195160 65552 195236 65558
rect 195573 65558 195574 65590
rect 195638 65590 195644 65622
rect 195976 65894 196052 65900
rect 195976 65830 195982 65894
rect 196046 65830 196052 65894
rect 195976 65622 196052 65830
rect 195976 65590 195982 65622
rect 195638 65558 195639 65590
rect 195573 65557 195639 65558
rect 195981 65558 195982 65590
rect 196046 65590 196052 65622
rect 196112 65894 196188 65900
rect 196112 65830 196118 65894
rect 196182 65830 196188 65894
rect 196661 65894 196727 65895
rect 196661 65862 196662 65894
rect 196112 65622 196188 65830
rect 196112 65590 196118 65622
rect 196046 65558 196047 65590
rect 195981 65557 196047 65558
rect 196117 65558 196118 65590
rect 196182 65590 196188 65622
rect 196656 65830 196662 65862
rect 196726 65862 196727 65894
rect 196726 65830 196732 65862
rect 196656 65622 196732 65830
rect 196182 65558 196183 65590
rect 196117 65557 196183 65558
rect 196656 65558 196662 65622
rect 196726 65558 196732 65622
rect 196656 65552 196732 65558
rect 22168 65486 22244 65492
rect 22168 65422 22174 65486
rect 22238 65422 22244 65486
rect 22445 65486 22511 65487
rect 22445 65454 22446 65486
rect 22168 65214 22244 65422
rect 22168 65182 22174 65214
rect 22173 65150 22174 65182
rect 22238 65182 22244 65214
rect 22440 65422 22446 65454
rect 22510 65454 22511 65486
rect 22984 65486 23060 65492
rect 22510 65422 22516 65454
rect 22440 65214 22516 65422
rect 22238 65150 22239 65182
rect 22173 65149 22239 65150
rect 22440 65150 22446 65214
rect 22510 65150 22516 65214
rect 22984 65422 22990 65486
rect 23054 65422 23060 65486
rect 23397 65486 23463 65487
rect 23397 65454 23398 65486
rect 22984 65214 23060 65422
rect 22984 65182 22990 65214
rect 22440 65144 22516 65150
rect 22989 65150 22990 65182
rect 23054 65182 23060 65214
rect 23392 65422 23398 65454
rect 23462 65454 23463 65486
rect 195029 65486 195095 65487
rect 195029 65454 195030 65486
rect 23462 65422 23468 65454
rect 23392 65214 23468 65422
rect 23054 65150 23055 65182
rect 22989 65149 23055 65150
rect 23392 65150 23398 65214
rect 23462 65150 23468 65214
rect 23392 65144 23468 65150
rect 195024 65422 195030 65454
rect 195094 65454 195095 65486
rect 195437 65486 195503 65487
rect 195437 65454 195438 65486
rect 195094 65422 195100 65454
rect 195024 65214 195100 65422
rect 195024 65150 195030 65214
rect 195094 65150 195100 65214
rect 195024 65144 195100 65150
rect 195432 65422 195438 65454
rect 195502 65454 195503 65486
rect 196248 65486 196324 65492
rect 195502 65422 195508 65454
rect 195432 65214 195508 65422
rect 195432 65150 195438 65214
rect 195502 65150 195508 65214
rect 196248 65422 196254 65486
rect 196318 65422 196324 65486
rect 196248 65214 196324 65422
rect 196248 65182 196254 65214
rect 195432 65144 195508 65150
rect 196253 65150 196254 65182
rect 196318 65182 196324 65214
rect 196318 65150 196319 65182
rect 196253 65149 196319 65150
rect 21765 65078 21831 65079
rect 21765 65046 21766 65078
rect 21760 65014 21766 65046
rect 21830 65046 21831 65078
rect 22581 65078 22647 65079
rect 22581 65046 22582 65078
rect 21830 65014 21836 65046
rect 21760 64806 21836 65014
rect 21760 64742 21766 64806
rect 21830 64742 21836 64806
rect 21760 64736 21836 64742
rect 22576 65014 22582 65046
rect 22646 65046 22647 65078
rect 23120 65078 23196 65084
rect 22646 65014 22652 65046
rect 22576 64806 22652 65014
rect 22576 64742 22582 64806
rect 22646 64742 22652 64806
rect 23120 65014 23126 65078
rect 23190 65014 23196 65078
rect 23533 65078 23599 65079
rect 23533 65046 23534 65078
rect 23120 64806 23196 65014
rect 23120 64774 23126 64806
rect 22576 64736 22652 64742
rect 23125 64742 23126 64774
rect 23190 64774 23196 64806
rect 23528 65014 23534 65046
rect 23598 65046 23599 65078
rect 195165 65078 195231 65079
rect 195165 65046 195166 65078
rect 23598 65014 23604 65046
rect 23528 64806 23604 65014
rect 23190 64742 23191 64774
rect 23125 64741 23191 64742
rect 23528 64742 23534 64806
rect 23598 64742 23604 64806
rect 23528 64736 23604 64742
rect 195160 65014 195166 65046
rect 195230 65046 195231 65078
rect 195568 65078 195644 65084
rect 195230 65014 195236 65046
rect 195160 64806 195236 65014
rect 195160 64742 195166 64806
rect 195230 64742 195236 64806
rect 195568 65014 195574 65078
rect 195638 65014 195644 65078
rect 195568 64806 195644 65014
rect 195568 64774 195574 64806
rect 195160 64736 195236 64742
rect 195573 64742 195574 64774
rect 195638 64774 195644 64806
rect 195840 65078 195916 65084
rect 195840 65014 195846 65078
rect 195910 65014 195916 65078
rect 195840 64806 195916 65014
rect 195840 64774 195846 64806
rect 195638 64742 195639 64774
rect 195573 64741 195639 64742
rect 195845 64742 195846 64774
rect 195910 64774 195916 64806
rect 196112 65078 196188 65084
rect 196112 65014 196118 65078
rect 196182 65014 196188 65078
rect 196112 64806 196188 65014
rect 196112 64774 196118 64806
rect 195910 64742 195911 64774
rect 195845 64741 195911 64742
rect 196117 64742 196118 64774
rect 196182 64774 196188 64806
rect 196656 65078 196732 65084
rect 196656 65014 196662 65078
rect 196726 65014 196732 65078
rect 196656 64806 196732 65014
rect 196656 64774 196662 64806
rect 196182 64742 196183 64774
rect 196117 64741 196183 64742
rect 196661 64742 196662 64774
rect 196726 64774 196732 64806
rect 196726 64742 196727 64774
rect 196661 64741 196727 64742
rect 22445 64670 22511 64671
rect 22445 64638 22446 64670
rect 22440 64606 22446 64638
rect 22510 64638 22511 64670
rect 22712 64670 22788 64676
rect 22510 64606 22516 64638
rect 21901 64398 21967 64399
rect 21901 64366 21902 64398
rect 952 64198 1230 64262
rect 1294 64198 1300 64262
rect 952 62630 1300 64198
rect 21896 64334 21902 64366
rect 21966 64366 21967 64398
rect 22440 64398 22516 64606
rect 21966 64334 21972 64366
rect 21896 64126 21972 64334
rect 22440 64334 22446 64398
rect 22510 64334 22516 64398
rect 22712 64606 22718 64670
rect 22782 64606 22788 64670
rect 22712 64398 22788 64606
rect 22712 64366 22718 64398
rect 22440 64328 22516 64334
rect 22717 64334 22718 64366
rect 22782 64366 22788 64398
rect 23120 64670 23196 64676
rect 23120 64606 23126 64670
rect 23190 64606 23196 64670
rect 23120 64398 23196 64606
rect 23120 64366 23126 64398
rect 22782 64334 22783 64366
rect 22717 64333 22783 64334
rect 23125 64334 23126 64366
rect 23190 64366 23196 64398
rect 23392 64670 23468 64676
rect 23392 64606 23398 64670
rect 23462 64606 23468 64670
rect 23392 64398 23468 64606
rect 195024 64670 195100 64676
rect 195024 64606 195030 64670
rect 195094 64606 195100 64670
rect 28565 64534 28631 64535
rect 28565 64502 28566 64534
rect 23392 64366 23398 64398
rect 23190 64334 23191 64366
rect 23125 64333 23191 64334
rect 23397 64334 23398 64366
rect 23462 64366 23468 64398
rect 28560 64470 28566 64502
rect 28630 64502 28631 64534
rect 28630 64470 28636 64502
rect 23462 64334 23463 64366
rect 23397 64333 23463 64334
rect 23125 64262 23191 64263
rect 23125 64230 23126 64262
rect 21896 64062 21902 64126
rect 21966 64062 21972 64126
rect 21896 64056 21972 64062
rect 23120 64198 23126 64230
rect 23190 64230 23191 64262
rect 23397 64262 23463 64263
rect 23397 64230 23398 64262
rect 23190 64198 23196 64230
rect 23120 63990 23196 64198
rect 23120 63926 23126 63990
rect 23190 63926 23196 63990
rect 23120 63920 23196 63926
rect 23392 64198 23398 64230
rect 23462 64230 23463 64262
rect 28560 64262 28636 64470
rect 195024 64398 195100 64606
rect 195024 64366 195030 64398
rect 195029 64334 195030 64366
rect 195094 64366 195100 64398
rect 195568 64670 195644 64676
rect 195568 64606 195574 64670
rect 195638 64606 195644 64670
rect 195568 64398 195644 64606
rect 195568 64366 195574 64398
rect 195094 64334 195095 64366
rect 195029 64333 195095 64334
rect 195573 64334 195574 64366
rect 195638 64366 195644 64398
rect 195976 64670 196052 64676
rect 195976 64606 195982 64670
rect 196046 64606 196052 64670
rect 195976 64398 196052 64606
rect 195976 64366 195982 64398
rect 195638 64334 195639 64366
rect 195573 64333 195639 64334
rect 195981 64334 195982 64366
rect 196046 64366 196052 64398
rect 196792 64398 196868 64404
rect 196046 64334 196047 64366
rect 195981 64333 196047 64334
rect 196792 64334 196798 64398
rect 196862 64334 196868 64398
rect 23462 64198 23468 64230
rect 23392 63990 23468 64198
rect 28560 64198 28566 64262
rect 28630 64198 28636 64262
rect 28560 64192 28636 64198
rect 195160 64262 195236 64268
rect 195160 64198 195166 64262
rect 195230 64198 195236 64262
rect 195573 64262 195639 64263
rect 195573 64230 195574 64262
rect 23392 63926 23398 63990
rect 23462 63926 23468 63990
rect 195160 63990 195236 64198
rect 195160 63958 195166 63990
rect 23392 63920 23468 63926
rect 195165 63926 195166 63958
rect 195230 63958 195236 63990
rect 195568 64198 195574 64230
rect 195638 64230 195639 64262
rect 195638 64198 195644 64230
rect 195568 63990 195644 64198
rect 196792 64126 196868 64334
rect 196792 64094 196798 64126
rect 196797 64062 196798 64094
rect 196862 64094 196868 64126
rect 217464 64398 217812 65966
rect 217464 64334 217470 64398
rect 217534 64334 217812 64398
rect 196862 64062 196863 64094
rect 196797 64061 196863 64062
rect 195230 63926 195231 63958
rect 195165 63925 195231 63926
rect 195568 63926 195574 63990
rect 195638 63926 195644 63990
rect 195568 63920 195644 63926
rect 22712 63854 22788 63860
rect 22712 63790 22718 63854
rect 22782 63790 22788 63854
rect 21896 63582 21972 63588
rect 21896 63518 21902 63582
rect 21966 63518 21972 63582
rect 22712 63582 22788 63790
rect 195976 63854 196052 63860
rect 195976 63790 195982 63854
rect 196046 63790 196052 63854
rect 22712 63550 22718 63582
rect 21896 63310 21972 63518
rect 22717 63518 22718 63550
rect 22782 63550 22788 63582
rect 28424 63718 28500 63724
rect 28424 63654 28430 63718
rect 28494 63654 28500 63718
rect 190133 63718 190199 63719
rect 190133 63686 190134 63718
rect 22782 63518 22783 63550
rect 22717 63517 22783 63518
rect 21896 63278 21902 63310
rect 21901 63246 21902 63278
rect 21966 63278 21972 63310
rect 28288 63446 28364 63452
rect 28288 63382 28294 63446
rect 28358 63382 28364 63446
rect 28424 63446 28500 63654
rect 28424 63414 28430 63446
rect 21966 63246 21967 63278
rect 21901 63245 21967 63246
rect 21901 63174 21967 63175
rect 21901 63142 21902 63174
rect 21896 63110 21902 63142
rect 21966 63142 21967 63174
rect 22309 63174 22375 63175
rect 22309 63142 22310 63174
rect 21966 63110 21972 63142
rect 21896 62902 21972 63110
rect 21896 62838 21902 62902
rect 21966 62838 21972 62902
rect 21896 62832 21972 62838
rect 22304 63110 22310 63142
rect 22374 63142 22375 63174
rect 22445 63174 22511 63175
rect 22445 63142 22446 63174
rect 22374 63110 22380 63142
rect 22304 62902 22380 63110
rect 22304 62838 22310 62902
rect 22374 62838 22380 62902
rect 22304 62832 22380 62838
rect 22440 63110 22446 63142
rect 22510 63142 22511 63174
rect 22510 63110 22516 63142
rect 22440 62902 22516 63110
rect 28288 63038 28364 63382
rect 28429 63382 28430 63414
rect 28494 63414 28500 63446
rect 190128 63654 190134 63686
rect 190198 63686 190199 63718
rect 190198 63654 190204 63686
rect 190128 63446 190204 63654
rect 195976 63582 196052 63790
rect 195976 63550 195982 63582
rect 195981 63518 195982 63550
rect 196046 63550 196052 63582
rect 196797 63582 196863 63583
rect 196797 63550 196798 63582
rect 196046 63518 196047 63550
rect 195981 63517 196047 63518
rect 196792 63518 196798 63550
rect 196862 63550 196863 63582
rect 196862 63518 196868 63550
rect 28494 63382 28495 63414
rect 28429 63381 28495 63382
rect 190128 63382 190134 63446
rect 190198 63382 190204 63446
rect 190128 63376 190204 63382
rect 28288 63006 28294 63038
rect 28293 62974 28294 63006
rect 28358 63006 28364 63038
rect 190128 63310 190204 63316
rect 190128 63246 190134 63310
rect 190198 63246 190204 63310
rect 190128 63038 190204 63246
rect 196792 63310 196868 63518
rect 196792 63246 196798 63310
rect 196862 63246 196868 63310
rect 196792 63240 196868 63246
rect 196117 63174 196183 63175
rect 196117 63142 196118 63174
rect 190128 63006 190134 63038
rect 28358 62974 28359 63006
rect 28293 62973 28359 62974
rect 190133 62974 190134 63006
rect 190198 63006 190204 63038
rect 196112 63110 196118 63142
rect 196182 63142 196183 63174
rect 196656 63174 196732 63180
rect 196182 63110 196188 63142
rect 190198 62974 190199 63006
rect 190133 62973 190199 62974
rect 22440 62838 22446 62902
rect 22510 62838 22516 62902
rect 190133 62902 190199 62903
rect 190133 62870 190134 62902
rect 22440 62832 22516 62838
rect 190128 62838 190134 62870
rect 190198 62870 190199 62902
rect 196112 62902 196188 63110
rect 190198 62838 190204 62870
rect 21765 62766 21831 62767
rect 21765 62734 21766 62766
rect 952 62566 1230 62630
rect 1294 62566 1300 62630
rect 952 60998 1300 62566
rect 21760 62702 21766 62734
rect 21830 62734 21831 62766
rect 22984 62766 23060 62772
rect 21830 62702 21836 62734
rect 21760 62494 21836 62702
rect 21760 62430 21766 62494
rect 21830 62430 21836 62494
rect 22984 62702 22990 62766
rect 23054 62702 23060 62766
rect 22984 62494 23060 62702
rect 22984 62462 22990 62494
rect 21760 62424 21836 62430
rect 22989 62430 22990 62462
rect 23054 62462 23060 62494
rect 23392 62766 23468 62772
rect 23392 62702 23398 62766
rect 23462 62702 23468 62766
rect 23392 62494 23468 62702
rect 190128 62630 190204 62838
rect 196112 62838 196118 62902
rect 196182 62838 196188 62902
rect 196656 63110 196662 63174
rect 196726 63110 196732 63174
rect 196656 62902 196732 63110
rect 196656 62870 196662 62902
rect 196112 62832 196188 62838
rect 196661 62838 196662 62870
rect 196726 62870 196732 62902
rect 196726 62838 196727 62870
rect 196661 62837 196727 62838
rect 190128 62566 190134 62630
rect 190198 62566 190204 62630
rect 190128 62560 190204 62566
rect 195024 62766 195100 62772
rect 195024 62702 195030 62766
rect 195094 62702 195100 62766
rect 23392 62462 23398 62494
rect 23054 62430 23055 62462
rect 22989 62429 23055 62430
rect 23397 62430 23398 62462
rect 23462 62462 23468 62494
rect 195024 62494 195100 62702
rect 195024 62462 195030 62494
rect 23462 62430 23463 62462
rect 23397 62429 23463 62430
rect 195029 62430 195030 62462
rect 195094 62462 195100 62494
rect 195432 62766 195508 62772
rect 195432 62702 195438 62766
rect 195502 62702 195508 62766
rect 195432 62494 195508 62702
rect 195432 62462 195438 62494
rect 195094 62430 195095 62462
rect 195029 62429 195095 62430
rect 195437 62430 195438 62462
rect 195502 62462 195508 62494
rect 196792 62766 196868 62772
rect 196792 62702 196798 62766
rect 196862 62702 196868 62766
rect 196792 62494 196868 62702
rect 196792 62462 196798 62494
rect 195502 62430 195503 62462
rect 195437 62429 195503 62430
rect 196797 62430 196798 62462
rect 196862 62462 196868 62494
rect 217464 62766 217812 64334
rect 217464 62702 217470 62766
rect 217534 62702 217812 62766
rect 196862 62430 196863 62462
rect 196797 62429 196863 62430
rect 21901 62358 21967 62359
rect 21901 62326 21902 62358
rect 21896 62294 21902 62326
rect 21966 62326 21967 62358
rect 22712 62358 22788 62364
rect 21966 62294 21972 62326
rect 21896 62086 21972 62294
rect 21896 62022 21902 62086
rect 21966 62022 21972 62086
rect 22712 62294 22718 62358
rect 22782 62294 22788 62358
rect 22712 62086 22788 62294
rect 22712 62054 22718 62086
rect 21896 62016 21972 62022
rect 22717 62022 22718 62054
rect 22782 62054 22788 62086
rect 23120 62358 23196 62364
rect 23120 62294 23126 62358
rect 23190 62294 23196 62358
rect 23397 62358 23463 62359
rect 23397 62326 23398 62358
rect 23120 62086 23196 62294
rect 23120 62054 23126 62086
rect 22782 62022 22783 62054
rect 22717 62021 22783 62022
rect 23125 62022 23126 62054
rect 23190 62054 23196 62086
rect 23392 62294 23398 62326
rect 23462 62326 23463 62358
rect 195024 62358 195100 62364
rect 23462 62294 23468 62326
rect 23392 62086 23468 62294
rect 23190 62022 23191 62054
rect 23125 62021 23191 62022
rect 23392 62022 23398 62086
rect 23462 62022 23468 62086
rect 195024 62294 195030 62358
rect 195094 62294 195100 62358
rect 195437 62358 195503 62359
rect 195437 62326 195438 62358
rect 195024 62086 195100 62294
rect 195024 62054 195030 62086
rect 23392 62016 23468 62022
rect 195029 62022 195030 62054
rect 195094 62054 195100 62086
rect 195432 62294 195438 62326
rect 195502 62326 195503 62358
rect 195976 62358 196052 62364
rect 195502 62294 195508 62326
rect 195432 62086 195508 62294
rect 195094 62022 195095 62054
rect 195029 62021 195095 62022
rect 195432 62022 195438 62086
rect 195502 62022 195508 62086
rect 195976 62294 195982 62358
rect 196046 62294 196052 62358
rect 196797 62358 196863 62359
rect 196797 62326 196798 62358
rect 195976 62086 196052 62294
rect 195976 62054 195982 62086
rect 195432 62016 195508 62022
rect 195981 62022 195982 62054
rect 196046 62054 196052 62086
rect 196792 62294 196798 62326
rect 196862 62326 196863 62358
rect 196862 62294 196868 62326
rect 196792 62086 196868 62294
rect 196046 62022 196047 62054
rect 195981 62021 196047 62022
rect 196792 62022 196798 62086
rect 196862 62022 196868 62086
rect 196792 62016 196868 62022
rect 21760 61950 21836 61956
rect 21760 61886 21766 61950
rect 21830 61886 21836 61950
rect 21760 61678 21836 61886
rect 21760 61646 21766 61678
rect 21765 61614 21766 61646
rect 21830 61646 21836 61678
rect 22168 61950 22244 61956
rect 22168 61886 22174 61950
rect 22238 61886 22244 61950
rect 22581 61950 22647 61951
rect 22581 61918 22582 61950
rect 22168 61678 22244 61886
rect 22168 61646 22174 61678
rect 21830 61614 21831 61646
rect 21765 61613 21831 61614
rect 22173 61614 22174 61646
rect 22238 61646 22244 61678
rect 22576 61886 22582 61918
rect 22646 61918 22647 61950
rect 22989 61950 23055 61951
rect 22989 61918 22990 61950
rect 22646 61886 22652 61918
rect 22576 61678 22652 61886
rect 22238 61614 22239 61646
rect 22173 61613 22239 61614
rect 22576 61614 22582 61678
rect 22646 61614 22652 61678
rect 22576 61608 22652 61614
rect 22984 61886 22990 61918
rect 23054 61918 23055 61950
rect 23528 61950 23604 61956
rect 23054 61886 23060 61918
rect 22984 61678 23060 61886
rect 22984 61614 22990 61678
rect 23054 61614 23060 61678
rect 23528 61886 23534 61950
rect 23598 61886 23604 61950
rect 195165 61950 195231 61951
rect 195165 61918 195166 61950
rect 23528 61678 23604 61886
rect 23528 61646 23534 61678
rect 22984 61608 23060 61614
rect 23533 61614 23534 61646
rect 23598 61646 23604 61678
rect 195160 61886 195166 61918
rect 195230 61918 195231 61950
rect 195568 61950 195644 61956
rect 195230 61886 195236 61918
rect 195160 61678 195236 61886
rect 23598 61614 23599 61646
rect 23533 61613 23599 61614
rect 195160 61614 195166 61678
rect 195230 61614 195236 61678
rect 195568 61886 195574 61950
rect 195638 61886 195644 61950
rect 196117 61950 196183 61951
rect 196117 61918 196118 61950
rect 195568 61678 195644 61886
rect 195568 61646 195574 61678
rect 195160 61608 195236 61614
rect 195573 61614 195574 61646
rect 195638 61646 195644 61678
rect 196112 61886 196118 61918
rect 196182 61918 196183 61950
rect 196253 61950 196319 61951
rect 196253 61918 196254 61950
rect 196182 61886 196188 61918
rect 196112 61678 196188 61886
rect 195638 61614 195639 61646
rect 195573 61613 195639 61614
rect 196112 61614 196118 61678
rect 196182 61614 196188 61678
rect 196112 61608 196188 61614
rect 196248 61886 196254 61918
rect 196318 61918 196319 61950
rect 196661 61950 196727 61951
rect 196661 61918 196662 61950
rect 196318 61886 196324 61918
rect 196248 61678 196324 61886
rect 196248 61614 196254 61678
rect 196318 61614 196324 61678
rect 196248 61608 196324 61614
rect 196656 61886 196662 61918
rect 196726 61918 196727 61950
rect 196726 61886 196732 61918
rect 196656 61678 196732 61886
rect 196656 61614 196662 61678
rect 196726 61614 196732 61678
rect 196656 61608 196732 61614
rect 21896 61542 21972 61548
rect 21896 61478 21902 61542
rect 21966 61478 21972 61542
rect 23125 61542 23191 61543
rect 23125 61510 23126 61542
rect 21896 61270 21972 61478
rect 21896 61238 21902 61270
rect 21901 61206 21902 61238
rect 21966 61238 21972 61270
rect 23120 61478 23126 61510
rect 23190 61510 23191 61542
rect 23533 61542 23599 61543
rect 23533 61510 23534 61542
rect 23190 61478 23196 61510
rect 23120 61270 23196 61478
rect 21966 61206 21967 61238
rect 21901 61205 21967 61206
rect 23120 61206 23126 61270
rect 23190 61206 23196 61270
rect 23120 61200 23196 61206
rect 23528 61478 23534 61510
rect 23598 61510 23599 61542
rect 195165 61542 195231 61543
rect 195165 61510 195166 61542
rect 23598 61478 23604 61510
rect 23528 61270 23604 61478
rect 23528 61206 23534 61270
rect 23598 61206 23604 61270
rect 23528 61200 23604 61206
rect 195160 61478 195166 61510
rect 195230 61510 195231 61542
rect 195573 61542 195639 61543
rect 195573 61510 195574 61542
rect 195230 61478 195236 61510
rect 195160 61270 195236 61478
rect 195160 61206 195166 61270
rect 195230 61206 195236 61270
rect 195160 61200 195236 61206
rect 195568 61478 195574 61510
rect 195638 61510 195639 61542
rect 195976 61542 196052 61548
rect 195638 61478 195644 61510
rect 195568 61270 195644 61478
rect 195568 61206 195574 61270
rect 195638 61206 195644 61270
rect 195976 61478 195982 61542
rect 196046 61478 196052 61542
rect 196661 61542 196727 61543
rect 196661 61510 196662 61542
rect 195976 61270 196052 61478
rect 195976 61238 195982 61270
rect 195568 61200 195644 61206
rect 195981 61206 195982 61238
rect 196046 61238 196052 61270
rect 196656 61478 196662 61510
rect 196726 61510 196727 61542
rect 196726 61478 196732 61510
rect 196656 61270 196732 61478
rect 196046 61206 196047 61238
rect 195981 61205 196047 61206
rect 196656 61206 196662 61270
rect 196726 61206 196732 61270
rect 196656 61200 196732 61206
rect 21901 61134 21967 61135
rect 21901 61102 21902 61134
rect 952 60934 1230 60998
rect 1294 60934 1300 60998
rect 952 59230 1300 60934
rect 21896 61070 21902 61102
rect 21966 61102 21967 61134
rect 22168 61134 22244 61140
rect 21966 61070 21972 61102
rect 21896 60862 21972 61070
rect 21896 60798 21902 60862
rect 21966 60798 21972 60862
rect 22168 61070 22174 61134
rect 22238 61070 22244 61134
rect 22717 61134 22783 61135
rect 22717 61102 22718 61134
rect 22168 60862 22244 61070
rect 22168 60830 22174 60862
rect 21896 60792 21972 60798
rect 22173 60798 22174 60830
rect 22238 60830 22244 60862
rect 22712 61070 22718 61102
rect 22782 61102 22783 61134
rect 22984 61134 23060 61140
rect 22782 61070 22788 61102
rect 22712 60862 22788 61070
rect 22238 60798 22239 60830
rect 22173 60797 22239 60798
rect 22712 60798 22718 60862
rect 22782 60798 22788 60862
rect 22984 61070 22990 61134
rect 23054 61070 23060 61134
rect 22984 60862 23060 61070
rect 22984 60830 22990 60862
rect 22712 60792 22788 60798
rect 22989 60798 22990 60830
rect 23054 60830 23060 60862
rect 23528 61134 23604 61140
rect 23528 61070 23534 61134
rect 23598 61070 23604 61134
rect 195029 61134 195095 61135
rect 195029 61102 195030 61134
rect 23528 60862 23604 61070
rect 23528 60830 23534 60862
rect 23054 60798 23055 60830
rect 22989 60797 23055 60798
rect 23533 60798 23534 60830
rect 23598 60830 23604 60862
rect 195024 61070 195030 61102
rect 195094 61102 195095 61134
rect 195432 61134 195508 61140
rect 195094 61070 195100 61102
rect 195024 60862 195100 61070
rect 23598 60798 23599 60830
rect 23533 60797 23599 60798
rect 195024 60798 195030 60862
rect 195094 60798 195100 60862
rect 195432 61070 195438 61134
rect 195502 61070 195508 61134
rect 196117 61134 196183 61135
rect 196117 61102 196118 61134
rect 195432 60862 195508 61070
rect 195432 60830 195438 60862
rect 195024 60792 195100 60798
rect 195437 60798 195438 60830
rect 195502 60830 195508 60862
rect 196112 61070 196118 61102
rect 196182 61102 196183 61134
rect 196656 61134 196732 61140
rect 196182 61070 196188 61102
rect 196112 60862 196188 61070
rect 195502 60798 195503 60830
rect 195437 60797 195503 60798
rect 196112 60798 196118 60862
rect 196182 60798 196188 60862
rect 196656 61070 196662 61134
rect 196726 61070 196732 61134
rect 196656 60862 196732 61070
rect 196656 60830 196662 60862
rect 196112 60792 196188 60798
rect 196661 60798 196662 60830
rect 196726 60830 196732 60862
rect 217464 61134 217812 62702
rect 217464 61070 217470 61134
rect 217534 61070 217812 61134
rect 196726 60798 196727 60830
rect 196661 60797 196727 60798
rect 22576 60726 22652 60732
rect 22576 60662 22582 60726
rect 22646 60662 22652 60726
rect 22989 60726 23055 60727
rect 22989 60694 22990 60726
rect 22576 60454 22652 60662
rect 22576 60422 22582 60454
rect 22581 60390 22582 60422
rect 22646 60422 22652 60454
rect 22984 60662 22990 60694
rect 23054 60694 23055 60726
rect 23533 60726 23599 60727
rect 23533 60694 23534 60726
rect 23054 60662 23060 60694
rect 22984 60454 23060 60662
rect 22646 60390 22647 60422
rect 22581 60389 22647 60390
rect 22984 60390 22990 60454
rect 23054 60390 23060 60454
rect 22984 60384 23060 60390
rect 23528 60662 23534 60694
rect 23598 60694 23599 60726
rect 195165 60726 195231 60727
rect 195165 60694 195166 60726
rect 23598 60662 23604 60694
rect 23528 60454 23604 60662
rect 23528 60390 23534 60454
rect 23598 60390 23604 60454
rect 23528 60384 23604 60390
rect 195160 60662 195166 60694
rect 195230 60694 195231 60726
rect 195437 60726 195503 60727
rect 195437 60694 195438 60726
rect 195230 60662 195236 60694
rect 195160 60454 195236 60662
rect 195160 60390 195166 60454
rect 195230 60390 195236 60454
rect 195160 60384 195236 60390
rect 195432 60662 195438 60694
rect 195502 60694 195503 60726
rect 195845 60726 195911 60727
rect 195845 60694 195846 60726
rect 195502 60662 195508 60694
rect 195432 60454 195508 60662
rect 195432 60390 195438 60454
rect 195502 60390 195508 60454
rect 195432 60384 195508 60390
rect 195840 60662 195846 60694
rect 195910 60694 195911 60726
rect 196248 60726 196324 60732
rect 195910 60662 195916 60694
rect 195840 60454 195916 60662
rect 195840 60390 195846 60454
rect 195910 60390 195916 60454
rect 196248 60662 196254 60726
rect 196318 60662 196324 60726
rect 196248 60454 196324 60662
rect 196248 60422 196254 60454
rect 195840 60384 195916 60390
rect 196253 60390 196254 60422
rect 196318 60422 196324 60454
rect 196318 60390 196319 60422
rect 196253 60389 196319 60390
rect 23120 60318 23196 60324
rect 23120 60254 23126 60318
rect 23190 60254 23196 60318
rect 23397 60318 23463 60319
rect 23397 60286 23398 60318
rect 23120 60046 23196 60254
rect 23120 60014 23126 60046
rect 23125 59982 23126 60014
rect 23190 60014 23196 60046
rect 23392 60254 23398 60286
rect 23462 60286 23463 60318
rect 28293 60318 28359 60319
rect 28293 60286 28294 60318
rect 23462 60254 23468 60286
rect 23392 60046 23468 60254
rect 23190 59982 23191 60014
rect 23125 59981 23191 59982
rect 23392 59982 23398 60046
rect 23462 59982 23468 60046
rect 23392 59976 23468 59982
rect 28288 60254 28294 60286
rect 28358 60286 28359 60318
rect 195024 60318 195100 60324
rect 28358 60254 28364 60286
rect 22581 59910 22647 59911
rect 22581 59878 22582 59910
rect 22576 59846 22582 59878
rect 22646 59878 22647 59910
rect 28288 59910 28364 60254
rect 195024 60254 195030 60318
rect 195094 60254 195100 60318
rect 195437 60318 195503 60319
rect 195437 60286 195438 60318
rect 195024 60046 195100 60254
rect 195024 60014 195030 60046
rect 195029 59982 195030 60014
rect 195094 60014 195100 60046
rect 195432 60254 195438 60286
rect 195502 60286 195503 60318
rect 195502 60254 195508 60286
rect 195432 60046 195508 60254
rect 195094 59982 195095 60014
rect 195029 59981 195095 59982
rect 195432 59982 195438 60046
rect 195502 59982 195508 60046
rect 195432 59976 195508 59982
rect 22646 59846 22652 59878
rect 21765 59638 21831 59639
rect 21765 59606 21766 59638
rect 21760 59574 21766 59606
rect 21830 59606 21831 59638
rect 22576 59638 22652 59846
rect 28288 59846 28294 59910
rect 28358 59846 28364 59910
rect 28288 59840 28364 59846
rect 21830 59574 21836 59606
rect 21760 59366 21836 59574
rect 22576 59574 22582 59638
rect 22646 59574 22652 59638
rect 22576 59568 22652 59574
rect 196656 59638 196732 59644
rect 196656 59574 196662 59638
rect 196726 59574 196732 59638
rect 21760 59302 21766 59366
rect 21830 59302 21836 59366
rect 28565 59366 28631 59367
rect 28565 59334 28566 59366
rect 21760 59296 21836 59302
rect 28560 59302 28566 59334
rect 28630 59334 28631 59366
rect 190264 59366 190340 59372
rect 28630 59302 28636 59334
rect 952 59166 1230 59230
rect 1294 59166 1300 59230
rect 952 57734 1300 59166
rect 21896 59230 21972 59236
rect 21896 59166 21902 59230
rect 21966 59166 21972 59230
rect 21896 58958 21972 59166
rect 21896 58926 21902 58958
rect 21901 58894 21902 58926
rect 21966 58926 21972 58958
rect 22576 59230 22652 59236
rect 22576 59166 22582 59230
rect 22646 59166 22652 59230
rect 22576 58958 22652 59166
rect 28560 59094 28636 59302
rect 28560 59030 28566 59094
rect 28630 59030 28636 59094
rect 190264 59302 190270 59366
rect 190334 59302 190340 59366
rect 196656 59366 196732 59574
rect 196656 59334 196662 59366
rect 190264 59094 190340 59302
rect 196661 59302 196662 59334
rect 196726 59334 196732 59366
rect 217464 59366 217812 61070
rect 196726 59302 196727 59334
rect 196661 59301 196727 59302
rect 217464 59302 217470 59366
rect 217534 59302 217812 59366
rect 195981 59230 196047 59231
rect 195981 59198 195982 59230
rect 190264 59062 190270 59094
rect 28560 59024 28636 59030
rect 190269 59030 190270 59062
rect 190334 59062 190340 59094
rect 195976 59166 195982 59198
rect 196046 59198 196047 59230
rect 196792 59230 196868 59236
rect 196046 59166 196052 59198
rect 190334 59030 190335 59062
rect 190269 59029 190335 59030
rect 22576 58926 22582 58958
rect 21966 58894 21967 58926
rect 21901 58893 21967 58894
rect 22581 58894 22582 58926
rect 22646 58926 22652 58958
rect 28565 58958 28631 58959
rect 28565 58926 28566 58958
rect 22646 58894 22647 58926
rect 22581 58893 22647 58894
rect 28560 58894 28566 58926
rect 28630 58926 28631 58958
rect 190128 58958 190204 58964
rect 28630 58894 28636 58926
rect 21760 58822 21836 58828
rect 21760 58758 21766 58822
rect 21830 58758 21836 58822
rect 21760 58550 21836 58758
rect 21760 58518 21766 58550
rect 21765 58486 21766 58518
rect 21830 58518 21836 58550
rect 22984 58822 23060 58828
rect 22984 58758 22990 58822
rect 23054 58758 23060 58822
rect 22984 58550 23060 58758
rect 22984 58518 22990 58550
rect 21830 58486 21831 58518
rect 21765 58485 21831 58486
rect 22989 58486 22990 58518
rect 23054 58518 23060 58550
rect 23528 58822 23604 58828
rect 23528 58758 23534 58822
rect 23598 58758 23604 58822
rect 23528 58550 23604 58758
rect 28560 58686 28636 58894
rect 28560 58622 28566 58686
rect 28630 58622 28636 58686
rect 190128 58894 190134 58958
rect 190198 58894 190204 58958
rect 190128 58686 190204 58894
rect 195976 58958 196052 59166
rect 195976 58894 195982 58958
rect 196046 58894 196052 58958
rect 196792 59166 196798 59230
rect 196862 59166 196868 59230
rect 196792 58958 196868 59166
rect 196792 58926 196798 58958
rect 195976 58888 196052 58894
rect 196797 58894 196798 58926
rect 196862 58926 196868 58958
rect 196862 58894 196863 58926
rect 196797 58893 196863 58894
rect 190128 58654 190134 58686
rect 28560 58616 28636 58622
rect 190133 58622 190134 58654
rect 190198 58654 190204 58686
rect 195160 58822 195236 58828
rect 195160 58758 195166 58822
rect 195230 58758 195236 58822
rect 190198 58622 190199 58654
rect 190133 58621 190199 58622
rect 23528 58518 23534 58550
rect 23054 58486 23055 58518
rect 22989 58485 23055 58486
rect 23533 58486 23534 58518
rect 23598 58518 23604 58550
rect 195160 58550 195236 58758
rect 195160 58518 195166 58550
rect 23598 58486 23599 58518
rect 23533 58485 23599 58486
rect 195165 58486 195166 58518
rect 195230 58518 195236 58550
rect 195432 58822 195508 58828
rect 195432 58758 195438 58822
rect 195502 58758 195508 58822
rect 196797 58822 196863 58823
rect 196797 58790 196798 58822
rect 195432 58550 195508 58758
rect 195432 58518 195438 58550
rect 195230 58486 195231 58518
rect 195165 58485 195231 58486
rect 195437 58486 195438 58518
rect 195502 58518 195508 58550
rect 196792 58758 196798 58790
rect 196862 58790 196863 58822
rect 196862 58758 196868 58790
rect 196792 58550 196868 58758
rect 195502 58486 195503 58518
rect 195437 58485 195503 58486
rect 196792 58486 196798 58550
rect 196862 58486 196868 58550
rect 196792 58480 196868 58486
rect 21896 58414 21972 58420
rect 21896 58350 21902 58414
rect 21966 58350 21972 58414
rect 22581 58414 22647 58415
rect 22581 58382 22582 58414
rect 21896 58142 21972 58350
rect 21896 58110 21902 58142
rect 21901 58078 21902 58110
rect 21966 58110 21972 58142
rect 22576 58350 22582 58382
rect 22646 58382 22647 58414
rect 22989 58414 23055 58415
rect 22989 58382 22990 58414
rect 22646 58350 22652 58382
rect 22576 58142 22652 58350
rect 21966 58078 21967 58110
rect 21901 58077 21967 58078
rect 22576 58078 22582 58142
rect 22646 58078 22652 58142
rect 22576 58072 22652 58078
rect 22984 58350 22990 58382
rect 23054 58382 23055 58414
rect 23533 58414 23599 58415
rect 23533 58382 23534 58414
rect 23054 58350 23060 58382
rect 22984 58142 23060 58350
rect 22984 58078 22990 58142
rect 23054 58078 23060 58142
rect 22984 58072 23060 58078
rect 23528 58350 23534 58382
rect 23598 58382 23599 58414
rect 195024 58414 195100 58420
rect 23598 58350 23604 58382
rect 23528 58142 23604 58350
rect 195024 58350 195030 58414
rect 195094 58350 195100 58414
rect 195437 58414 195503 58415
rect 195437 58382 195438 58414
rect 23528 58078 23534 58142
rect 23598 58078 23604 58142
rect 28429 58142 28495 58143
rect 28429 58110 28430 58142
rect 23528 58072 23604 58078
rect 28424 58078 28430 58110
rect 28494 58110 28495 58142
rect 195024 58142 195100 58350
rect 195024 58110 195030 58142
rect 28494 58078 28500 58110
rect 21901 58006 21967 58007
rect 21901 57974 21902 58006
rect 952 57670 1230 57734
rect 1294 57670 1300 57734
rect 952 55966 1300 57670
rect 21896 57942 21902 57974
rect 21966 57974 21967 58006
rect 22989 58006 23055 58007
rect 22989 57974 22990 58006
rect 21966 57942 21972 57974
rect 21896 57734 21972 57942
rect 21896 57670 21902 57734
rect 21966 57670 21972 57734
rect 21896 57664 21972 57670
rect 22984 57942 22990 57974
rect 23054 57974 23055 58006
rect 23392 58006 23468 58012
rect 23054 57942 23060 57974
rect 22984 57734 23060 57942
rect 22984 57670 22990 57734
rect 23054 57670 23060 57734
rect 23392 57942 23398 58006
rect 23462 57942 23468 58006
rect 23392 57734 23468 57942
rect 28424 57870 28500 58078
rect 195029 58078 195030 58110
rect 195094 58110 195100 58142
rect 195432 58350 195438 58382
rect 195502 58382 195503 58414
rect 195976 58414 196052 58420
rect 195502 58350 195508 58382
rect 195432 58142 195508 58350
rect 195094 58078 195095 58110
rect 195029 58077 195095 58078
rect 195432 58078 195438 58142
rect 195502 58078 195508 58142
rect 195976 58350 195982 58414
rect 196046 58350 196052 58414
rect 195976 58142 196052 58350
rect 195976 58110 195982 58142
rect 195432 58072 195508 58078
rect 195981 58078 195982 58110
rect 196046 58110 196052 58142
rect 196112 58414 196188 58420
rect 196112 58350 196118 58414
rect 196182 58350 196188 58414
rect 196661 58414 196727 58415
rect 196661 58382 196662 58414
rect 196112 58142 196188 58350
rect 196112 58110 196118 58142
rect 196046 58078 196047 58110
rect 195981 58077 196047 58078
rect 196117 58078 196118 58110
rect 196182 58110 196188 58142
rect 196656 58350 196662 58382
rect 196726 58382 196727 58414
rect 196726 58350 196732 58382
rect 196656 58142 196732 58350
rect 196182 58078 196183 58110
rect 196117 58077 196183 58078
rect 196656 58078 196662 58142
rect 196726 58078 196732 58142
rect 196656 58072 196732 58078
rect 195029 58006 195095 58007
rect 195029 57974 195030 58006
rect 28424 57806 28430 57870
rect 28494 57806 28500 57870
rect 28424 57800 28500 57806
rect 195024 57942 195030 57974
rect 195094 57974 195095 58006
rect 195568 58006 195644 58012
rect 195094 57942 195100 57974
rect 23392 57702 23398 57734
rect 22984 57664 23060 57670
rect 23397 57670 23398 57702
rect 23462 57702 23468 57734
rect 195024 57734 195100 57942
rect 23462 57670 23463 57702
rect 23397 57669 23463 57670
rect 195024 57670 195030 57734
rect 195094 57670 195100 57734
rect 195568 57942 195574 58006
rect 195638 57942 195644 58006
rect 196389 58006 196455 58007
rect 196389 57974 196390 58006
rect 195568 57734 195644 57942
rect 195568 57702 195574 57734
rect 195024 57664 195100 57670
rect 195573 57670 195574 57702
rect 195638 57702 195644 57734
rect 196384 57942 196390 57974
rect 196454 57974 196455 58006
rect 196792 58006 196868 58012
rect 196454 57942 196460 57974
rect 196384 57734 196460 57942
rect 195638 57670 195639 57702
rect 195573 57669 195639 57670
rect 196384 57670 196390 57734
rect 196454 57670 196460 57734
rect 196792 57942 196798 58006
rect 196862 57942 196868 58006
rect 196792 57734 196868 57942
rect 196792 57702 196798 57734
rect 196384 57664 196460 57670
rect 196797 57670 196798 57702
rect 196862 57702 196868 57734
rect 196862 57670 196863 57702
rect 196797 57669 196863 57670
rect 21760 57598 21836 57604
rect 21760 57534 21766 57598
rect 21830 57534 21836 57598
rect 21760 57326 21836 57534
rect 21760 57294 21766 57326
rect 21765 57262 21766 57294
rect 21830 57294 21836 57326
rect 22168 57598 22244 57604
rect 22168 57534 22174 57598
rect 22238 57534 22244 57598
rect 22168 57326 22244 57534
rect 22168 57294 22174 57326
rect 21830 57262 21831 57294
rect 21765 57261 21831 57262
rect 22173 57262 22174 57294
rect 22238 57294 22244 57326
rect 22576 57598 22652 57604
rect 22576 57534 22582 57598
rect 22646 57534 22652 57598
rect 22989 57598 23055 57599
rect 22989 57566 22990 57598
rect 22576 57326 22652 57534
rect 22576 57294 22582 57326
rect 22238 57262 22239 57294
rect 22173 57261 22239 57262
rect 22581 57262 22582 57294
rect 22646 57294 22652 57326
rect 22984 57534 22990 57566
rect 23054 57566 23055 57598
rect 23533 57598 23599 57599
rect 23533 57566 23534 57598
rect 23054 57534 23060 57566
rect 22984 57326 23060 57534
rect 22646 57262 22647 57294
rect 22581 57261 22647 57262
rect 22984 57262 22990 57326
rect 23054 57262 23060 57326
rect 22984 57256 23060 57262
rect 23528 57534 23534 57566
rect 23598 57566 23599 57598
rect 195165 57598 195231 57599
rect 195165 57566 195166 57598
rect 23598 57534 23604 57566
rect 23528 57326 23604 57534
rect 23528 57262 23534 57326
rect 23598 57262 23604 57326
rect 23528 57256 23604 57262
rect 195160 57534 195166 57566
rect 195230 57566 195231 57598
rect 195437 57598 195503 57599
rect 195437 57566 195438 57598
rect 195230 57534 195236 57566
rect 195160 57326 195236 57534
rect 195160 57262 195166 57326
rect 195230 57262 195236 57326
rect 195160 57256 195236 57262
rect 195432 57534 195438 57566
rect 195502 57566 195503 57598
rect 196117 57598 196183 57599
rect 196117 57566 196118 57598
rect 195502 57534 195508 57566
rect 195432 57326 195508 57534
rect 195432 57262 195438 57326
rect 195502 57262 195508 57326
rect 195432 57256 195508 57262
rect 196112 57534 196118 57566
rect 196182 57566 196183 57598
rect 196248 57598 196324 57604
rect 196182 57534 196188 57566
rect 196112 57326 196188 57534
rect 196112 57262 196118 57326
rect 196182 57262 196188 57326
rect 196248 57534 196254 57598
rect 196318 57534 196324 57598
rect 196661 57598 196727 57599
rect 196661 57566 196662 57598
rect 196248 57326 196324 57534
rect 196248 57294 196254 57326
rect 196112 57256 196188 57262
rect 196253 57262 196254 57294
rect 196318 57294 196324 57326
rect 196656 57534 196662 57566
rect 196726 57566 196727 57598
rect 217464 57598 217812 59302
rect 196726 57534 196732 57566
rect 196656 57326 196732 57534
rect 196318 57262 196319 57294
rect 196253 57261 196319 57262
rect 196656 57262 196662 57326
rect 196726 57262 196732 57326
rect 196656 57256 196732 57262
rect 217464 57534 217470 57598
rect 217534 57534 217812 57598
rect 21765 57190 21831 57191
rect 21765 57158 21766 57190
rect 21760 57126 21766 57158
rect 21830 57158 21831 57190
rect 23125 57190 23191 57191
rect 23125 57158 23126 57190
rect 21830 57126 21836 57158
rect 21760 56918 21836 57126
rect 21760 56854 21766 56918
rect 21830 56854 21836 56918
rect 21760 56848 21836 56854
rect 23120 57126 23126 57158
rect 23190 57158 23191 57190
rect 23533 57190 23599 57191
rect 23533 57158 23534 57190
rect 23190 57126 23196 57158
rect 23120 56918 23196 57126
rect 23120 56854 23126 56918
rect 23190 56854 23196 56918
rect 23120 56848 23196 56854
rect 23528 57126 23534 57158
rect 23598 57158 23599 57190
rect 195165 57190 195231 57191
rect 195165 57158 195166 57190
rect 23598 57126 23604 57158
rect 23528 56918 23604 57126
rect 23528 56854 23534 56918
rect 23598 56854 23604 56918
rect 23528 56848 23604 56854
rect 195160 57126 195166 57158
rect 195230 57158 195231 57190
rect 195432 57190 195508 57196
rect 195230 57126 195236 57158
rect 195160 56918 195236 57126
rect 195160 56854 195166 56918
rect 195230 56854 195236 56918
rect 195432 57126 195438 57190
rect 195502 57126 195508 57190
rect 195845 57190 195911 57191
rect 195845 57158 195846 57190
rect 195432 56918 195508 57126
rect 195432 56886 195438 56918
rect 195160 56848 195236 56854
rect 195437 56854 195438 56886
rect 195502 56886 195508 56918
rect 195840 57126 195846 57158
rect 195910 57158 195911 57190
rect 196112 57190 196188 57196
rect 195910 57126 195916 57158
rect 195840 56918 195916 57126
rect 195502 56854 195503 56886
rect 195437 56853 195503 56854
rect 195840 56854 195846 56918
rect 195910 56854 195916 56918
rect 196112 57126 196118 57190
rect 196182 57126 196188 57190
rect 196112 56918 196188 57126
rect 196112 56886 196118 56918
rect 195840 56848 195916 56854
rect 196117 56854 196118 56886
rect 196182 56886 196188 56918
rect 196792 57190 196868 57196
rect 196792 57126 196798 57190
rect 196862 57126 196868 57190
rect 196792 56918 196868 57126
rect 196792 56886 196798 56918
rect 196182 56854 196183 56886
rect 196117 56853 196183 56854
rect 196797 56854 196798 56886
rect 196862 56886 196868 56918
rect 196862 56854 196863 56886
rect 196797 56853 196863 56854
rect 22168 56782 22244 56788
rect 22168 56718 22174 56782
rect 22238 56718 22244 56782
rect 22717 56782 22783 56783
rect 22717 56750 22718 56782
rect 22168 56510 22244 56718
rect 22168 56478 22174 56510
rect 22173 56446 22174 56478
rect 22238 56478 22244 56510
rect 22712 56718 22718 56750
rect 22782 56750 22783 56782
rect 22984 56782 23060 56788
rect 22782 56718 22788 56750
rect 22712 56510 22788 56718
rect 22238 56446 22239 56478
rect 22173 56445 22239 56446
rect 22712 56446 22718 56510
rect 22782 56446 22788 56510
rect 22984 56718 22990 56782
rect 23054 56718 23060 56782
rect 22984 56510 23060 56718
rect 22984 56478 22990 56510
rect 22712 56440 22788 56446
rect 22989 56446 22990 56478
rect 23054 56478 23060 56510
rect 23528 56782 23604 56788
rect 23528 56718 23534 56782
rect 23598 56718 23604 56782
rect 23528 56510 23604 56718
rect 195160 56782 195236 56788
rect 195160 56718 195166 56782
rect 195230 56718 195236 56782
rect 195437 56782 195503 56783
rect 195437 56750 195438 56782
rect 190269 56646 190335 56647
rect 190269 56614 190270 56646
rect 23528 56478 23534 56510
rect 23054 56446 23055 56478
rect 22989 56445 23055 56446
rect 23533 56446 23534 56478
rect 23598 56478 23604 56510
rect 190264 56582 190270 56614
rect 190334 56614 190335 56646
rect 190334 56582 190340 56614
rect 23598 56446 23599 56478
rect 23533 56445 23599 56446
rect 22989 56374 23055 56375
rect 22989 56342 22990 56374
rect 22984 56310 22990 56342
rect 23054 56342 23055 56374
rect 23533 56374 23599 56375
rect 23533 56342 23534 56374
rect 23054 56310 23060 56342
rect 22984 56102 23060 56310
rect 22984 56038 22990 56102
rect 23054 56038 23060 56102
rect 22984 56032 23060 56038
rect 23528 56310 23534 56342
rect 23598 56342 23599 56374
rect 190264 56374 190340 56582
rect 195160 56510 195236 56718
rect 195160 56478 195166 56510
rect 195165 56446 195166 56478
rect 195230 56478 195236 56510
rect 195432 56718 195438 56750
rect 195502 56750 195503 56782
rect 196248 56782 196324 56788
rect 195502 56718 195508 56750
rect 195432 56510 195508 56718
rect 195230 56446 195231 56478
rect 195165 56445 195231 56446
rect 195432 56446 195438 56510
rect 195502 56446 195508 56510
rect 196248 56718 196254 56782
rect 196318 56718 196324 56782
rect 196248 56510 196324 56718
rect 196248 56478 196254 56510
rect 195432 56440 195508 56446
rect 196253 56446 196254 56478
rect 196318 56478 196324 56510
rect 196318 56446 196319 56478
rect 196253 56445 196319 56446
rect 23598 56310 23604 56342
rect 23528 56102 23604 56310
rect 190264 56310 190270 56374
rect 190334 56310 190340 56374
rect 190264 56304 190340 56310
rect 195160 56374 195236 56380
rect 195160 56310 195166 56374
rect 195230 56310 195236 56374
rect 23528 56038 23534 56102
rect 23598 56038 23604 56102
rect 195160 56102 195236 56310
rect 195160 56070 195166 56102
rect 23528 56032 23604 56038
rect 195165 56038 195166 56070
rect 195230 56070 195236 56102
rect 195568 56374 195644 56380
rect 195568 56310 195574 56374
rect 195638 56310 195644 56374
rect 195568 56102 195644 56310
rect 195568 56070 195574 56102
rect 195230 56038 195231 56070
rect 195165 56037 195231 56038
rect 195573 56038 195574 56070
rect 195638 56070 195644 56102
rect 195638 56038 195639 56070
rect 195573 56037 195639 56038
rect 952 55902 1230 55966
rect 1294 55902 1300 55966
rect 952 54198 1300 55902
rect 22712 55966 22788 55972
rect 22712 55902 22718 55966
rect 22782 55902 22788 55966
rect 22989 55966 23055 55967
rect 22989 55934 22990 55966
rect 21760 55694 21836 55700
rect 21760 55630 21766 55694
rect 21830 55630 21836 55694
rect 22712 55694 22788 55902
rect 22712 55662 22718 55694
rect 21760 55422 21836 55630
rect 22717 55630 22718 55662
rect 22782 55662 22788 55694
rect 22984 55902 22990 55934
rect 23054 55934 23055 55966
rect 23397 55966 23463 55967
rect 23397 55934 23398 55966
rect 23054 55902 23060 55934
rect 22984 55694 23060 55902
rect 22782 55630 22783 55662
rect 22717 55629 22783 55630
rect 22984 55630 22990 55694
rect 23054 55630 23060 55694
rect 22984 55624 23060 55630
rect 23392 55902 23398 55934
rect 23462 55934 23463 55966
rect 195029 55966 195095 55967
rect 195029 55934 195030 55966
rect 23462 55902 23468 55934
rect 23392 55694 23468 55902
rect 195024 55902 195030 55934
rect 195094 55934 195095 55966
rect 195437 55966 195503 55967
rect 195437 55934 195438 55966
rect 195094 55902 195100 55934
rect 23392 55630 23398 55694
rect 23462 55630 23468 55694
rect 23392 55624 23468 55630
rect 28288 55830 28364 55836
rect 28288 55766 28294 55830
rect 28358 55766 28364 55830
rect 28288 55558 28364 55766
rect 195024 55694 195100 55902
rect 195024 55630 195030 55694
rect 195094 55630 195100 55694
rect 195024 55624 195100 55630
rect 195432 55902 195438 55934
rect 195502 55934 195503 55966
rect 195981 55966 196047 55967
rect 195981 55934 195982 55966
rect 195502 55902 195508 55934
rect 195432 55694 195508 55902
rect 195432 55630 195438 55694
rect 195502 55630 195508 55694
rect 195432 55624 195508 55630
rect 195976 55902 195982 55934
rect 196046 55934 196047 55966
rect 196117 55966 196183 55967
rect 196117 55934 196118 55966
rect 196046 55902 196052 55934
rect 195976 55694 196052 55902
rect 195976 55630 195982 55694
rect 196046 55630 196052 55694
rect 195976 55624 196052 55630
rect 196112 55902 196118 55934
rect 196182 55934 196183 55966
rect 217464 55966 217812 57534
rect 196182 55902 196188 55934
rect 196112 55694 196188 55902
rect 217464 55902 217470 55966
rect 217534 55902 217812 55966
rect 196112 55630 196118 55694
rect 196182 55630 196188 55694
rect 196112 55624 196188 55630
rect 196656 55694 196732 55700
rect 196656 55630 196662 55694
rect 196726 55630 196732 55694
rect 28288 55526 28294 55558
rect 28293 55494 28294 55526
rect 28358 55526 28364 55558
rect 28358 55494 28359 55526
rect 28293 55493 28359 55494
rect 21760 55390 21766 55422
rect 21765 55358 21766 55390
rect 21830 55390 21836 55422
rect 28288 55422 28364 55428
rect 21830 55358 21831 55390
rect 21765 55357 21831 55358
rect 28288 55358 28294 55422
rect 28358 55358 28364 55422
rect 190133 55422 190199 55423
rect 190133 55390 190134 55422
rect 21765 55286 21831 55287
rect 21765 55254 21766 55286
rect 21760 55222 21766 55254
rect 21830 55254 21831 55286
rect 22581 55286 22647 55287
rect 22581 55254 22582 55286
rect 21830 55222 21836 55254
rect 21760 55014 21836 55222
rect 21760 54950 21766 55014
rect 21830 54950 21836 55014
rect 21760 54944 21836 54950
rect 22576 55222 22582 55254
rect 22646 55254 22647 55286
rect 22646 55222 22652 55254
rect 22576 55014 22652 55222
rect 28288 55150 28364 55358
rect 28288 55118 28294 55150
rect 28293 55086 28294 55118
rect 28358 55118 28364 55150
rect 190128 55358 190134 55390
rect 190198 55390 190199 55422
rect 196656 55422 196732 55630
rect 196656 55390 196662 55422
rect 190198 55358 190204 55390
rect 190128 55150 190204 55358
rect 196661 55358 196662 55390
rect 196726 55390 196732 55422
rect 196726 55358 196727 55390
rect 196661 55357 196727 55358
rect 196117 55286 196183 55287
rect 196117 55254 196118 55286
rect 28358 55086 28359 55118
rect 28293 55085 28359 55086
rect 190128 55086 190134 55150
rect 190198 55086 190204 55150
rect 190128 55080 190204 55086
rect 196112 55222 196118 55254
rect 196182 55254 196183 55286
rect 196661 55286 196727 55287
rect 196661 55254 196662 55286
rect 196182 55222 196188 55254
rect 22576 54950 22582 55014
rect 22646 54950 22652 55014
rect 28565 55014 28631 55015
rect 28565 54982 28566 55014
rect 22576 54944 22652 54950
rect 28560 54950 28566 54982
rect 28630 54982 28631 55014
rect 190264 55014 190340 55020
rect 28630 54950 28636 54982
rect 21901 54878 21967 54879
rect 21901 54846 21902 54878
rect 21896 54814 21902 54846
rect 21966 54846 21967 54878
rect 21966 54814 21972 54846
rect 21896 54606 21972 54814
rect 21896 54542 21902 54606
rect 21966 54542 21972 54606
rect 21896 54536 21972 54542
rect 28288 54742 28364 54748
rect 28288 54678 28294 54742
rect 28358 54678 28364 54742
rect 952 54134 1230 54198
rect 1294 54134 1300 54198
rect 21760 54470 21836 54476
rect 21760 54406 21766 54470
rect 21830 54406 21836 54470
rect 22445 54470 22511 54471
rect 22445 54438 22446 54470
rect 21760 54198 21836 54406
rect 21760 54166 21766 54198
rect 952 52566 1300 54134
rect 21765 54134 21766 54166
rect 21830 54166 21836 54198
rect 22440 54406 22446 54438
rect 22510 54438 22511 54470
rect 23120 54470 23196 54476
rect 22510 54406 22516 54438
rect 22440 54198 22516 54406
rect 21830 54134 21831 54166
rect 21765 54133 21831 54134
rect 22440 54134 22446 54198
rect 22510 54134 22516 54198
rect 23120 54406 23126 54470
rect 23190 54406 23196 54470
rect 23397 54470 23463 54471
rect 23397 54438 23398 54470
rect 23120 54198 23196 54406
rect 23120 54166 23126 54198
rect 22440 54128 22516 54134
rect 23125 54134 23126 54166
rect 23190 54166 23196 54198
rect 23392 54406 23398 54438
rect 23462 54438 23463 54470
rect 28288 54470 28364 54678
rect 28560 54742 28636 54950
rect 28560 54678 28566 54742
rect 28630 54678 28636 54742
rect 190264 54950 190270 55014
rect 190334 54950 190340 55014
rect 190264 54742 190340 54950
rect 196112 55014 196188 55222
rect 196112 54950 196118 55014
rect 196182 54950 196188 55014
rect 196112 54944 196188 54950
rect 196656 55222 196662 55254
rect 196726 55254 196727 55286
rect 196726 55222 196732 55254
rect 196656 55014 196732 55222
rect 196656 54950 196662 55014
rect 196726 54950 196732 55014
rect 196656 54944 196732 54950
rect 190264 54710 190270 54742
rect 28560 54672 28636 54678
rect 190269 54678 190270 54710
rect 190334 54710 190340 54742
rect 196792 54878 196868 54884
rect 196792 54814 196798 54878
rect 196862 54814 196868 54878
rect 190334 54678 190335 54710
rect 190269 54677 190335 54678
rect 196792 54606 196868 54814
rect 196792 54574 196798 54606
rect 196797 54542 196798 54574
rect 196862 54574 196868 54606
rect 196862 54542 196863 54574
rect 196797 54541 196863 54542
rect 28288 54438 28294 54470
rect 23462 54406 23468 54438
rect 23392 54198 23468 54406
rect 28293 54406 28294 54438
rect 28358 54438 28364 54470
rect 195160 54470 195236 54476
rect 28358 54406 28359 54438
rect 28293 54405 28359 54406
rect 195160 54406 195166 54470
rect 195230 54406 195236 54470
rect 195573 54470 195639 54471
rect 195573 54438 195574 54470
rect 23190 54134 23191 54166
rect 23125 54133 23191 54134
rect 23392 54134 23398 54198
rect 23462 54134 23468 54198
rect 195160 54198 195236 54406
rect 195160 54166 195166 54198
rect 23392 54128 23468 54134
rect 195165 54134 195166 54166
rect 195230 54166 195236 54198
rect 195568 54406 195574 54438
rect 195638 54438 195639 54470
rect 195840 54470 195916 54476
rect 195638 54406 195644 54438
rect 195568 54198 195644 54406
rect 195230 54134 195231 54166
rect 195165 54133 195231 54134
rect 195568 54134 195574 54198
rect 195638 54134 195644 54198
rect 195840 54406 195846 54470
rect 195910 54406 195916 54470
rect 196389 54470 196455 54471
rect 196389 54438 196390 54470
rect 195840 54198 195916 54406
rect 195840 54166 195846 54198
rect 195568 54128 195644 54134
rect 195845 54134 195846 54166
rect 195910 54166 195916 54198
rect 196384 54406 196390 54438
rect 196454 54438 196455 54470
rect 196797 54470 196863 54471
rect 196797 54438 196798 54470
rect 196454 54406 196460 54438
rect 196384 54198 196460 54406
rect 195910 54134 195911 54166
rect 195845 54133 195911 54134
rect 196384 54134 196390 54198
rect 196454 54134 196460 54198
rect 196384 54128 196460 54134
rect 196792 54406 196798 54438
rect 196862 54438 196863 54470
rect 196862 54406 196868 54438
rect 196792 54198 196868 54406
rect 196792 54134 196798 54198
rect 196862 54134 196868 54198
rect 196792 54128 196868 54134
rect 217464 54334 217812 55902
rect 217464 54270 217470 54334
rect 217534 54270 217812 54334
rect 21896 54062 21972 54068
rect 21896 53998 21902 54062
rect 21966 53998 21972 54062
rect 21896 53790 21972 53998
rect 21896 53758 21902 53790
rect 21901 53726 21902 53758
rect 21966 53758 21972 53790
rect 22304 54062 22380 54068
rect 22304 53998 22310 54062
rect 22374 53998 22380 54062
rect 22304 53790 22380 53998
rect 22304 53758 22310 53790
rect 21966 53726 21967 53758
rect 21901 53725 21967 53726
rect 22309 53726 22310 53758
rect 22374 53758 22380 53790
rect 22712 54062 22788 54068
rect 22712 53998 22718 54062
rect 22782 53998 22788 54062
rect 22712 53790 22788 53998
rect 22712 53758 22718 53790
rect 22374 53726 22375 53758
rect 22309 53725 22375 53726
rect 22717 53726 22718 53758
rect 22782 53758 22788 53790
rect 22984 54062 23060 54068
rect 22984 53998 22990 54062
rect 23054 53998 23060 54062
rect 22984 53790 23060 53998
rect 22984 53758 22990 53790
rect 22782 53726 22783 53758
rect 22717 53725 22783 53726
rect 22989 53726 22990 53758
rect 23054 53758 23060 53790
rect 23392 54062 23468 54068
rect 23392 53998 23398 54062
rect 23462 53998 23468 54062
rect 195165 54062 195231 54063
rect 195165 54030 195166 54062
rect 23392 53790 23468 53998
rect 23392 53758 23398 53790
rect 23054 53726 23055 53758
rect 22989 53725 23055 53726
rect 23397 53726 23398 53758
rect 23462 53758 23468 53790
rect 195160 53998 195166 54030
rect 195230 54030 195231 54062
rect 195573 54062 195639 54063
rect 195573 54030 195574 54062
rect 195230 53998 195236 54030
rect 195160 53790 195236 53998
rect 23462 53726 23463 53758
rect 23397 53725 23463 53726
rect 195160 53726 195166 53790
rect 195230 53726 195236 53790
rect 195160 53720 195236 53726
rect 195568 53998 195574 54030
rect 195638 54030 195639 54062
rect 196792 54062 196868 54068
rect 195638 53998 195644 54030
rect 195568 53790 195644 53998
rect 195568 53726 195574 53790
rect 195638 53726 195644 53790
rect 196792 53998 196798 54062
rect 196862 53998 196868 54062
rect 196792 53790 196868 53998
rect 196792 53758 196798 53790
rect 195568 53720 195644 53726
rect 196797 53726 196798 53758
rect 196862 53758 196868 53790
rect 196862 53726 196863 53758
rect 196797 53725 196863 53726
rect 21901 53654 21967 53655
rect 21901 53622 21902 53654
rect 21896 53590 21902 53622
rect 21966 53622 21967 53654
rect 23120 53654 23196 53660
rect 21966 53590 21972 53622
rect 21896 53382 21972 53590
rect 21896 53318 21902 53382
rect 21966 53318 21972 53382
rect 23120 53590 23126 53654
rect 23190 53590 23196 53654
rect 23120 53382 23196 53590
rect 23120 53350 23126 53382
rect 21896 53312 21972 53318
rect 23125 53318 23126 53350
rect 23190 53350 23196 53382
rect 23392 53654 23468 53660
rect 23392 53590 23398 53654
rect 23462 53590 23468 53654
rect 195029 53654 195095 53655
rect 195029 53622 195030 53654
rect 23392 53382 23468 53590
rect 23392 53350 23398 53382
rect 23190 53318 23191 53350
rect 23125 53317 23191 53318
rect 23397 53318 23398 53350
rect 23462 53350 23468 53382
rect 195024 53590 195030 53622
rect 195094 53622 195095 53654
rect 195568 53654 195644 53660
rect 195094 53590 195100 53622
rect 195024 53382 195100 53590
rect 23462 53318 23463 53350
rect 23397 53317 23463 53318
rect 195024 53318 195030 53382
rect 195094 53318 195100 53382
rect 195568 53590 195574 53654
rect 195638 53590 195644 53654
rect 196389 53654 196455 53655
rect 196389 53622 196390 53654
rect 195568 53382 195644 53590
rect 195568 53350 195574 53382
rect 195024 53312 195100 53318
rect 195573 53318 195574 53350
rect 195638 53350 195644 53382
rect 196384 53590 196390 53622
rect 196454 53622 196455 53654
rect 196797 53654 196863 53655
rect 196797 53622 196798 53654
rect 196454 53590 196460 53622
rect 196384 53382 196460 53590
rect 195638 53318 195639 53350
rect 195573 53317 195639 53318
rect 196384 53318 196390 53382
rect 196454 53318 196460 53382
rect 196384 53312 196460 53318
rect 196792 53590 196798 53622
rect 196862 53622 196863 53654
rect 196862 53590 196868 53622
rect 196792 53382 196868 53590
rect 196792 53318 196798 53382
rect 196862 53318 196868 53382
rect 196792 53312 196868 53318
rect 21760 53246 21836 53252
rect 21760 53182 21766 53246
rect 21830 53182 21836 53246
rect 22445 53246 22511 53247
rect 22445 53214 22446 53246
rect 21760 52974 21836 53182
rect 21760 52942 21766 52974
rect 21765 52910 21766 52942
rect 21830 52942 21836 52974
rect 22440 53182 22446 53214
rect 22510 53214 22511 53246
rect 22989 53246 23055 53247
rect 22989 53214 22990 53246
rect 22510 53182 22516 53214
rect 22440 52974 22516 53182
rect 21830 52910 21831 52942
rect 21765 52909 21831 52910
rect 22440 52910 22446 52974
rect 22510 52910 22516 52974
rect 22440 52904 22516 52910
rect 22984 53182 22990 53214
rect 23054 53214 23055 53246
rect 23533 53246 23599 53247
rect 23533 53214 23534 53246
rect 23054 53182 23060 53214
rect 22984 52974 23060 53182
rect 22984 52910 22990 52974
rect 23054 52910 23060 52974
rect 22984 52904 23060 52910
rect 23528 53182 23534 53214
rect 23598 53214 23599 53246
rect 195165 53246 195231 53247
rect 195165 53214 195166 53246
rect 23598 53182 23604 53214
rect 23528 52974 23604 53182
rect 23528 52910 23534 52974
rect 23598 52910 23604 52974
rect 23528 52904 23604 52910
rect 195160 53182 195166 53214
rect 195230 53214 195231 53246
rect 195437 53246 195503 53247
rect 195437 53214 195438 53246
rect 195230 53182 195236 53214
rect 195160 52974 195236 53182
rect 195160 52910 195166 52974
rect 195230 52910 195236 52974
rect 195160 52904 195236 52910
rect 195432 53182 195438 53214
rect 195502 53214 195503 53246
rect 195845 53246 195911 53247
rect 195845 53214 195846 53246
rect 195502 53182 195508 53214
rect 195432 52974 195508 53182
rect 195432 52910 195438 52974
rect 195502 52910 195508 52974
rect 195432 52904 195508 52910
rect 195840 53182 195846 53214
rect 195910 53214 195911 53246
rect 196389 53246 196455 53247
rect 196389 53214 196390 53246
rect 195910 53182 195916 53214
rect 195840 52974 195916 53182
rect 195840 52910 195846 52974
rect 195910 52910 195916 52974
rect 195840 52904 195916 52910
rect 196384 53182 196390 53214
rect 196454 53214 196455 53246
rect 196656 53246 196732 53252
rect 196454 53182 196460 53214
rect 196384 52974 196460 53182
rect 196384 52910 196390 52974
rect 196454 52910 196460 52974
rect 196656 53182 196662 53246
rect 196726 53182 196732 53246
rect 196656 52974 196732 53182
rect 196656 52942 196662 52974
rect 196384 52904 196460 52910
rect 196661 52910 196662 52942
rect 196726 52942 196732 52974
rect 196726 52910 196727 52942
rect 196661 52909 196727 52910
rect 952 52502 1230 52566
rect 1294 52502 1300 52566
rect 22304 52838 22380 52844
rect 22304 52774 22310 52838
rect 22374 52774 22380 52838
rect 22304 52566 22380 52774
rect 22304 52534 22310 52566
rect 952 50934 1300 52502
rect 22309 52502 22310 52534
rect 22374 52534 22380 52566
rect 22984 52838 23060 52844
rect 22984 52774 22990 52838
rect 23054 52774 23060 52838
rect 22984 52566 23060 52774
rect 22984 52534 22990 52566
rect 22374 52502 22375 52534
rect 22309 52501 22375 52502
rect 22989 52502 22990 52534
rect 23054 52534 23060 52566
rect 23392 52838 23468 52844
rect 23392 52774 23398 52838
rect 23462 52774 23468 52838
rect 195165 52838 195231 52839
rect 195165 52806 195166 52838
rect 23392 52566 23468 52774
rect 23392 52534 23398 52566
rect 23054 52502 23055 52534
rect 22989 52501 23055 52502
rect 23397 52502 23398 52534
rect 23462 52534 23468 52566
rect 195160 52774 195166 52806
rect 195230 52806 195231 52838
rect 195432 52838 195508 52844
rect 195230 52774 195236 52806
rect 195160 52566 195236 52774
rect 23462 52502 23463 52534
rect 23397 52501 23463 52502
rect 195160 52502 195166 52566
rect 195230 52502 195236 52566
rect 195432 52774 195438 52838
rect 195502 52774 195508 52838
rect 195432 52566 195508 52774
rect 195432 52534 195438 52566
rect 195160 52496 195236 52502
rect 195437 52502 195438 52534
rect 195502 52534 195508 52566
rect 195976 52838 196052 52844
rect 195976 52774 195982 52838
rect 196046 52774 196052 52838
rect 195976 52566 196052 52774
rect 195976 52534 195982 52566
rect 195502 52502 195503 52534
rect 195437 52501 195503 52502
rect 195981 52502 195982 52534
rect 196046 52534 196052 52566
rect 196112 52838 196188 52844
rect 196112 52774 196118 52838
rect 196182 52774 196188 52838
rect 196112 52566 196188 52774
rect 196112 52534 196118 52566
rect 196046 52502 196047 52534
rect 195981 52501 196047 52502
rect 196117 52502 196118 52534
rect 196182 52534 196188 52566
rect 196384 52838 196460 52844
rect 196384 52774 196390 52838
rect 196454 52774 196460 52838
rect 196384 52566 196460 52774
rect 196384 52534 196390 52566
rect 196182 52502 196183 52534
rect 196117 52501 196183 52502
rect 196389 52502 196390 52534
rect 196454 52534 196460 52566
rect 217464 52702 217812 54270
rect 217464 52638 217470 52702
rect 217534 52638 217812 52702
rect 196454 52502 196455 52534
rect 196389 52501 196455 52502
rect 22989 52430 23055 52431
rect 22989 52398 22990 52430
rect 22984 52366 22990 52398
rect 23054 52398 23055 52430
rect 23397 52430 23463 52431
rect 23397 52398 23398 52430
rect 23054 52366 23060 52398
rect 22984 52158 23060 52366
rect 22984 52094 22990 52158
rect 23054 52094 23060 52158
rect 22984 52088 23060 52094
rect 23392 52366 23398 52398
rect 23462 52398 23463 52430
rect 195160 52430 195236 52436
rect 23462 52366 23468 52398
rect 23392 52158 23468 52366
rect 23392 52094 23398 52158
rect 23462 52094 23468 52158
rect 195160 52366 195166 52430
rect 195230 52366 195236 52430
rect 195160 52158 195236 52366
rect 195160 52126 195166 52158
rect 23392 52088 23468 52094
rect 195165 52094 195166 52126
rect 195230 52126 195236 52158
rect 195432 52430 195508 52436
rect 195432 52366 195438 52430
rect 195502 52366 195508 52430
rect 195432 52158 195508 52366
rect 195432 52126 195438 52158
rect 195230 52094 195231 52126
rect 195165 52093 195231 52094
rect 195437 52094 195438 52126
rect 195502 52126 195508 52158
rect 195502 52094 195503 52126
rect 195437 52093 195503 52094
rect 22440 52022 22516 52028
rect 22440 51958 22446 52022
rect 22510 51958 22516 52022
rect 21896 51750 21972 51756
rect 21896 51686 21902 51750
rect 21966 51686 21972 51750
rect 22440 51750 22516 51958
rect 22440 51718 22446 51750
rect 21896 51478 21972 51686
rect 22445 51686 22446 51718
rect 22510 51718 22516 51750
rect 23120 52022 23196 52028
rect 23120 51958 23126 52022
rect 23190 51958 23196 52022
rect 23120 51750 23196 51958
rect 23120 51718 23126 51750
rect 22510 51686 22511 51718
rect 22445 51685 22511 51686
rect 23125 51686 23126 51718
rect 23190 51718 23196 51750
rect 23528 52022 23604 52028
rect 23528 51958 23534 52022
rect 23598 51958 23604 52022
rect 23528 51750 23604 51958
rect 195160 52022 195236 52028
rect 195160 51958 195166 52022
rect 195230 51958 195236 52022
rect 195437 52022 195503 52023
rect 195437 51990 195438 52022
rect 23528 51718 23534 51750
rect 23190 51686 23191 51718
rect 23125 51685 23191 51686
rect 23533 51686 23534 51718
rect 23598 51718 23604 51750
rect 28288 51886 28364 51892
rect 28288 51822 28294 51886
rect 28358 51822 28364 51886
rect 23598 51686 23599 51718
rect 23533 51685 23599 51686
rect 28288 51614 28364 51822
rect 195160 51750 195236 51958
rect 195160 51718 195166 51750
rect 195165 51686 195166 51718
rect 195230 51718 195236 51750
rect 195432 51958 195438 51990
rect 195502 51990 195503 52022
rect 195845 52022 195911 52023
rect 195845 51990 195846 52022
rect 195502 51958 195508 51990
rect 195432 51750 195508 51958
rect 195230 51686 195231 51718
rect 195165 51685 195231 51686
rect 195432 51686 195438 51750
rect 195502 51686 195508 51750
rect 195432 51680 195508 51686
rect 195840 51958 195846 51990
rect 195910 51990 195911 52022
rect 195910 51958 195916 51990
rect 195840 51750 195916 51958
rect 195840 51686 195846 51750
rect 195910 51686 195916 51750
rect 196661 51750 196727 51751
rect 196661 51718 196662 51750
rect 195840 51680 195916 51686
rect 196656 51686 196662 51718
rect 196726 51718 196727 51750
rect 196726 51686 196732 51718
rect 28288 51582 28294 51614
rect 28293 51550 28294 51582
rect 28358 51582 28364 51614
rect 28358 51550 28359 51582
rect 28293 51549 28359 51550
rect 21896 51446 21902 51478
rect 21901 51414 21902 51446
rect 21966 51446 21972 51478
rect 28288 51478 28364 51484
rect 21966 51414 21967 51446
rect 21901 51413 21967 51414
rect 28288 51414 28294 51478
rect 28358 51414 28364 51478
rect 21760 51342 21836 51348
rect 21760 51278 21766 51342
rect 21830 51278 21836 51342
rect 21760 51070 21836 51278
rect 21760 51038 21766 51070
rect 21765 51006 21766 51038
rect 21830 51038 21836 51070
rect 22712 51342 22788 51348
rect 22712 51278 22718 51342
rect 22782 51278 22788 51342
rect 22712 51070 22788 51278
rect 28288 51206 28364 51414
rect 28288 51174 28294 51206
rect 28293 51142 28294 51174
rect 28358 51174 28364 51206
rect 190264 51478 190340 51484
rect 190264 51414 190270 51478
rect 190334 51414 190340 51478
rect 190264 51206 190340 51414
rect 196656 51478 196732 51686
rect 196656 51414 196662 51478
rect 196726 51414 196732 51478
rect 196656 51408 196732 51414
rect 195981 51342 196047 51343
rect 195981 51310 195982 51342
rect 190264 51174 190270 51206
rect 28358 51142 28359 51174
rect 28293 51141 28359 51142
rect 190269 51142 190270 51174
rect 190334 51174 190340 51206
rect 195976 51278 195982 51310
rect 196046 51310 196047 51342
rect 196656 51342 196732 51348
rect 196046 51278 196052 51310
rect 190334 51142 190335 51174
rect 190269 51141 190335 51142
rect 22712 51038 22718 51070
rect 21830 51006 21831 51038
rect 21765 51005 21831 51006
rect 22717 51006 22718 51038
rect 22782 51038 22788 51070
rect 195976 51070 196052 51278
rect 22782 51006 22783 51038
rect 22717 51005 22783 51006
rect 195976 51006 195982 51070
rect 196046 51006 196052 51070
rect 196656 51278 196662 51342
rect 196726 51278 196732 51342
rect 196656 51070 196732 51278
rect 196656 51038 196662 51070
rect 195976 51000 196052 51006
rect 196661 51006 196662 51038
rect 196726 51038 196732 51070
rect 196726 51006 196727 51038
rect 196661 51005 196727 51006
rect 952 50870 1230 50934
rect 1294 50870 1300 50934
rect 952 49302 1300 50870
rect 21760 50934 21836 50940
rect 21760 50870 21766 50934
rect 21830 50870 21836 50934
rect 21760 50662 21836 50870
rect 21760 50630 21766 50662
rect 21765 50598 21766 50630
rect 21830 50630 21836 50662
rect 196656 50934 196732 50940
rect 196656 50870 196662 50934
rect 196726 50870 196732 50934
rect 196656 50662 196732 50870
rect 196656 50630 196662 50662
rect 21830 50598 21831 50630
rect 21765 50597 21831 50598
rect 196661 50598 196662 50630
rect 196726 50630 196732 50662
rect 217464 50798 217812 52638
rect 217464 50734 217470 50798
rect 217534 50734 217812 50798
rect 196726 50598 196727 50630
rect 196661 50597 196727 50598
rect 21901 50526 21967 50527
rect 21901 50494 21902 50526
rect 21896 50462 21902 50494
rect 21966 50494 21967 50526
rect 22717 50526 22783 50527
rect 22717 50494 22718 50526
rect 21966 50462 21972 50494
rect 21896 50254 21972 50462
rect 21896 50190 21902 50254
rect 21966 50190 21972 50254
rect 21896 50184 21972 50190
rect 22712 50462 22718 50494
rect 22782 50494 22783 50526
rect 22989 50526 23055 50527
rect 22989 50494 22990 50526
rect 22782 50462 22788 50494
rect 22712 50254 22788 50462
rect 22712 50190 22718 50254
rect 22782 50190 22788 50254
rect 22712 50184 22788 50190
rect 22984 50462 22990 50494
rect 23054 50494 23055 50526
rect 23397 50526 23463 50527
rect 23397 50494 23398 50526
rect 23054 50462 23060 50494
rect 22984 50254 23060 50462
rect 22984 50190 22990 50254
rect 23054 50190 23060 50254
rect 22984 50184 23060 50190
rect 23392 50462 23398 50494
rect 23462 50494 23463 50526
rect 195024 50526 195100 50532
rect 23462 50462 23468 50494
rect 23392 50254 23468 50462
rect 195024 50462 195030 50526
rect 195094 50462 195100 50526
rect 195437 50526 195503 50527
rect 195437 50494 195438 50526
rect 23392 50190 23398 50254
rect 23462 50190 23468 50254
rect 23392 50184 23468 50190
rect 28288 50254 28364 50260
rect 28288 50190 28294 50254
rect 28358 50190 28364 50254
rect 195024 50254 195100 50462
rect 195024 50222 195030 50254
rect 21760 50118 21836 50124
rect 21760 50054 21766 50118
rect 21830 50054 21836 50118
rect 22309 50118 22375 50119
rect 22309 50086 22310 50118
rect 21760 49846 21836 50054
rect 21760 49814 21766 49846
rect 21765 49782 21766 49814
rect 21830 49814 21836 49846
rect 22304 50054 22310 50086
rect 22374 50086 22375 50118
rect 22984 50118 23060 50124
rect 22374 50054 22380 50086
rect 22304 49846 22380 50054
rect 21830 49782 21831 49814
rect 21765 49781 21831 49782
rect 22304 49782 22310 49846
rect 22374 49782 22380 49846
rect 22984 50054 22990 50118
rect 23054 50054 23060 50118
rect 23397 50118 23463 50119
rect 23397 50086 23398 50118
rect 22984 49846 23060 50054
rect 22984 49814 22990 49846
rect 22304 49776 22380 49782
rect 22989 49782 22990 49814
rect 23054 49814 23060 49846
rect 23392 50054 23398 50086
rect 23462 50086 23463 50118
rect 23462 50054 23468 50086
rect 23392 49846 23468 50054
rect 28288 49982 28364 50190
rect 195029 50190 195030 50222
rect 195094 50222 195100 50254
rect 195432 50462 195438 50494
rect 195502 50494 195503 50526
rect 195976 50526 196052 50532
rect 195502 50462 195508 50494
rect 195432 50254 195508 50462
rect 195094 50190 195095 50222
rect 195029 50189 195095 50190
rect 195432 50190 195438 50254
rect 195502 50190 195508 50254
rect 195976 50462 195982 50526
rect 196046 50462 196052 50526
rect 195976 50254 196052 50462
rect 195976 50222 195982 50254
rect 195432 50184 195508 50190
rect 195981 50190 195982 50222
rect 196046 50222 196052 50254
rect 196792 50526 196868 50532
rect 196792 50462 196798 50526
rect 196862 50462 196868 50526
rect 196792 50254 196868 50462
rect 196792 50222 196798 50254
rect 196046 50190 196047 50222
rect 195981 50189 196047 50190
rect 196797 50190 196798 50222
rect 196862 50222 196868 50254
rect 196862 50190 196863 50222
rect 196797 50189 196863 50190
rect 195029 50118 195095 50119
rect 195029 50086 195030 50118
rect 28288 49950 28294 49982
rect 28293 49918 28294 49950
rect 28358 49950 28364 49982
rect 195024 50054 195030 50086
rect 195094 50086 195095 50118
rect 195432 50118 195508 50124
rect 195094 50054 195100 50086
rect 28358 49918 28359 49950
rect 28293 49917 28359 49918
rect 23054 49782 23055 49814
rect 22989 49781 23055 49782
rect 23392 49782 23398 49846
rect 23462 49782 23468 49846
rect 23392 49776 23468 49782
rect 195024 49846 195100 50054
rect 195024 49782 195030 49846
rect 195094 49782 195100 49846
rect 195432 50054 195438 50118
rect 195502 50054 195508 50118
rect 196389 50118 196455 50119
rect 196389 50086 196390 50118
rect 195432 49846 195508 50054
rect 195432 49814 195438 49846
rect 195024 49776 195100 49782
rect 195437 49782 195438 49814
rect 195502 49814 195508 49846
rect 196384 50054 196390 50086
rect 196454 50086 196455 50118
rect 196797 50118 196863 50119
rect 196797 50086 196798 50118
rect 196454 50054 196460 50086
rect 196384 49846 196460 50054
rect 195502 49782 195503 49814
rect 195437 49781 195503 49782
rect 196384 49782 196390 49846
rect 196454 49782 196460 49846
rect 196384 49776 196460 49782
rect 196792 50054 196798 50086
rect 196862 50086 196863 50118
rect 196862 50054 196868 50086
rect 196792 49846 196868 50054
rect 196792 49782 196798 49846
rect 196862 49782 196868 49846
rect 196792 49776 196868 49782
rect 21765 49710 21831 49711
rect 21765 49678 21766 49710
rect 21760 49646 21766 49678
rect 21830 49678 21831 49710
rect 22173 49710 22239 49711
rect 22173 49678 22174 49710
rect 21830 49646 21836 49678
rect 21760 49438 21836 49646
rect 21760 49374 21766 49438
rect 21830 49374 21836 49438
rect 21760 49368 21836 49374
rect 22168 49646 22174 49678
rect 22238 49678 22239 49710
rect 22712 49710 22788 49716
rect 22238 49646 22244 49678
rect 22168 49438 22244 49646
rect 22168 49374 22174 49438
rect 22238 49374 22244 49438
rect 22712 49646 22718 49710
rect 22782 49646 22788 49710
rect 22989 49710 23055 49711
rect 22989 49678 22990 49710
rect 22712 49438 22788 49646
rect 22712 49406 22718 49438
rect 22168 49368 22244 49374
rect 22717 49374 22718 49406
rect 22782 49406 22788 49438
rect 22984 49646 22990 49678
rect 23054 49678 23055 49710
rect 23392 49710 23468 49716
rect 23054 49646 23060 49678
rect 22984 49438 23060 49646
rect 22782 49374 22783 49406
rect 22717 49373 22783 49374
rect 22984 49374 22990 49438
rect 23054 49374 23060 49438
rect 23392 49646 23398 49710
rect 23462 49646 23468 49710
rect 23392 49438 23468 49646
rect 23392 49406 23398 49438
rect 22984 49368 23060 49374
rect 23397 49374 23398 49406
rect 23462 49406 23468 49438
rect 195024 49710 195100 49716
rect 195024 49646 195030 49710
rect 195094 49646 195100 49710
rect 195437 49710 195503 49711
rect 195437 49678 195438 49710
rect 195024 49438 195100 49646
rect 195024 49406 195030 49438
rect 23462 49374 23463 49406
rect 23397 49373 23463 49374
rect 195029 49374 195030 49406
rect 195094 49406 195100 49438
rect 195432 49646 195438 49678
rect 195502 49678 195503 49710
rect 195845 49710 195911 49711
rect 195845 49678 195846 49710
rect 195502 49646 195508 49678
rect 195432 49438 195508 49646
rect 195094 49374 195095 49406
rect 195029 49373 195095 49374
rect 195432 49374 195438 49438
rect 195502 49374 195508 49438
rect 195432 49368 195508 49374
rect 195840 49646 195846 49678
rect 195910 49678 195911 49710
rect 196661 49710 196727 49711
rect 196661 49678 196662 49710
rect 195910 49646 195916 49678
rect 195840 49438 195916 49646
rect 195840 49374 195846 49438
rect 195910 49374 195916 49438
rect 195840 49368 195916 49374
rect 196656 49646 196662 49678
rect 196726 49678 196727 49710
rect 196726 49646 196732 49678
rect 196656 49438 196732 49646
rect 196656 49374 196662 49438
rect 196726 49374 196732 49438
rect 196656 49368 196732 49374
rect 952 49238 1230 49302
rect 1294 49238 1300 49302
rect 21901 49302 21967 49303
rect 21901 49270 21902 49302
rect 952 47670 1300 49238
rect 21896 49238 21902 49270
rect 21966 49270 21967 49302
rect 22309 49302 22375 49303
rect 22309 49270 22310 49302
rect 21966 49238 21972 49270
rect 21896 49030 21972 49238
rect 21896 48966 21902 49030
rect 21966 48966 21972 49030
rect 21896 48960 21972 48966
rect 22304 49238 22310 49270
rect 22374 49270 22375 49302
rect 23120 49302 23196 49308
rect 22374 49238 22380 49270
rect 22304 49030 22380 49238
rect 22304 48966 22310 49030
rect 22374 48966 22380 49030
rect 23120 49238 23126 49302
rect 23190 49238 23196 49302
rect 23397 49302 23463 49303
rect 23397 49270 23398 49302
rect 23120 49030 23196 49238
rect 23120 48998 23126 49030
rect 22304 48960 22380 48966
rect 23125 48966 23126 48998
rect 23190 48998 23196 49030
rect 23392 49238 23398 49270
rect 23462 49270 23463 49302
rect 195029 49302 195095 49303
rect 195029 49270 195030 49302
rect 23462 49238 23468 49270
rect 23392 49030 23468 49238
rect 23190 48966 23191 48998
rect 23125 48965 23191 48966
rect 23392 48966 23398 49030
rect 23462 48966 23468 49030
rect 23392 48960 23468 48966
rect 195024 49238 195030 49270
rect 195094 49270 195095 49302
rect 195568 49302 195644 49308
rect 195094 49238 195100 49270
rect 195024 49030 195100 49238
rect 195024 48966 195030 49030
rect 195094 48966 195100 49030
rect 195568 49238 195574 49302
rect 195638 49238 195644 49302
rect 195568 49030 195644 49238
rect 195568 48998 195574 49030
rect 195024 48960 195100 48966
rect 195573 48966 195574 48998
rect 195638 48998 195644 49030
rect 196384 49302 196460 49308
rect 196384 49238 196390 49302
rect 196454 49238 196460 49302
rect 196797 49302 196863 49303
rect 196797 49270 196798 49302
rect 196384 49030 196460 49238
rect 196384 48998 196390 49030
rect 195638 48966 195639 48998
rect 195573 48965 195639 48966
rect 196389 48966 196390 48998
rect 196454 48998 196460 49030
rect 196792 49238 196798 49270
rect 196862 49270 196863 49302
rect 196862 49238 196868 49270
rect 196792 49030 196868 49238
rect 196454 48966 196455 48998
rect 196389 48965 196455 48966
rect 196792 48966 196798 49030
rect 196862 48966 196868 49030
rect 196792 48960 196868 48966
rect 217464 49166 217812 50734
rect 217464 49102 217470 49166
rect 217534 49102 217812 49166
rect 22168 48894 22244 48900
rect 22168 48830 22174 48894
rect 22238 48830 22244 48894
rect 22989 48894 23055 48895
rect 22989 48862 22990 48894
rect 22168 48622 22244 48830
rect 22168 48590 22174 48622
rect 22173 48558 22174 48590
rect 22238 48590 22244 48622
rect 22984 48830 22990 48862
rect 23054 48862 23055 48894
rect 23528 48894 23604 48900
rect 23054 48830 23060 48862
rect 22984 48622 23060 48830
rect 22238 48558 22239 48590
rect 22173 48557 22239 48558
rect 22984 48558 22990 48622
rect 23054 48558 23060 48622
rect 23528 48830 23534 48894
rect 23598 48830 23604 48894
rect 195165 48894 195231 48895
rect 195165 48862 195166 48894
rect 23528 48622 23604 48830
rect 23528 48590 23534 48622
rect 22984 48552 23060 48558
rect 23533 48558 23534 48590
rect 23598 48590 23604 48622
rect 195160 48830 195166 48862
rect 195230 48862 195231 48894
rect 195437 48894 195503 48895
rect 195437 48862 195438 48894
rect 195230 48830 195236 48862
rect 195160 48622 195236 48830
rect 23598 48558 23599 48590
rect 23533 48557 23599 48558
rect 195160 48558 195166 48622
rect 195230 48558 195236 48622
rect 195160 48552 195236 48558
rect 195432 48830 195438 48862
rect 195502 48862 195503 48894
rect 195845 48894 195911 48895
rect 195845 48862 195846 48894
rect 195502 48830 195508 48862
rect 195432 48622 195508 48830
rect 195432 48558 195438 48622
rect 195502 48558 195508 48622
rect 195432 48552 195508 48558
rect 195840 48830 195846 48862
rect 195910 48862 195911 48894
rect 196248 48894 196324 48900
rect 195910 48830 195916 48862
rect 195840 48622 195916 48830
rect 195840 48558 195846 48622
rect 195910 48558 195916 48622
rect 196248 48830 196254 48894
rect 196318 48830 196324 48894
rect 196248 48622 196324 48830
rect 196248 48590 196254 48622
rect 195840 48552 195916 48558
rect 196253 48558 196254 48590
rect 196318 48590 196324 48622
rect 196318 48558 196319 48590
rect 196253 48557 196319 48558
rect 21896 48486 21972 48492
rect 21896 48422 21902 48486
rect 21966 48422 21972 48486
rect 21896 48214 21972 48422
rect 21896 48182 21902 48214
rect 21901 48150 21902 48182
rect 21966 48182 21972 48214
rect 22304 48486 22380 48492
rect 22304 48422 22310 48486
rect 22374 48422 22380 48486
rect 22581 48486 22647 48487
rect 22581 48454 22582 48486
rect 22304 48214 22380 48422
rect 22304 48182 22310 48214
rect 21966 48150 21967 48182
rect 21901 48149 21967 48150
rect 22309 48150 22310 48182
rect 22374 48182 22380 48214
rect 22576 48422 22582 48454
rect 22646 48454 22647 48486
rect 23125 48486 23191 48487
rect 23125 48454 23126 48486
rect 22646 48422 22652 48454
rect 22576 48214 22652 48422
rect 22374 48150 22375 48182
rect 22309 48149 22375 48150
rect 22576 48150 22582 48214
rect 22646 48150 22652 48214
rect 22576 48144 22652 48150
rect 23120 48422 23126 48454
rect 23190 48454 23191 48486
rect 23533 48486 23599 48487
rect 23533 48454 23534 48486
rect 23190 48422 23196 48454
rect 23120 48214 23196 48422
rect 23120 48150 23126 48214
rect 23190 48150 23196 48214
rect 23120 48144 23196 48150
rect 23528 48422 23534 48454
rect 23598 48454 23599 48486
rect 195024 48486 195100 48492
rect 23598 48422 23604 48454
rect 23528 48214 23604 48422
rect 23528 48150 23534 48214
rect 23598 48150 23604 48214
rect 195024 48422 195030 48486
rect 195094 48422 195100 48486
rect 195573 48486 195639 48487
rect 195573 48454 195574 48486
rect 195024 48214 195100 48422
rect 195024 48182 195030 48214
rect 23528 48144 23604 48150
rect 195029 48150 195030 48182
rect 195094 48182 195100 48214
rect 195568 48422 195574 48454
rect 195638 48454 195639 48486
rect 195845 48486 195911 48487
rect 195845 48454 195846 48486
rect 195638 48422 195644 48454
rect 195568 48214 195644 48422
rect 195094 48150 195095 48182
rect 195029 48149 195095 48150
rect 195568 48150 195574 48214
rect 195638 48150 195644 48214
rect 195568 48144 195644 48150
rect 195840 48422 195846 48454
rect 195910 48454 195911 48486
rect 196112 48486 196188 48492
rect 195910 48422 195916 48454
rect 195840 48214 195916 48422
rect 195840 48150 195846 48214
rect 195910 48150 195916 48214
rect 196112 48422 196118 48486
rect 196182 48422 196188 48486
rect 196112 48214 196188 48422
rect 196112 48182 196118 48214
rect 195840 48144 195916 48150
rect 196117 48150 196118 48182
rect 196182 48182 196188 48214
rect 196792 48486 196868 48492
rect 196792 48422 196798 48486
rect 196862 48422 196868 48486
rect 196792 48214 196868 48422
rect 196792 48182 196798 48214
rect 196182 48150 196183 48182
rect 196117 48149 196183 48150
rect 196797 48150 196798 48182
rect 196862 48182 196868 48214
rect 196862 48150 196863 48182
rect 196797 48149 196863 48150
rect 22717 48078 22783 48079
rect 22717 48046 22718 48078
rect 22712 48014 22718 48046
rect 22782 48046 22783 48078
rect 22984 48078 23060 48084
rect 22782 48014 22788 48046
rect 952 47606 1230 47670
rect 1294 47606 1300 47670
rect 952 46038 1300 47606
rect 21896 47806 21972 47812
rect 21896 47742 21902 47806
rect 21966 47742 21972 47806
rect 21896 47534 21972 47742
rect 22712 47806 22788 48014
rect 22712 47742 22718 47806
rect 22782 47742 22788 47806
rect 22984 48014 22990 48078
rect 23054 48014 23060 48078
rect 22984 47806 23060 48014
rect 22984 47774 22990 47806
rect 22712 47736 22788 47742
rect 22989 47742 22990 47774
rect 23054 47774 23060 47806
rect 23528 48078 23604 48084
rect 23528 48014 23534 48078
rect 23598 48014 23604 48078
rect 23528 47806 23604 48014
rect 23528 47774 23534 47806
rect 23054 47742 23055 47774
rect 22989 47741 23055 47742
rect 23533 47742 23534 47774
rect 23598 47774 23604 47806
rect 195160 48078 195236 48084
rect 195160 48014 195166 48078
rect 195230 48014 195236 48078
rect 195160 47806 195236 48014
rect 195160 47774 195166 47806
rect 23598 47742 23599 47774
rect 23533 47741 23599 47742
rect 195165 47742 195166 47774
rect 195230 47774 195236 47806
rect 195432 48078 195508 48084
rect 195432 48014 195438 48078
rect 195502 48014 195508 48078
rect 195432 47806 195508 48014
rect 195432 47774 195438 47806
rect 195230 47742 195231 47774
rect 195165 47741 195231 47742
rect 195437 47742 195438 47774
rect 195502 47774 195508 47806
rect 196248 48078 196324 48084
rect 196248 48014 196254 48078
rect 196318 48014 196324 48078
rect 196248 47806 196324 48014
rect 196248 47774 196254 47806
rect 195502 47742 195503 47774
rect 195437 47741 195503 47742
rect 196253 47742 196254 47774
rect 196318 47774 196324 47806
rect 196656 47806 196732 47812
rect 196318 47742 196319 47774
rect 196253 47741 196319 47742
rect 196656 47742 196662 47806
rect 196726 47742 196732 47806
rect 22989 47670 23055 47671
rect 22989 47638 22990 47670
rect 21896 47502 21902 47534
rect 21901 47470 21902 47502
rect 21966 47502 21972 47534
rect 22984 47606 22990 47638
rect 23054 47638 23055 47670
rect 23528 47670 23604 47676
rect 23054 47606 23060 47638
rect 21966 47470 21967 47502
rect 21901 47469 21967 47470
rect 22984 47398 23060 47606
rect 22984 47334 22990 47398
rect 23054 47334 23060 47398
rect 23528 47606 23534 47670
rect 23598 47606 23604 47670
rect 195165 47670 195231 47671
rect 195165 47638 195166 47670
rect 23528 47398 23604 47606
rect 23528 47366 23534 47398
rect 22984 47328 23060 47334
rect 23533 47334 23534 47366
rect 23598 47366 23604 47398
rect 195160 47606 195166 47638
rect 195230 47638 195231 47670
rect 195437 47670 195503 47671
rect 195437 47638 195438 47670
rect 195230 47606 195236 47638
rect 195160 47398 195236 47606
rect 23598 47334 23599 47366
rect 23533 47333 23599 47334
rect 195160 47334 195166 47398
rect 195230 47334 195236 47398
rect 195160 47328 195236 47334
rect 195432 47606 195438 47638
rect 195502 47638 195503 47670
rect 195502 47606 195508 47638
rect 195432 47398 195508 47606
rect 196656 47534 196732 47742
rect 196656 47502 196662 47534
rect 196661 47470 196662 47502
rect 196726 47502 196732 47534
rect 217464 47534 217812 49102
rect 196726 47470 196727 47502
rect 196661 47469 196727 47470
rect 217464 47470 217470 47534
rect 217534 47470 217812 47534
rect 195432 47334 195438 47398
rect 195502 47334 195508 47398
rect 195432 47328 195508 47334
rect 22440 47262 22516 47268
rect 22440 47198 22446 47262
rect 22510 47198 22516 47262
rect 21901 46990 21967 46991
rect 21901 46958 21902 46990
rect 21896 46926 21902 46958
rect 21966 46958 21967 46990
rect 22440 46990 22516 47198
rect 22440 46958 22446 46990
rect 21966 46926 21972 46958
rect 21896 46718 21972 46926
rect 22445 46926 22446 46958
rect 22510 46958 22516 46990
rect 28288 47126 28364 47132
rect 28288 47062 28294 47126
rect 28358 47062 28364 47126
rect 22510 46926 22511 46958
rect 22445 46925 22511 46926
rect 22309 46854 22375 46855
rect 22309 46822 22310 46854
rect 21896 46654 21902 46718
rect 21966 46654 21972 46718
rect 21896 46648 21972 46654
rect 22304 46790 22310 46822
rect 22374 46822 22375 46854
rect 28288 46854 28364 47062
rect 196797 46990 196863 46991
rect 196797 46958 196798 46990
rect 28288 46822 28294 46854
rect 22374 46790 22380 46822
rect 22304 46724 22380 46790
rect 28293 46790 28294 46822
rect 28358 46822 28364 46854
rect 196792 46926 196798 46958
rect 196862 46958 196863 46990
rect 196862 46926 196868 46958
rect 28358 46790 28359 46822
rect 28293 46789 28359 46790
rect 22304 46718 22516 46724
rect 22304 46654 22446 46718
rect 22510 46654 22516 46718
rect 22304 46648 22516 46654
rect 196792 46718 196868 46926
rect 196792 46654 196798 46718
rect 196862 46654 196868 46718
rect 196792 46648 196868 46654
rect 21760 46582 21836 46588
rect 21760 46518 21766 46582
rect 21830 46518 21836 46582
rect 21760 46310 21836 46518
rect 21760 46278 21766 46310
rect 21765 46246 21766 46278
rect 21830 46278 21836 46310
rect 22576 46582 22652 46588
rect 22576 46518 22582 46582
rect 22646 46518 22652 46582
rect 22989 46582 23055 46583
rect 22989 46550 22990 46582
rect 22576 46310 22652 46518
rect 22576 46278 22582 46310
rect 21830 46246 21831 46278
rect 21765 46245 21831 46246
rect 22581 46246 22582 46278
rect 22646 46278 22652 46310
rect 22984 46518 22990 46550
rect 23054 46550 23055 46582
rect 23528 46582 23604 46588
rect 23054 46518 23060 46550
rect 22984 46310 23060 46518
rect 22646 46246 22647 46278
rect 22581 46245 22647 46246
rect 22984 46246 22990 46310
rect 23054 46246 23060 46310
rect 23528 46518 23534 46582
rect 23598 46518 23604 46582
rect 195165 46582 195231 46583
rect 195165 46550 195166 46582
rect 23528 46310 23604 46518
rect 195160 46518 195166 46550
rect 195230 46550 195231 46582
rect 195437 46582 195503 46583
rect 195437 46550 195438 46582
rect 195230 46518 195236 46550
rect 23528 46278 23534 46310
rect 22984 46240 23060 46246
rect 23533 46246 23534 46278
rect 23598 46278 23604 46310
rect 190133 46310 190199 46311
rect 190133 46278 190134 46310
rect 23598 46246 23599 46278
rect 23533 46245 23599 46246
rect 190128 46246 190134 46278
rect 190198 46278 190199 46310
rect 195160 46310 195236 46518
rect 190198 46246 190204 46278
rect 21901 46174 21967 46175
rect 21901 46142 21902 46174
rect 952 45974 1230 46038
rect 1294 45974 1300 46038
rect 952 44134 1300 45974
rect 21896 46110 21902 46142
rect 21966 46142 21967 46174
rect 23120 46174 23196 46180
rect 21966 46110 21972 46142
rect 21896 45902 21972 46110
rect 21896 45838 21902 45902
rect 21966 45838 21972 45902
rect 23120 46110 23126 46174
rect 23190 46110 23196 46174
rect 23397 46174 23463 46175
rect 23397 46142 23398 46174
rect 23120 45902 23196 46110
rect 23120 45870 23126 45902
rect 21896 45832 21972 45838
rect 23125 45838 23126 45870
rect 23190 45870 23196 45902
rect 23392 46110 23398 46142
rect 23462 46142 23463 46174
rect 23462 46110 23468 46142
rect 23392 45902 23468 46110
rect 190128 46038 190204 46246
rect 195160 46246 195166 46310
rect 195230 46246 195236 46310
rect 195160 46240 195236 46246
rect 195432 46518 195438 46550
rect 195502 46550 195503 46582
rect 196253 46582 196319 46583
rect 196253 46550 196254 46582
rect 195502 46518 195508 46550
rect 195432 46310 195508 46518
rect 195432 46246 195438 46310
rect 195502 46246 195508 46310
rect 195432 46240 195508 46246
rect 196248 46518 196254 46550
rect 196318 46550 196319 46582
rect 196656 46582 196732 46588
rect 196318 46518 196324 46550
rect 196248 46310 196324 46518
rect 196248 46246 196254 46310
rect 196318 46246 196324 46310
rect 196656 46518 196662 46582
rect 196726 46518 196732 46582
rect 196656 46310 196732 46518
rect 196656 46278 196662 46310
rect 196248 46240 196324 46246
rect 196661 46246 196662 46278
rect 196726 46278 196732 46310
rect 196726 46246 196727 46278
rect 196661 46245 196727 46246
rect 190128 45974 190134 46038
rect 190198 45974 190204 46038
rect 190128 45968 190204 45974
rect 195024 46174 195100 46180
rect 195024 46110 195030 46174
rect 195094 46110 195100 46174
rect 23190 45838 23191 45870
rect 23125 45837 23191 45838
rect 23392 45838 23398 45902
rect 23462 45838 23468 45902
rect 195024 45902 195100 46110
rect 195024 45870 195030 45902
rect 23392 45832 23468 45838
rect 195029 45838 195030 45870
rect 195094 45870 195100 45902
rect 195568 46174 195644 46180
rect 195568 46110 195574 46174
rect 195638 46110 195644 46174
rect 196797 46174 196863 46175
rect 196797 46142 196798 46174
rect 195568 45902 195644 46110
rect 195568 45870 195574 45902
rect 195094 45838 195095 45870
rect 195029 45837 195095 45838
rect 195573 45838 195574 45870
rect 195638 45870 195644 45902
rect 196792 46110 196798 46142
rect 196862 46142 196863 46174
rect 196862 46110 196868 46142
rect 196792 45902 196868 46110
rect 195638 45838 195639 45870
rect 195573 45837 195639 45838
rect 196792 45838 196798 45902
rect 196862 45838 196868 45902
rect 196792 45832 196868 45838
rect 217464 46038 217812 47470
rect 217464 45974 217470 46038
rect 217534 45974 217812 46038
rect 21901 45766 21967 45767
rect 21901 45734 21902 45766
rect 21896 45702 21902 45734
rect 21966 45734 21967 45766
rect 22168 45766 22244 45772
rect 21966 45702 21972 45734
rect 14693 45630 14759 45631
rect 14693 45598 14694 45630
rect 14688 45566 14694 45598
rect 14758 45598 14759 45630
rect 14758 45566 14764 45598
rect 952 44070 1230 44134
rect 1294 44070 1300 44134
rect 952 42502 1300 44070
rect 952 42438 1230 42502
rect 1294 42438 1300 42502
rect 952 40870 1300 42438
rect 14552 44134 14628 44140
rect 14552 44070 14558 44134
rect 14622 44070 14628 44134
rect 14552 41550 14628 44070
rect 14688 42910 14764 45566
rect 21896 45494 21972 45702
rect 21896 45430 21902 45494
rect 21966 45430 21972 45494
rect 22168 45702 22174 45766
rect 22238 45702 22244 45766
rect 23125 45766 23191 45767
rect 23125 45734 23126 45766
rect 22168 45494 22244 45702
rect 22168 45462 22174 45494
rect 21896 45424 21972 45430
rect 22173 45430 22174 45462
rect 22238 45462 22244 45494
rect 23120 45702 23126 45734
rect 23190 45734 23191 45766
rect 23528 45766 23604 45772
rect 23190 45702 23196 45734
rect 23120 45494 23196 45702
rect 22238 45430 22239 45462
rect 22173 45429 22239 45430
rect 23120 45430 23126 45494
rect 23190 45430 23196 45494
rect 23528 45702 23534 45766
rect 23598 45702 23604 45766
rect 23528 45494 23604 45702
rect 23528 45462 23534 45494
rect 23120 45424 23196 45430
rect 23533 45430 23534 45462
rect 23598 45462 23604 45494
rect 195160 45766 195236 45772
rect 195160 45702 195166 45766
rect 195230 45702 195236 45766
rect 195573 45766 195639 45767
rect 195573 45734 195574 45766
rect 195160 45494 195236 45702
rect 195160 45462 195166 45494
rect 23598 45430 23599 45462
rect 23533 45429 23599 45430
rect 195165 45430 195166 45462
rect 195230 45462 195236 45494
rect 195568 45702 195574 45734
rect 195638 45734 195639 45766
rect 195840 45766 195916 45772
rect 195638 45702 195644 45734
rect 195568 45494 195644 45702
rect 195230 45430 195231 45462
rect 195165 45429 195231 45430
rect 195568 45430 195574 45494
rect 195638 45430 195644 45494
rect 195840 45702 195846 45766
rect 195910 45702 195916 45766
rect 195840 45494 195916 45702
rect 195840 45462 195846 45494
rect 195568 45424 195644 45430
rect 195845 45430 195846 45462
rect 195910 45462 195916 45494
rect 196656 45766 196732 45772
rect 196656 45702 196662 45766
rect 196726 45702 196732 45766
rect 196656 45494 196732 45702
rect 196656 45462 196662 45494
rect 195910 45430 195911 45462
rect 195845 45429 195911 45430
rect 196661 45430 196662 45462
rect 196726 45462 196732 45494
rect 196726 45430 196727 45462
rect 196661 45429 196727 45430
rect 21896 45358 21972 45364
rect 21896 45294 21902 45358
rect 21966 45294 21972 45358
rect 21896 45086 21972 45294
rect 21896 45054 21902 45086
rect 21901 45022 21902 45054
rect 21966 45054 21972 45086
rect 22712 45358 22788 45364
rect 22712 45294 22718 45358
rect 22782 45294 22788 45358
rect 22989 45358 23055 45359
rect 22989 45326 22990 45358
rect 22712 45086 22788 45294
rect 22712 45054 22718 45086
rect 21966 45022 21967 45054
rect 21901 45021 21967 45022
rect 22717 45022 22718 45054
rect 22782 45054 22788 45086
rect 22984 45294 22990 45326
rect 23054 45326 23055 45358
rect 23533 45358 23599 45359
rect 23533 45326 23534 45358
rect 23054 45294 23060 45326
rect 22984 45086 23060 45294
rect 22782 45022 22783 45054
rect 22717 45021 22783 45022
rect 22984 45022 22990 45086
rect 23054 45022 23060 45086
rect 22984 45016 23060 45022
rect 23528 45294 23534 45326
rect 23598 45326 23599 45358
rect 195165 45358 195231 45359
rect 195165 45326 195166 45358
rect 23598 45294 23604 45326
rect 23528 45086 23604 45294
rect 23528 45022 23534 45086
rect 23598 45022 23604 45086
rect 23528 45016 23604 45022
rect 195160 45294 195166 45326
rect 195230 45326 195231 45358
rect 195432 45358 195508 45364
rect 195230 45294 195236 45326
rect 195160 45086 195236 45294
rect 195160 45022 195166 45086
rect 195230 45022 195236 45086
rect 195432 45294 195438 45358
rect 195502 45294 195508 45358
rect 195845 45358 195911 45359
rect 195845 45326 195846 45358
rect 195432 45086 195508 45294
rect 195432 45054 195438 45086
rect 195160 45016 195236 45022
rect 195437 45022 195438 45054
rect 195502 45054 195508 45086
rect 195840 45294 195846 45326
rect 195910 45326 195911 45358
rect 196112 45358 196188 45364
rect 195910 45294 195916 45326
rect 195840 45086 195916 45294
rect 195502 45022 195503 45054
rect 195437 45021 195503 45022
rect 195840 45022 195846 45086
rect 195910 45022 195916 45086
rect 196112 45294 196118 45358
rect 196182 45294 196188 45358
rect 196661 45358 196727 45359
rect 196661 45326 196662 45358
rect 196112 45086 196188 45294
rect 196112 45054 196118 45086
rect 195840 45016 195916 45022
rect 196117 45022 196118 45054
rect 196182 45054 196188 45086
rect 196656 45294 196662 45326
rect 196726 45326 196727 45358
rect 196726 45294 196732 45326
rect 196656 45086 196732 45294
rect 196182 45022 196183 45054
rect 196117 45021 196183 45022
rect 196656 45022 196662 45086
rect 196726 45022 196732 45086
rect 196656 45016 196732 45022
rect 21896 44950 21972 44956
rect 21896 44886 21902 44950
rect 21966 44886 21972 44950
rect 22309 44950 22375 44951
rect 22309 44918 22310 44950
rect 21896 44678 21972 44886
rect 21896 44646 21902 44678
rect 21901 44614 21902 44646
rect 21966 44646 21972 44678
rect 22304 44886 22310 44918
rect 22374 44918 22375 44950
rect 23120 44950 23196 44956
rect 22374 44886 22380 44918
rect 22304 44678 22380 44886
rect 21966 44614 21967 44646
rect 21901 44613 21967 44614
rect 22304 44614 22310 44678
rect 22374 44614 22380 44678
rect 23120 44886 23126 44950
rect 23190 44886 23196 44950
rect 23120 44678 23196 44886
rect 23120 44646 23126 44678
rect 22304 44608 22380 44614
rect 23125 44614 23126 44646
rect 23190 44646 23196 44678
rect 23392 44950 23468 44956
rect 23392 44886 23398 44950
rect 23462 44886 23468 44950
rect 23392 44678 23468 44886
rect 23392 44646 23398 44678
rect 23190 44614 23191 44646
rect 23125 44613 23191 44614
rect 23397 44614 23398 44646
rect 23462 44646 23468 44678
rect 195024 44950 195100 44956
rect 195024 44886 195030 44950
rect 195094 44886 195100 44950
rect 195437 44950 195503 44951
rect 195437 44918 195438 44950
rect 195024 44678 195100 44886
rect 195024 44646 195030 44678
rect 23462 44614 23463 44646
rect 23397 44613 23463 44614
rect 195029 44614 195030 44646
rect 195094 44646 195100 44678
rect 195432 44886 195438 44918
rect 195502 44918 195503 44950
rect 196389 44950 196455 44951
rect 196389 44918 196390 44950
rect 195502 44886 195508 44918
rect 195432 44678 195508 44886
rect 195094 44614 195095 44646
rect 195029 44613 195095 44614
rect 195432 44614 195438 44678
rect 195502 44614 195508 44678
rect 195432 44608 195508 44614
rect 196384 44886 196390 44918
rect 196454 44918 196455 44950
rect 196797 44950 196863 44951
rect 196797 44918 196798 44950
rect 196454 44886 196460 44918
rect 196384 44678 196460 44886
rect 196384 44614 196390 44678
rect 196454 44614 196460 44678
rect 196384 44608 196460 44614
rect 196792 44886 196798 44918
rect 196862 44918 196863 44950
rect 196862 44886 196868 44918
rect 196792 44678 196868 44886
rect 196792 44614 196798 44678
rect 196862 44614 196868 44678
rect 196792 44608 196868 44614
rect 21760 44542 21836 44548
rect 21760 44478 21766 44542
rect 21830 44478 21836 44542
rect 21760 44270 21836 44478
rect 21760 44238 21766 44270
rect 21765 44206 21766 44238
rect 21830 44238 21836 44270
rect 22168 44542 22244 44548
rect 22168 44478 22174 44542
rect 22238 44478 22244 44542
rect 22168 44270 22244 44478
rect 22168 44238 22174 44270
rect 21830 44206 21831 44238
rect 21765 44205 21831 44206
rect 22173 44206 22174 44238
rect 22238 44238 22244 44270
rect 22576 44542 22652 44548
rect 22576 44478 22582 44542
rect 22646 44478 22652 44542
rect 22989 44542 23055 44543
rect 22989 44510 22990 44542
rect 22576 44270 22652 44478
rect 22576 44238 22582 44270
rect 22238 44206 22239 44238
rect 22173 44205 22239 44206
rect 22581 44206 22582 44238
rect 22646 44238 22652 44270
rect 22984 44478 22990 44510
rect 23054 44510 23055 44542
rect 23528 44542 23604 44548
rect 23054 44478 23060 44510
rect 22984 44270 23060 44478
rect 22646 44206 22647 44238
rect 22581 44205 22647 44206
rect 22984 44206 22990 44270
rect 23054 44206 23060 44270
rect 23528 44478 23534 44542
rect 23598 44478 23604 44542
rect 195165 44542 195231 44543
rect 195165 44510 195166 44542
rect 23528 44270 23604 44478
rect 23528 44238 23534 44270
rect 22984 44200 23060 44206
rect 23533 44206 23534 44238
rect 23598 44238 23604 44270
rect 195160 44478 195166 44510
rect 195230 44510 195231 44542
rect 195568 44542 195644 44548
rect 195230 44478 195236 44510
rect 195160 44270 195236 44478
rect 23598 44206 23599 44238
rect 23533 44205 23599 44206
rect 195160 44206 195166 44270
rect 195230 44206 195236 44270
rect 195568 44478 195574 44542
rect 195638 44478 195644 44542
rect 195568 44270 195644 44478
rect 195568 44238 195574 44270
rect 195160 44200 195236 44206
rect 195573 44206 195574 44238
rect 195638 44238 195644 44270
rect 196248 44542 196324 44548
rect 196248 44478 196254 44542
rect 196318 44478 196324 44542
rect 196661 44542 196727 44543
rect 196661 44510 196662 44542
rect 196248 44270 196324 44478
rect 196248 44238 196254 44270
rect 195638 44206 195639 44238
rect 195573 44205 195639 44206
rect 196253 44206 196254 44238
rect 196318 44238 196324 44270
rect 196656 44478 196662 44510
rect 196726 44510 196727 44542
rect 196726 44478 196732 44510
rect 196656 44270 196732 44478
rect 196318 44206 196319 44238
rect 196253 44205 196319 44206
rect 196656 44206 196662 44270
rect 196726 44206 196732 44270
rect 196656 44200 196732 44206
rect 217464 44270 217812 45974
rect 217464 44206 217470 44270
rect 217534 44206 217812 44270
rect 22440 44134 22516 44140
rect 22440 44070 22446 44134
rect 22510 44070 22516 44134
rect 23125 44134 23191 44135
rect 23125 44102 23126 44134
rect 22440 43862 22516 44070
rect 22440 43830 22446 43862
rect 22445 43798 22446 43830
rect 22510 43830 22516 43862
rect 23120 44070 23126 44102
rect 23190 44102 23191 44134
rect 23533 44134 23599 44135
rect 23533 44102 23534 44134
rect 23190 44070 23196 44102
rect 23120 43862 23196 44070
rect 22510 43798 22511 43830
rect 22445 43797 22511 43798
rect 23120 43798 23126 43862
rect 23190 43798 23196 43862
rect 23120 43792 23196 43798
rect 23528 44070 23534 44102
rect 23598 44102 23599 44134
rect 195024 44134 195100 44140
rect 23598 44070 23604 44102
rect 23528 43862 23604 44070
rect 23528 43798 23534 43862
rect 23598 43798 23604 43862
rect 195024 44070 195030 44134
rect 195094 44070 195100 44134
rect 195573 44134 195639 44135
rect 195573 44102 195574 44134
rect 195024 43862 195100 44070
rect 195024 43830 195030 43862
rect 23528 43792 23604 43798
rect 195029 43798 195030 43830
rect 195094 43830 195100 43862
rect 195568 44070 195574 44102
rect 195638 44102 195639 44134
rect 195976 44134 196052 44140
rect 195638 44070 195644 44102
rect 195568 43862 195644 44070
rect 195094 43798 195095 43830
rect 195029 43797 195095 43798
rect 195568 43798 195574 43862
rect 195638 43798 195644 43862
rect 195976 44070 195982 44134
rect 196046 44070 196052 44134
rect 195976 43862 196052 44070
rect 195976 43830 195982 43862
rect 195568 43792 195644 43798
rect 195981 43798 195982 43830
rect 196046 43830 196052 43862
rect 196384 44134 196460 44140
rect 196384 44070 196390 44134
rect 196454 44070 196460 44134
rect 196384 43862 196460 44070
rect 196384 43830 196390 43862
rect 196046 43798 196047 43830
rect 195981 43797 196047 43798
rect 196389 43798 196390 43830
rect 196454 43830 196460 43862
rect 196454 43798 196455 43830
rect 196389 43797 196455 43798
rect 22989 43726 23055 43727
rect 22989 43694 22990 43726
rect 22984 43662 22990 43694
rect 23054 43694 23055 43726
rect 23397 43726 23463 43727
rect 23397 43694 23398 43726
rect 23054 43662 23060 43694
rect 22984 43454 23060 43662
rect 22984 43390 22990 43454
rect 23054 43390 23060 43454
rect 22984 43384 23060 43390
rect 23392 43662 23398 43694
rect 23462 43694 23463 43726
rect 195029 43726 195095 43727
rect 195029 43694 195030 43726
rect 23462 43662 23468 43694
rect 23392 43454 23468 43662
rect 195024 43662 195030 43694
rect 195094 43694 195095 43726
rect 195573 43726 195639 43727
rect 195573 43694 195574 43726
rect 195094 43662 195100 43694
rect 23392 43390 23398 43454
rect 23462 43390 23468 43454
rect 190133 43454 190199 43455
rect 190133 43422 190134 43454
rect 23392 43384 23468 43390
rect 190128 43390 190134 43422
rect 190198 43422 190199 43454
rect 195024 43454 195100 43662
rect 190198 43390 190204 43422
rect 22440 43318 22516 43324
rect 22440 43254 22446 43318
rect 22510 43254 22516 43318
rect 21765 43046 21831 43047
rect 21765 43014 21766 43046
rect 14688 42846 14694 42910
rect 14758 42846 14764 42910
rect 14688 42840 14764 42846
rect 21760 42982 21766 43014
rect 21830 43014 21831 43046
rect 22440 43046 22516 43254
rect 28293 43182 28359 43183
rect 28293 43150 28294 43182
rect 22440 43014 22446 43046
rect 21830 42982 21836 43014
rect 14552 41518 14558 41550
rect 14557 41486 14558 41518
rect 14622 41518 14628 41550
rect 14688 42774 14764 42780
rect 14688 42710 14694 42774
rect 14758 42710 14764 42774
rect 14622 41486 14623 41518
rect 14557 41485 14623 41486
rect 14557 41278 14623 41279
rect 14557 41246 14558 41278
rect 952 40806 1230 40870
rect 1294 40806 1300 40870
rect 952 39238 1300 40806
rect 952 39174 1230 39238
rect 1294 39174 1300 39238
rect 952 37470 1300 39174
rect 14552 41214 14558 41246
rect 14622 41246 14623 41278
rect 14622 41214 14628 41246
rect 14552 38694 14628 41214
rect 14688 40054 14764 42710
rect 21760 42774 21836 42982
rect 22445 42982 22446 43014
rect 22510 43014 22516 43046
rect 28288 43118 28294 43150
rect 28358 43150 28359 43182
rect 190128 43182 190204 43390
rect 195024 43390 195030 43454
rect 195094 43390 195100 43454
rect 195024 43384 195100 43390
rect 195568 43662 195574 43694
rect 195638 43694 195639 43726
rect 195638 43662 195644 43694
rect 195568 43454 195644 43662
rect 195568 43390 195574 43454
rect 195638 43390 195644 43454
rect 195568 43384 195644 43390
rect 196389 43318 196455 43319
rect 196389 43286 196390 43318
rect 196384 43254 196390 43286
rect 196454 43286 196455 43318
rect 196454 43254 196460 43286
rect 28358 43118 28364 43150
rect 22510 42982 22511 43014
rect 22445 42981 22511 42982
rect 21760 42710 21766 42774
rect 21830 42710 21836 42774
rect 21760 42704 21836 42710
rect 22440 42910 22516 42916
rect 22440 42846 22446 42910
rect 22510 42846 22516 42910
rect 21760 42638 21836 42644
rect 21760 42574 21766 42638
rect 21830 42574 21836 42638
rect 22440 42638 22516 42846
rect 28288 42910 28364 43118
rect 190128 43118 190134 43182
rect 190198 43118 190204 43182
rect 190128 43112 190204 43118
rect 190264 43182 190340 43188
rect 190264 43118 190270 43182
rect 190334 43118 190340 43182
rect 28288 42846 28294 42910
rect 28358 42846 28364 42910
rect 28288 42840 28364 42846
rect 28560 42910 28636 42916
rect 28560 42846 28566 42910
rect 28630 42846 28636 42910
rect 190264 42910 190340 43118
rect 196384 43046 196460 43254
rect 196384 42982 196390 43046
rect 196454 42982 196460 43046
rect 196661 43046 196727 43047
rect 196661 43014 196662 43046
rect 196384 42976 196460 42982
rect 196656 42982 196662 43014
rect 196726 43014 196727 43046
rect 196726 42982 196732 43014
rect 190264 42878 190270 42910
rect 28288 42774 28364 42780
rect 28288 42710 28294 42774
rect 28358 42710 28364 42774
rect 22440 42606 22446 42638
rect 21760 42366 21836 42574
rect 22445 42574 22446 42606
rect 22510 42606 22516 42638
rect 22717 42638 22783 42639
rect 22717 42606 22718 42638
rect 22510 42574 22511 42606
rect 22445 42573 22511 42574
rect 22712 42574 22718 42606
rect 22782 42606 22783 42638
rect 22782 42574 22788 42606
rect 21760 42334 21766 42366
rect 21765 42302 21766 42334
rect 21830 42334 21836 42366
rect 22712 42366 22788 42574
rect 28288 42502 28364 42710
rect 28288 42470 28294 42502
rect 28293 42438 28294 42470
rect 28358 42470 28364 42502
rect 28560 42502 28636 42846
rect 190269 42846 190270 42878
rect 190334 42878 190340 42910
rect 190334 42846 190335 42878
rect 190269 42845 190335 42846
rect 190269 42774 190335 42775
rect 190269 42742 190270 42774
rect 28560 42470 28566 42502
rect 28358 42438 28359 42470
rect 28293 42437 28359 42438
rect 28565 42438 28566 42470
rect 28630 42470 28636 42502
rect 190264 42710 190270 42742
rect 190334 42742 190335 42774
rect 196656 42774 196732 42982
rect 190334 42710 190340 42742
rect 190264 42502 190340 42710
rect 196656 42710 196662 42774
rect 196726 42710 196732 42774
rect 196656 42704 196732 42710
rect 28630 42438 28631 42470
rect 28565 42437 28631 42438
rect 190264 42438 190270 42502
rect 190334 42438 190340 42502
rect 190264 42432 190340 42438
rect 196384 42638 196460 42644
rect 196384 42574 196390 42638
rect 196454 42574 196460 42638
rect 21830 42302 21831 42334
rect 21765 42301 21831 42302
rect 22712 42302 22718 42366
rect 22782 42302 22788 42366
rect 196384 42366 196460 42574
rect 196384 42334 196390 42366
rect 22712 42296 22788 42302
rect 196389 42302 196390 42334
rect 196454 42334 196460 42366
rect 196656 42638 196732 42644
rect 196656 42574 196662 42638
rect 196726 42574 196732 42638
rect 196656 42366 196732 42574
rect 196656 42334 196662 42366
rect 196454 42302 196455 42334
rect 196389 42301 196455 42302
rect 196661 42302 196662 42334
rect 196726 42334 196732 42366
rect 217464 42638 217812 44206
rect 217464 42574 217470 42638
rect 217534 42574 217812 42638
rect 196726 42302 196727 42334
rect 196661 42301 196727 42302
rect 21765 42230 21831 42231
rect 21765 42198 21766 42230
rect 21760 42166 21766 42198
rect 21830 42198 21831 42230
rect 23120 42230 23196 42236
rect 21830 42166 21836 42198
rect 21760 41958 21836 42166
rect 21760 41894 21766 41958
rect 21830 41894 21836 41958
rect 23120 42166 23126 42230
rect 23190 42166 23196 42230
rect 23533 42230 23599 42231
rect 23533 42198 23534 42230
rect 23120 41958 23196 42166
rect 23120 41926 23126 41958
rect 21760 41888 21836 41894
rect 23125 41894 23126 41926
rect 23190 41926 23196 41958
rect 23528 42166 23534 42198
rect 23598 42198 23599 42230
rect 195165 42230 195231 42231
rect 195165 42198 195166 42230
rect 23598 42166 23604 42198
rect 23528 41958 23604 42166
rect 23190 41894 23191 41926
rect 23125 41893 23191 41894
rect 23528 41894 23534 41958
rect 23598 41894 23604 41958
rect 23528 41888 23604 41894
rect 195160 42166 195166 42198
rect 195230 42198 195231 42230
rect 195568 42230 195644 42236
rect 195230 42166 195236 42198
rect 195160 41958 195236 42166
rect 195160 41894 195166 41958
rect 195230 41894 195236 41958
rect 195568 42166 195574 42230
rect 195638 42166 195644 42230
rect 196661 42230 196727 42231
rect 196661 42198 196662 42230
rect 195568 41958 195644 42166
rect 195568 41926 195574 41958
rect 195160 41888 195236 41894
rect 195573 41894 195574 41926
rect 195638 41926 195644 41958
rect 196656 42166 196662 42198
rect 196726 42198 196727 42230
rect 196726 42166 196732 42198
rect 196656 41958 196732 42166
rect 195638 41894 195639 41926
rect 195573 41893 195639 41894
rect 196656 41894 196662 41958
rect 196726 41894 196732 41958
rect 196656 41888 196732 41894
rect 21901 41822 21967 41823
rect 21901 41790 21902 41822
rect 21896 41758 21902 41790
rect 21966 41790 21967 41822
rect 22445 41822 22511 41823
rect 22445 41790 22446 41822
rect 21966 41758 21972 41790
rect 21896 41550 21972 41758
rect 21896 41486 21902 41550
rect 21966 41486 21972 41550
rect 21896 41480 21972 41486
rect 22440 41758 22446 41790
rect 22510 41790 22511 41822
rect 22712 41822 22788 41828
rect 22510 41758 22516 41790
rect 22440 41550 22516 41758
rect 22440 41486 22446 41550
rect 22510 41486 22516 41550
rect 22712 41758 22718 41822
rect 22782 41758 22788 41822
rect 22989 41822 23055 41823
rect 22989 41790 22990 41822
rect 22712 41550 22788 41758
rect 22712 41518 22718 41550
rect 22440 41480 22516 41486
rect 22717 41486 22718 41518
rect 22782 41518 22788 41550
rect 22984 41758 22990 41790
rect 23054 41790 23055 41822
rect 23392 41822 23468 41828
rect 23054 41758 23060 41790
rect 22984 41550 23060 41758
rect 22782 41486 22783 41518
rect 22717 41485 22783 41486
rect 22984 41486 22990 41550
rect 23054 41486 23060 41550
rect 23392 41758 23398 41822
rect 23462 41758 23468 41822
rect 23392 41550 23468 41758
rect 195024 41822 195100 41828
rect 195024 41758 195030 41822
rect 195094 41758 195100 41822
rect 195437 41822 195503 41823
rect 195437 41790 195438 41822
rect 23392 41518 23398 41550
rect 22984 41480 23060 41486
rect 23397 41486 23398 41518
rect 23462 41518 23468 41550
rect 28288 41550 28364 41556
rect 23462 41486 23463 41518
rect 23397 41485 23463 41486
rect 28288 41486 28294 41550
rect 28358 41486 28364 41550
rect 21901 41414 21967 41415
rect 21901 41382 21902 41414
rect 21896 41350 21902 41382
rect 21966 41382 21967 41414
rect 22309 41414 22375 41415
rect 22309 41382 22310 41414
rect 21966 41350 21972 41382
rect 21896 41142 21972 41350
rect 21896 41078 21902 41142
rect 21966 41078 21972 41142
rect 21896 41072 21972 41078
rect 22304 41350 22310 41382
rect 22374 41382 22375 41414
rect 23125 41414 23191 41415
rect 23125 41382 23126 41414
rect 22374 41350 22380 41382
rect 22304 41142 22380 41350
rect 22304 41078 22310 41142
rect 22374 41078 22380 41142
rect 22304 41072 22380 41078
rect 23120 41350 23126 41382
rect 23190 41382 23191 41414
rect 23397 41414 23463 41415
rect 23397 41382 23398 41414
rect 23190 41350 23196 41382
rect 23120 41142 23196 41350
rect 23120 41078 23126 41142
rect 23190 41078 23196 41142
rect 23120 41072 23196 41078
rect 23392 41350 23398 41382
rect 23462 41382 23463 41414
rect 23462 41350 23468 41382
rect 23392 41142 23468 41350
rect 28288 41278 28364 41486
rect 28288 41246 28294 41278
rect 28293 41214 28294 41246
rect 28358 41246 28364 41278
rect 190128 41550 190204 41556
rect 190128 41486 190134 41550
rect 190198 41486 190204 41550
rect 195024 41550 195100 41758
rect 195024 41518 195030 41550
rect 190128 41278 190204 41486
rect 195029 41486 195030 41518
rect 195094 41518 195100 41550
rect 195432 41758 195438 41790
rect 195502 41790 195503 41822
rect 196792 41822 196868 41828
rect 195502 41758 195508 41790
rect 195432 41550 195508 41758
rect 195094 41486 195095 41518
rect 195029 41485 195095 41486
rect 195432 41486 195438 41550
rect 195502 41486 195508 41550
rect 196792 41758 196798 41822
rect 196862 41758 196868 41822
rect 196792 41550 196868 41758
rect 196792 41518 196798 41550
rect 195432 41480 195508 41486
rect 196797 41486 196798 41518
rect 196862 41518 196868 41550
rect 196862 41486 196863 41518
rect 196797 41485 196863 41486
rect 190128 41246 190134 41278
rect 28358 41214 28359 41246
rect 28293 41213 28359 41214
rect 190133 41214 190134 41246
rect 190198 41246 190204 41278
rect 195160 41414 195236 41420
rect 195160 41350 195166 41414
rect 195230 41350 195236 41414
rect 195573 41414 195639 41415
rect 195573 41382 195574 41414
rect 190198 41214 190199 41246
rect 190133 41213 190199 41214
rect 23392 41078 23398 41142
rect 23462 41078 23468 41142
rect 195160 41142 195236 41350
rect 195160 41110 195166 41142
rect 23392 41072 23468 41078
rect 195165 41078 195166 41110
rect 195230 41110 195236 41142
rect 195568 41350 195574 41382
rect 195638 41382 195639 41414
rect 195840 41414 195916 41420
rect 195638 41350 195644 41382
rect 195568 41142 195644 41350
rect 195230 41078 195231 41110
rect 195165 41077 195231 41078
rect 195568 41078 195574 41142
rect 195638 41078 195644 41142
rect 195840 41350 195846 41414
rect 195910 41350 195916 41414
rect 196389 41414 196455 41415
rect 196389 41382 196390 41414
rect 195840 41142 195916 41350
rect 195840 41110 195846 41142
rect 195568 41072 195644 41078
rect 195845 41078 195846 41110
rect 195910 41110 195916 41142
rect 196384 41350 196390 41382
rect 196454 41382 196455 41414
rect 196797 41414 196863 41415
rect 196797 41382 196798 41414
rect 196454 41350 196460 41382
rect 196384 41142 196460 41350
rect 195910 41078 195911 41110
rect 195845 41077 195911 41078
rect 196384 41078 196390 41142
rect 196454 41078 196460 41142
rect 196384 41072 196460 41078
rect 196792 41350 196798 41382
rect 196862 41382 196863 41414
rect 196862 41350 196868 41382
rect 196792 41142 196868 41350
rect 196792 41078 196798 41142
rect 196862 41078 196868 41142
rect 196792 41072 196868 41078
rect 21896 41006 21972 41012
rect 21896 40942 21902 41006
rect 21966 40942 21972 41006
rect 22581 41006 22647 41007
rect 22581 40974 22582 41006
rect 21896 40734 21972 40942
rect 21896 40702 21902 40734
rect 21901 40670 21902 40702
rect 21966 40702 21972 40734
rect 22576 40942 22582 40974
rect 22646 40974 22647 41006
rect 22989 41006 23055 41007
rect 22989 40974 22990 41006
rect 22646 40942 22652 40974
rect 22576 40734 22652 40942
rect 21966 40670 21967 40702
rect 21901 40669 21967 40670
rect 22576 40670 22582 40734
rect 22646 40670 22652 40734
rect 22576 40664 22652 40670
rect 22984 40942 22990 40974
rect 23054 40974 23055 41006
rect 23533 41006 23599 41007
rect 23533 40974 23534 41006
rect 23054 40942 23060 40974
rect 22984 40734 23060 40942
rect 22984 40670 22990 40734
rect 23054 40670 23060 40734
rect 22984 40664 23060 40670
rect 23528 40942 23534 40974
rect 23598 40974 23599 41006
rect 195165 41006 195231 41007
rect 195165 40974 195166 41006
rect 23598 40942 23604 40974
rect 23528 40734 23604 40942
rect 23528 40670 23534 40734
rect 23598 40670 23604 40734
rect 23528 40664 23604 40670
rect 195160 40942 195166 40974
rect 195230 40974 195231 41006
rect 195432 41006 195508 41012
rect 195230 40942 195236 40974
rect 195160 40734 195236 40942
rect 195160 40670 195166 40734
rect 195230 40670 195236 40734
rect 195432 40942 195438 41006
rect 195502 40942 195508 41006
rect 196661 41006 196727 41007
rect 196661 40974 196662 41006
rect 195432 40734 195508 40942
rect 195432 40702 195438 40734
rect 195160 40664 195236 40670
rect 195437 40670 195438 40702
rect 195502 40702 195508 40734
rect 196656 40942 196662 40974
rect 196726 40974 196727 41006
rect 196726 40942 196732 40974
rect 196656 40734 196732 40942
rect 195502 40670 195503 40702
rect 195437 40669 195503 40670
rect 196656 40670 196662 40734
rect 196726 40670 196732 40734
rect 196656 40664 196732 40670
rect 217464 40870 217812 42574
rect 217464 40806 217470 40870
rect 217534 40806 217812 40870
rect 21901 40598 21967 40599
rect 21901 40566 21902 40598
rect 21896 40534 21902 40566
rect 21966 40566 21967 40598
rect 22309 40598 22375 40599
rect 22309 40566 22310 40598
rect 21966 40534 21972 40566
rect 21896 40326 21972 40534
rect 21896 40262 21902 40326
rect 21966 40262 21972 40326
rect 21896 40256 21972 40262
rect 22304 40534 22310 40566
rect 22374 40566 22375 40598
rect 23120 40598 23196 40604
rect 22374 40534 22380 40566
rect 22304 40326 22380 40534
rect 22304 40262 22310 40326
rect 22374 40262 22380 40326
rect 23120 40534 23126 40598
rect 23190 40534 23196 40598
rect 23120 40326 23196 40534
rect 23120 40294 23126 40326
rect 22304 40256 22380 40262
rect 23125 40262 23126 40294
rect 23190 40294 23196 40326
rect 23392 40598 23468 40604
rect 23392 40534 23398 40598
rect 23462 40534 23468 40598
rect 23392 40326 23468 40534
rect 23392 40294 23398 40326
rect 23190 40262 23191 40294
rect 23125 40261 23191 40262
rect 23397 40262 23398 40294
rect 23462 40294 23468 40326
rect 195024 40598 195100 40604
rect 195024 40534 195030 40598
rect 195094 40534 195100 40598
rect 195437 40598 195503 40599
rect 195437 40566 195438 40598
rect 195024 40326 195100 40534
rect 195024 40294 195030 40326
rect 23462 40262 23463 40294
rect 23397 40261 23463 40262
rect 195029 40262 195030 40294
rect 195094 40294 195100 40326
rect 195432 40534 195438 40566
rect 195502 40566 195503 40598
rect 196389 40598 196455 40599
rect 196389 40566 196390 40598
rect 195502 40534 195508 40566
rect 195432 40326 195508 40534
rect 195094 40262 195095 40294
rect 195029 40261 195095 40262
rect 195432 40262 195438 40326
rect 195502 40262 195508 40326
rect 195432 40256 195508 40262
rect 196384 40534 196390 40566
rect 196454 40566 196455 40598
rect 196792 40598 196868 40604
rect 196454 40534 196460 40566
rect 196384 40326 196460 40534
rect 196384 40262 196390 40326
rect 196454 40262 196460 40326
rect 196792 40534 196798 40598
rect 196862 40534 196868 40598
rect 196792 40326 196868 40534
rect 196792 40294 196798 40326
rect 196384 40256 196460 40262
rect 196797 40262 196798 40294
rect 196862 40294 196868 40326
rect 196862 40262 196863 40294
rect 196797 40261 196863 40262
rect 22173 40190 22239 40191
rect 22173 40158 22174 40190
rect 14688 40022 14694 40054
rect 14693 39990 14694 40022
rect 14758 40022 14764 40054
rect 22168 40126 22174 40158
rect 22238 40158 22239 40190
rect 22445 40190 22511 40191
rect 22445 40158 22446 40190
rect 22238 40126 22244 40158
rect 14758 39990 14759 40022
rect 14693 39989 14759 39990
rect 14552 38630 14558 38694
rect 14622 38630 14628 38694
rect 14552 38624 14628 38630
rect 14688 39918 14764 39924
rect 14688 39854 14694 39918
rect 14758 39854 14764 39918
rect 952 37406 1230 37470
rect 1294 37406 1300 37470
rect 952 35702 1300 37406
rect 14552 38558 14628 38564
rect 14552 38494 14558 38558
rect 14622 38494 14628 38558
rect 14552 35838 14628 38494
rect 14688 37198 14764 39854
rect 22168 39918 22244 40126
rect 22168 39854 22174 39918
rect 22238 39854 22244 39918
rect 22168 39848 22244 39854
rect 22440 40126 22446 40158
rect 22510 40158 22511 40190
rect 22989 40190 23055 40191
rect 22989 40158 22990 40190
rect 22510 40126 22516 40158
rect 22440 39918 22516 40126
rect 22440 39854 22446 39918
rect 22510 39854 22516 39918
rect 22440 39848 22516 39854
rect 22984 40126 22990 40158
rect 23054 40158 23055 40190
rect 23533 40190 23599 40191
rect 23533 40158 23534 40190
rect 23054 40126 23060 40158
rect 22984 39918 23060 40126
rect 22984 39854 22990 39918
rect 23054 39854 23060 39918
rect 22984 39848 23060 39854
rect 23528 40126 23534 40158
rect 23598 40158 23599 40190
rect 195160 40190 195236 40196
rect 23598 40126 23604 40158
rect 23528 39918 23604 40126
rect 195160 40126 195166 40190
rect 195230 40126 195236 40190
rect 23528 39854 23534 39918
rect 23598 39854 23604 39918
rect 23528 39848 23604 39854
rect 28288 40054 28364 40060
rect 28288 39990 28294 40054
rect 28358 39990 28364 40054
rect 190133 40054 190199 40055
rect 190133 40022 190134 40054
rect 22984 39782 23060 39788
rect 22984 39718 22990 39782
rect 23054 39718 23060 39782
rect 22984 39510 23060 39718
rect 22984 39478 22990 39510
rect 22989 39446 22990 39478
rect 23054 39478 23060 39510
rect 23392 39782 23468 39788
rect 23392 39718 23398 39782
rect 23462 39718 23468 39782
rect 28288 39782 28364 39990
rect 28288 39750 28294 39782
rect 23392 39510 23468 39718
rect 28293 39718 28294 39750
rect 28358 39750 28364 39782
rect 190128 39990 190134 40022
rect 190198 40022 190199 40054
rect 190198 39990 190204 40022
rect 190128 39782 190204 39990
rect 195160 39918 195236 40126
rect 195160 39886 195166 39918
rect 195165 39854 195166 39886
rect 195230 39886 195236 39918
rect 195568 40190 195644 40196
rect 195568 40126 195574 40190
rect 195638 40126 195644 40190
rect 195568 39918 195644 40126
rect 195568 39886 195574 39918
rect 195230 39854 195231 39886
rect 195165 39853 195231 39854
rect 195573 39854 195574 39886
rect 195638 39886 195644 39918
rect 195840 40190 195916 40196
rect 195840 40126 195846 40190
rect 195910 40126 195916 40190
rect 196253 40190 196319 40191
rect 196253 40158 196254 40190
rect 195840 39918 195916 40126
rect 195840 39886 195846 39918
rect 195638 39854 195639 39886
rect 195573 39853 195639 39854
rect 195845 39854 195846 39886
rect 195910 39886 195916 39918
rect 196248 40126 196254 40158
rect 196318 40158 196319 40190
rect 196318 40126 196324 40158
rect 196248 39918 196324 40126
rect 195910 39854 195911 39886
rect 195845 39853 195911 39854
rect 196248 39854 196254 39918
rect 196318 39854 196324 39918
rect 196248 39848 196324 39854
rect 28358 39718 28359 39750
rect 28293 39717 28359 39718
rect 190128 39718 190134 39782
rect 190198 39718 190204 39782
rect 195165 39782 195231 39783
rect 195165 39750 195166 39782
rect 190128 39712 190204 39718
rect 195160 39718 195166 39750
rect 195230 39750 195231 39782
rect 195573 39782 195639 39783
rect 195573 39750 195574 39782
rect 195230 39718 195236 39750
rect 23392 39478 23398 39510
rect 23054 39446 23055 39478
rect 22989 39445 23055 39446
rect 23397 39446 23398 39478
rect 23462 39478 23468 39510
rect 195160 39510 195236 39718
rect 23462 39446 23463 39478
rect 23397 39445 23463 39446
rect 195160 39446 195166 39510
rect 195230 39446 195236 39510
rect 195160 39440 195236 39446
rect 195568 39718 195574 39750
rect 195638 39750 195639 39782
rect 195638 39718 195644 39750
rect 195568 39510 195644 39718
rect 195568 39446 195574 39510
rect 195638 39446 195644 39510
rect 195568 39440 195644 39446
rect 22168 39374 22244 39380
rect 22168 39310 22174 39374
rect 22238 39310 22244 39374
rect 22445 39374 22511 39375
rect 22445 39342 22446 39374
rect 21765 39102 21831 39103
rect 21765 39070 21766 39102
rect 21760 39038 21766 39070
rect 21830 39070 21831 39102
rect 22168 39102 22244 39310
rect 22168 39070 22174 39102
rect 21830 39038 21836 39070
rect 21760 38830 21836 39038
rect 22173 39038 22174 39070
rect 22238 39070 22244 39102
rect 22440 39310 22446 39342
rect 22510 39342 22511 39374
rect 22989 39374 23055 39375
rect 22989 39342 22990 39374
rect 22510 39310 22516 39342
rect 22440 39102 22516 39310
rect 22238 39038 22239 39070
rect 22173 39037 22239 39038
rect 22440 39038 22446 39102
rect 22510 39038 22516 39102
rect 22440 39032 22516 39038
rect 22984 39310 22990 39342
rect 23054 39342 23055 39374
rect 23397 39374 23463 39375
rect 23397 39342 23398 39374
rect 23054 39310 23060 39342
rect 22984 39102 23060 39310
rect 22984 39038 22990 39102
rect 23054 39038 23060 39102
rect 22984 39032 23060 39038
rect 23392 39310 23398 39342
rect 23462 39342 23463 39374
rect 195160 39374 195236 39380
rect 23462 39310 23468 39342
rect 23392 39102 23468 39310
rect 23392 39038 23398 39102
rect 23462 39038 23468 39102
rect 195160 39310 195166 39374
rect 195230 39310 195236 39374
rect 195160 39102 195236 39310
rect 195160 39070 195166 39102
rect 23392 39032 23468 39038
rect 195165 39038 195166 39070
rect 195230 39070 195236 39102
rect 195432 39374 195508 39380
rect 195432 39310 195438 39374
rect 195502 39310 195508 39374
rect 195432 39102 195508 39310
rect 195432 39070 195438 39102
rect 195230 39038 195231 39070
rect 195165 39037 195231 39038
rect 195437 39038 195438 39070
rect 195502 39070 195508 39102
rect 196248 39374 196324 39380
rect 196248 39310 196254 39374
rect 196318 39310 196324 39374
rect 196248 39102 196324 39310
rect 196248 39070 196254 39102
rect 195502 39038 195503 39070
rect 195437 39037 195503 39038
rect 196253 39038 196254 39070
rect 196318 39070 196324 39102
rect 196656 39102 196732 39108
rect 196318 39038 196319 39070
rect 196253 39037 196319 39038
rect 196656 39038 196662 39102
rect 196726 39038 196732 39102
rect 190133 38966 190199 38967
rect 190133 38934 190134 38966
rect 190128 38902 190134 38934
rect 190198 38934 190199 38966
rect 190198 38902 190204 38934
rect 21760 38766 21766 38830
rect 21830 38766 21836 38830
rect 21760 38760 21836 38766
rect 28288 38830 28364 38836
rect 28288 38766 28294 38830
rect 28358 38766 28364 38830
rect 21896 38694 21972 38700
rect 21896 38630 21902 38694
rect 21966 38630 21972 38694
rect 21896 38422 21972 38630
rect 21896 38390 21902 38422
rect 21901 38358 21902 38390
rect 21966 38390 21972 38422
rect 22576 38694 22652 38700
rect 22576 38630 22582 38694
rect 22646 38630 22652 38694
rect 22576 38422 22652 38630
rect 28288 38558 28364 38766
rect 28288 38526 28294 38558
rect 28293 38494 28294 38526
rect 28358 38526 28364 38558
rect 190128 38558 190204 38902
rect 190269 38830 190335 38831
rect 190269 38798 190270 38830
rect 28358 38494 28359 38526
rect 28293 38493 28359 38494
rect 190128 38494 190134 38558
rect 190198 38494 190204 38558
rect 190128 38488 190204 38494
rect 190264 38766 190270 38798
rect 190334 38798 190335 38830
rect 196656 38830 196732 39038
rect 196656 38798 196662 38830
rect 190334 38766 190340 38798
rect 190264 38558 190340 38766
rect 196661 38766 196662 38798
rect 196726 38798 196732 38830
rect 217464 39102 217812 40806
rect 217464 39038 217470 39102
rect 217534 39038 217812 39102
rect 196726 38766 196727 38798
rect 196661 38765 196727 38766
rect 195845 38694 195911 38695
rect 195845 38662 195846 38694
rect 190264 38494 190270 38558
rect 190334 38494 190340 38558
rect 190264 38488 190340 38494
rect 195840 38630 195846 38662
rect 195910 38662 195911 38694
rect 196661 38694 196727 38695
rect 196661 38662 196662 38694
rect 195910 38630 195916 38662
rect 22576 38390 22582 38422
rect 21966 38358 21967 38390
rect 21901 38357 21967 38358
rect 22581 38358 22582 38390
rect 22646 38390 22652 38422
rect 195840 38422 195916 38630
rect 22646 38358 22647 38390
rect 22581 38357 22647 38358
rect 195840 38358 195846 38422
rect 195910 38358 195916 38422
rect 195840 38352 195916 38358
rect 196656 38630 196662 38662
rect 196726 38662 196727 38694
rect 196726 38630 196732 38662
rect 196656 38422 196732 38630
rect 196656 38358 196662 38422
rect 196726 38358 196732 38422
rect 196656 38352 196732 38358
rect 21901 38286 21967 38287
rect 21901 38254 21902 38286
rect 21896 38222 21902 38254
rect 21966 38254 21967 38286
rect 22984 38286 23060 38292
rect 21966 38222 21972 38254
rect 21896 38014 21972 38222
rect 21896 37950 21902 38014
rect 21966 37950 21972 38014
rect 22984 38222 22990 38286
rect 23054 38222 23060 38286
rect 23397 38286 23463 38287
rect 23397 38254 23398 38286
rect 22984 38014 23060 38222
rect 22984 37982 22990 38014
rect 21896 37944 21972 37950
rect 22989 37950 22990 37982
rect 23054 37982 23060 38014
rect 23392 38222 23398 38254
rect 23462 38254 23463 38286
rect 195160 38286 195236 38292
rect 23462 38222 23468 38254
rect 23392 38014 23468 38222
rect 23054 37950 23055 37982
rect 22989 37949 23055 37950
rect 23392 37950 23398 38014
rect 23462 37950 23468 38014
rect 195160 38222 195166 38286
rect 195230 38222 195236 38286
rect 195160 38014 195236 38222
rect 195160 37982 195166 38014
rect 23392 37944 23468 37950
rect 195165 37950 195166 37982
rect 195230 37982 195236 38014
rect 195432 38286 195508 38292
rect 195432 38222 195438 38286
rect 195502 38222 195508 38286
rect 196797 38286 196863 38287
rect 196797 38254 196798 38286
rect 195432 38014 195508 38222
rect 195432 37982 195438 38014
rect 195230 37950 195231 37982
rect 195165 37949 195231 37950
rect 195437 37950 195438 37982
rect 195502 37982 195508 38014
rect 196792 38222 196798 38254
rect 196862 38254 196863 38286
rect 196862 38222 196868 38254
rect 196792 38014 196868 38222
rect 195502 37950 195503 37982
rect 195437 37949 195503 37950
rect 196792 37950 196798 38014
rect 196862 37950 196868 38014
rect 196792 37944 196868 37950
rect 21760 37878 21836 37884
rect 21760 37814 21766 37878
rect 21830 37814 21836 37878
rect 21760 37606 21836 37814
rect 21760 37574 21766 37606
rect 21765 37542 21766 37574
rect 21830 37574 21836 37606
rect 22168 37878 22244 37884
rect 22168 37814 22174 37878
rect 22238 37814 22244 37878
rect 22581 37878 22647 37879
rect 22581 37846 22582 37878
rect 22168 37606 22244 37814
rect 22168 37574 22174 37606
rect 21830 37542 21831 37574
rect 21765 37541 21831 37542
rect 22173 37542 22174 37574
rect 22238 37574 22244 37606
rect 22576 37814 22582 37846
rect 22646 37846 22647 37878
rect 22989 37878 23055 37879
rect 22989 37846 22990 37878
rect 22646 37814 22652 37846
rect 22576 37606 22652 37814
rect 22238 37542 22239 37574
rect 22173 37541 22239 37542
rect 22576 37542 22582 37606
rect 22646 37542 22652 37606
rect 22576 37536 22652 37542
rect 22984 37814 22990 37846
rect 23054 37846 23055 37878
rect 23528 37878 23604 37884
rect 23054 37814 23060 37846
rect 22984 37606 23060 37814
rect 22984 37542 22990 37606
rect 23054 37542 23060 37606
rect 23528 37814 23534 37878
rect 23598 37814 23604 37878
rect 195165 37878 195231 37879
rect 195165 37846 195166 37878
rect 23528 37606 23604 37814
rect 195160 37814 195166 37846
rect 195230 37846 195231 37878
rect 195437 37878 195503 37879
rect 195437 37846 195438 37878
rect 195230 37814 195236 37846
rect 23528 37574 23534 37606
rect 22984 37536 23060 37542
rect 23533 37542 23534 37574
rect 23598 37574 23604 37606
rect 190133 37606 190199 37607
rect 190133 37574 190134 37606
rect 23598 37542 23599 37574
rect 23533 37541 23599 37542
rect 190128 37542 190134 37574
rect 190198 37574 190199 37606
rect 195160 37606 195236 37814
rect 190198 37542 190204 37574
rect 14688 37166 14694 37198
rect 14693 37134 14694 37166
rect 14758 37166 14764 37198
rect 21896 37470 21972 37476
rect 21896 37406 21902 37470
rect 21966 37406 21972 37470
rect 21896 37198 21972 37406
rect 21896 37166 21902 37198
rect 14758 37134 14759 37166
rect 14693 37133 14759 37134
rect 21901 37134 21902 37166
rect 21966 37166 21972 37198
rect 22712 37470 22788 37476
rect 22712 37406 22718 37470
rect 22782 37406 22788 37470
rect 22989 37470 23055 37471
rect 22989 37438 22990 37470
rect 22712 37198 22788 37406
rect 22712 37166 22718 37198
rect 21966 37134 21967 37166
rect 21901 37133 21967 37134
rect 22717 37134 22718 37166
rect 22782 37166 22788 37198
rect 22984 37406 22990 37438
rect 23054 37438 23055 37470
rect 23397 37470 23463 37471
rect 23397 37438 23398 37470
rect 23054 37406 23060 37438
rect 22984 37198 23060 37406
rect 22782 37134 22783 37166
rect 22717 37133 22783 37134
rect 22984 37134 22990 37198
rect 23054 37134 23060 37198
rect 22984 37128 23060 37134
rect 23392 37406 23398 37438
rect 23462 37438 23463 37470
rect 23462 37406 23468 37438
rect 23392 37198 23468 37406
rect 190128 37334 190204 37542
rect 195160 37542 195166 37606
rect 195230 37542 195236 37606
rect 195160 37536 195236 37542
rect 195432 37814 195438 37846
rect 195502 37846 195503 37878
rect 196248 37878 196324 37884
rect 195502 37814 195508 37846
rect 195432 37606 195508 37814
rect 195432 37542 195438 37606
rect 195502 37542 195508 37606
rect 196248 37814 196254 37878
rect 196318 37814 196324 37878
rect 196661 37878 196727 37879
rect 196661 37846 196662 37878
rect 196248 37606 196324 37814
rect 196248 37574 196254 37606
rect 195432 37536 195508 37542
rect 196253 37542 196254 37574
rect 196318 37574 196324 37606
rect 196656 37814 196662 37846
rect 196726 37846 196727 37878
rect 196726 37814 196732 37846
rect 196656 37606 196732 37814
rect 196318 37542 196319 37574
rect 196253 37541 196319 37542
rect 196656 37542 196662 37606
rect 196726 37542 196732 37606
rect 196656 37536 196732 37542
rect 217464 37606 217812 39038
rect 217464 37542 217470 37606
rect 217534 37542 217812 37606
rect 190128 37270 190134 37334
rect 190198 37270 190204 37334
rect 190128 37264 190204 37270
rect 195024 37470 195100 37476
rect 195024 37406 195030 37470
rect 195094 37406 195100 37470
rect 23392 37134 23398 37198
rect 23462 37134 23468 37198
rect 195024 37198 195100 37406
rect 195024 37166 195030 37198
rect 23392 37128 23468 37134
rect 195029 37134 195030 37166
rect 195094 37166 195100 37198
rect 195568 37470 195644 37476
rect 195568 37406 195574 37470
rect 195638 37406 195644 37470
rect 195568 37198 195644 37406
rect 195568 37166 195574 37198
rect 195094 37134 195095 37166
rect 195029 37133 195095 37134
rect 195573 37134 195574 37166
rect 195638 37166 195644 37198
rect 196792 37470 196868 37476
rect 196792 37406 196798 37470
rect 196862 37406 196868 37470
rect 196792 37198 196868 37406
rect 196792 37166 196798 37198
rect 195638 37134 195639 37166
rect 195573 37133 195639 37134
rect 196797 37134 196798 37166
rect 196862 37166 196868 37198
rect 196862 37134 196863 37166
rect 196797 37133 196863 37134
rect 14693 37062 14759 37063
rect 14693 37030 14694 37062
rect 14552 35806 14558 35838
rect 14557 35774 14558 35806
rect 14622 35806 14628 35838
rect 14688 36998 14694 37030
rect 14758 37030 14759 37062
rect 21901 37062 21967 37063
rect 21901 37030 21902 37062
rect 14758 36998 14764 37030
rect 14622 35774 14623 35806
rect 14557 35773 14623 35774
rect 952 35638 1230 35702
rect 1294 35638 1300 35702
rect 952 34070 1300 35638
rect 14688 34478 14764 36998
rect 21896 36998 21902 37030
rect 21966 37030 21967 37062
rect 22309 37062 22375 37063
rect 22309 37030 22310 37062
rect 21966 36998 21972 37030
rect 21896 36790 21972 36998
rect 21896 36726 21902 36790
rect 21966 36726 21972 36790
rect 21896 36720 21972 36726
rect 22304 36998 22310 37030
rect 22374 37030 22375 37062
rect 22984 37062 23060 37068
rect 22374 36998 22380 37030
rect 22304 36790 22380 36998
rect 22304 36726 22310 36790
rect 22374 36726 22380 36790
rect 22984 36998 22990 37062
rect 23054 36998 23060 37062
rect 22984 36790 23060 36998
rect 22984 36758 22990 36790
rect 22304 36720 22380 36726
rect 22989 36726 22990 36758
rect 23054 36758 23060 36790
rect 23528 37062 23604 37068
rect 23528 36998 23534 37062
rect 23598 36998 23604 37062
rect 23528 36790 23604 36998
rect 23528 36758 23534 36790
rect 23054 36726 23055 36758
rect 22989 36725 23055 36726
rect 23533 36726 23534 36758
rect 23598 36758 23604 36790
rect 195160 37062 195236 37068
rect 195160 36998 195166 37062
rect 195230 36998 195236 37062
rect 195573 37062 195639 37063
rect 195573 37030 195574 37062
rect 195160 36790 195236 36998
rect 195160 36758 195166 36790
rect 23598 36726 23599 36758
rect 23533 36725 23599 36726
rect 195165 36726 195166 36758
rect 195230 36758 195236 36790
rect 195568 36998 195574 37030
rect 195638 37030 195639 37062
rect 196797 37062 196863 37063
rect 196797 37030 196798 37062
rect 195638 36998 195644 37030
rect 195568 36790 195644 36998
rect 195230 36726 195231 36758
rect 195165 36725 195231 36726
rect 195568 36726 195574 36790
rect 195638 36726 195644 36790
rect 195568 36720 195644 36726
rect 196792 36998 196798 37030
rect 196862 37030 196863 37062
rect 196862 36998 196868 37030
rect 196792 36790 196868 36998
rect 196792 36726 196798 36790
rect 196862 36726 196868 36790
rect 196792 36720 196868 36726
rect 21896 36654 21972 36660
rect 21896 36590 21902 36654
rect 21966 36590 21972 36654
rect 22581 36654 22647 36655
rect 22581 36622 22582 36654
rect 21896 36382 21972 36590
rect 21896 36350 21902 36382
rect 21901 36318 21902 36350
rect 21966 36350 21972 36382
rect 22576 36590 22582 36622
rect 22646 36622 22647 36654
rect 22984 36654 23060 36660
rect 22646 36590 22652 36622
rect 22576 36382 22652 36590
rect 21966 36318 21967 36350
rect 21901 36317 21967 36318
rect 22576 36318 22582 36382
rect 22646 36318 22652 36382
rect 22984 36590 22990 36654
rect 23054 36590 23060 36654
rect 23533 36654 23599 36655
rect 23533 36622 23534 36654
rect 22984 36382 23060 36590
rect 22984 36350 22990 36382
rect 22576 36312 22652 36318
rect 22989 36318 22990 36350
rect 23054 36350 23060 36382
rect 23528 36590 23534 36622
rect 23598 36622 23599 36654
rect 195165 36654 195231 36655
rect 195165 36622 195166 36654
rect 23598 36590 23604 36622
rect 23528 36382 23604 36590
rect 23054 36318 23055 36350
rect 22989 36317 23055 36318
rect 23528 36318 23534 36382
rect 23598 36318 23604 36382
rect 23528 36312 23604 36318
rect 195160 36590 195166 36622
rect 195230 36622 195231 36654
rect 195432 36654 195508 36660
rect 195230 36590 195236 36622
rect 195160 36382 195236 36590
rect 195160 36318 195166 36382
rect 195230 36318 195236 36382
rect 195432 36590 195438 36654
rect 195502 36590 195508 36654
rect 195432 36382 195508 36590
rect 195432 36350 195438 36382
rect 195160 36312 195236 36318
rect 195437 36318 195438 36350
rect 195502 36350 195508 36382
rect 196792 36654 196868 36660
rect 196792 36590 196798 36654
rect 196862 36590 196868 36654
rect 196792 36382 196868 36590
rect 196792 36350 196798 36382
rect 195502 36318 195503 36350
rect 195437 36317 195503 36318
rect 196797 36318 196798 36350
rect 196862 36350 196868 36382
rect 196862 36318 196863 36350
rect 196797 36317 196863 36318
rect 22445 36246 22511 36247
rect 22445 36214 22446 36246
rect 22440 36182 22446 36214
rect 22510 36214 22511 36246
rect 22712 36246 22788 36252
rect 22510 36182 22516 36214
rect 22440 35974 22516 36182
rect 22440 35910 22446 35974
rect 22510 35910 22516 35974
rect 22712 36182 22718 36246
rect 22782 36182 22788 36246
rect 22712 35974 22788 36182
rect 22712 35942 22718 35974
rect 22440 35904 22516 35910
rect 22717 35910 22718 35942
rect 22782 35942 22788 35974
rect 23120 36246 23196 36252
rect 23120 36182 23126 36246
rect 23190 36182 23196 36246
rect 23120 35974 23196 36182
rect 23120 35942 23126 35974
rect 22782 35910 22783 35942
rect 22717 35909 22783 35910
rect 23125 35910 23126 35942
rect 23190 35942 23196 35974
rect 23392 36246 23468 36252
rect 23392 36182 23398 36246
rect 23462 36182 23468 36246
rect 23392 35974 23468 36182
rect 195024 36246 195100 36252
rect 195024 36182 195030 36246
rect 195094 36182 195100 36246
rect 195437 36246 195503 36247
rect 195437 36214 195438 36246
rect 28293 36110 28359 36111
rect 28293 36078 28294 36110
rect 23392 35942 23398 35974
rect 23190 35910 23191 35942
rect 23125 35909 23191 35910
rect 23397 35910 23398 35942
rect 23462 35942 23468 35974
rect 28288 36046 28294 36078
rect 28358 36078 28359 36110
rect 28358 36046 28364 36078
rect 23462 35910 23463 35942
rect 23397 35909 23463 35910
rect 22989 35838 23055 35839
rect 22989 35806 22990 35838
rect 22984 35774 22990 35806
rect 23054 35806 23055 35838
rect 23533 35838 23599 35839
rect 23533 35806 23534 35838
rect 23054 35774 23060 35806
rect 18501 35702 18567 35703
rect 18501 35670 18502 35702
rect 14688 34414 14694 34478
rect 14758 34414 14764 34478
rect 14688 34408 14764 34414
rect 18496 35638 18502 35670
rect 18566 35670 18567 35702
rect 18566 35638 18572 35670
rect 16597 34206 16663 34207
rect 16597 34174 16598 34206
rect 952 34006 1230 34070
rect 1294 34006 1300 34070
rect 952 32438 1300 34006
rect 952 32374 1230 32438
rect 1294 32374 1300 32438
rect 952 30806 1300 32374
rect 16592 34142 16598 34174
rect 16662 34174 16663 34206
rect 16662 34142 16668 34174
rect 16592 31622 16668 34142
rect 18496 34070 18572 35638
rect 22984 35566 23060 35774
rect 22984 35502 22990 35566
rect 23054 35502 23060 35566
rect 22984 35496 23060 35502
rect 23528 35774 23534 35806
rect 23598 35806 23599 35838
rect 28288 35838 28364 36046
rect 195024 35974 195100 36182
rect 195024 35942 195030 35974
rect 195029 35910 195030 35942
rect 195094 35942 195100 35974
rect 195432 36182 195438 36214
rect 195502 36214 195503 36246
rect 196389 36246 196455 36247
rect 196389 36214 196390 36246
rect 195502 36182 195508 36214
rect 195432 35974 195508 36182
rect 195094 35910 195095 35942
rect 195029 35909 195095 35910
rect 195432 35910 195438 35974
rect 195502 35910 195508 35974
rect 195432 35904 195508 35910
rect 196384 36182 196390 36214
rect 196454 36214 196455 36246
rect 196454 36182 196460 36214
rect 196384 35974 196460 36182
rect 196384 35910 196390 35974
rect 196454 35910 196460 35974
rect 196384 35904 196460 35910
rect 23598 35774 23604 35806
rect 23528 35566 23604 35774
rect 28288 35774 28294 35838
rect 28358 35774 28364 35838
rect 28288 35768 28364 35774
rect 195160 35838 195236 35844
rect 195160 35774 195166 35838
rect 195230 35774 195236 35838
rect 195437 35838 195503 35839
rect 195437 35806 195438 35838
rect 23528 35502 23534 35566
rect 23598 35502 23604 35566
rect 195160 35566 195236 35774
rect 195160 35534 195166 35566
rect 23528 35496 23604 35502
rect 195165 35502 195166 35534
rect 195230 35534 195236 35566
rect 195432 35774 195438 35806
rect 195502 35806 195503 35838
rect 217464 35838 217812 37542
rect 195502 35774 195508 35806
rect 195432 35566 195508 35774
rect 195230 35502 195231 35534
rect 195165 35501 195231 35502
rect 195432 35502 195438 35566
rect 195502 35502 195508 35566
rect 195432 35496 195508 35502
rect 217464 35774 217470 35838
rect 217534 35774 217812 35838
rect 22304 35430 22380 35436
rect 22304 35366 22310 35430
rect 22374 35366 22380 35430
rect 21901 35158 21967 35159
rect 21901 35126 21902 35158
rect 21896 35094 21902 35126
rect 21966 35126 21967 35158
rect 22304 35158 22380 35366
rect 22304 35126 22310 35158
rect 21966 35094 21972 35126
rect 21896 34886 21972 35094
rect 22309 35094 22310 35126
rect 22374 35126 22380 35158
rect 22440 35430 22516 35436
rect 22440 35366 22446 35430
rect 22510 35366 22516 35430
rect 22440 35158 22516 35366
rect 22440 35126 22446 35158
rect 22374 35094 22375 35126
rect 22309 35093 22375 35094
rect 22445 35094 22446 35126
rect 22510 35126 22516 35158
rect 22984 35430 23060 35436
rect 22984 35366 22990 35430
rect 23054 35366 23060 35430
rect 22984 35158 23060 35366
rect 22984 35126 22990 35158
rect 22510 35094 22511 35126
rect 22445 35093 22511 35094
rect 22989 35094 22990 35126
rect 23054 35126 23060 35158
rect 23392 35430 23468 35436
rect 23392 35366 23398 35430
rect 23462 35366 23468 35430
rect 195165 35430 195231 35431
rect 195165 35398 195166 35430
rect 23392 35158 23468 35366
rect 195160 35366 195166 35398
rect 195230 35398 195231 35430
rect 195432 35430 195508 35436
rect 195230 35366 195236 35398
rect 190269 35294 190335 35295
rect 190269 35262 190270 35294
rect 23392 35126 23398 35158
rect 23054 35094 23055 35126
rect 22989 35093 23055 35094
rect 23397 35094 23398 35126
rect 23462 35126 23468 35158
rect 190264 35230 190270 35262
rect 190334 35262 190335 35294
rect 190334 35230 190340 35262
rect 23462 35094 23463 35126
rect 23397 35093 23463 35094
rect 190264 35022 190340 35230
rect 195160 35158 195236 35366
rect 195160 35094 195166 35158
rect 195230 35094 195236 35158
rect 195432 35366 195438 35430
rect 195502 35366 195508 35430
rect 195432 35158 195508 35366
rect 195432 35126 195438 35158
rect 195160 35088 195236 35094
rect 195437 35094 195438 35126
rect 195502 35126 195508 35158
rect 195976 35430 196052 35436
rect 195976 35366 195982 35430
rect 196046 35366 196052 35430
rect 195976 35158 196052 35366
rect 195976 35126 195982 35158
rect 195502 35094 195503 35126
rect 195437 35093 195503 35094
rect 195981 35094 195982 35126
rect 196046 35126 196052 35158
rect 196112 35430 196188 35436
rect 196112 35366 196118 35430
rect 196182 35366 196188 35430
rect 196112 35158 196188 35366
rect 196112 35126 196118 35158
rect 196046 35094 196047 35126
rect 195981 35093 196047 35094
rect 196117 35094 196118 35126
rect 196182 35126 196188 35158
rect 196792 35158 196868 35164
rect 196182 35094 196183 35126
rect 196117 35093 196183 35094
rect 196792 35094 196798 35158
rect 196862 35094 196868 35158
rect 190264 34958 190270 35022
rect 190334 34958 190340 35022
rect 190264 34952 190340 34958
rect 21896 34822 21902 34886
rect 21966 34822 21972 34886
rect 21896 34816 21972 34822
rect 28424 34886 28500 34892
rect 28424 34822 28430 34886
rect 28494 34822 28500 34886
rect 21760 34750 21836 34756
rect 21760 34686 21766 34750
rect 21830 34686 21836 34750
rect 21760 34478 21836 34686
rect 21760 34446 21766 34478
rect 21765 34414 21766 34446
rect 21830 34446 21836 34478
rect 22168 34750 22244 34756
rect 22168 34686 22174 34750
rect 22238 34686 22244 34750
rect 22581 34750 22647 34751
rect 22581 34718 22582 34750
rect 22168 34478 22244 34686
rect 22168 34446 22174 34478
rect 21830 34414 21831 34446
rect 21765 34413 21831 34414
rect 22173 34414 22174 34446
rect 22238 34446 22244 34478
rect 22576 34686 22582 34718
rect 22646 34718 22647 34750
rect 22646 34686 22652 34718
rect 22576 34478 22652 34686
rect 28424 34614 28500 34822
rect 28424 34582 28430 34614
rect 28429 34550 28430 34582
rect 28494 34582 28500 34614
rect 190128 34886 190204 34892
rect 190128 34822 190134 34886
rect 190198 34822 190204 34886
rect 196792 34886 196868 35094
rect 196792 34854 196798 34886
rect 190128 34614 190204 34822
rect 196797 34822 196798 34854
rect 196862 34854 196868 34886
rect 196862 34822 196863 34854
rect 196797 34821 196863 34822
rect 195845 34750 195911 34751
rect 195845 34718 195846 34750
rect 190128 34582 190134 34614
rect 28494 34550 28495 34582
rect 28429 34549 28495 34550
rect 190133 34550 190134 34582
rect 190198 34582 190204 34614
rect 195840 34686 195846 34718
rect 195910 34718 195911 34750
rect 196661 34750 196727 34751
rect 196661 34718 196662 34750
rect 195910 34686 195916 34718
rect 190198 34550 190199 34582
rect 190133 34549 190199 34550
rect 22238 34414 22239 34446
rect 22173 34413 22239 34414
rect 22576 34414 22582 34478
rect 22646 34414 22652 34478
rect 22576 34408 22652 34414
rect 28288 34478 28364 34484
rect 28288 34414 28294 34478
rect 28358 34414 28364 34478
rect 190133 34478 190199 34479
rect 190133 34446 190134 34478
rect 21765 34342 21831 34343
rect 21765 34310 21766 34342
rect 18496 34006 18502 34070
rect 18566 34006 18572 34070
rect 18496 34000 18572 34006
rect 21760 34278 21766 34310
rect 21830 34310 21831 34342
rect 21830 34278 21836 34310
rect 21760 34070 21836 34278
rect 28288 34206 28364 34414
rect 190128 34414 190134 34446
rect 190198 34446 190199 34478
rect 195840 34478 195916 34686
rect 190198 34414 190204 34446
rect 28288 34174 28294 34206
rect 28293 34142 28294 34174
rect 28358 34174 28364 34206
rect 28424 34206 28500 34212
rect 28358 34142 28359 34174
rect 28293 34141 28359 34142
rect 28424 34142 28430 34206
rect 28494 34142 28500 34206
rect 21760 34006 21766 34070
rect 21830 34006 21836 34070
rect 21760 34000 21836 34006
rect 18224 33934 18300 33940
rect 18224 33870 18230 33934
rect 18294 33870 18300 33934
rect 18224 33254 18300 33870
rect 18224 33222 18230 33254
rect 18229 33190 18230 33222
rect 18294 33222 18300 33254
rect 18904 33934 18980 33940
rect 18904 33870 18910 33934
rect 18974 33870 18980 33934
rect 18904 33254 18980 33870
rect 18904 33222 18910 33254
rect 18294 33190 18295 33222
rect 18229 33189 18295 33190
rect 18909 33190 18910 33222
rect 18974 33222 18980 33254
rect 19312 33934 19388 33940
rect 19312 33870 19318 33934
rect 19382 33870 19388 33934
rect 19312 33254 19388 33870
rect 21760 33934 21836 33940
rect 21760 33870 21766 33934
rect 21830 33870 21836 33934
rect 21760 33662 21836 33870
rect 21760 33630 21766 33662
rect 21765 33598 21766 33630
rect 21830 33630 21836 33662
rect 22168 33934 22244 33940
rect 22168 33870 22174 33934
rect 22238 33870 22244 33934
rect 22168 33662 22244 33870
rect 22168 33630 22174 33662
rect 21830 33598 21831 33630
rect 21765 33597 21831 33598
rect 22173 33598 22174 33630
rect 22238 33630 22244 33662
rect 22576 33934 22652 33940
rect 22576 33870 22582 33934
rect 22646 33870 22652 33934
rect 22576 33662 22652 33870
rect 22576 33630 22582 33662
rect 22238 33598 22239 33630
rect 22173 33597 22239 33598
rect 22581 33598 22582 33630
rect 22646 33630 22652 33662
rect 22984 33934 23060 33940
rect 22984 33870 22990 33934
rect 23054 33870 23060 33934
rect 22984 33662 23060 33870
rect 22984 33630 22990 33662
rect 22646 33598 22647 33630
rect 22581 33597 22647 33598
rect 22989 33598 22990 33630
rect 23054 33630 23060 33662
rect 23528 33934 23604 33940
rect 23528 33870 23534 33934
rect 23598 33870 23604 33934
rect 28424 33934 28500 34142
rect 190128 34206 190204 34414
rect 195840 34414 195846 34478
rect 195910 34414 195916 34478
rect 195840 34408 195916 34414
rect 196656 34686 196662 34718
rect 196726 34718 196727 34750
rect 196726 34686 196732 34718
rect 196656 34478 196732 34686
rect 196656 34414 196662 34478
rect 196726 34414 196732 34478
rect 196656 34408 196732 34414
rect 196661 34342 196727 34343
rect 196661 34310 196662 34342
rect 190128 34142 190134 34206
rect 190198 34142 190204 34206
rect 190128 34136 190204 34142
rect 196656 34278 196662 34310
rect 196726 34310 196727 34342
rect 196726 34278 196732 34310
rect 196656 34070 196732 34278
rect 196656 34006 196662 34070
rect 196726 34006 196732 34070
rect 196656 34000 196732 34006
rect 217464 34206 217812 35774
rect 217464 34142 217470 34206
rect 217534 34142 217812 34206
rect 28424 33902 28430 33934
rect 23528 33662 23604 33870
rect 28429 33870 28430 33902
rect 28494 33902 28500 33934
rect 195160 33934 195236 33940
rect 28494 33870 28495 33902
rect 28429 33869 28495 33870
rect 195160 33870 195166 33934
rect 195230 33870 195236 33934
rect 195437 33934 195503 33935
rect 195437 33902 195438 33934
rect 23528 33630 23534 33662
rect 23054 33598 23055 33630
rect 22989 33597 23055 33598
rect 23533 33598 23534 33630
rect 23598 33630 23604 33662
rect 195160 33662 195236 33870
rect 195160 33630 195166 33662
rect 23598 33598 23599 33630
rect 23533 33597 23599 33598
rect 195165 33598 195166 33630
rect 195230 33630 195236 33662
rect 195432 33870 195438 33902
rect 195502 33902 195503 33934
rect 196389 33934 196455 33935
rect 196389 33902 196390 33934
rect 195502 33870 195508 33902
rect 195432 33662 195508 33870
rect 195230 33598 195231 33630
rect 195165 33597 195231 33598
rect 195432 33598 195438 33662
rect 195502 33598 195508 33662
rect 195432 33592 195508 33598
rect 196384 33870 196390 33902
rect 196454 33902 196455 33934
rect 196656 33934 196732 33940
rect 196454 33870 196460 33902
rect 196384 33662 196460 33870
rect 196384 33598 196390 33662
rect 196454 33598 196460 33662
rect 196656 33870 196662 33934
rect 196726 33870 196732 33934
rect 196656 33662 196732 33870
rect 196656 33630 196662 33662
rect 196384 33592 196460 33598
rect 196661 33598 196662 33630
rect 196726 33630 196732 33662
rect 198832 33934 198908 33940
rect 198832 33870 198838 33934
rect 198902 33870 198908 33934
rect 199109 33934 199175 33935
rect 199109 33902 199110 33934
rect 196726 33598 196727 33630
rect 196661 33597 196727 33598
rect 21765 33526 21831 33527
rect 21765 33494 21766 33526
rect 19312 33222 19318 33254
rect 18974 33190 18975 33222
rect 18909 33189 18975 33190
rect 19317 33190 19318 33222
rect 19382 33222 19388 33254
rect 21760 33462 21766 33494
rect 21830 33494 21831 33526
rect 22581 33526 22647 33527
rect 22581 33494 22582 33526
rect 21830 33462 21836 33494
rect 21760 33254 21836 33462
rect 19382 33190 19383 33222
rect 19317 33189 19383 33190
rect 21760 33190 21766 33254
rect 21830 33190 21836 33254
rect 21760 33184 21836 33190
rect 22576 33462 22582 33494
rect 22646 33494 22647 33526
rect 23120 33526 23196 33532
rect 22646 33462 22652 33494
rect 22576 33254 22652 33462
rect 22576 33190 22582 33254
rect 22646 33190 22652 33254
rect 23120 33462 23126 33526
rect 23190 33462 23196 33526
rect 23120 33254 23196 33462
rect 23120 33222 23126 33254
rect 22576 33184 22652 33190
rect 23125 33190 23126 33222
rect 23190 33222 23196 33254
rect 23528 33526 23604 33532
rect 23528 33462 23534 33526
rect 23598 33462 23604 33526
rect 195165 33526 195231 33527
rect 195165 33494 195166 33526
rect 23528 33254 23604 33462
rect 23528 33222 23534 33254
rect 23190 33190 23191 33222
rect 23125 33189 23191 33190
rect 23533 33190 23534 33222
rect 23598 33222 23604 33254
rect 195160 33462 195166 33494
rect 195230 33494 195231 33526
rect 195568 33526 195644 33532
rect 195230 33462 195236 33494
rect 195160 33254 195236 33462
rect 23598 33190 23599 33222
rect 23533 33189 23599 33190
rect 195160 33190 195166 33254
rect 195230 33190 195236 33254
rect 195568 33462 195574 33526
rect 195638 33462 195644 33526
rect 196117 33526 196183 33527
rect 196117 33494 196118 33526
rect 195568 33254 195644 33462
rect 195568 33222 195574 33254
rect 195160 33184 195236 33190
rect 195573 33190 195574 33222
rect 195638 33222 195644 33254
rect 196112 33462 196118 33494
rect 196182 33494 196183 33526
rect 196384 33526 196460 33532
rect 196182 33462 196188 33494
rect 196112 33254 196188 33462
rect 195638 33190 195639 33222
rect 195573 33189 195639 33190
rect 196112 33190 196118 33254
rect 196182 33190 196188 33254
rect 196384 33462 196390 33526
rect 196454 33462 196460 33526
rect 196661 33526 196727 33527
rect 196661 33494 196662 33526
rect 196384 33254 196460 33462
rect 196384 33222 196390 33254
rect 196112 33184 196188 33190
rect 196389 33190 196390 33222
rect 196454 33222 196460 33254
rect 196656 33462 196662 33494
rect 196726 33494 196727 33526
rect 196726 33462 196732 33494
rect 196656 33254 196732 33462
rect 196454 33190 196455 33222
rect 196389 33189 196455 33190
rect 196656 33190 196662 33254
rect 196726 33190 196732 33254
rect 198832 33254 198908 33870
rect 198832 33222 198838 33254
rect 196656 33184 196732 33190
rect 198837 33190 198838 33222
rect 198902 33222 198908 33254
rect 199104 33870 199110 33902
rect 199174 33902 199175 33934
rect 200469 33934 200535 33935
rect 200469 33902 200470 33934
rect 199174 33870 199180 33902
rect 199104 33254 199180 33870
rect 198902 33190 198903 33222
rect 198837 33189 198903 33190
rect 199104 33190 199110 33254
rect 199174 33190 199180 33254
rect 199104 33184 199180 33190
rect 200464 33870 200470 33902
rect 200534 33902 200535 33934
rect 200534 33870 200540 33902
rect 200464 33254 200540 33870
rect 200464 33190 200470 33254
rect 200534 33190 200540 33254
rect 200464 33184 200540 33190
rect 18093 33118 18159 33119
rect 18093 33086 18094 33118
rect 18088 33054 18094 33086
rect 18158 33086 18159 33118
rect 18773 33118 18839 33119
rect 18773 33086 18774 33118
rect 18158 33054 18164 33086
rect 18088 32438 18164 33054
rect 18088 32374 18094 32438
rect 18158 32374 18164 32438
rect 18088 32368 18164 32374
rect 18768 33054 18774 33086
rect 18838 33086 18839 33118
rect 19453 33118 19519 33119
rect 19453 33086 19454 33118
rect 18838 33054 18844 33086
rect 18768 32444 18844 33054
rect 19448 33054 19454 33086
rect 19518 33086 19519 33118
rect 21896 33118 21972 33124
rect 19518 33054 19524 33086
rect 18768 32438 18980 32444
rect 18768 32374 18910 32438
rect 18974 32374 18980 32438
rect 18768 32368 18980 32374
rect 19448 32438 19524 33054
rect 21896 33054 21902 33118
rect 21966 33054 21972 33118
rect 22445 33118 22511 33119
rect 22445 33086 22446 33118
rect 21896 32846 21972 33054
rect 21896 32814 21902 32846
rect 21901 32782 21902 32814
rect 21966 32814 21972 32846
rect 22440 33054 22446 33086
rect 22510 33086 22511 33118
rect 22989 33118 23055 33119
rect 22989 33086 22990 33118
rect 22510 33054 22516 33086
rect 22440 32846 22516 33054
rect 21966 32782 21967 32814
rect 21901 32781 21967 32782
rect 22440 32782 22446 32846
rect 22510 32782 22516 32846
rect 22440 32776 22516 32782
rect 22984 33054 22990 33086
rect 23054 33086 23055 33118
rect 23397 33118 23463 33119
rect 23397 33086 23398 33118
rect 23054 33054 23060 33086
rect 22984 32846 23060 33054
rect 22984 32782 22990 32846
rect 23054 32782 23060 32846
rect 22984 32776 23060 32782
rect 23392 33054 23398 33086
rect 23462 33086 23463 33118
rect 195024 33118 195100 33124
rect 23462 33054 23468 33086
rect 23392 32846 23468 33054
rect 23392 32782 23398 32846
rect 23462 32782 23468 32846
rect 195024 33054 195030 33118
rect 195094 33054 195100 33118
rect 195024 32846 195100 33054
rect 195024 32814 195030 32846
rect 23392 32776 23468 32782
rect 195029 32782 195030 32814
rect 195094 32814 195100 32846
rect 195568 33118 195644 33124
rect 195568 33054 195574 33118
rect 195638 33054 195644 33118
rect 195568 32846 195644 33054
rect 195568 32814 195574 32846
rect 195094 32782 195095 32814
rect 195029 32781 195095 32782
rect 195573 32782 195574 32814
rect 195638 32814 195644 32846
rect 195976 33118 196052 33124
rect 195976 33054 195982 33118
rect 196046 33054 196052 33118
rect 195976 32846 196052 33054
rect 195976 32814 195982 32846
rect 195638 32782 195639 32814
rect 195573 32781 195639 32782
rect 195981 32782 195982 32814
rect 196046 32814 196052 32846
rect 196112 33118 196188 33124
rect 196112 33054 196118 33118
rect 196182 33054 196188 33118
rect 196112 32846 196188 33054
rect 196112 32814 196118 32846
rect 196046 32782 196047 32814
rect 195981 32781 196047 32782
rect 196117 32782 196118 32814
rect 196182 32814 196188 32846
rect 196792 33118 196868 33124
rect 196792 33054 196798 33118
rect 196862 33054 196868 33118
rect 196792 32846 196868 33054
rect 196792 32814 196798 32846
rect 196182 32782 196183 32814
rect 196117 32781 196183 32782
rect 196797 32782 196798 32814
rect 196862 32814 196868 32846
rect 199104 33118 199180 33124
rect 199104 33054 199110 33118
rect 199174 33054 199180 33118
rect 199789 33118 199855 33119
rect 199789 33086 199790 33118
rect 196862 32782 196863 32814
rect 196797 32781 196863 32782
rect 21901 32710 21967 32711
rect 21901 32678 21902 32710
rect 19448 32374 19454 32438
rect 19518 32374 19524 32438
rect 19448 32368 19524 32374
rect 21896 32646 21902 32678
rect 21966 32678 21967 32710
rect 23125 32710 23191 32711
rect 23125 32678 23126 32710
rect 21966 32646 21972 32678
rect 21896 32438 21972 32646
rect 21896 32374 21902 32438
rect 21966 32374 21972 32438
rect 21896 32368 21972 32374
rect 23120 32646 23126 32678
rect 23190 32678 23191 32710
rect 23397 32710 23463 32711
rect 23397 32678 23398 32710
rect 23190 32646 23196 32678
rect 23120 32438 23196 32646
rect 23120 32374 23126 32438
rect 23190 32374 23196 32438
rect 23120 32368 23196 32374
rect 23392 32646 23398 32678
rect 23462 32678 23463 32710
rect 195160 32710 195236 32716
rect 23462 32646 23468 32678
rect 23392 32438 23468 32646
rect 23392 32374 23398 32438
rect 23462 32374 23468 32438
rect 195160 32646 195166 32710
rect 195230 32646 195236 32710
rect 195160 32438 195236 32646
rect 195160 32406 195166 32438
rect 23392 32368 23468 32374
rect 195165 32374 195166 32406
rect 195230 32406 195236 32438
rect 195432 32710 195508 32716
rect 195432 32646 195438 32710
rect 195502 32646 195508 32710
rect 195981 32710 196047 32711
rect 195981 32678 195982 32710
rect 195432 32438 195508 32646
rect 195432 32406 195438 32438
rect 195230 32374 195231 32406
rect 195165 32373 195231 32374
rect 195437 32374 195438 32406
rect 195502 32406 195508 32438
rect 195976 32646 195982 32678
rect 196046 32678 196047 32710
rect 196389 32710 196455 32711
rect 196389 32678 196390 32710
rect 196046 32646 196052 32678
rect 195976 32438 196052 32646
rect 195502 32374 195503 32406
rect 195437 32373 195503 32374
rect 195976 32374 195982 32438
rect 196046 32374 196052 32438
rect 195976 32368 196052 32374
rect 196384 32646 196390 32678
rect 196454 32678 196455 32710
rect 196797 32710 196863 32711
rect 196797 32678 196798 32710
rect 196454 32646 196460 32678
rect 196384 32438 196460 32646
rect 196384 32374 196390 32438
rect 196454 32374 196460 32438
rect 196384 32368 196460 32374
rect 196792 32646 196798 32678
rect 196862 32678 196863 32710
rect 196862 32646 196868 32678
rect 196792 32438 196868 32646
rect 196792 32374 196798 32438
rect 196862 32374 196868 32438
rect 199104 32438 199180 33054
rect 199104 32406 199110 32438
rect 196792 32368 196868 32374
rect 199109 32374 199110 32406
rect 199174 32406 199180 32438
rect 199784 33054 199790 33086
rect 199854 33086 199855 33118
rect 200469 33118 200535 33119
rect 200469 33086 200470 33118
rect 199854 33054 199860 33086
rect 199784 32444 199860 33054
rect 200464 33054 200470 33086
rect 200534 33086 200535 33118
rect 200534 33054 200540 33086
rect 199784 32438 199996 32444
rect 199174 32374 199175 32406
rect 199109 32373 199175 32374
rect 199784 32374 199926 32438
rect 199990 32374 199996 32438
rect 199784 32368 199996 32374
rect 200464 32438 200540 33054
rect 200464 32374 200470 32438
rect 200534 32374 200540 32438
rect 200464 32368 200540 32374
rect 217464 32574 217812 34142
rect 217464 32510 217470 32574
rect 217534 32510 217812 32574
rect 18093 32302 18159 32303
rect 18093 32270 18094 32302
rect 16592 31558 16598 31622
rect 16662 31558 16668 31622
rect 16592 31552 16668 31558
rect 18088 32238 18094 32270
rect 18158 32270 18159 32302
rect 18909 32302 18975 32303
rect 18909 32270 18910 32302
rect 18158 32238 18164 32270
rect 18088 31622 18164 32238
rect 18088 31558 18094 31622
rect 18158 31558 18164 31622
rect 18088 31552 18164 31558
rect 18904 32238 18910 32270
rect 18974 32270 18975 32302
rect 19448 32302 19524 32308
rect 18974 32238 18980 32270
rect 18904 31622 18980 32238
rect 18904 31558 18910 31622
rect 18974 31558 18980 31622
rect 19448 32238 19454 32302
rect 19518 32238 19524 32302
rect 19448 31622 19524 32238
rect 19448 31590 19454 31622
rect 18904 31552 18980 31558
rect 19453 31558 19454 31590
rect 19518 31590 19524 31622
rect 19856 32302 19932 32308
rect 19856 32238 19862 32302
rect 19926 32238 19932 32302
rect 22173 32302 22239 32303
rect 22173 32270 22174 32302
rect 19856 31622 19932 32238
rect 22168 32238 22174 32270
rect 22238 32270 22239 32302
rect 22712 32302 22788 32308
rect 22238 32238 22244 32270
rect 22168 32030 22244 32238
rect 22168 31966 22174 32030
rect 22238 31966 22244 32030
rect 22712 32238 22718 32302
rect 22782 32238 22788 32302
rect 22712 32030 22788 32238
rect 22712 31998 22718 32030
rect 22168 31960 22244 31966
rect 22717 31966 22718 31998
rect 22782 31998 22788 32030
rect 22984 32302 23060 32308
rect 22984 32238 22990 32302
rect 23054 32238 23060 32302
rect 23533 32302 23599 32303
rect 23533 32270 23534 32302
rect 22984 32030 23060 32238
rect 22984 31998 22990 32030
rect 22782 31966 22783 31998
rect 22717 31965 22783 31966
rect 22989 31966 22990 31998
rect 23054 31998 23060 32030
rect 23528 32238 23534 32270
rect 23598 32270 23599 32302
rect 195165 32302 195231 32303
rect 195165 32270 195166 32302
rect 23598 32238 23604 32270
rect 23528 32030 23604 32238
rect 23054 31966 23055 31998
rect 22989 31965 23055 31966
rect 23528 31966 23534 32030
rect 23598 31966 23604 32030
rect 23528 31960 23604 31966
rect 195160 32238 195166 32270
rect 195230 32270 195231 32302
rect 195437 32302 195503 32303
rect 195437 32270 195438 32302
rect 195230 32238 195236 32270
rect 195160 32030 195236 32238
rect 195160 31966 195166 32030
rect 195230 31966 195236 32030
rect 195160 31960 195236 31966
rect 195432 32238 195438 32270
rect 195502 32270 195503 32302
rect 196112 32302 196188 32308
rect 195502 32238 195508 32270
rect 195432 32030 195508 32238
rect 195432 31966 195438 32030
rect 195502 31966 195508 32030
rect 196112 32238 196118 32302
rect 196182 32238 196188 32302
rect 196112 32030 196188 32238
rect 196112 31998 196118 32030
rect 195432 31960 195508 31966
rect 196117 31966 196118 31998
rect 196182 31998 196188 32030
rect 198968 32302 199044 32308
rect 198968 32238 198974 32302
rect 199038 32238 199044 32302
rect 199245 32302 199311 32303
rect 199245 32270 199246 32302
rect 196182 31966 196183 31998
rect 196117 31965 196183 31966
rect 19856 31590 19862 31622
rect 19518 31558 19519 31590
rect 19453 31557 19519 31558
rect 19861 31558 19862 31590
rect 19926 31590 19932 31622
rect 21896 31894 21972 31900
rect 21896 31830 21902 31894
rect 21966 31830 21972 31894
rect 21896 31622 21972 31830
rect 21896 31590 21902 31622
rect 19926 31558 19927 31590
rect 19861 31557 19927 31558
rect 21901 31558 21902 31590
rect 21966 31590 21972 31622
rect 22304 31894 22380 31900
rect 22304 31830 22310 31894
rect 22374 31830 22380 31894
rect 22304 31622 22380 31830
rect 22304 31590 22310 31622
rect 21966 31558 21967 31590
rect 21901 31557 21967 31558
rect 22309 31558 22310 31590
rect 22374 31590 22380 31622
rect 22440 31894 22516 31900
rect 22440 31830 22446 31894
rect 22510 31830 22516 31894
rect 22440 31622 22516 31830
rect 22440 31590 22446 31622
rect 22374 31558 22375 31590
rect 22309 31557 22375 31558
rect 22445 31558 22446 31590
rect 22510 31590 22516 31622
rect 23120 31894 23196 31900
rect 23120 31830 23126 31894
rect 23190 31830 23196 31894
rect 23397 31894 23463 31895
rect 23397 31862 23398 31894
rect 23120 31622 23196 31830
rect 23120 31590 23126 31622
rect 22510 31558 22511 31590
rect 22445 31557 22511 31558
rect 23125 31558 23126 31590
rect 23190 31590 23196 31622
rect 23392 31830 23398 31862
rect 23462 31862 23463 31894
rect 195024 31894 195100 31900
rect 23462 31830 23468 31862
rect 23392 31622 23468 31830
rect 23190 31558 23191 31590
rect 23125 31557 23191 31558
rect 23392 31558 23398 31622
rect 23462 31558 23468 31622
rect 195024 31830 195030 31894
rect 195094 31830 195100 31894
rect 195437 31894 195503 31895
rect 195437 31862 195438 31894
rect 195024 31622 195100 31830
rect 195024 31590 195030 31622
rect 23392 31552 23468 31558
rect 195029 31558 195030 31590
rect 195094 31590 195100 31622
rect 195432 31830 195438 31862
rect 195502 31862 195503 31894
rect 196384 31894 196460 31900
rect 195502 31830 195508 31862
rect 195432 31622 195508 31830
rect 195094 31558 195095 31590
rect 195029 31557 195095 31558
rect 195432 31558 195438 31622
rect 195502 31558 195508 31622
rect 196384 31830 196390 31894
rect 196454 31830 196460 31894
rect 196661 31894 196727 31895
rect 196661 31862 196662 31894
rect 196384 31622 196460 31830
rect 196384 31590 196390 31622
rect 195432 31552 195508 31558
rect 196389 31558 196390 31590
rect 196454 31590 196460 31622
rect 196656 31830 196662 31862
rect 196726 31862 196727 31894
rect 196726 31830 196732 31862
rect 196656 31622 196732 31830
rect 196454 31558 196455 31590
rect 196389 31557 196455 31558
rect 196656 31558 196662 31622
rect 196726 31558 196732 31622
rect 198968 31622 199044 32238
rect 198968 31590 198974 31622
rect 196656 31552 196732 31558
rect 198973 31558 198974 31590
rect 199038 31590 199044 31622
rect 199240 32238 199246 32270
rect 199310 32270 199311 32302
rect 200464 32302 200540 32308
rect 199310 32238 199316 32270
rect 199240 31622 199316 32238
rect 199038 31558 199039 31590
rect 198973 31557 199039 31558
rect 199240 31558 199246 31622
rect 199310 31558 199316 31622
rect 200464 32238 200470 32302
rect 200534 32238 200540 32302
rect 201829 32302 201895 32303
rect 201829 32270 201830 32302
rect 200464 31622 200540 32238
rect 200464 31590 200470 31622
rect 199240 31552 199316 31558
rect 200469 31558 200470 31590
rect 200534 31590 200540 31622
rect 201824 32238 201830 32270
rect 201894 32270 201895 32302
rect 201894 32238 201900 32270
rect 201824 31622 201900 32238
rect 200534 31558 200535 31590
rect 200469 31557 200535 31558
rect 201824 31558 201830 31622
rect 201894 31558 201900 31622
rect 201824 31552 201900 31558
rect 952 30742 1230 30806
rect 1294 30742 1300 30806
rect 952 29174 1300 30742
rect 18904 31486 18980 31492
rect 18904 31422 18910 31486
rect 18974 31422 18980 31486
rect 19317 31486 19383 31487
rect 19317 31454 19318 31486
rect 2108 30356 2174 30357
rect 2108 30292 2109 30356
rect 2173 30292 2174 30356
rect 2108 30291 2174 30292
rect 952 29110 1230 29174
rect 1294 29110 1300 29174
rect 952 27542 1300 29110
rect 952 27478 1230 27542
rect 1294 27478 1300 27542
rect 1904 28086 1980 28092
rect 1904 28022 1910 28086
rect 1974 28022 1980 28086
rect 1904 27542 1980 28022
rect 1904 27510 1910 27542
rect 952 25638 1300 27478
rect 1909 27478 1910 27510
rect 1974 27510 1980 27542
rect 1974 27478 1975 27510
rect 1909 27477 1975 27478
rect 952 25574 1230 25638
rect 1294 25574 1300 25638
rect 952 24006 1300 25574
rect 952 23942 1230 24006
rect 1294 23942 1300 24006
rect 952 22374 1300 23942
rect 2111 22950 2171 30291
rect 18904 30126 18980 31422
rect 18904 30094 18910 30126
rect 18909 30062 18910 30094
rect 18974 30094 18980 30126
rect 19312 31422 19318 31454
rect 19382 31454 19383 31486
rect 22576 31486 22652 31492
rect 19382 31422 19388 31454
rect 19312 30126 19388 31422
rect 22576 31422 22582 31486
rect 22646 31422 22652 31486
rect 22989 31486 23055 31487
rect 22989 31454 22990 31486
rect 21765 31214 21831 31215
rect 21765 31182 21766 31214
rect 21760 31150 21766 31182
rect 21830 31182 21831 31214
rect 22576 31214 22652 31422
rect 22576 31182 22582 31214
rect 21830 31150 21836 31182
rect 21760 30942 21836 31150
rect 22581 31150 22582 31182
rect 22646 31182 22652 31214
rect 22984 31422 22990 31454
rect 23054 31454 23055 31486
rect 23528 31486 23604 31492
rect 23054 31422 23060 31454
rect 22984 31214 23060 31422
rect 22646 31150 22647 31182
rect 22581 31149 22647 31150
rect 22984 31150 22990 31214
rect 23054 31150 23060 31214
rect 23528 31422 23534 31486
rect 23598 31422 23604 31486
rect 195165 31486 195231 31487
rect 195165 31454 195166 31486
rect 23528 31214 23604 31422
rect 195160 31422 195166 31454
rect 195230 31454 195231 31486
rect 195437 31486 195503 31487
rect 195437 31454 195438 31486
rect 195230 31422 195236 31454
rect 28565 31350 28631 31351
rect 28565 31318 28566 31350
rect 23528 31182 23534 31214
rect 22984 31144 23060 31150
rect 23533 31150 23534 31182
rect 23598 31182 23604 31214
rect 28560 31286 28566 31318
rect 28630 31318 28631 31350
rect 190133 31350 190199 31351
rect 190133 31318 190134 31350
rect 28630 31286 28636 31318
rect 23598 31150 23599 31182
rect 23533 31149 23599 31150
rect 21760 30878 21766 30942
rect 21830 30878 21836 30942
rect 21760 30872 21836 30878
rect 22984 31078 23060 31084
rect 22984 31014 22990 31078
rect 23054 31014 23060 31078
rect 23533 31078 23599 31079
rect 23533 31046 23534 31078
rect 22984 30806 23060 31014
rect 22984 30774 22990 30806
rect 22989 30742 22990 30774
rect 23054 30774 23060 30806
rect 23528 31014 23534 31046
rect 23598 31046 23599 31078
rect 28560 31078 28636 31286
rect 23598 31014 23604 31046
rect 23528 30806 23604 31014
rect 28560 31014 28566 31078
rect 28630 31014 28636 31078
rect 28560 31008 28636 31014
rect 190128 31286 190134 31318
rect 190198 31318 190199 31350
rect 190198 31286 190204 31318
rect 190128 31078 190204 31286
rect 195160 31214 195236 31422
rect 195160 31150 195166 31214
rect 195230 31150 195236 31214
rect 195160 31144 195236 31150
rect 195432 31422 195438 31454
rect 195502 31454 195503 31486
rect 195845 31486 195911 31487
rect 195845 31454 195846 31486
rect 195502 31422 195508 31454
rect 195432 31214 195508 31422
rect 195432 31150 195438 31214
rect 195502 31150 195508 31214
rect 195432 31144 195508 31150
rect 195840 31422 195846 31454
rect 195910 31454 195911 31486
rect 196248 31486 196324 31492
rect 195910 31422 195916 31454
rect 195840 31214 195916 31422
rect 195840 31150 195846 31214
rect 195910 31150 195916 31214
rect 196248 31422 196254 31486
rect 196318 31422 196324 31486
rect 196248 31214 196324 31422
rect 198832 31486 198908 31492
rect 198832 31422 198838 31486
rect 198902 31422 198908 31486
rect 199109 31486 199175 31487
rect 199109 31454 199110 31486
rect 196248 31182 196254 31214
rect 195840 31144 195916 31150
rect 196253 31150 196254 31182
rect 196318 31182 196324 31214
rect 196656 31214 196732 31220
rect 196318 31150 196319 31182
rect 196253 31149 196319 31150
rect 196656 31150 196662 31214
rect 196726 31150 196732 31214
rect 190128 31014 190134 31078
rect 190198 31014 190204 31078
rect 190128 31008 190204 31014
rect 195024 31078 195100 31084
rect 195024 31014 195030 31078
rect 195094 31014 195100 31078
rect 23054 30742 23055 30774
rect 22989 30741 23055 30742
rect 23528 30742 23534 30806
rect 23598 30742 23604 30806
rect 195024 30806 195100 31014
rect 195024 30774 195030 30806
rect 23528 30736 23604 30742
rect 195029 30742 195030 30774
rect 195094 30774 195100 30806
rect 195568 31078 195644 31084
rect 195568 31014 195574 31078
rect 195638 31014 195644 31078
rect 195568 30806 195644 31014
rect 196656 30942 196732 31150
rect 198832 31078 198908 31422
rect 198832 31046 198838 31078
rect 198837 31014 198838 31046
rect 198902 31046 198908 31078
rect 199104 31422 199110 31454
rect 199174 31454 199175 31486
rect 199784 31486 199860 31492
rect 199174 31422 199180 31454
rect 198902 31014 198903 31046
rect 198837 31013 198903 31014
rect 196656 30910 196662 30942
rect 196661 30878 196662 30910
rect 196726 30910 196732 30942
rect 196726 30878 196727 30910
rect 196661 30877 196727 30878
rect 195568 30774 195574 30806
rect 195094 30742 195095 30774
rect 195029 30741 195095 30742
rect 195573 30742 195574 30774
rect 195638 30774 195644 30806
rect 195638 30742 195639 30774
rect 195573 30741 195639 30742
rect 22032 30670 22108 30676
rect 22032 30606 22038 30670
rect 22102 30606 22108 30670
rect 21765 30398 21831 30399
rect 21765 30366 21766 30398
rect 18974 30062 18975 30094
rect 18909 30061 18975 30062
rect 19312 30062 19318 30126
rect 19382 30062 19388 30126
rect 19312 30056 19388 30062
rect 21760 30334 21766 30366
rect 21830 30366 21831 30398
rect 21830 30334 21836 30366
rect 21760 30126 21836 30334
rect 22032 30262 22108 30606
rect 22168 30670 22244 30676
rect 22168 30606 22174 30670
rect 22238 30606 22244 30670
rect 22581 30670 22647 30671
rect 22581 30638 22582 30670
rect 22168 30398 22244 30606
rect 22168 30366 22174 30398
rect 22173 30334 22174 30366
rect 22238 30366 22244 30398
rect 22576 30606 22582 30638
rect 22646 30638 22647 30670
rect 196248 30670 196324 30676
rect 22646 30606 22652 30638
rect 22576 30398 22652 30606
rect 196248 30606 196254 30670
rect 196318 30606 196324 30670
rect 22238 30334 22239 30366
rect 22173 30333 22239 30334
rect 22576 30334 22582 30398
rect 22646 30334 22652 30398
rect 22576 30328 22652 30334
rect 190128 30534 190204 30540
rect 190128 30470 190134 30534
rect 190198 30470 190204 30534
rect 22032 30230 22038 30262
rect 22037 30198 22038 30230
rect 22102 30230 22108 30262
rect 190128 30262 190204 30470
rect 196248 30398 196324 30606
rect 196248 30366 196254 30398
rect 196253 30334 196254 30366
rect 196318 30366 196324 30398
rect 196656 30398 196732 30404
rect 196318 30334 196319 30366
rect 196253 30333 196319 30334
rect 196656 30334 196662 30398
rect 196726 30334 196732 30398
rect 190128 30230 190134 30262
rect 22102 30198 22103 30230
rect 22037 30197 22103 30198
rect 190133 30198 190134 30230
rect 190198 30230 190204 30262
rect 190198 30198 190199 30230
rect 190133 30197 190199 30198
rect 21760 30062 21766 30126
rect 21830 30062 21836 30126
rect 196656 30126 196732 30334
rect 196656 30094 196662 30126
rect 21760 30056 21836 30062
rect 196661 30062 196662 30094
rect 196726 30094 196732 30126
rect 199104 30126 199180 31422
rect 196726 30062 196727 30094
rect 196661 30061 196727 30062
rect 199104 30062 199110 30126
rect 199174 30062 199180 30126
rect 199784 31422 199790 31486
rect 199854 31422 199860 31486
rect 199784 30126 199860 31422
rect 199784 30094 199790 30126
rect 199104 30056 199180 30062
rect 199789 30062 199790 30094
rect 199854 30094 199860 30126
rect 217464 30670 217812 32510
rect 217464 30606 217470 30670
rect 217534 30606 217812 30670
rect 199854 30062 199855 30094
rect 199789 30061 199855 30062
rect 18229 29990 18295 29991
rect 18229 29958 18230 29990
rect 18224 29926 18230 29958
rect 18294 29958 18295 29990
rect 18773 29990 18839 29991
rect 18773 29958 18774 29990
rect 18294 29926 18300 29958
rect 18224 29310 18300 29926
rect 18224 29246 18230 29310
rect 18294 29246 18300 29310
rect 18224 29240 18300 29246
rect 18768 29926 18774 29958
rect 18838 29958 18839 29990
rect 19312 29990 19388 29996
rect 18838 29926 18844 29958
rect 18768 29316 18844 29926
rect 19312 29926 19318 29990
rect 19382 29926 19388 29990
rect 19861 29990 19927 29991
rect 19861 29958 19862 29990
rect 18768 29310 18980 29316
rect 18768 29246 18910 29310
rect 18974 29246 18980 29310
rect 19312 29310 19388 29926
rect 19312 29278 19318 29310
rect 18768 29240 18980 29246
rect 19317 29246 19318 29278
rect 19382 29278 19388 29310
rect 19856 29926 19862 29958
rect 19926 29958 19927 29990
rect 21896 29990 21972 29996
rect 19926 29926 19932 29958
rect 19856 29310 19932 29926
rect 21896 29926 21902 29990
rect 21966 29926 21972 29990
rect 21896 29718 21972 29926
rect 21896 29686 21902 29718
rect 21901 29654 21902 29686
rect 21966 29686 21972 29718
rect 22440 29990 22516 29996
rect 22440 29926 22446 29990
rect 22510 29926 22516 29990
rect 23125 29990 23191 29991
rect 23125 29958 23126 29990
rect 22440 29718 22516 29926
rect 22440 29686 22446 29718
rect 21966 29654 21967 29686
rect 21901 29653 21967 29654
rect 22445 29654 22446 29686
rect 22510 29686 22516 29718
rect 23120 29926 23126 29958
rect 23190 29958 23191 29990
rect 23392 29990 23468 29996
rect 23190 29926 23196 29958
rect 23120 29718 23196 29926
rect 22510 29654 22511 29686
rect 22445 29653 22511 29654
rect 23120 29654 23126 29718
rect 23190 29654 23196 29718
rect 23392 29926 23398 29990
rect 23462 29926 23468 29990
rect 195165 29990 195231 29991
rect 195165 29958 195166 29990
rect 23392 29718 23468 29926
rect 23392 29686 23398 29718
rect 23120 29648 23196 29654
rect 23397 29654 23398 29686
rect 23462 29686 23468 29718
rect 195160 29926 195166 29958
rect 195230 29958 195231 29990
rect 195432 29990 195508 29996
rect 195230 29926 195236 29958
rect 195160 29718 195236 29926
rect 23462 29654 23463 29686
rect 23397 29653 23463 29654
rect 195160 29654 195166 29718
rect 195230 29654 195236 29718
rect 195432 29926 195438 29990
rect 195502 29926 195508 29990
rect 195845 29990 195911 29991
rect 195845 29958 195846 29990
rect 195432 29718 195508 29926
rect 195432 29686 195438 29718
rect 195160 29648 195236 29654
rect 195437 29654 195438 29686
rect 195502 29686 195508 29718
rect 195840 29926 195846 29958
rect 195910 29958 195911 29990
rect 196792 29990 196868 29996
rect 195910 29926 195916 29958
rect 195840 29718 195916 29926
rect 195502 29654 195503 29686
rect 195437 29653 195503 29654
rect 195840 29654 195846 29718
rect 195910 29654 195916 29718
rect 196792 29926 196798 29990
rect 196862 29926 196868 29990
rect 196792 29718 196868 29926
rect 196792 29686 196798 29718
rect 195840 29648 195916 29654
rect 196797 29654 196798 29686
rect 196862 29686 196868 29718
rect 199104 29990 199180 29996
rect 199104 29926 199110 29990
rect 199174 29926 199180 29990
rect 199381 29990 199447 29991
rect 199381 29958 199382 29990
rect 199104 29718 199180 29926
rect 199104 29686 199110 29718
rect 196862 29654 196863 29686
rect 196797 29653 196863 29654
rect 199109 29654 199110 29686
rect 199174 29686 199180 29718
rect 199376 29926 199382 29958
rect 199446 29958 199447 29990
rect 199784 29990 199996 29996
rect 199446 29926 199452 29958
rect 199174 29654 199175 29686
rect 199109 29653 199175 29654
rect 21901 29582 21967 29583
rect 21901 29550 21902 29582
rect 19382 29246 19383 29278
rect 19317 29245 19383 29246
rect 19856 29246 19862 29310
rect 19926 29246 19932 29310
rect 19856 29240 19932 29246
rect 21896 29518 21902 29550
rect 21966 29550 21967 29582
rect 22309 29582 22375 29583
rect 22309 29550 22310 29582
rect 21966 29518 21972 29550
rect 21896 29310 21972 29518
rect 21896 29246 21902 29310
rect 21966 29246 21972 29310
rect 21896 29240 21972 29246
rect 22304 29518 22310 29550
rect 22374 29550 22375 29582
rect 22717 29582 22783 29583
rect 22717 29550 22718 29582
rect 22374 29518 22380 29550
rect 22304 29310 22380 29518
rect 22304 29246 22310 29310
rect 22374 29246 22380 29310
rect 22304 29240 22380 29246
rect 22712 29518 22718 29550
rect 22782 29550 22783 29582
rect 22989 29582 23055 29583
rect 22989 29550 22990 29582
rect 22782 29518 22788 29550
rect 22712 29310 22788 29518
rect 22712 29246 22718 29310
rect 22782 29246 22788 29310
rect 22712 29240 22788 29246
rect 22984 29518 22990 29550
rect 23054 29550 23055 29582
rect 23397 29582 23463 29583
rect 23397 29550 23398 29582
rect 23054 29518 23060 29550
rect 22984 29310 23060 29518
rect 22984 29246 22990 29310
rect 23054 29246 23060 29310
rect 22984 29240 23060 29246
rect 23392 29518 23398 29550
rect 23462 29550 23463 29582
rect 195160 29582 195236 29588
rect 23462 29518 23468 29550
rect 23392 29310 23468 29518
rect 23392 29246 23398 29310
rect 23462 29246 23468 29310
rect 195160 29518 195166 29582
rect 195230 29518 195236 29582
rect 195160 29310 195236 29518
rect 195160 29278 195166 29310
rect 23392 29240 23468 29246
rect 195165 29246 195166 29278
rect 195230 29278 195236 29310
rect 195432 29582 195508 29588
rect 195432 29518 195438 29582
rect 195502 29518 195508 29582
rect 195432 29310 195508 29518
rect 195432 29278 195438 29310
rect 195230 29246 195231 29278
rect 195165 29245 195231 29246
rect 195437 29246 195438 29278
rect 195502 29278 195508 29310
rect 195840 29582 195916 29588
rect 195840 29518 195846 29582
rect 195910 29518 195916 29582
rect 195840 29310 195916 29518
rect 195840 29278 195846 29310
rect 195502 29246 195503 29278
rect 195437 29245 195503 29246
rect 195845 29246 195846 29278
rect 195910 29278 195916 29310
rect 196656 29582 196732 29588
rect 196656 29518 196662 29582
rect 196726 29518 196732 29582
rect 196656 29310 196732 29518
rect 196656 29278 196662 29310
rect 195910 29246 195911 29278
rect 195845 29245 195911 29246
rect 196661 29246 196662 29278
rect 196726 29278 196732 29310
rect 199376 29310 199452 29926
rect 196726 29246 196727 29278
rect 196661 29245 196727 29246
rect 199376 29246 199382 29310
rect 199446 29246 199452 29310
rect 199784 29926 199926 29990
rect 199990 29926 199996 29990
rect 200605 29990 200671 29991
rect 200605 29958 200606 29990
rect 199784 29920 199996 29926
rect 200600 29926 200606 29958
rect 200670 29958 200671 29990
rect 200670 29926 200676 29958
rect 199784 29310 199860 29920
rect 199784 29278 199790 29310
rect 199376 29240 199452 29246
rect 199789 29246 199790 29278
rect 199854 29278 199860 29310
rect 200600 29310 200676 29926
rect 199854 29246 199855 29278
rect 199789 29245 199855 29246
rect 200600 29246 200606 29310
rect 200670 29246 200676 29310
rect 200600 29240 200676 29246
rect 18224 29174 18300 29180
rect 18224 29110 18230 29174
rect 18294 29110 18300 29174
rect 18224 28494 18300 29110
rect 18904 29174 18980 29180
rect 18904 29110 18910 29174
rect 18974 29110 18980 29174
rect 18904 28630 18980 29110
rect 18904 28598 18910 28630
rect 18909 28566 18910 28598
rect 18974 28598 18980 28630
rect 19448 29174 19524 29180
rect 19448 29110 19454 29174
rect 19518 29110 19524 29174
rect 18974 28566 18975 28598
rect 18909 28565 18975 28566
rect 18224 28462 18230 28494
rect 18229 28430 18230 28462
rect 18294 28462 18300 28494
rect 19448 28494 19524 29110
rect 21760 29174 21836 29180
rect 21760 29110 21766 29174
rect 21830 29110 21836 29174
rect 22581 29174 22647 29175
rect 22581 29142 22582 29174
rect 21760 28902 21836 29110
rect 21760 28870 21766 28902
rect 21765 28838 21766 28870
rect 21830 28870 21836 28902
rect 22576 29110 22582 29142
rect 22646 29142 22647 29174
rect 23120 29174 23196 29180
rect 22646 29110 22652 29142
rect 22576 28902 22652 29110
rect 21830 28838 21831 28870
rect 21765 28837 21831 28838
rect 22576 28838 22582 28902
rect 22646 28838 22652 28902
rect 23120 29110 23126 29174
rect 23190 29110 23196 29174
rect 23533 29174 23599 29175
rect 23533 29142 23534 29174
rect 23120 28902 23196 29110
rect 23120 28870 23126 28902
rect 22576 28832 22652 28838
rect 23125 28838 23126 28870
rect 23190 28870 23196 28902
rect 23528 29110 23534 29142
rect 23598 29142 23599 29174
rect 195160 29174 195236 29180
rect 23598 29110 23604 29142
rect 23528 28902 23604 29110
rect 23190 28838 23191 28870
rect 23125 28837 23191 28838
rect 23528 28838 23534 28902
rect 23598 28838 23604 28902
rect 195160 29110 195166 29174
rect 195230 29110 195236 29174
rect 195437 29174 195503 29175
rect 195437 29142 195438 29174
rect 195160 28902 195236 29110
rect 195160 28870 195166 28902
rect 23528 28832 23604 28838
rect 195165 28838 195166 28870
rect 195230 28870 195236 28902
rect 195432 29110 195438 29142
rect 195502 29142 195503 29174
rect 195845 29174 195911 29175
rect 195845 29142 195846 29174
rect 195502 29110 195508 29142
rect 195432 28902 195508 29110
rect 195230 28838 195231 28870
rect 195165 28837 195231 28838
rect 195432 28838 195438 28902
rect 195502 28838 195508 28902
rect 195432 28832 195508 28838
rect 195840 29110 195846 29142
rect 195910 29142 195911 29174
rect 196248 29174 196324 29180
rect 195910 29110 195916 29142
rect 195840 28902 195916 29110
rect 195840 28838 195846 28902
rect 195910 28838 195916 28902
rect 196248 29110 196254 29174
rect 196318 29110 196324 29174
rect 196661 29174 196727 29175
rect 196661 29142 196662 29174
rect 196248 28902 196324 29110
rect 196248 28870 196254 28902
rect 195840 28832 195916 28838
rect 196253 28838 196254 28870
rect 196318 28870 196324 28902
rect 196656 29110 196662 29142
rect 196726 29142 196727 29174
rect 198837 29174 198903 29175
rect 198837 29142 198838 29174
rect 196726 29110 196732 29142
rect 196656 28902 196732 29110
rect 196318 28838 196319 28870
rect 196253 28837 196319 28838
rect 196656 28838 196662 28902
rect 196726 28838 196732 28902
rect 196656 28832 196732 28838
rect 198832 29110 198838 29142
rect 198902 29142 198903 29174
rect 199240 29174 199316 29180
rect 198902 29110 198908 29142
rect 19448 28462 19454 28494
rect 18294 28430 18295 28462
rect 18229 28429 18295 28430
rect 19453 28430 19454 28462
rect 19518 28462 19524 28494
rect 21896 28766 21972 28772
rect 21896 28702 21902 28766
rect 21966 28702 21972 28766
rect 21896 28494 21972 28702
rect 21896 28462 21902 28494
rect 19518 28430 19519 28462
rect 19453 28429 19519 28430
rect 21901 28430 21902 28462
rect 21966 28462 21972 28494
rect 22304 28766 22380 28772
rect 22304 28702 22310 28766
rect 22374 28702 22380 28766
rect 22304 28494 22380 28702
rect 22304 28462 22310 28494
rect 21966 28430 21967 28462
rect 21901 28429 21967 28430
rect 22309 28430 22310 28462
rect 22374 28462 22380 28494
rect 22712 28766 22788 28772
rect 22712 28702 22718 28766
rect 22782 28702 22788 28766
rect 22989 28766 23055 28767
rect 22989 28734 22990 28766
rect 22712 28494 22788 28702
rect 22712 28462 22718 28494
rect 22374 28430 22375 28462
rect 22309 28429 22375 28430
rect 22717 28430 22718 28462
rect 22782 28462 22788 28494
rect 22984 28702 22990 28734
rect 23054 28734 23055 28766
rect 23392 28766 23468 28772
rect 23054 28702 23060 28734
rect 22984 28494 23060 28702
rect 22782 28430 22783 28462
rect 22717 28429 22783 28430
rect 22984 28430 22990 28494
rect 23054 28430 23060 28494
rect 23392 28702 23398 28766
rect 23462 28702 23468 28766
rect 195029 28766 195095 28767
rect 195029 28734 195030 28766
rect 23392 28494 23468 28702
rect 23392 28462 23398 28494
rect 22984 28424 23060 28430
rect 23397 28430 23398 28462
rect 23462 28462 23468 28494
rect 195024 28702 195030 28734
rect 195094 28734 195095 28766
rect 195437 28766 195503 28767
rect 195437 28734 195438 28766
rect 195094 28702 195100 28734
rect 195024 28494 195100 28702
rect 23462 28430 23463 28462
rect 23397 28429 23463 28430
rect 195024 28430 195030 28494
rect 195094 28430 195100 28494
rect 195024 28424 195100 28430
rect 195432 28702 195438 28734
rect 195502 28734 195503 28766
rect 196792 28766 196868 28772
rect 195502 28702 195508 28734
rect 195432 28494 195508 28702
rect 195432 28430 195438 28494
rect 195502 28430 195508 28494
rect 196792 28702 196798 28766
rect 196862 28702 196868 28766
rect 196792 28494 196868 28702
rect 196792 28462 196798 28494
rect 195432 28424 195508 28430
rect 196797 28430 196798 28462
rect 196862 28462 196868 28494
rect 198832 28494 198908 29110
rect 196862 28430 196863 28462
rect 196797 28429 196863 28430
rect 198832 28430 198838 28494
rect 198902 28430 198908 28494
rect 199240 29110 199246 29174
rect 199310 29110 199316 29174
rect 199240 28494 199316 29110
rect 199240 28462 199246 28494
rect 198832 28424 198908 28430
rect 199245 28430 199246 28462
rect 199310 28462 199316 28494
rect 200464 29174 200540 29180
rect 200464 29110 200470 29174
rect 200534 29110 200540 29174
rect 200464 28494 200540 29110
rect 200464 28462 200470 28494
rect 199310 28430 199311 28462
rect 199245 28429 199311 28430
rect 200469 28430 200470 28462
rect 200534 28462 200540 28494
rect 217464 29038 217812 30606
rect 217464 28974 217470 29038
rect 217534 28974 217812 29038
rect 200534 28430 200535 28462
rect 200469 28429 200535 28430
rect 18088 28358 18164 28364
rect 18088 28294 18094 28358
rect 18158 28294 18164 28358
rect 18365 28358 18431 28359
rect 18365 28326 18366 28358
rect 18088 27678 18164 28294
rect 18360 28294 18366 28326
rect 18430 28326 18431 28358
rect 19045 28358 19111 28359
rect 19045 28326 19046 28358
rect 18430 28294 18436 28326
rect 18360 28086 18436 28294
rect 18360 28022 18366 28086
rect 18430 28022 18436 28086
rect 18360 28016 18436 28022
rect 19040 28294 19046 28326
rect 19110 28326 19111 28358
rect 19312 28358 19388 28364
rect 19110 28294 19116 28326
rect 18088 27646 18094 27678
rect 18093 27614 18094 27646
rect 18158 27646 18164 27678
rect 19040 27678 19116 28294
rect 19312 28294 19318 28358
rect 19382 28294 19388 28358
rect 19312 28086 19388 28294
rect 19312 28054 19318 28086
rect 19317 28022 19318 28054
rect 19382 28054 19388 28086
rect 19448 28358 19524 28364
rect 19448 28294 19454 28358
rect 19518 28294 19524 28358
rect 19861 28358 19927 28359
rect 19861 28326 19862 28358
rect 19382 28022 19383 28054
rect 19317 28021 19383 28022
rect 18158 27614 18159 27646
rect 18093 27613 18159 27614
rect 19040 27614 19046 27678
rect 19110 27614 19116 27678
rect 19448 27678 19524 28294
rect 19448 27646 19454 27678
rect 19040 27608 19116 27614
rect 19453 27614 19454 27646
rect 19518 27646 19524 27678
rect 19856 28294 19862 28326
rect 19926 28326 19927 28358
rect 21901 28358 21967 28359
rect 21901 28326 21902 28358
rect 19926 28294 19932 28326
rect 19856 27678 19932 28294
rect 21896 28294 21902 28326
rect 21966 28326 21967 28358
rect 22445 28358 22511 28359
rect 22445 28326 22446 28358
rect 21966 28294 21972 28326
rect 21896 28086 21972 28294
rect 21896 28022 21902 28086
rect 21966 28022 21972 28086
rect 21896 28016 21972 28022
rect 22440 28294 22446 28326
rect 22510 28326 22511 28358
rect 22984 28358 23060 28364
rect 22510 28294 22516 28326
rect 22440 28086 22516 28294
rect 22440 28022 22446 28086
rect 22510 28022 22516 28086
rect 22984 28294 22990 28358
rect 23054 28294 23060 28358
rect 23397 28358 23463 28359
rect 23397 28326 23398 28358
rect 22984 28086 23060 28294
rect 22984 28054 22990 28086
rect 22440 28016 22516 28022
rect 22989 28022 22990 28054
rect 23054 28054 23060 28086
rect 23392 28294 23398 28326
rect 23462 28326 23463 28358
rect 195160 28358 195236 28364
rect 23462 28294 23468 28326
rect 23392 28086 23468 28294
rect 23054 28022 23055 28054
rect 22989 28021 23055 28022
rect 23392 28022 23398 28086
rect 23462 28022 23468 28086
rect 195160 28294 195166 28358
rect 195230 28294 195236 28358
rect 195160 28086 195236 28294
rect 195160 28054 195166 28086
rect 23392 28016 23468 28022
rect 195165 28022 195166 28054
rect 195230 28054 195236 28086
rect 195432 28358 195508 28364
rect 195432 28294 195438 28358
rect 195502 28294 195508 28358
rect 196389 28358 196455 28359
rect 196389 28326 196390 28358
rect 195432 28086 195508 28294
rect 195432 28054 195438 28086
rect 195230 28022 195231 28054
rect 195165 28021 195231 28022
rect 195437 28022 195438 28054
rect 195502 28054 195508 28086
rect 196384 28294 196390 28326
rect 196454 28326 196455 28358
rect 196797 28358 196863 28359
rect 196797 28326 196798 28358
rect 196454 28294 196460 28326
rect 196384 28086 196460 28294
rect 195502 28022 195503 28054
rect 195437 28021 195503 28022
rect 196384 28022 196390 28086
rect 196454 28022 196460 28086
rect 196384 28016 196460 28022
rect 196792 28294 196798 28326
rect 196862 28326 196863 28358
rect 198968 28358 199044 28364
rect 196862 28294 196868 28326
rect 196792 28086 196868 28294
rect 196792 28022 196798 28086
rect 196862 28022 196868 28086
rect 196792 28016 196868 28022
rect 198968 28294 198974 28358
rect 199038 28294 199044 28358
rect 199381 28358 199447 28359
rect 199381 28326 199382 28358
rect 21765 27950 21831 27951
rect 21765 27918 21766 27950
rect 19518 27614 19519 27646
rect 19453 27613 19519 27614
rect 19856 27614 19862 27678
rect 19926 27614 19932 27678
rect 19856 27608 19932 27614
rect 21760 27886 21766 27918
rect 21830 27918 21831 27950
rect 22173 27950 22239 27951
rect 22173 27918 22174 27950
rect 21830 27886 21836 27918
rect 21760 27678 21836 27886
rect 21760 27614 21766 27678
rect 21830 27614 21836 27678
rect 21760 27608 21836 27614
rect 22168 27886 22174 27918
rect 22238 27918 22239 27950
rect 22581 27950 22647 27951
rect 22581 27918 22582 27950
rect 22238 27886 22244 27918
rect 22168 27678 22244 27886
rect 22168 27614 22174 27678
rect 22238 27614 22244 27678
rect 22168 27608 22244 27614
rect 22576 27886 22582 27918
rect 22646 27918 22647 27950
rect 23125 27950 23191 27951
rect 23125 27918 23126 27950
rect 22646 27886 22652 27918
rect 22576 27678 22652 27886
rect 22576 27614 22582 27678
rect 22646 27614 22652 27678
rect 22576 27608 22652 27614
rect 23120 27886 23126 27918
rect 23190 27918 23191 27950
rect 23392 27950 23468 27956
rect 23190 27886 23196 27918
rect 23120 27678 23196 27886
rect 23120 27614 23126 27678
rect 23190 27614 23196 27678
rect 23392 27886 23398 27950
rect 23462 27886 23468 27950
rect 195165 27950 195231 27951
rect 195165 27918 195166 27950
rect 23392 27678 23468 27886
rect 23392 27646 23398 27678
rect 23120 27608 23196 27614
rect 23397 27614 23398 27646
rect 23462 27646 23468 27678
rect 195160 27886 195166 27918
rect 195230 27918 195231 27950
rect 195432 27950 195508 27956
rect 195230 27886 195236 27918
rect 195160 27678 195236 27886
rect 23462 27614 23463 27646
rect 23397 27613 23463 27614
rect 195160 27614 195166 27678
rect 195230 27614 195236 27678
rect 195432 27886 195438 27950
rect 195502 27886 195508 27950
rect 195432 27678 195508 27886
rect 195432 27646 195438 27678
rect 195160 27608 195236 27614
rect 195437 27614 195438 27646
rect 195502 27646 195508 27678
rect 195976 27950 196052 27956
rect 195976 27886 195982 27950
rect 196046 27886 196052 27950
rect 195976 27678 196052 27886
rect 195976 27646 195982 27678
rect 195502 27614 195503 27646
rect 195437 27613 195503 27614
rect 195981 27614 195982 27646
rect 196046 27646 196052 27678
rect 196792 27950 196868 27956
rect 196792 27886 196798 27950
rect 196862 27886 196868 27950
rect 196792 27678 196868 27886
rect 196792 27646 196798 27678
rect 196046 27614 196047 27646
rect 195981 27613 196047 27614
rect 196797 27614 196798 27646
rect 196862 27646 196868 27678
rect 198968 27678 199044 28294
rect 198968 27646 198974 27678
rect 196862 27614 196863 27646
rect 196797 27613 196863 27614
rect 198973 27614 198974 27646
rect 199038 27646 199044 27678
rect 199376 28294 199382 28326
rect 199446 28326 199447 28358
rect 200464 28358 200540 28364
rect 199446 28294 199452 28326
rect 199376 27678 199452 28294
rect 199038 27614 199039 27646
rect 198973 27613 199039 27614
rect 199376 27614 199382 27678
rect 199446 27614 199452 27678
rect 200464 28294 200470 28358
rect 200534 28294 200540 28358
rect 200464 27678 200540 28294
rect 200464 27646 200470 27678
rect 199376 27608 199452 27614
rect 200469 27614 200470 27646
rect 200534 27646 200540 27678
rect 200534 27614 200535 27646
rect 200469 27613 200535 27614
rect 19453 27542 19519 27543
rect 19453 27510 19454 27542
rect 19448 27478 19454 27510
rect 19518 27510 19519 27542
rect 19720 27542 19796 27548
rect 19518 27478 19524 27510
rect 19448 26182 19524 27478
rect 19448 26118 19454 26182
rect 19518 26118 19524 26182
rect 19720 27478 19726 27542
rect 19790 27478 19796 27542
rect 22309 27542 22375 27543
rect 22309 27510 22310 27542
rect 19720 26182 19796 27478
rect 22304 27478 22310 27510
rect 22374 27510 22375 27542
rect 23120 27542 23196 27548
rect 22374 27478 22380 27510
rect 21901 27270 21967 27271
rect 21901 27238 21902 27270
rect 21896 27206 21902 27238
rect 21966 27238 21967 27270
rect 22304 27270 22380 27478
rect 21966 27206 21972 27238
rect 21896 26998 21972 27206
rect 22304 27206 22310 27270
rect 22374 27206 22380 27270
rect 23120 27478 23126 27542
rect 23190 27478 23196 27542
rect 23397 27542 23463 27543
rect 23397 27510 23398 27542
rect 23120 27270 23196 27478
rect 23120 27238 23126 27270
rect 22304 27200 22380 27206
rect 23125 27206 23126 27238
rect 23190 27238 23196 27270
rect 23392 27478 23398 27510
rect 23462 27510 23463 27542
rect 195024 27542 195100 27548
rect 23462 27478 23468 27510
rect 23392 27270 23468 27478
rect 23190 27206 23191 27238
rect 23125 27205 23191 27206
rect 23392 27206 23398 27270
rect 23462 27206 23468 27270
rect 195024 27478 195030 27542
rect 195094 27478 195100 27542
rect 195437 27542 195503 27543
rect 195437 27510 195438 27542
rect 195024 27270 195100 27478
rect 195024 27238 195030 27270
rect 23392 27200 23468 27206
rect 195029 27206 195030 27238
rect 195094 27238 195100 27270
rect 195432 27478 195438 27510
rect 195502 27510 195503 27542
rect 196389 27542 196455 27543
rect 196389 27510 196390 27542
rect 195502 27478 195508 27510
rect 195432 27270 195508 27478
rect 195094 27206 195095 27238
rect 195029 27205 195095 27206
rect 195432 27206 195438 27270
rect 195502 27206 195508 27270
rect 195432 27200 195508 27206
rect 196384 27478 196390 27510
rect 196454 27510 196455 27542
rect 200464 27542 200540 27548
rect 196454 27478 196460 27510
rect 196384 27270 196460 27478
rect 200464 27478 200470 27542
rect 200534 27478 200540 27542
rect 198968 27406 199044 27412
rect 198968 27342 198974 27406
rect 199038 27342 199044 27406
rect 196384 27206 196390 27270
rect 196454 27206 196460 27270
rect 196797 27270 196863 27271
rect 196797 27238 196798 27270
rect 196384 27200 196460 27206
rect 196792 27206 196798 27238
rect 196862 27238 196863 27270
rect 196862 27206 196868 27238
rect 21896 26934 21902 26998
rect 21966 26934 21972 26998
rect 21896 26928 21972 26934
rect 23120 27134 23196 27140
rect 23120 27070 23126 27134
rect 23190 27070 23196 27134
rect 23120 26862 23196 27070
rect 23120 26830 23126 26862
rect 23125 26798 23126 26830
rect 23190 26830 23196 26862
rect 23528 27134 23604 27140
rect 23528 27070 23534 27134
rect 23598 27070 23604 27134
rect 195165 27134 195231 27135
rect 195165 27102 195166 27134
rect 23528 26862 23604 27070
rect 23528 26830 23534 26862
rect 23190 26798 23191 26830
rect 23125 26797 23191 26798
rect 23533 26798 23534 26830
rect 23598 26830 23604 26862
rect 195160 27070 195166 27102
rect 195230 27102 195231 27134
rect 195568 27134 195644 27140
rect 195230 27070 195236 27102
rect 195160 26862 195236 27070
rect 23598 26798 23599 26830
rect 23533 26797 23599 26798
rect 195160 26798 195166 26862
rect 195230 26798 195236 26862
rect 195568 27070 195574 27134
rect 195638 27070 195644 27134
rect 195568 26862 195644 27070
rect 196792 26998 196868 27206
rect 196792 26934 196798 26998
rect 196862 26934 196868 26998
rect 196792 26928 196868 26934
rect 195568 26830 195574 26862
rect 195160 26792 195236 26798
rect 195573 26798 195574 26830
rect 195638 26830 195644 26862
rect 195638 26798 195639 26830
rect 195573 26797 195639 26798
rect 22173 26726 22239 26727
rect 22173 26694 22174 26726
rect 22168 26662 22174 26694
rect 22238 26694 22239 26726
rect 22440 26726 22516 26732
rect 22238 26662 22244 26694
rect 19720 26150 19726 26182
rect 19448 26112 19524 26118
rect 19725 26118 19726 26150
rect 19790 26150 19796 26182
rect 21896 26454 21972 26460
rect 21896 26390 21902 26454
rect 21966 26390 21972 26454
rect 21896 26182 21972 26390
rect 22168 26454 22244 26662
rect 22168 26390 22174 26454
rect 22238 26390 22244 26454
rect 22440 26662 22446 26726
rect 22510 26662 22516 26726
rect 22440 26454 22516 26662
rect 196384 26726 196460 26732
rect 196384 26662 196390 26726
rect 196454 26662 196460 26726
rect 28565 26590 28631 26591
rect 28565 26558 28566 26590
rect 22440 26422 22446 26454
rect 22168 26384 22244 26390
rect 22445 26390 22446 26422
rect 22510 26422 22516 26454
rect 28560 26526 28566 26558
rect 28630 26558 28631 26590
rect 190264 26590 190340 26596
rect 28630 26526 28636 26558
rect 22510 26390 22511 26422
rect 22445 26389 22511 26390
rect 28560 26318 28636 26526
rect 28560 26254 28566 26318
rect 28630 26254 28636 26318
rect 190264 26526 190270 26590
rect 190334 26526 190340 26590
rect 190264 26318 190340 26526
rect 196384 26454 196460 26662
rect 196384 26422 196390 26454
rect 196389 26390 196390 26422
rect 196454 26422 196460 26454
rect 196797 26454 196863 26455
rect 196797 26422 196798 26454
rect 196454 26390 196455 26422
rect 196389 26389 196455 26390
rect 196792 26390 196798 26422
rect 196862 26422 196863 26454
rect 196862 26390 196868 26422
rect 190264 26286 190270 26318
rect 28560 26248 28636 26254
rect 190269 26254 190270 26286
rect 190334 26286 190340 26318
rect 190334 26254 190335 26286
rect 190269 26253 190335 26254
rect 21896 26150 21902 26182
rect 19790 26118 19791 26150
rect 19725 26117 19791 26118
rect 21901 26118 21902 26150
rect 21966 26150 21972 26182
rect 28424 26182 28500 26188
rect 21966 26118 21967 26150
rect 21901 26117 21967 26118
rect 28424 26118 28430 26182
rect 28494 26118 28500 26182
rect 190269 26182 190335 26183
rect 190269 26150 190270 26182
rect 18632 26046 18708 26052
rect 18632 25982 18638 26046
rect 18702 25982 18708 26046
rect 21765 26046 21831 26047
rect 21765 26014 21766 26046
rect 18632 25366 18708 25982
rect 21760 25982 21766 26014
rect 21830 26014 21831 26046
rect 22168 26046 22244 26052
rect 21830 25982 21836 26014
rect 19448 25910 19524 25916
rect 19448 25846 19454 25910
rect 19518 25846 19524 25910
rect 18632 25334 18638 25366
rect 18637 25302 18638 25334
rect 18702 25334 18708 25366
rect 18768 25638 18844 25644
rect 18768 25574 18774 25638
rect 18838 25574 18844 25638
rect 19317 25638 19383 25639
rect 19317 25606 19318 25638
rect 18768 25366 18844 25574
rect 18768 25334 18774 25366
rect 18702 25302 18703 25334
rect 18637 25301 18703 25302
rect 18773 25302 18774 25334
rect 18838 25334 18844 25366
rect 19312 25574 19318 25606
rect 19382 25606 19383 25638
rect 19382 25574 19388 25606
rect 19312 25366 19388 25574
rect 18838 25302 18839 25334
rect 18773 25301 18839 25302
rect 19312 25302 19318 25366
rect 19382 25302 19388 25366
rect 19448 25366 19524 25846
rect 19720 25910 19796 25916
rect 19720 25846 19726 25910
rect 19790 25846 19796 25910
rect 19720 25502 19796 25846
rect 21760 25774 21836 25982
rect 21760 25710 21766 25774
rect 21830 25710 21836 25774
rect 22168 25982 22174 26046
rect 22238 25982 22244 26046
rect 22168 25774 22244 25982
rect 22168 25742 22174 25774
rect 21760 25704 21836 25710
rect 22173 25710 22174 25742
rect 22238 25742 22244 25774
rect 22576 26046 22652 26052
rect 22576 25982 22582 26046
rect 22646 25982 22652 26046
rect 22576 25774 22652 25982
rect 28424 25910 28500 26118
rect 28424 25878 28430 25910
rect 28429 25846 28430 25878
rect 28494 25878 28500 25910
rect 190264 26118 190270 26150
rect 190334 26150 190335 26182
rect 196792 26182 196868 26390
rect 190334 26118 190340 26150
rect 190264 25910 190340 26118
rect 196792 26118 196798 26182
rect 196862 26118 196868 26182
rect 198968 26182 199044 27342
rect 198968 26150 198974 26182
rect 196792 26112 196868 26118
rect 198973 26118 198974 26150
rect 199038 26150 199044 26182
rect 200464 26182 200540 27478
rect 200464 26150 200470 26182
rect 199038 26118 199039 26150
rect 198973 26117 199039 26118
rect 200469 26118 200470 26150
rect 200534 26150 200540 26182
rect 217464 27406 217812 28974
rect 217464 27342 217470 27406
rect 217534 27342 217812 27406
rect 200534 26118 200535 26150
rect 200469 26117 200535 26118
rect 196253 26046 196319 26047
rect 196253 26014 196254 26046
rect 28494 25846 28495 25878
rect 28429 25845 28495 25846
rect 190264 25846 190270 25910
rect 190334 25846 190340 25910
rect 190264 25840 190340 25846
rect 196248 25982 196254 26014
rect 196318 26014 196319 26046
rect 196656 26046 196732 26052
rect 196318 25982 196324 26014
rect 22576 25742 22582 25774
rect 22238 25710 22239 25742
rect 22173 25709 22239 25710
rect 22581 25710 22582 25742
rect 22646 25742 22652 25774
rect 28288 25774 28364 25780
rect 22646 25710 22647 25742
rect 22581 25709 22647 25710
rect 28288 25710 28294 25774
rect 28358 25710 28364 25774
rect 19720 25470 19726 25502
rect 19725 25438 19726 25470
rect 19790 25470 19796 25502
rect 21896 25638 21972 25644
rect 21896 25574 21902 25638
rect 21966 25574 21972 25638
rect 23125 25638 23191 25639
rect 23125 25606 23126 25638
rect 19790 25438 19791 25470
rect 19725 25437 19791 25438
rect 19448 25334 19454 25366
rect 19312 25296 19388 25302
rect 19453 25302 19454 25334
rect 19518 25334 19524 25366
rect 21896 25366 21972 25574
rect 21896 25334 21902 25366
rect 19518 25302 19519 25334
rect 19453 25301 19519 25302
rect 21901 25302 21902 25334
rect 21966 25334 21972 25366
rect 23120 25574 23126 25606
rect 23190 25606 23191 25638
rect 23392 25638 23468 25644
rect 23190 25574 23196 25606
rect 23120 25366 23196 25574
rect 21966 25302 21967 25334
rect 21901 25301 21967 25302
rect 23120 25302 23126 25366
rect 23190 25302 23196 25366
rect 23392 25574 23398 25638
rect 23462 25574 23468 25638
rect 23392 25366 23468 25574
rect 28288 25502 28364 25710
rect 196248 25774 196324 25982
rect 196248 25710 196254 25774
rect 196318 25710 196324 25774
rect 196656 25982 196662 26046
rect 196726 25982 196732 26046
rect 196656 25774 196732 25982
rect 199648 26046 199724 26052
rect 199648 25982 199654 26046
rect 199718 25982 199724 26046
rect 196656 25742 196662 25774
rect 196248 25704 196324 25710
rect 196661 25710 196662 25742
rect 196726 25742 196732 25774
rect 199376 25910 199452 25916
rect 199376 25846 199382 25910
rect 199446 25846 199452 25910
rect 196726 25710 196727 25742
rect 196661 25709 196727 25710
rect 28288 25470 28294 25502
rect 28293 25438 28294 25470
rect 28358 25470 28364 25502
rect 195024 25638 195100 25644
rect 195024 25574 195030 25638
rect 195094 25574 195100 25638
rect 28358 25438 28359 25470
rect 28293 25437 28359 25438
rect 23392 25334 23398 25366
rect 23120 25296 23196 25302
rect 23397 25302 23398 25334
rect 23462 25334 23468 25366
rect 195024 25366 195100 25574
rect 195024 25334 195030 25366
rect 23462 25302 23463 25334
rect 23397 25301 23463 25302
rect 195029 25302 195030 25334
rect 195094 25334 195100 25366
rect 195432 25638 195508 25644
rect 195432 25574 195438 25638
rect 195502 25574 195508 25638
rect 196661 25638 196727 25639
rect 196661 25606 196662 25638
rect 195432 25366 195508 25574
rect 195432 25334 195438 25366
rect 195094 25302 195095 25334
rect 195029 25301 195095 25302
rect 195437 25302 195438 25334
rect 195502 25334 195508 25366
rect 196656 25574 196662 25606
rect 196726 25606 196727 25638
rect 196726 25574 196732 25606
rect 196656 25366 196732 25574
rect 195502 25302 195503 25334
rect 195437 25301 195503 25302
rect 196656 25302 196662 25366
rect 196726 25302 196732 25366
rect 199376 25366 199452 25846
rect 199376 25334 199382 25366
rect 196656 25296 196732 25302
rect 199381 25302 199382 25334
rect 199446 25334 199452 25366
rect 199648 25366 199724 25982
rect 199648 25334 199654 25366
rect 199446 25302 199447 25334
rect 199381 25301 199447 25302
rect 199653 25302 199654 25334
rect 199718 25334 199724 25366
rect 200192 26046 200268 26052
rect 200192 25982 200198 26046
rect 200262 25982 200268 26046
rect 201285 26046 201351 26047
rect 201285 26014 201286 26046
rect 200192 25366 200268 25982
rect 200192 25334 200198 25366
rect 199718 25302 199719 25334
rect 199653 25301 199719 25302
rect 200197 25302 200198 25334
rect 200262 25334 200268 25366
rect 201280 25982 201286 26014
rect 201350 26014 201351 26046
rect 201350 25982 201356 26014
rect 201280 25366 201356 25982
rect 200262 25302 200263 25334
rect 200197 25301 200263 25302
rect 201280 25302 201286 25366
rect 201350 25302 201356 25366
rect 201280 25296 201356 25302
rect 217464 25774 217812 27342
rect 217464 25710 217470 25774
rect 217534 25710 217812 25774
rect 17136 25230 17212 25236
rect 17136 25166 17142 25230
rect 17206 25166 17212 25230
rect 17136 24006 17212 25166
rect 17136 23974 17142 24006
rect 17141 23942 17142 23974
rect 17206 23974 17212 24006
rect 17544 25230 17620 25236
rect 17544 25166 17550 25230
rect 17614 25166 17620 25230
rect 21901 25230 21967 25231
rect 21901 25198 21902 25230
rect 17206 23942 17207 23974
rect 17141 23941 17207 23942
rect 15237 23870 15303 23871
rect 15237 23838 15238 23870
rect 15232 23806 15238 23838
rect 15302 23838 15303 23870
rect 15302 23806 15308 23838
rect 2108 22949 2174 22950
rect 2108 22885 2109 22949
rect 2173 22885 2174 22949
rect 2108 22884 2174 22885
rect 952 22310 1230 22374
rect 1294 22310 1300 22374
rect 952 20742 1300 22310
rect 952 20678 1230 20742
rect 1294 20678 1300 20742
rect 952 18974 1300 20678
rect 15096 22510 15172 22516
rect 15096 22446 15102 22510
rect 15166 22446 15172 22510
rect 2725 20606 2791 20607
rect 2725 20574 2726 20606
rect 2720 20542 2726 20574
rect 2790 20574 2791 20606
rect 2790 20542 2796 20574
rect 2720 19790 2796 20542
rect 2720 19726 2726 19790
rect 2790 19726 2796 19790
rect 15096 19790 15172 22446
rect 15232 21150 15308 23806
rect 17544 22646 17620 25166
rect 17544 22614 17550 22646
rect 17549 22582 17550 22614
rect 17614 22614 17620 22646
rect 21896 25166 21902 25198
rect 21966 25198 21967 25230
rect 23397 25230 23463 25231
rect 23397 25198 23398 25230
rect 21966 25166 21972 25198
rect 17614 22582 17615 22614
rect 17549 22581 17615 22582
rect 21896 22374 21972 25166
rect 23392 25166 23398 25198
rect 23462 25198 23463 25230
rect 195024 25230 195100 25236
rect 23462 25166 23468 25198
rect 23392 24822 23468 25166
rect 23392 24758 23398 24822
rect 23462 24758 23468 24822
rect 23392 24752 23468 24758
rect 195024 25166 195030 25230
rect 195094 25166 195100 25230
rect 199381 25230 199447 25231
rect 199381 25198 199382 25230
rect 29925 24686 29991 24687
rect 29925 24654 29926 24686
rect 29920 24622 29926 24654
rect 29990 24654 29991 24686
rect 29990 24622 29996 24654
rect 21896 22310 21902 22374
rect 21966 22310 21972 22374
rect 21896 22304 21972 22310
rect 23120 24550 23196 24556
rect 23120 24486 23126 24550
rect 23190 24486 23196 24550
rect 15232 21086 15238 21150
rect 15302 21086 15308 21150
rect 15232 21080 15308 21086
rect 21760 22238 21836 22244
rect 21760 22174 21766 22238
rect 21830 22174 21836 22238
rect 15237 21014 15303 21015
rect 15237 20982 15238 21014
rect 15096 19758 15102 19790
rect 2720 19720 2796 19726
rect 15101 19726 15102 19758
rect 15166 19758 15172 19790
rect 15232 20950 15238 20982
rect 15302 20982 15303 21014
rect 15302 20950 15308 20982
rect 15166 19726 15167 19758
rect 15101 19725 15167 19726
rect 15101 19654 15167 19655
rect 15101 19622 15102 19654
rect 952 18910 1230 18974
rect 1294 18910 1300 18974
rect 952 17342 1300 18910
rect 952 17278 1230 17342
rect 1294 17278 1300 17342
rect 952 15574 1300 17278
rect 15096 19590 15102 19622
rect 15166 19622 15167 19654
rect 15166 19590 15172 19622
rect 15096 16934 15172 19590
rect 15232 18430 15308 20950
rect 20541 20878 20607 20879
rect 20541 20846 20542 20878
rect 15232 18366 15238 18430
rect 15302 18366 15308 18430
rect 15232 18360 15308 18366
rect 20536 20814 20542 20846
rect 20606 20846 20607 20878
rect 20606 20814 20612 20846
rect 15237 18158 15303 18159
rect 15237 18126 15238 18158
rect 15096 16870 15102 16934
rect 15166 16870 15172 16934
rect 15096 16864 15172 16870
rect 15232 18094 15238 18126
rect 15302 18126 15303 18158
rect 20536 18158 20612 20814
rect 21760 19518 21836 22174
rect 23120 21014 23196 24486
rect 29376 24414 29452 24420
rect 29376 24350 29382 24414
rect 29446 24350 29452 24414
rect 29376 23734 29452 24350
rect 29376 23702 29382 23734
rect 29381 23670 29382 23702
rect 29446 23702 29452 23734
rect 29446 23670 29447 23702
rect 29381 23669 29447 23670
rect 29653 23598 29719 23599
rect 29653 23566 29654 23598
rect 23120 20982 23126 21014
rect 23125 20950 23126 20982
rect 23190 20982 23196 21014
rect 29648 23534 29654 23566
rect 29718 23566 29719 23598
rect 29718 23534 29724 23566
rect 23190 20950 23191 20982
rect 23125 20949 23191 20950
rect 21760 19486 21766 19518
rect 21765 19454 21766 19486
rect 21830 19486 21836 19518
rect 21830 19454 21831 19486
rect 21765 19453 21831 19454
rect 21765 19382 21831 19383
rect 21765 19350 21766 19382
rect 15302 18094 15308 18126
rect 952 15510 1230 15574
rect 1294 15510 1300 15574
rect 952 13942 1300 15510
rect 15096 16798 15172 16804
rect 15096 16734 15102 16798
rect 15166 16734 15172 16798
rect 15096 14078 15172 16734
rect 15232 15574 15308 18094
rect 20536 18094 20542 18158
rect 20606 18094 20612 18158
rect 20536 18088 20612 18094
rect 21760 19318 21766 19350
rect 21830 19350 21831 19382
rect 21830 19318 21836 19350
rect 20405 18022 20471 18023
rect 20405 17990 20406 18022
rect 15232 15510 15238 15574
rect 15302 15510 15308 15574
rect 15232 15504 15308 15510
rect 20400 17958 20406 17990
rect 20470 17990 20471 18022
rect 20470 17958 20476 17990
rect 15096 14046 15102 14078
rect 15101 14014 15102 14046
rect 15166 14046 15172 14078
rect 15232 15438 15308 15444
rect 15232 15374 15238 15438
rect 15302 15374 15308 15438
rect 15166 14014 15167 14046
rect 15101 14013 15167 14014
rect 952 13878 1230 13942
rect 1294 13878 1300 13942
rect 952 12310 1300 13878
rect 15232 12718 15308 15374
rect 20400 15302 20476 17958
rect 21760 16798 21836 19318
rect 29648 18974 29724 23534
rect 29920 22238 29996 24622
rect 30600 24414 30676 24420
rect 30600 24350 30606 24414
rect 30670 24350 30676 24414
rect 30600 23734 30676 24350
rect 39304 24414 39380 24420
rect 39304 24350 39310 24414
rect 39374 24350 39380 24414
rect 30600 23702 30606 23734
rect 30605 23670 30606 23702
rect 30670 23702 30676 23734
rect 32232 24278 32308 24284
rect 32232 24214 32238 24278
rect 32302 24214 32308 24278
rect 32917 24278 32983 24279
rect 32917 24246 32918 24278
rect 32232 23734 32308 24214
rect 32232 23702 32238 23734
rect 30670 23670 30671 23702
rect 30605 23669 30671 23670
rect 32237 23670 32238 23702
rect 32302 23702 32308 23734
rect 32912 24214 32918 24246
rect 32982 24246 32983 24278
rect 33456 24278 33532 24284
rect 32982 24214 32988 24246
rect 32912 23734 32988 24214
rect 32302 23670 32303 23702
rect 32237 23669 32303 23670
rect 32912 23670 32918 23734
rect 32982 23670 32988 23734
rect 33456 24214 33462 24278
rect 33526 24214 33532 24278
rect 34141 24278 34207 24279
rect 34141 24246 34142 24278
rect 33456 23734 33532 24214
rect 33456 23702 33462 23734
rect 32912 23664 32988 23670
rect 33461 23670 33462 23702
rect 33526 23702 33532 23734
rect 34136 24214 34142 24246
rect 34206 24246 34207 24278
rect 35501 24278 35567 24279
rect 35501 24246 35502 24278
rect 34206 24214 34212 24246
rect 34136 23734 34212 24214
rect 33526 23670 33527 23702
rect 33461 23669 33527 23670
rect 34136 23670 34142 23734
rect 34206 23670 34212 23734
rect 34136 23664 34212 23670
rect 35496 24214 35502 24246
rect 35566 24246 35567 24278
rect 37128 24278 37204 24284
rect 35566 24214 35572 24246
rect 35496 23734 35572 24214
rect 35496 23670 35502 23734
rect 35566 23670 35572 23734
rect 37128 24214 37134 24278
rect 37198 24214 37204 24278
rect 37128 23734 37204 24214
rect 37128 23702 37134 23734
rect 35496 23664 35572 23670
rect 37133 23670 37134 23702
rect 37198 23702 37204 23734
rect 38488 24278 38564 24284
rect 38488 24214 38494 24278
rect 38558 24214 38564 24278
rect 38488 23734 38564 24214
rect 38488 23702 38494 23734
rect 37198 23670 37199 23702
rect 37133 23669 37199 23670
rect 38493 23670 38494 23702
rect 38558 23702 38564 23734
rect 39304 23734 39380 24350
rect 58072 24414 58148 24420
rect 58072 24350 58078 24414
rect 58142 24350 58148 24414
rect 39304 23702 39310 23734
rect 38558 23670 38559 23702
rect 38493 23669 38559 23670
rect 39309 23670 39310 23702
rect 39374 23702 39380 23734
rect 40936 24278 41012 24284
rect 40936 24214 40942 24278
rect 41006 24214 41012 24278
rect 41621 24278 41687 24279
rect 41621 24246 41622 24278
rect 40936 23734 41012 24214
rect 40936 23702 40942 23734
rect 39374 23670 39375 23702
rect 39309 23669 39375 23670
rect 40941 23670 40942 23702
rect 41006 23702 41012 23734
rect 41616 24214 41622 24246
rect 41686 24246 41687 24278
rect 42845 24278 42911 24279
rect 42845 24246 42846 24278
rect 41686 24214 41692 24246
rect 41616 23734 41692 24214
rect 41006 23670 41007 23702
rect 40941 23669 41007 23670
rect 41616 23670 41622 23734
rect 41686 23670 41692 23734
rect 41616 23664 41692 23670
rect 42840 24214 42846 24246
rect 42910 24246 42911 24278
rect 44608 24278 44684 24284
rect 42910 24214 42916 24246
rect 42840 23734 42916 24214
rect 42840 23670 42846 23734
rect 42910 23670 42916 23734
rect 44608 24214 44614 24278
rect 44678 24214 44684 24278
rect 45429 24278 45495 24279
rect 45429 24246 45430 24278
rect 44608 23734 44684 24214
rect 44608 23702 44614 23734
rect 42840 23664 42916 23670
rect 44613 23670 44614 23702
rect 44678 23702 44684 23734
rect 45424 24214 45430 24246
rect 45494 24246 45495 24278
rect 47192 24278 47268 24284
rect 45494 24214 45500 24246
rect 45424 23734 45500 24214
rect 44678 23670 44679 23702
rect 44613 23669 44679 23670
rect 45424 23670 45430 23734
rect 45494 23670 45500 23734
rect 47192 24214 47198 24278
rect 47262 24214 47268 24278
rect 47192 23734 47268 24214
rect 47192 23702 47198 23734
rect 45424 23664 45500 23670
rect 47197 23670 47198 23702
rect 47262 23702 47268 23734
rect 48008 24278 48084 24284
rect 48008 24214 48014 24278
rect 48078 24214 48084 24278
rect 48008 23734 48084 24214
rect 48008 23702 48014 23734
rect 47262 23670 47263 23702
rect 47197 23669 47263 23670
rect 48013 23670 48014 23702
rect 48078 23702 48084 23734
rect 49640 24278 49716 24284
rect 49640 24214 49646 24278
rect 49710 24214 49716 24278
rect 50461 24278 50527 24279
rect 50461 24246 50462 24278
rect 49640 23734 49716 24214
rect 49640 23702 49646 23734
rect 48078 23670 48079 23702
rect 48013 23669 48079 23670
rect 49645 23670 49646 23702
rect 49710 23702 49716 23734
rect 50456 24214 50462 24246
rect 50526 24246 50527 24278
rect 50864 24278 50940 24284
rect 50526 24214 50532 24246
rect 50456 23734 50532 24214
rect 49710 23670 49711 23702
rect 49645 23669 49711 23670
rect 50456 23670 50462 23734
rect 50526 23670 50532 23734
rect 50864 24214 50870 24278
rect 50934 24214 50940 24278
rect 51685 24278 51751 24279
rect 51685 24246 51686 24278
rect 50864 23734 50940 24214
rect 50864 23702 50870 23734
rect 50456 23664 50532 23670
rect 50869 23670 50870 23702
rect 50934 23702 50940 23734
rect 51680 24214 51686 24246
rect 51750 24246 51751 24278
rect 52909 24278 52975 24279
rect 52909 24246 52910 24278
rect 51750 24214 51756 24246
rect 51680 23734 51756 24214
rect 50934 23670 50935 23702
rect 50869 23669 50935 23670
rect 51680 23670 51686 23734
rect 51750 23670 51756 23734
rect 51680 23664 51756 23670
rect 52904 24214 52910 24246
rect 52974 24246 52975 24278
rect 54672 24278 54748 24284
rect 52974 24214 52980 24246
rect 52904 23734 52980 24214
rect 52904 23670 52910 23734
rect 52974 23670 52980 23734
rect 54672 24214 54678 24278
rect 54742 24214 54748 24278
rect 55357 24278 55423 24279
rect 55357 24246 55358 24278
rect 54672 23734 54748 24214
rect 54672 23702 54678 23734
rect 52904 23664 52980 23670
rect 54677 23670 54678 23702
rect 54742 23702 54748 23734
rect 55352 24214 55358 24246
rect 55422 24246 55423 24278
rect 56581 24278 56647 24279
rect 56581 24246 56582 24278
rect 55422 24214 55428 24246
rect 55352 23734 55428 24214
rect 54742 23670 54743 23702
rect 54677 23669 54743 23670
rect 55352 23670 55358 23734
rect 55422 23670 55428 23734
rect 55352 23664 55428 23670
rect 56576 24214 56582 24246
rect 56646 24246 56647 24278
rect 56646 24214 56652 24246
rect 56576 23734 56652 24214
rect 56576 23670 56582 23734
rect 56646 23670 56652 23734
rect 58072 23734 58148 24350
rect 114240 24414 114316 24420
rect 114240 24350 114246 24414
rect 114310 24350 114316 24414
rect 58072 23702 58078 23734
rect 56576 23664 56652 23670
rect 58077 23670 58078 23702
rect 58142 23702 58148 23734
rect 59704 24278 59780 24284
rect 59704 24214 59710 24278
rect 59774 24214 59780 24278
rect 60389 24278 60455 24279
rect 60389 24246 60390 24278
rect 59704 23734 59780 24214
rect 59704 23702 59710 23734
rect 58142 23670 58143 23702
rect 58077 23669 58143 23670
rect 59709 23670 59710 23702
rect 59774 23702 59780 23734
rect 60384 24214 60390 24246
rect 60454 24246 60455 24278
rect 61613 24278 61679 24279
rect 61613 24246 61614 24278
rect 60454 24214 60460 24246
rect 60384 23734 60460 24214
rect 59774 23670 59775 23702
rect 59709 23669 59775 23670
rect 60384 23670 60390 23734
rect 60454 23670 60460 23734
rect 60384 23664 60460 23670
rect 61608 24214 61614 24246
rect 61678 24246 61679 24278
rect 62152 24278 62228 24284
rect 61678 24214 61684 24246
rect 61608 23734 61684 24214
rect 61608 23670 61614 23734
rect 61678 23670 61684 23734
rect 62152 24214 62158 24278
rect 62222 24214 62228 24278
rect 62837 24278 62903 24279
rect 62837 24246 62838 24278
rect 62152 23734 62228 24214
rect 62152 23702 62158 23734
rect 61608 23664 61684 23670
rect 62157 23670 62158 23702
rect 62222 23702 62228 23734
rect 62832 24214 62838 24246
rect 62902 24246 62903 24278
rect 64061 24278 64127 24279
rect 64061 24246 64062 24278
rect 62902 24214 62908 24246
rect 62832 23734 62908 24214
rect 62222 23670 62223 23702
rect 62157 23669 62223 23670
rect 62832 23670 62838 23734
rect 62902 23670 62908 23734
rect 62832 23664 62908 23670
rect 64056 24214 64062 24246
rect 64126 24246 64127 24278
rect 66645 24278 66711 24279
rect 66645 24246 66646 24278
rect 64126 24214 64132 24246
rect 64056 23734 64132 24214
rect 64056 23670 64062 23734
rect 64126 23670 64132 23734
rect 64056 23664 64132 23670
rect 66640 24214 66646 24246
rect 66710 24246 66711 24278
rect 67869 24278 67935 24279
rect 67869 24246 67870 24278
rect 66710 24214 66716 24246
rect 66640 23734 66716 24214
rect 66640 23670 66646 23734
rect 66710 23670 66716 23734
rect 66640 23664 66716 23670
rect 67864 24214 67870 24246
rect 67934 24246 67935 24278
rect 68408 24278 68484 24284
rect 67934 24214 67940 24246
rect 67864 23734 67940 24214
rect 67864 23670 67870 23734
rect 67934 23670 67940 23734
rect 68408 24214 68414 24278
rect 68478 24214 68484 24278
rect 69093 24278 69159 24279
rect 69093 24246 69094 24278
rect 68408 23734 68484 24214
rect 68408 23702 68414 23734
rect 67864 23664 67940 23670
rect 68413 23670 68414 23702
rect 68478 23702 68484 23734
rect 69088 24214 69094 24246
rect 69158 24246 69159 24278
rect 69632 24278 69708 24284
rect 69158 24214 69164 24246
rect 69088 23734 69164 24214
rect 68478 23670 68479 23702
rect 68413 23669 68479 23670
rect 69088 23670 69094 23734
rect 69158 23670 69164 23734
rect 69632 24214 69638 24278
rect 69702 24214 69708 24278
rect 70317 24278 70383 24279
rect 70317 24246 70318 24278
rect 69632 23734 69708 24214
rect 69632 23702 69638 23734
rect 69088 23664 69164 23670
rect 69637 23670 69638 23702
rect 69702 23702 69708 23734
rect 70312 24214 70318 24246
rect 70382 24246 70383 24278
rect 70856 24278 70932 24284
rect 70382 24214 70388 24246
rect 70312 23734 70388 24214
rect 69702 23670 69703 23702
rect 69637 23669 69703 23670
rect 70312 23670 70318 23734
rect 70382 23670 70388 23734
rect 70856 24214 70862 24278
rect 70926 24214 70932 24278
rect 71677 24278 71743 24279
rect 71677 24246 71678 24278
rect 70856 23734 70932 24214
rect 70856 23702 70862 23734
rect 70312 23664 70388 23670
rect 70861 23670 70862 23702
rect 70926 23702 70932 23734
rect 71672 24214 71678 24246
rect 71742 24246 71743 24278
rect 73440 24278 73516 24284
rect 71742 24214 71748 24246
rect 71672 23734 71748 24214
rect 70926 23670 70927 23702
rect 70861 23669 70927 23670
rect 71672 23670 71678 23734
rect 71742 23670 71748 23734
rect 73440 24214 73446 24278
rect 73510 24214 73516 24278
rect 73440 23734 73516 24214
rect 73440 23702 73446 23734
rect 71672 23664 71748 23670
rect 73445 23670 73446 23702
rect 73510 23702 73516 23734
rect 74664 24278 74740 24284
rect 74664 24214 74670 24278
rect 74734 24214 74740 24278
rect 74664 23734 74740 24214
rect 74664 23702 74670 23734
rect 73510 23670 73511 23702
rect 73445 23669 73511 23670
rect 74669 23670 74670 23702
rect 74734 23702 74740 23734
rect 75208 24278 75284 24284
rect 75208 24214 75214 24278
rect 75278 24214 75284 24278
rect 75208 23734 75284 24214
rect 75208 23702 75214 23734
rect 74734 23670 74735 23702
rect 74669 23669 74735 23670
rect 75213 23670 75214 23702
rect 75278 23702 75284 23734
rect 75888 24278 75964 24284
rect 75888 24214 75894 24278
rect 75958 24214 75964 24278
rect 76573 24278 76639 24279
rect 76573 24246 76574 24278
rect 75888 23734 75964 24214
rect 75888 23702 75894 23734
rect 75278 23670 75279 23702
rect 75213 23669 75279 23670
rect 75893 23670 75894 23702
rect 75958 23702 75964 23734
rect 76568 24214 76574 24246
rect 76638 24246 76639 24278
rect 78336 24278 78412 24284
rect 76638 24214 76644 24246
rect 76568 23734 76644 24214
rect 75958 23670 75959 23702
rect 75893 23669 75959 23670
rect 76568 23670 76574 23734
rect 76638 23670 76644 23734
rect 78336 24214 78342 24278
rect 78406 24214 78412 24278
rect 78336 23734 78412 24214
rect 78336 23702 78342 23734
rect 76568 23664 76644 23670
rect 78341 23670 78342 23702
rect 78406 23702 78412 23734
rect 79560 24278 79636 24284
rect 79560 24214 79566 24278
rect 79630 24214 79636 24278
rect 79560 23734 79636 24214
rect 79560 23702 79566 23734
rect 78406 23670 78407 23702
rect 78341 23669 78407 23670
rect 79565 23670 79566 23702
rect 79630 23702 79636 23734
rect 80512 24278 80588 24284
rect 80512 24214 80518 24278
rect 80582 24214 80588 24278
rect 80512 23734 80588 24214
rect 80512 23702 80518 23734
rect 79630 23670 79631 23702
rect 79565 23669 79631 23670
rect 80517 23670 80518 23702
rect 80582 23702 80588 23734
rect 82008 24278 82084 24284
rect 82008 24214 82014 24278
rect 82078 24214 82084 24278
rect 82008 23734 82084 24214
rect 82008 23702 82014 23734
rect 80582 23670 80583 23702
rect 80517 23669 80583 23670
rect 82013 23670 82014 23702
rect 82078 23702 82084 23734
rect 83368 24278 83444 24284
rect 83368 24214 83374 24278
rect 83438 24214 83444 24278
rect 83368 23734 83444 24214
rect 83368 23702 83374 23734
rect 82078 23670 82079 23702
rect 82013 23669 82079 23670
rect 83373 23670 83374 23702
rect 83438 23702 83444 23734
rect 84592 24278 84668 24284
rect 84592 24214 84598 24278
rect 84662 24214 84668 24278
rect 85685 24278 85751 24279
rect 85685 24246 85686 24278
rect 84592 23734 84668 24214
rect 84592 23702 84598 23734
rect 83438 23670 83439 23702
rect 83373 23669 83439 23670
rect 84597 23670 84598 23702
rect 84662 23702 84668 23734
rect 85680 24214 85686 24246
rect 85750 24246 85751 24278
rect 86501 24278 86567 24279
rect 86501 24246 86502 24278
rect 85750 24214 85756 24246
rect 85680 23734 85756 24214
rect 84662 23670 84663 23702
rect 84597 23669 84663 23670
rect 85680 23670 85686 23734
rect 85750 23670 85756 23734
rect 85680 23664 85756 23670
rect 86496 24214 86502 24246
rect 86566 24246 86567 24278
rect 88400 24278 88476 24284
rect 86566 24214 86572 24246
rect 86496 23734 86572 24214
rect 86496 23670 86502 23734
rect 86566 23670 86572 23734
rect 88400 24214 88406 24278
rect 88470 24214 88476 24278
rect 89085 24278 89151 24279
rect 89085 24246 89086 24278
rect 88400 23734 88476 24214
rect 88400 23702 88406 23734
rect 86496 23664 86572 23670
rect 88405 23670 88406 23702
rect 88470 23702 88476 23734
rect 89080 24214 89086 24246
rect 89150 24246 89151 24278
rect 89765 24278 89831 24279
rect 89765 24246 89766 24278
rect 89150 24214 89156 24246
rect 89080 23734 89156 24214
rect 88470 23670 88471 23702
rect 88405 23669 88471 23670
rect 89080 23670 89086 23734
rect 89150 23670 89156 23734
rect 89080 23664 89156 23670
rect 89760 24214 89766 24246
rect 89830 24246 89831 24278
rect 92072 24278 92148 24284
rect 89830 24214 89836 24246
rect 89760 23734 89836 24214
rect 89760 23670 89766 23734
rect 89830 23670 89836 23734
rect 92072 24214 92078 24278
rect 92142 24214 92148 24278
rect 92072 23734 92148 24214
rect 92072 23702 92078 23734
rect 89760 23664 89836 23670
rect 92077 23670 92078 23702
rect 92142 23702 92148 23734
rect 94656 24278 94732 24284
rect 94656 24214 94662 24278
rect 94726 24214 94732 24278
rect 95341 24278 95407 24279
rect 95341 24246 95342 24278
rect 94656 23734 94732 24214
rect 94656 23702 94662 23734
rect 92142 23670 92143 23702
rect 92077 23669 92143 23670
rect 94661 23670 94662 23702
rect 94726 23702 94732 23734
rect 95336 24214 95342 24246
rect 95406 24246 95407 24278
rect 95744 24278 95820 24284
rect 95406 24214 95412 24246
rect 95336 23734 95412 24214
rect 94726 23670 94727 23702
rect 94661 23669 94727 23670
rect 95336 23670 95342 23734
rect 95406 23670 95412 23734
rect 95744 24214 95750 24278
rect 95814 24214 95820 24278
rect 95744 23734 95820 24214
rect 95744 23702 95750 23734
rect 95336 23664 95412 23670
rect 95749 23670 95750 23702
rect 95814 23702 95820 23734
rect 97104 24278 97180 24284
rect 97104 24214 97110 24278
rect 97174 24214 97180 24278
rect 97789 24278 97855 24279
rect 97789 24246 97790 24278
rect 97104 23734 97180 24214
rect 97104 23702 97110 23734
rect 95814 23670 95815 23702
rect 95749 23669 95815 23670
rect 97109 23670 97110 23702
rect 97174 23702 97180 23734
rect 97784 24214 97790 24246
rect 97854 24246 97855 24278
rect 100776 24278 100852 24284
rect 97854 24214 97860 24246
rect 97784 23734 97860 24214
rect 97174 23670 97175 23702
rect 97109 23669 97175 23670
rect 97784 23670 97790 23734
rect 97854 23670 97860 23734
rect 100776 24214 100782 24278
rect 100846 24214 100852 24278
rect 101597 24278 101663 24279
rect 101597 24246 101598 24278
rect 100776 23734 100852 24214
rect 100776 23702 100782 23734
rect 97784 23664 97860 23670
rect 100781 23670 100782 23702
rect 100846 23702 100852 23734
rect 101592 24214 101598 24246
rect 101662 24246 101663 24278
rect 102136 24278 102212 24284
rect 101662 24214 101668 24246
rect 101592 23734 101668 24214
rect 100846 23670 100847 23702
rect 100781 23669 100847 23670
rect 101592 23670 101598 23734
rect 101662 23670 101668 23734
rect 102136 24214 102142 24278
rect 102206 24214 102212 24278
rect 102136 23734 102212 24214
rect 102136 23702 102142 23734
rect 101592 23664 101668 23670
rect 102141 23670 102142 23702
rect 102206 23702 102212 23734
rect 103360 24278 103436 24284
rect 103360 24214 103366 24278
rect 103430 24214 103436 24278
rect 104045 24278 104111 24279
rect 104045 24246 104046 24278
rect 103360 23734 103436 24214
rect 103360 23702 103366 23734
rect 102206 23670 102207 23702
rect 102141 23669 102207 23670
rect 103365 23670 103366 23702
rect 103430 23702 103436 23734
rect 104040 24214 104046 24246
rect 104110 24246 104111 24278
rect 104584 24278 104660 24284
rect 104110 24214 104116 24246
rect 104040 23734 104116 24214
rect 103430 23670 103431 23702
rect 103365 23669 103431 23670
rect 104040 23670 104046 23734
rect 104110 23670 104116 23734
rect 104584 24214 104590 24278
rect 104654 24214 104660 24278
rect 105269 24278 105335 24279
rect 105269 24246 105270 24278
rect 104584 23734 104660 24214
rect 104584 23702 104590 23734
rect 104040 23664 104116 23670
rect 104589 23670 104590 23702
rect 104654 23702 104660 23734
rect 105264 24214 105270 24246
rect 105334 24246 105335 24278
rect 109616 24278 109692 24284
rect 105334 24214 105340 24246
rect 105264 23734 105340 24214
rect 104654 23670 104655 23702
rect 104589 23669 104655 23670
rect 105264 23670 105270 23734
rect 105334 23670 105340 23734
rect 109616 24214 109622 24278
rect 109686 24214 109692 24278
rect 110301 24278 110367 24279
rect 110301 24246 110302 24278
rect 109616 23734 109692 24214
rect 109616 23702 109622 23734
rect 105264 23664 105340 23670
rect 109621 23670 109622 23702
rect 109686 23702 109692 23734
rect 110296 24214 110302 24246
rect 110366 24246 110367 24278
rect 110840 24278 110916 24284
rect 110366 24214 110372 24246
rect 110296 23734 110372 24214
rect 109686 23670 109687 23702
rect 109621 23669 109687 23670
rect 110296 23670 110302 23734
rect 110366 23670 110372 23734
rect 110840 24214 110846 24278
rect 110910 24214 110916 24278
rect 111525 24278 111591 24279
rect 111525 24246 111526 24278
rect 110840 23734 110916 24214
rect 110840 23702 110846 23734
rect 110296 23664 110372 23670
rect 110845 23670 110846 23702
rect 110910 23702 110916 23734
rect 111520 24214 111526 24246
rect 111590 24246 111591 24278
rect 112749 24278 112815 24279
rect 112749 24246 112750 24278
rect 111590 24214 111596 24246
rect 111520 23734 111596 24214
rect 110910 23670 110911 23702
rect 110845 23669 110911 23670
rect 111520 23670 111526 23734
rect 111590 23670 111596 23734
rect 111520 23664 111596 23670
rect 112744 24214 112750 24246
rect 112814 24246 112815 24278
rect 113288 24278 113364 24284
rect 112814 24214 112820 24246
rect 112744 23734 112820 24214
rect 112744 23670 112750 23734
rect 112814 23670 112820 23734
rect 113288 24214 113294 24278
rect 113358 24214 113364 24278
rect 113288 23734 113364 24214
rect 113288 23702 113294 23734
rect 112744 23664 112820 23670
rect 113293 23670 113294 23702
rect 113358 23702 113364 23734
rect 114240 23734 114316 24350
rect 136680 24414 136756 24420
rect 136680 24350 136686 24414
rect 136750 24350 136756 24414
rect 115333 24278 115399 24279
rect 115333 24246 115334 24278
rect 114240 23702 114246 23734
rect 113358 23670 113359 23702
rect 113293 23669 113359 23670
rect 114245 23670 114246 23702
rect 114310 23702 114316 23734
rect 115328 24214 115334 24246
rect 115398 24246 115399 24278
rect 117096 24278 117172 24284
rect 115398 24214 115404 24246
rect 115328 23734 115404 24214
rect 114310 23670 114311 23702
rect 114245 23669 114311 23670
rect 115328 23670 115334 23734
rect 115398 23670 115404 23734
rect 117096 24214 117102 24278
rect 117166 24214 117172 24278
rect 117096 23734 117172 24214
rect 117096 23702 117102 23734
rect 115328 23664 115404 23670
rect 117101 23670 117102 23702
rect 117166 23702 117172 23734
rect 117640 24278 117716 24284
rect 117640 24214 117646 24278
rect 117710 24214 117716 24278
rect 119005 24278 119071 24279
rect 119005 24246 119006 24278
rect 117640 23734 117716 24214
rect 117640 23702 117646 23734
rect 117166 23670 117167 23702
rect 117101 23669 117167 23670
rect 117645 23670 117646 23702
rect 117710 23702 117716 23734
rect 119000 24214 119006 24246
rect 119070 24246 119071 24278
rect 120229 24278 120295 24279
rect 120229 24246 120230 24278
rect 119070 24214 119076 24246
rect 119000 23734 119076 24214
rect 117710 23670 117711 23702
rect 117645 23669 117711 23670
rect 119000 23670 119006 23734
rect 119070 23670 119076 23734
rect 119000 23664 119076 23670
rect 120224 24214 120230 24246
rect 120294 24246 120295 24278
rect 121992 24278 122068 24284
rect 120294 24214 120300 24246
rect 120224 23734 120300 24214
rect 120224 23670 120230 23734
rect 120294 23670 120300 23734
rect 121992 24214 121998 24278
rect 122062 24214 122068 24278
rect 121992 23734 122068 24214
rect 121992 23702 121998 23734
rect 120224 23664 120300 23670
rect 121997 23670 121998 23702
rect 122062 23702 122068 23734
rect 122944 24278 123020 24284
rect 122944 24214 122950 24278
rect 123014 24214 123020 24278
rect 122944 23734 123020 24214
rect 122944 23702 122950 23734
rect 122062 23670 122063 23702
rect 121997 23669 122063 23670
rect 122949 23670 122950 23702
rect 123014 23702 123020 23734
rect 123896 24278 123972 24284
rect 123896 24214 123902 24278
rect 123966 24214 123972 24278
rect 123896 23734 123972 24214
rect 123896 23702 123902 23734
rect 123014 23670 123015 23702
rect 122949 23669 123015 23670
rect 123901 23670 123902 23702
rect 123966 23702 123972 23734
rect 124440 24278 124516 24284
rect 124440 24214 124446 24278
rect 124510 24214 124516 24278
rect 124440 23734 124516 24214
rect 124440 23702 124446 23734
rect 123966 23670 123967 23702
rect 123901 23669 123967 23670
rect 124445 23670 124446 23702
rect 124510 23702 124516 23734
rect 125800 24278 125876 24284
rect 125800 24214 125806 24278
rect 125870 24214 125876 24278
rect 125800 23734 125876 24214
rect 125800 23702 125806 23734
rect 124510 23670 124511 23702
rect 124445 23669 124511 23670
rect 125805 23670 125806 23702
rect 125870 23702 125876 23734
rect 127024 24278 127100 24284
rect 127024 24214 127030 24278
rect 127094 24214 127100 24278
rect 128933 24278 128999 24279
rect 128933 24246 128934 24278
rect 127024 23734 127100 24214
rect 127024 23702 127030 23734
rect 125870 23670 125871 23702
rect 125805 23669 125871 23670
rect 127029 23670 127030 23702
rect 127094 23702 127100 23734
rect 128928 24214 128934 24246
rect 128998 24246 128999 24278
rect 130293 24278 130359 24279
rect 130293 24246 130294 24278
rect 128998 24214 129004 24246
rect 128928 23734 129004 24214
rect 127094 23670 127095 23702
rect 127029 23669 127095 23670
rect 128928 23670 128934 23734
rect 128998 23670 129004 23734
rect 128928 23664 129004 23670
rect 130288 24214 130294 24246
rect 130358 24246 130359 24278
rect 131648 24278 131724 24284
rect 130358 24214 130364 24246
rect 130288 23734 130364 24214
rect 130288 23670 130294 23734
rect 130358 23670 130364 23734
rect 131648 24214 131654 24278
rect 131718 24214 131724 24278
rect 131648 23734 131724 24214
rect 131648 23702 131654 23734
rect 130288 23664 130364 23670
rect 131653 23670 131654 23702
rect 131718 23702 131724 23734
rect 133280 24278 133356 24284
rect 133280 24214 133286 24278
rect 133350 24214 133356 24278
rect 133280 23734 133356 24214
rect 133280 23702 133286 23734
rect 131718 23670 131719 23702
rect 131653 23669 131719 23670
rect 133285 23670 133286 23702
rect 133350 23702 133356 23734
rect 134504 24278 134580 24284
rect 134504 24214 134510 24278
rect 134574 24214 134580 24278
rect 135189 24278 135255 24279
rect 135189 24246 135190 24278
rect 134504 23734 134580 24214
rect 134504 23702 134510 23734
rect 133350 23670 133351 23702
rect 133285 23669 133351 23670
rect 134509 23670 134510 23702
rect 134574 23702 134580 23734
rect 135184 24214 135190 24246
rect 135254 24246 135255 24278
rect 135728 24278 135804 24284
rect 135254 24214 135260 24246
rect 135184 23734 135260 24214
rect 134574 23670 134575 23702
rect 134509 23669 134575 23670
rect 135184 23670 135190 23734
rect 135254 23670 135260 23734
rect 135728 24214 135734 24278
rect 135798 24214 135804 24278
rect 135728 23734 135804 24214
rect 135728 23702 135734 23734
rect 135184 23664 135260 23670
rect 135733 23670 135734 23702
rect 135798 23702 135804 23734
rect 136680 23734 136756 24350
rect 145384 24414 145460 24420
rect 145384 24350 145390 24414
rect 145454 24350 145460 24414
rect 136680 23702 136686 23734
rect 135798 23670 135799 23702
rect 135733 23669 135799 23670
rect 136685 23670 136686 23702
rect 136750 23702 136756 23734
rect 138176 24278 138252 24284
rect 138176 24214 138182 24278
rect 138246 24214 138252 24278
rect 138176 23734 138252 24214
rect 138176 23702 138182 23734
rect 136750 23670 136751 23702
rect 136685 23669 136751 23670
rect 138181 23670 138182 23702
rect 138246 23702 138252 23734
rect 139536 24278 139612 24284
rect 139536 24214 139542 24278
rect 139606 24214 139612 24278
rect 140221 24278 140287 24279
rect 140221 24246 140222 24278
rect 139536 23734 139612 24214
rect 139536 23702 139542 23734
rect 138246 23670 138247 23702
rect 138181 23669 138247 23670
rect 139541 23670 139542 23702
rect 139606 23702 139612 23734
rect 140216 24214 140222 24246
rect 140286 24246 140287 24278
rect 141853 24278 141919 24279
rect 141853 24246 141854 24278
rect 140286 24214 140292 24246
rect 140216 23734 140292 24214
rect 139606 23670 139607 23702
rect 139541 23669 139607 23670
rect 140216 23670 140222 23734
rect 140286 23670 140292 23734
rect 140216 23664 140292 23670
rect 141848 24214 141854 24246
rect 141918 24246 141919 24278
rect 143208 24278 143284 24284
rect 141918 24214 141924 24246
rect 141848 23734 141924 24214
rect 141848 23670 141854 23734
rect 141918 23670 141924 23734
rect 143208 24214 143214 24278
rect 143278 24214 143284 24278
rect 144029 24278 144095 24279
rect 144029 24246 144030 24278
rect 143208 23734 143284 24214
rect 143208 23702 143214 23734
rect 141848 23664 141924 23670
rect 143213 23670 143214 23702
rect 143278 23702 143284 23734
rect 144024 24214 144030 24246
rect 144094 24246 144095 24278
rect 144094 24214 144100 24246
rect 144024 23734 144100 24214
rect 143278 23670 143279 23702
rect 143213 23669 143279 23670
rect 144024 23670 144030 23734
rect 144094 23670 144100 23734
rect 145384 23734 145460 24350
rect 179112 24414 179188 24420
rect 179112 24350 179118 24414
rect 179182 24350 179188 24414
rect 195024 24414 195100 25166
rect 199376 25166 199382 25198
rect 199446 25198 199447 25230
rect 199920 25230 199996 25236
rect 199446 25166 199452 25198
rect 199376 24958 199452 25166
rect 199376 24894 199382 24958
rect 199446 24894 199452 24958
rect 199920 25166 199926 25230
rect 199990 25166 199996 25230
rect 201149 25230 201215 25231
rect 201149 25198 201150 25230
rect 199920 24958 199996 25166
rect 199920 24926 199926 24958
rect 199376 24888 199452 24894
rect 199925 24894 199926 24926
rect 199990 24926 199996 24958
rect 201144 25166 201150 25198
rect 201214 25198 201215 25230
rect 204005 25230 204071 25231
rect 204005 25198 204006 25230
rect 201214 25166 201220 25198
rect 199990 24894 199991 24926
rect 199925 24893 199991 24894
rect 195024 24382 195030 24414
rect 146477 24278 146543 24279
rect 146477 24246 146478 24278
rect 145384 23702 145390 23734
rect 144024 23664 144100 23670
rect 145389 23670 145390 23702
rect 145454 23702 145460 23734
rect 146472 24214 146478 24246
rect 146542 24246 146543 24278
rect 147016 24278 147092 24284
rect 146542 24214 146548 24246
rect 146472 23734 146548 24214
rect 145454 23670 145455 23702
rect 145389 23669 145455 23670
rect 146472 23670 146478 23734
rect 146542 23670 146548 23734
rect 147016 24214 147022 24278
rect 147086 24214 147092 24278
rect 147701 24278 147767 24279
rect 147701 24246 147702 24278
rect 147016 23734 147092 24214
rect 147016 23702 147022 23734
rect 146472 23664 146548 23670
rect 147021 23670 147022 23702
rect 147086 23702 147092 23734
rect 147696 24214 147702 24246
rect 147766 24246 147767 24278
rect 149061 24278 149127 24279
rect 149061 24246 149062 24278
rect 147766 24214 147772 24246
rect 147696 23734 147772 24214
rect 147086 23670 147087 23702
rect 147021 23669 147087 23670
rect 147696 23670 147702 23734
rect 147766 23670 147772 23734
rect 147696 23664 147772 23670
rect 149056 24214 149062 24246
rect 149126 24246 149127 24278
rect 150416 24278 150492 24284
rect 149126 24214 149132 24246
rect 149056 23734 149132 24214
rect 149056 23670 149062 23734
rect 149126 23670 149132 23734
rect 150416 24214 150422 24278
rect 150486 24214 150492 24278
rect 150416 23734 150492 24214
rect 150416 23702 150422 23734
rect 149056 23664 149132 23670
rect 150421 23670 150422 23702
rect 150486 23702 150492 23734
rect 152048 24278 152124 24284
rect 152048 24214 152054 24278
rect 152118 24214 152124 24278
rect 152733 24278 152799 24279
rect 152733 24246 152734 24278
rect 152048 23734 152124 24214
rect 152048 23702 152054 23734
rect 150486 23670 150487 23702
rect 150421 23669 150487 23670
rect 152053 23670 152054 23702
rect 152118 23702 152124 23734
rect 152728 24214 152734 24246
rect 152798 24246 152799 24278
rect 153272 24278 153348 24284
rect 152798 24214 152804 24246
rect 152728 23734 152804 24214
rect 152118 23670 152119 23702
rect 152053 23669 152119 23670
rect 152728 23670 152734 23734
rect 152798 23670 152804 23734
rect 153272 24214 153278 24278
rect 153342 24214 153348 24278
rect 153272 23734 153348 24214
rect 153272 23702 153278 23734
rect 152728 23664 152804 23670
rect 153277 23670 153278 23702
rect 153342 23702 153348 23734
rect 154496 24278 154572 24284
rect 154496 24214 154502 24278
rect 154566 24214 154572 24278
rect 155181 24278 155247 24279
rect 155181 24246 155182 24278
rect 154496 23734 154572 24214
rect 154496 23702 154502 23734
rect 153342 23670 153343 23702
rect 153277 23669 153343 23670
rect 154501 23670 154502 23702
rect 154566 23702 154572 23734
rect 155176 24214 155182 24246
rect 155246 24246 155247 24278
rect 155720 24278 155796 24284
rect 155246 24214 155252 24246
rect 155176 23734 155252 24214
rect 154566 23670 154567 23702
rect 154501 23669 154567 23670
rect 155176 23670 155182 23734
rect 155246 23670 155252 23734
rect 155720 24214 155726 24278
rect 155790 24214 155796 24278
rect 155720 23734 155796 24214
rect 155720 23702 155726 23734
rect 155176 23664 155252 23670
rect 155725 23670 155726 23702
rect 155790 23702 155796 23734
rect 156944 24278 157020 24284
rect 156944 24214 156950 24278
rect 157014 24214 157020 24278
rect 156944 23734 157020 24214
rect 156944 23702 156950 23734
rect 155790 23670 155791 23702
rect 155725 23669 155791 23670
rect 156949 23670 156950 23702
rect 157014 23702 157020 23734
rect 158168 24278 158244 24284
rect 158168 24214 158174 24278
rect 158238 24214 158244 24278
rect 158168 23734 158244 24214
rect 158168 23702 158174 23734
rect 157014 23670 157015 23702
rect 156949 23669 157015 23670
rect 158173 23670 158174 23702
rect 158238 23702 158244 23734
rect 159528 24278 159604 24284
rect 159528 24214 159534 24278
rect 159598 24214 159604 24278
rect 160213 24278 160279 24279
rect 160213 24246 160214 24278
rect 159528 23734 159604 24214
rect 159528 23702 159534 23734
rect 158238 23670 158239 23702
rect 158173 23669 158239 23670
rect 159533 23670 159534 23702
rect 159598 23702 159604 23734
rect 160208 24214 160214 24246
rect 160278 24246 160279 24278
rect 160752 24278 160828 24284
rect 160278 24214 160284 24246
rect 160208 23734 160284 24214
rect 159598 23670 159599 23702
rect 159533 23669 159599 23670
rect 160208 23670 160214 23734
rect 160278 23670 160284 23734
rect 160752 24214 160758 24278
rect 160822 24214 160828 24278
rect 161437 24278 161503 24279
rect 161437 24246 161438 24278
rect 160752 23734 160828 24214
rect 160752 23702 160758 23734
rect 160208 23664 160284 23670
rect 160757 23670 160758 23702
rect 160822 23702 160828 23734
rect 161432 24214 161438 24246
rect 161502 24246 161503 24278
rect 163200 24278 163276 24284
rect 161502 24214 161508 24246
rect 161432 23734 161508 24214
rect 160822 23670 160823 23702
rect 160757 23669 160823 23670
rect 161432 23670 161438 23734
rect 161502 23670 161508 23734
rect 163200 24214 163206 24278
rect 163270 24214 163276 24278
rect 163200 23734 163276 24214
rect 163200 23702 163206 23734
rect 161432 23664 161508 23670
rect 163205 23670 163206 23702
rect 163270 23702 163276 23734
rect 164424 24278 164500 24284
rect 164424 24214 164430 24278
rect 164494 24214 164500 24278
rect 164424 23734 164500 24214
rect 164424 23702 164430 23734
rect 163270 23670 163271 23702
rect 163205 23669 163271 23670
rect 164429 23670 164430 23702
rect 164494 23702 164500 23734
rect 165376 24278 165452 24284
rect 165376 24214 165382 24278
rect 165446 24214 165452 24278
rect 165376 23734 165452 24214
rect 165376 23702 165382 23734
rect 164494 23670 164495 23702
rect 164429 23669 164495 23670
rect 165381 23670 165382 23702
rect 165446 23702 165452 23734
rect 166872 24278 166948 24284
rect 166872 24214 166878 24278
rect 166942 24214 166948 24278
rect 166872 23734 166948 24214
rect 166872 23702 166878 23734
rect 165446 23670 165447 23702
rect 165381 23669 165447 23670
rect 166877 23670 166878 23702
rect 166942 23702 166948 23734
rect 168232 24278 168308 24284
rect 168232 24214 168238 24278
rect 168302 24214 168308 24278
rect 168232 23734 168308 24214
rect 168232 23702 168238 23734
rect 166942 23670 166943 23702
rect 166877 23669 166943 23670
rect 168237 23670 168238 23702
rect 168302 23702 168308 23734
rect 169456 24278 169532 24284
rect 169456 24214 169462 24278
rect 169526 24214 169532 24278
rect 170549 24278 170615 24279
rect 170549 24246 170550 24278
rect 169456 23734 169532 24214
rect 169456 23702 169462 23734
rect 168302 23670 168303 23702
rect 168237 23669 168303 23670
rect 169461 23670 169462 23702
rect 169526 23702 169532 23734
rect 170544 24214 170550 24246
rect 170614 24246 170615 24278
rect 171365 24278 171431 24279
rect 171365 24246 171366 24278
rect 170614 24214 170620 24246
rect 170544 23734 170620 24214
rect 169526 23670 169527 23702
rect 169461 23669 169527 23670
rect 170544 23670 170550 23734
rect 170614 23670 170620 23734
rect 170544 23664 170620 23670
rect 171360 24214 171366 24246
rect 171430 24246 171431 24278
rect 171904 24278 171980 24284
rect 171430 24214 171436 24246
rect 171360 23734 171436 24214
rect 171360 23670 171366 23734
rect 171430 23670 171436 23734
rect 171904 24214 171910 24278
rect 171974 24214 171980 24278
rect 171904 23734 171980 24214
rect 171904 23702 171910 23734
rect 171360 23664 171436 23670
rect 171909 23670 171910 23702
rect 171974 23702 171980 23734
rect 173264 24278 173340 24284
rect 173264 24214 173270 24278
rect 173334 24214 173340 24278
rect 175173 24278 175239 24279
rect 175173 24246 175174 24278
rect 173264 23734 173340 24214
rect 173264 23702 173270 23734
rect 171974 23670 171975 23702
rect 171909 23669 171975 23670
rect 173269 23670 173270 23702
rect 173334 23702 173340 23734
rect 175168 24214 175174 24246
rect 175238 24246 175239 24278
rect 176936 24278 177012 24284
rect 175238 24214 175244 24246
rect 175168 23734 175244 24214
rect 173334 23670 173335 23702
rect 173269 23669 173335 23670
rect 175168 23670 175174 23734
rect 175238 23670 175244 23734
rect 176936 24214 176942 24278
rect 177006 24214 177012 24278
rect 176936 23734 177012 24214
rect 176936 23702 176942 23734
rect 175168 23664 175244 23670
rect 176941 23670 176942 23702
rect 177006 23702 177012 23734
rect 178160 24278 178236 24284
rect 178160 24214 178166 24278
rect 178230 24214 178236 24278
rect 178160 23734 178236 24214
rect 178160 23702 178166 23734
rect 177006 23670 177007 23702
rect 176941 23669 177007 23670
rect 178165 23670 178166 23702
rect 178230 23702 178236 23734
rect 179112 23734 179188 24350
rect 195029 24350 195030 24382
rect 195094 24382 195100 24414
rect 195094 24350 195095 24382
rect 195029 24349 195095 24350
rect 180205 24278 180271 24279
rect 180205 24246 180206 24278
rect 179112 23702 179118 23734
rect 178230 23670 178231 23702
rect 178165 23669 178231 23670
rect 179117 23670 179118 23702
rect 179182 23702 179188 23734
rect 180200 24214 180206 24246
rect 180270 24246 180271 24278
rect 181429 24278 181495 24279
rect 181429 24246 181430 24278
rect 180270 24214 180276 24246
rect 180200 23734 180276 24214
rect 179182 23670 179183 23702
rect 179117 23669 179183 23670
rect 180200 23670 180206 23734
rect 180270 23670 180276 23734
rect 180200 23664 180276 23670
rect 181424 24214 181430 24246
rect 181494 24246 181495 24278
rect 183192 24278 183268 24284
rect 181494 24214 181500 24246
rect 181424 23734 181500 24214
rect 181424 23670 181430 23734
rect 181494 23670 181500 23734
rect 183192 24214 183198 24278
rect 183262 24214 183268 24278
rect 183192 23734 183268 24214
rect 183192 23702 183198 23734
rect 181424 23664 181500 23670
rect 183197 23670 183198 23702
rect 183262 23702 183268 23734
rect 185640 24278 185716 24284
rect 185640 24214 185646 24278
rect 185710 24214 185716 24278
rect 186461 24278 186527 24279
rect 186461 24246 186462 24278
rect 185640 23734 185716 24214
rect 185640 23702 185646 23734
rect 183262 23670 183263 23702
rect 183197 23669 183263 23670
rect 185645 23670 185646 23702
rect 185710 23702 185716 23734
rect 186456 24214 186462 24246
rect 186526 24246 186527 24278
rect 187685 24278 187751 24279
rect 187685 24246 187686 24278
rect 186526 24214 186532 24246
rect 186456 23734 186532 24214
rect 185710 23670 185711 23702
rect 185645 23669 185711 23670
rect 186456 23670 186462 23734
rect 186526 23670 186532 23734
rect 186456 23664 186532 23670
rect 187680 24214 187686 24246
rect 187750 24246 187751 24278
rect 188909 24278 188975 24279
rect 188909 24246 188910 24278
rect 187750 24214 187756 24246
rect 187680 23734 187756 24214
rect 187680 23670 187686 23734
rect 187750 23670 187756 23734
rect 187680 23664 187756 23670
rect 188904 24214 188910 24246
rect 188974 24246 188975 24278
rect 188974 24214 188980 24246
rect 188904 23734 188980 24214
rect 188904 23670 188910 23734
rect 188974 23670 188980 23734
rect 188904 23664 188980 23670
rect 34685 23598 34751 23599
rect 34685 23566 34686 23598
rect 29920 22174 29926 22238
rect 29990 22174 29996 22238
rect 29920 22168 29996 22174
rect 34680 23534 34686 23566
rect 34750 23566 34751 23598
rect 39717 23598 39783 23599
rect 39717 23566 39718 23598
rect 34750 23534 34756 23566
rect 29920 22102 29996 22108
rect 29920 22038 29926 22102
rect 29990 22038 29996 22102
rect 29920 19654 29996 22038
rect 29920 19622 29926 19654
rect 29925 19590 29926 19622
rect 29990 19622 29996 19654
rect 30056 19654 30132 19660
rect 29990 19590 29991 19622
rect 29925 19589 29991 19590
rect 30056 19590 30062 19654
rect 30126 19590 30132 19654
rect 29648 18910 29654 18974
rect 29718 18910 29724 18974
rect 29648 18904 29724 18910
rect 29789 18838 29855 18839
rect 29789 18806 29790 18838
rect 29784 18774 29790 18806
rect 29854 18806 29855 18838
rect 29854 18774 29860 18806
rect 29784 18158 29860 18774
rect 29784 18094 29790 18158
rect 29854 18094 29860 18158
rect 29784 18088 29860 18094
rect 29920 18022 29996 18028
rect 29920 17958 29926 18022
rect 29990 17958 29996 18022
rect 28973 17614 29039 17615
rect 28973 17582 28974 17614
rect 21760 16734 21766 16798
rect 21830 16734 21836 16798
rect 21760 16728 21836 16734
rect 28968 17550 28974 17582
rect 29038 17582 29039 17614
rect 29038 17550 29044 17582
rect 20400 15238 20406 15302
rect 20470 15238 20476 15302
rect 20400 15232 20476 15238
rect 21760 16526 21836 16532
rect 21760 16462 21766 16526
rect 21830 16462 21836 16526
rect 21760 13942 21836 16462
rect 21760 13910 21766 13942
rect 21765 13878 21766 13910
rect 21830 13910 21836 13942
rect 21896 15166 21972 15172
rect 21896 15102 21902 15166
rect 21966 15102 21972 15166
rect 21830 13878 21831 13910
rect 21765 13877 21831 13878
rect 20405 13806 20471 13807
rect 20405 13774 20406 13806
rect 15232 12686 15238 12718
rect 15237 12654 15238 12686
rect 15302 12686 15308 12718
rect 20400 13742 20406 13774
rect 20470 13774 20471 13806
rect 20470 13742 20476 13774
rect 15302 12654 15303 12686
rect 15237 12653 15303 12654
rect 952 12246 1230 12310
rect 1294 12246 1300 12310
rect 2040 12582 2116 12588
rect 2040 12518 2046 12582
rect 2110 12518 2116 12582
rect 2040 12310 2116 12518
rect 2040 12278 2046 12310
rect 952 10678 1300 12246
rect 2045 12246 2046 12278
rect 2110 12278 2116 12310
rect 2110 12246 2111 12278
rect 2045 12245 2111 12246
rect 20400 11086 20476 13742
rect 21896 12446 21972 15102
rect 21896 12414 21902 12446
rect 21901 12382 21902 12414
rect 21966 12414 21972 12446
rect 21966 12382 21967 12414
rect 21901 12381 21967 12382
rect 20400 11022 20406 11086
rect 20470 11022 20476 11086
rect 20400 11016 20476 11022
rect 952 10614 1230 10678
rect 1294 10614 1300 10678
rect 952 9046 1300 10614
rect 952 8982 1230 9046
rect 1294 8982 1300 9046
rect 952 7142 1300 8982
rect 952 7078 1230 7142
rect 1294 7078 1300 7142
rect 952 5510 1300 7078
rect 952 5446 1230 5510
rect 1294 5446 1300 5510
rect 952 3878 1300 5446
rect 952 3814 1230 3878
rect 1294 3814 1300 3878
rect 952 2246 1300 3814
rect 16869 3606 16935 3607
rect 16869 3574 16870 3606
rect 16864 3542 16870 3574
rect 16934 3574 16935 3606
rect 16934 3542 16940 3574
rect 16461 2654 16527 2655
rect 16461 2622 16462 2654
rect 952 2182 1230 2246
rect 1294 2182 1300 2246
rect 952 1294 1300 2182
rect 16456 2590 16462 2622
rect 16526 2622 16527 2654
rect 16526 2590 16532 2622
rect 3677 1838 3743 1839
rect 3677 1806 3678 1838
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 1300 1294
rect 952 1158 1300 1230
rect 3672 1774 3678 1806
rect 3742 1806 3743 1838
rect 5445 1838 5511 1839
rect 5445 1806 5446 1838
rect 3742 1774 3748 1806
rect 3672 1294 3748 1774
rect 3672 1230 3678 1294
rect 3742 1230 3748 1294
rect 3672 1224 3748 1230
rect 5440 1774 5446 1806
rect 5510 1806 5511 1838
rect 6941 1838 7007 1839
rect 6941 1806 6942 1838
rect 5510 1774 5516 1806
rect 5440 1294 5516 1774
rect 5440 1230 5446 1294
rect 5510 1230 5516 1294
rect 5440 1224 5516 1230
rect 6936 1774 6942 1806
rect 7006 1806 7007 1838
rect 8709 1838 8775 1839
rect 8709 1806 8710 1838
rect 7006 1774 7012 1806
rect 6936 1294 7012 1774
rect 6936 1230 6942 1294
rect 7006 1230 7012 1294
rect 6936 1224 7012 1230
rect 8704 1774 8710 1806
rect 8774 1806 8775 1838
rect 10477 1838 10543 1839
rect 10477 1806 10478 1838
rect 8774 1774 8780 1806
rect 8704 1294 8780 1774
rect 8704 1230 8710 1294
rect 8774 1230 8780 1294
rect 8704 1224 8780 1230
rect 10472 1774 10478 1806
rect 10542 1806 10543 1838
rect 12109 1838 12175 1839
rect 12109 1806 12110 1838
rect 10542 1774 10548 1806
rect 10472 1294 10548 1774
rect 10472 1230 10478 1294
rect 10542 1230 10548 1294
rect 10472 1224 10548 1230
rect 12104 1774 12110 1806
rect 12174 1806 12175 1838
rect 13741 1838 13807 1839
rect 13741 1806 13742 1838
rect 12174 1774 12180 1806
rect 12104 1294 12180 1774
rect 12104 1230 12110 1294
rect 12174 1230 12180 1294
rect 12104 1224 12180 1230
rect 13736 1774 13742 1806
rect 13806 1806 13807 1838
rect 15509 1838 15575 1839
rect 15509 1806 15510 1838
rect 13806 1774 13812 1806
rect 13736 1294 13812 1774
rect 13736 1230 13742 1294
rect 13806 1230 13812 1294
rect 13736 1224 13812 1230
rect 15504 1774 15510 1806
rect 15574 1806 15575 1838
rect 15574 1774 15580 1806
rect 15504 1294 15580 1774
rect 15504 1230 15510 1294
rect 15574 1230 15580 1294
rect 15504 1224 15580 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 1300 1158
rect 952 1022 1300 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 1300 1022
rect 952 952 1300 958
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 620 614
rect 272 478 620 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 620 478
rect 272 342 620 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 620 342
rect 272 272 620 278
rect 16456 0 16532 2590
rect 16864 614 16940 3542
rect 17685 2654 17751 2655
rect 17685 2622 17686 2654
rect 17680 2590 17686 2622
rect 17750 2622 17751 2654
rect 18773 2654 18839 2655
rect 18773 2622 18774 2654
rect 17750 2590 17756 2622
rect 17141 1838 17207 1839
rect 17141 1806 17142 1838
rect 17136 1774 17142 1806
rect 17206 1806 17207 1838
rect 17206 1774 17212 1806
rect 17136 1294 17212 1774
rect 17136 1230 17142 1294
rect 17206 1230 17212 1294
rect 17136 1224 17212 1230
rect 16864 550 16870 614
rect 16934 550 16940 614
rect 16864 544 16940 550
rect 17680 0 17756 2590
rect 18768 2590 18774 2622
rect 18838 2622 18839 2654
rect 19997 2654 20063 2655
rect 19997 2622 19998 2654
rect 18838 2590 18844 2622
rect 18768 0 18844 2590
rect 19992 2590 19998 2622
rect 20062 2622 20063 2654
rect 21085 2654 21151 2655
rect 21085 2622 21086 2654
rect 20062 2590 20068 2622
rect 19045 1838 19111 1839
rect 19045 1806 19046 1838
rect 19040 1774 19046 1806
rect 19110 1806 19111 1838
rect 19110 1774 19116 1806
rect 19040 1294 19116 1774
rect 19040 1230 19046 1294
rect 19110 1230 19116 1294
rect 19040 1224 19116 1230
rect 19992 0 20068 2590
rect 21080 2590 21086 2622
rect 21150 2622 21151 2654
rect 22309 2654 22375 2655
rect 22309 2622 22310 2654
rect 21150 2590 21156 2622
rect 20405 1838 20471 1839
rect 20405 1806 20406 1838
rect 20400 1774 20406 1806
rect 20470 1806 20471 1838
rect 20470 1774 20476 1806
rect 20400 1294 20476 1774
rect 20400 1230 20406 1294
rect 20470 1230 20476 1294
rect 20400 1224 20476 1230
rect 21080 0 21156 2590
rect 22304 2590 22310 2622
rect 22374 2622 22375 2654
rect 23533 2654 23599 2655
rect 23533 2622 23534 2654
rect 22374 2590 22380 2622
rect 22173 1838 22239 1839
rect 22173 1806 22174 1838
rect 22168 1774 22174 1806
rect 22238 1806 22239 1838
rect 22238 1774 22244 1806
rect 22168 1294 22244 1774
rect 22168 1230 22174 1294
rect 22238 1230 22244 1294
rect 22168 1224 22244 1230
rect 22304 0 22380 2590
rect 23528 2590 23534 2622
rect 23598 2622 23599 2654
rect 24621 2654 24687 2655
rect 24621 2622 24622 2654
rect 23598 2590 23604 2622
rect 23528 0 23604 2590
rect 24616 2590 24622 2622
rect 24686 2622 24687 2654
rect 25981 2654 26047 2655
rect 25981 2622 25982 2654
rect 24686 2590 24692 2622
rect 23941 1838 24007 1839
rect 23941 1806 23942 1838
rect 23936 1774 23942 1806
rect 24006 1806 24007 1838
rect 24006 1774 24012 1806
rect 23936 1294 24012 1774
rect 23936 1230 23942 1294
rect 24006 1230 24012 1294
rect 23936 1224 24012 1230
rect 24616 0 24692 2590
rect 25976 2590 25982 2622
rect 26046 2622 26047 2654
rect 27069 2654 27135 2655
rect 27069 2622 27070 2654
rect 26046 2590 26052 2622
rect 25437 1838 25503 1839
rect 25437 1806 25438 1838
rect 25432 1774 25438 1806
rect 25502 1806 25503 1838
rect 25502 1774 25508 1806
rect 25432 1294 25508 1774
rect 25432 1230 25438 1294
rect 25502 1230 25508 1294
rect 25432 1224 25508 1230
rect 25976 0 26052 2590
rect 27064 2590 27070 2622
rect 27134 2622 27135 2654
rect 28293 2654 28359 2655
rect 28293 2622 28294 2654
rect 27134 2590 27140 2622
rect 27064 0 27140 2590
rect 28288 2590 28294 2622
rect 28358 2622 28359 2654
rect 28358 2590 28364 2622
rect 27205 1838 27271 1839
rect 27205 1806 27206 1838
rect 27200 1774 27206 1806
rect 27270 1806 27271 1838
rect 27270 1774 27276 1806
rect 27200 1294 27276 1774
rect 27200 1230 27206 1294
rect 27270 1230 27276 1294
rect 27200 1224 27276 1230
rect 28288 0 28364 2590
rect 28837 1838 28903 1839
rect 28837 1806 28838 1838
rect 28832 1774 28838 1806
rect 28902 1806 28903 1838
rect 28902 1774 28908 1806
rect 28832 1294 28908 1774
rect 28832 1230 28838 1294
rect 28902 1230 28908 1294
rect 28832 1224 28908 1230
rect 28968 0 29044 17550
rect 29784 17478 29860 17484
rect 29784 17414 29790 17478
rect 29854 17414 29860 17478
rect 29784 17070 29860 17414
rect 29784 17038 29790 17070
rect 29789 17006 29790 17038
rect 29854 17038 29860 17070
rect 29854 17006 29855 17038
rect 29789 17005 29855 17006
rect 29789 16934 29855 16935
rect 29789 16902 29790 16934
rect 29784 16870 29790 16902
rect 29854 16902 29855 16934
rect 29854 16870 29860 16902
rect 29653 16390 29719 16391
rect 29653 16358 29654 16390
rect 29648 16326 29654 16358
rect 29718 16358 29719 16390
rect 29718 16326 29724 16358
rect 29240 15846 29316 15852
rect 29240 15782 29246 15846
rect 29310 15782 29316 15846
rect 29240 14078 29316 15782
rect 29512 15574 29588 15580
rect 29512 15510 29518 15574
rect 29582 15510 29588 15574
rect 29512 15166 29588 15510
rect 29648 15574 29724 16326
rect 29784 16254 29860 16870
rect 29920 16526 29996 17958
rect 30056 17886 30132 19590
rect 34680 18974 34756 23534
rect 39712 23534 39718 23566
rect 39782 23566 39783 23598
rect 45424 23598 45500 23604
rect 39782 23534 39788 23566
rect 35088 22102 35164 22108
rect 35088 22038 35094 22102
rect 35158 22038 35164 22102
rect 34680 18910 34686 18974
rect 34750 18910 34756 18974
rect 34680 18904 34756 18910
rect 34952 19654 35028 19660
rect 34952 19590 34958 19654
rect 35022 19590 35028 19654
rect 35088 19654 35164 22038
rect 35088 19622 35094 19654
rect 34685 18838 34751 18839
rect 34685 18806 34686 18838
rect 34680 18774 34686 18806
rect 34750 18806 34751 18838
rect 34750 18774 34756 18806
rect 34680 18158 34756 18774
rect 34680 18094 34686 18158
rect 34750 18094 34756 18158
rect 34680 18088 34756 18094
rect 30056 17854 30062 17886
rect 30061 17822 30062 17854
rect 30126 17854 30132 17886
rect 34816 18022 34892 18028
rect 34816 17958 34822 18022
rect 34886 17958 34892 18022
rect 30126 17822 30127 17854
rect 30061 17821 30127 17822
rect 34549 17614 34615 17615
rect 34549 17582 34550 17614
rect 29920 16494 29926 16526
rect 29925 16462 29926 16494
rect 29990 16494 29996 16526
rect 34544 17550 34550 17582
rect 34614 17582 34615 17614
rect 34614 17550 34620 17582
rect 29990 16462 29991 16494
rect 29925 16461 29991 16462
rect 29784 16190 29790 16254
rect 29854 16190 29860 16254
rect 29784 16184 29860 16190
rect 29648 15510 29654 15574
rect 29718 15510 29724 15574
rect 29648 15504 29724 15510
rect 29512 15134 29518 15166
rect 29517 15102 29518 15134
rect 29582 15134 29588 15166
rect 29582 15102 29583 15134
rect 29517 15101 29583 15102
rect 29240 14046 29246 14078
rect 29245 14014 29246 14046
rect 29310 14046 29316 14078
rect 29310 14014 29311 14046
rect 29245 14013 29311 14014
rect 29245 2654 29311 2655
rect 29245 2622 29246 2654
rect 29240 2590 29246 2622
rect 29310 2622 29311 2654
rect 30605 2654 30671 2655
rect 30605 2622 30606 2654
rect 29310 2590 29316 2622
rect 29240 0 29316 2590
rect 30600 2590 30606 2622
rect 30670 2622 30671 2654
rect 31693 2654 31759 2655
rect 31693 2622 31694 2654
rect 30670 2590 30676 2622
rect 30469 1838 30535 1839
rect 30469 1806 30470 1838
rect 30464 1774 30470 1806
rect 30534 1806 30535 1838
rect 30534 1774 30540 1806
rect 30464 1294 30540 1774
rect 30464 1230 30470 1294
rect 30534 1230 30540 1294
rect 30464 1224 30540 1230
rect 30600 0 30676 2590
rect 31688 2590 31694 2622
rect 31758 2622 31759 2654
rect 32781 2654 32847 2655
rect 32781 2622 32782 2654
rect 31758 2590 31764 2622
rect 31688 0 31764 2590
rect 32776 2590 32782 2622
rect 32846 2622 32847 2654
rect 34005 2654 34071 2655
rect 34005 2622 34006 2654
rect 32846 2590 32852 2622
rect 32373 1838 32439 1839
rect 32373 1806 32374 1838
rect 32368 1774 32374 1806
rect 32438 1806 32439 1838
rect 32438 1774 32444 1806
rect 32368 1294 32444 1774
rect 32368 1230 32374 1294
rect 32438 1230 32444 1294
rect 32368 1224 32444 1230
rect 32776 0 32852 2590
rect 34000 2590 34006 2622
rect 34070 2622 34071 2654
rect 34070 2590 34076 2622
rect 33869 1838 33935 1839
rect 33869 1806 33870 1838
rect 33864 1774 33870 1806
rect 33934 1806 33935 1838
rect 33934 1774 33940 1806
rect 33864 1294 33940 1774
rect 33864 1230 33870 1294
rect 33934 1230 33940 1294
rect 33864 1224 33940 1230
rect 34000 0 34076 2590
rect 34544 0 34620 17550
rect 34816 16526 34892 17958
rect 34952 17886 35028 19590
rect 35093 19590 35094 19622
rect 35158 19622 35164 19654
rect 35158 19590 35159 19622
rect 35093 19589 35159 19590
rect 39712 18974 39788 23534
rect 45424 23534 45430 23598
rect 45494 23534 45500 23598
rect 49373 23598 49439 23599
rect 49373 23566 49374 23598
rect 39984 22102 40060 22108
rect 39984 22038 39990 22102
rect 40054 22038 40060 22102
rect 39712 18910 39718 18974
rect 39782 18910 39788 18974
rect 39712 18904 39788 18910
rect 39848 19654 39924 19660
rect 39848 19590 39854 19654
rect 39918 19590 39924 19654
rect 39984 19654 40060 22038
rect 39984 19622 39990 19654
rect 39717 18838 39783 18839
rect 39717 18806 39718 18838
rect 39712 18774 39718 18806
rect 39782 18806 39783 18838
rect 39782 18774 39788 18806
rect 39712 18158 39788 18774
rect 39712 18094 39718 18158
rect 39782 18094 39788 18158
rect 39712 18088 39788 18094
rect 34952 17854 34958 17886
rect 34957 17822 34958 17854
rect 35022 17854 35028 17886
rect 39712 18022 39788 18028
rect 39712 17958 39718 18022
rect 39782 17958 39788 18022
rect 35022 17822 35023 17854
rect 34957 17821 35023 17822
rect 34952 17614 35028 17620
rect 34952 17550 34958 17614
rect 35022 17550 35028 17614
rect 39445 17614 39511 17615
rect 39445 17582 39446 17614
rect 34952 17070 35028 17550
rect 34952 17038 34958 17070
rect 34957 17006 34958 17038
rect 35022 17038 35028 17070
rect 39440 17550 39446 17582
rect 39510 17582 39511 17614
rect 39510 17550 39516 17582
rect 35022 17006 35023 17038
rect 34957 17005 35023 17006
rect 34957 16934 35023 16935
rect 34957 16902 34958 16934
rect 34816 16494 34822 16526
rect 34821 16462 34822 16494
rect 34886 16494 34892 16526
rect 34952 16870 34958 16902
rect 35022 16902 35023 16934
rect 35022 16870 35028 16902
rect 34886 16462 34887 16494
rect 34821 16461 34887 16462
rect 34821 16390 34887 16391
rect 34821 16358 34822 16390
rect 34816 16326 34822 16358
rect 34886 16358 34887 16390
rect 34886 16326 34892 16358
rect 34816 15574 34892 16326
rect 34952 16254 35028 16870
rect 34952 16190 34958 16254
rect 35022 16190 35028 16254
rect 34952 16184 35028 16190
rect 34816 15510 34822 15574
rect 34886 15510 34892 15574
rect 34816 15504 34892 15510
rect 35093 2654 35159 2655
rect 35093 2622 35094 2654
rect 35088 2590 35094 2622
rect 35158 2622 35159 2654
rect 36453 2654 36519 2655
rect 36453 2622 36454 2654
rect 35158 2590 35164 2622
rect 35088 0 35164 2590
rect 36448 2590 36454 2622
rect 36518 2622 36519 2654
rect 37541 2654 37607 2655
rect 37541 2622 37542 2654
rect 36518 2590 36524 2622
rect 35501 1838 35567 1839
rect 35501 1806 35502 1838
rect 35496 1774 35502 1806
rect 35566 1806 35567 1838
rect 35566 1774 35572 1806
rect 35496 1294 35572 1774
rect 35496 1230 35502 1294
rect 35566 1230 35572 1294
rect 35496 1224 35572 1230
rect 36448 0 36524 2590
rect 37536 2590 37542 2622
rect 37606 2622 37607 2654
rect 38629 2654 38695 2655
rect 38629 2622 38630 2654
rect 37606 2590 37612 2622
rect 37269 1838 37335 1839
rect 37269 1806 37270 1838
rect 37264 1774 37270 1806
rect 37334 1806 37335 1838
rect 37334 1774 37340 1806
rect 37264 1294 37340 1774
rect 37264 1230 37270 1294
rect 37334 1230 37340 1294
rect 37264 1224 37340 1230
rect 37536 0 37612 2590
rect 38624 2590 38630 2622
rect 38694 2622 38695 2654
rect 38694 2590 38700 2622
rect 38624 0 38700 2590
rect 38901 1838 38967 1839
rect 38901 1806 38902 1838
rect 38896 1774 38902 1806
rect 38966 1806 38967 1838
rect 38966 1774 38972 1806
rect 38896 1294 38972 1774
rect 38896 1230 38902 1294
rect 38966 1230 38972 1294
rect 38896 1224 38972 1230
rect 39440 0 39516 17550
rect 39712 16526 39788 17958
rect 39848 17886 39924 19590
rect 39989 19590 39990 19622
rect 40054 19622 40060 19654
rect 44880 22102 44956 22108
rect 44880 22038 44886 22102
rect 44950 22038 44956 22102
rect 44880 19654 44956 22038
rect 44880 19622 44886 19654
rect 40054 19590 40055 19622
rect 39989 19589 40055 19590
rect 44885 19590 44886 19622
rect 44950 19622 44956 19654
rect 45016 19654 45092 19660
rect 44950 19590 44951 19622
rect 44885 19589 44951 19590
rect 45016 19590 45022 19654
rect 45086 19590 45092 19654
rect 44749 18838 44815 18839
rect 44749 18806 44750 18838
rect 44744 18774 44750 18806
rect 44814 18806 44815 18838
rect 44814 18774 44820 18806
rect 44744 18158 44820 18774
rect 44744 18094 44750 18158
rect 44814 18094 44820 18158
rect 44744 18088 44820 18094
rect 39848 17854 39854 17886
rect 39853 17822 39854 17854
rect 39918 17854 39924 17886
rect 44880 18022 44956 18028
rect 44880 17958 44886 18022
rect 44950 17958 44956 18022
rect 39918 17822 39919 17854
rect 39853 17821 39919 17822
rect 39848 17614 39924 17620
rect 39848 17550 39854 17614
rect 39918 17550 39924 17614
rect 44205 17614 44271 17615
rect 44205 17582 44206 17614
rect 39848 17070 39924 17550
rect 39848 17038 39854 17070
rect 39853 17006 39854 17038
rect 39918 17038 39924 17070
rect 44200 17550 44206 17582
rect 44270 17582 44271 17614
rect 44270 17550 44276 17582
rect 39918 17006 39919 17038
rect 39853 17005 39919 17006
rect 39853 16934 39919 16935
rect 39853 16902 39854 16934
rect 39712 16494 39718 16526
rect 39717 16462 39718 16494
rect 39782 16494 39788 16526
rect 39848 16870 39854 16902
rect 39918 16902 39919 16934
rect 39918 16870 39924 16902
rect 39782 16462 39783 16494
rect 39717 16461 39783 16462
rect 39717 16390 39783 16391
rect 39717 16358 39718 16390
rect 39712 16326 39718 16358
rect 39782 16358 39783 16390
rect 39782 16326 39788 16358
rect 39712 15574 39788 16326
rect 39848 16254 39924 16870
rect 39848 16190 39854 16254
rect 39918 16190 39924 16254
rect 39848 16184 39924 16190
rect 39712 15510 39718 15574
rect 39782 15510 39788 15574
rect 39712 15504 39788 15510
rect 39853 2654 39919 2655
rect 39853 2622 39854 2654
rect 39848 2590 39854 2622
rect 39918 2622 39919 2654
rect 40941 2654 41007 2655
rect 40941 2622 40942 2654
rect 39918 2590 39924 2622
rect 39848 0 39924 2590
rect 40936 2590 40942 2622
rect 41006 2622 41007 2654
rect 42301 2654 42367 2655
rect 42301 2622 42302 2654
rect 41006 2590 41012 2622
rect 40805 1838 40871 1839
rect 40805 1806 40806 1838
rect 40800 1774 40806 1806
rect 40870 1806 40871 1838
rect 40870 1774 40876 1806
rect 40800 1294 40876 1774
rect 40800 1230 40806 1294
rect 40870 1230 40876 1294
rect 40800 1224 40876 1230
rect 40936 0 41012 2590
rect 42296 2590 42302 2622
rect 42366 2622 42367 2654
rect 43389 2654 43455 2655
rect 43389 2622 43390 2654
rect 42366 2590 42372 2622
rect 42296 0 42372 2590
rect 43384 2590 43390 2622
rect 43454 2622 43455 2654
rect 43454 2590 43460 2622
rect 42437 1838 42503 1839
rect 42437 1806 42438 1838
rect 42432 1774 42438 1806
rect 42502 1806 42503 1838
rect 42502 1774 42508 1806
rect 42432 1294 42508 1774
rect 42432 1230 42438 1294
rect 42502 1230 42508 1294
rect 42432 1224 42508 1230
rect 43384 0 43460 2590
rect 43933 1838 43999 1839
rect 43933 1806 43934 1838
rect 43928 1774 43934 1806
rect 43998 1806 43999 1838
rect 43998 1774 44004 1806
rect 43928 1294 44004 1774
rect 43928 1230 43934 1294
rect 43998 1230 44004 1294
rect 43928 1224 44004 1230
rect 44200 0 44276 17550
rect 44744 17478 44820 17484
rect 44744 17414 44750 17478
rect 44814 17414 44820 17478
rect 44744 17070 44820 17414
rect 44744 17038 44750 17070
rect 44749 17006 44750 17038
rect 44814 17038 44820 17070
rect 44814 17006 44815 17038
rect 44749 17005 44815 17006
rect 44613 16934 44679 16935
rect 44613 16902 44614 16934
rect 44608 16870 44614 16902
rect 44678 16902 44679 16934
rect 44678 16870 44684 16902
rect 44608 16254 44684 16870
rect 44880 16526 44956 17958
rect 45016 17886 45092 19590
rect 45424 18974 45500 23534
rect 45424 18942 45430 18974
rect 45429 18910 45430 18942
rect 45494 18942 45500 18974
rect 49368 23534 49374 23566
rect 49438 23566 49439 23598
rect 54269 23598 54335 23599
rect 54269 23566 54270 23598
rect 49438 23534 49444 23566
rect 49368 18974 49444 23534
rect 54264 23534 54270 23566
rect 54334 23566 54335 23598
rect 60792 23598 60868 23604
rect 54334 23534 54340 23566
rect 50048 22102 50124 22108
rect 50048 22038 50054 22102
rect 50118 22038 50124 22102
rect 45494 18910 45495 18942
rect 45429 18909 45495 18910
rect 49368 18910 49374 18974
rect 49438 18910 49444 18974
rect 49368 18904 49444 18910
rect 49912 19654 49988 19660
rect 49912 19590 49918 19654
rect 49982 19590 49988 19654
rect 50048 19654 50124 22038
rect 50048 19622 50054 19654
rect 49645 18838 49711 18839
rect 49645 18806 49646 18838
rect 49640 18774 49646 18806
rect 49710 18806 49711 18838
rect 49710 18774 49716 18806
rect 49640 18158 49716 18774
rect 49640 18094 49646 18158
rect 49710 18094 49716 18158
rect 49640 18088 49716 18094
rect 45016 17854 45022 17886
rect 45021 17822 45022 17854
rect 45086 17854 45092 17886
rect 49776 18022 49852 18028
rect 49776 17958 49782 18022
rect 49846 17958 49852 18022
rect 45086 17822 45087 17854
rect 45021 17821 45087 17822
rect 49509 17614 49575 17615
rect 49509 17582 49510 17614
rect 44880 16494 44886 16526
rect 44885 16462 44886 16494
rect 44950 16494 44956 16526
rect 49504 17550 49510 17582
rect 49574 17582 49575 17614
rect 49574 17550 49580 17582
rect 44950 16462 44951 16494
rect 44885 16461 44951 16462
rect 44749 16390 44815 16391
rect 44749 16358 44750 16390
rect 44608 16190 44614 16254
rect 44678 16190 44684 16254
rect 44608 16184 44684 16190
rect 44744 16326 44750 16358
rect 44814 16358 44815 16390
rect 44814 16326 44820 16358
rect 44744 15574 44820 16326
rect 44744 15510 44750 15574
rect 44814 15510 44820 15574
rect 44744 15504 44820 15510
rect 44613 2654 44679 2655
rect 44613 2622 44614 2654
rect 44608 2590 44614 2622
rect 44678 2622 44679 2654
rect 45837 2654 45903 2655
rect 45837 2622 45838 2654
rect 44678 2590 44684 2622
rect 44608 0 44684 2590
rect 45832 2590 45838 2622
rect 45902 2622 45903 2654
rect 46925 2654 46991 2655
rect 46925 2622 46926 2654
rect 45902 2590 45908 2622
rect 45701 1838 45767 1839
rect 45701 1806 45702 1838
rect 45696 1774 45702 1806
rect 45766 1806 45767 1838
rect 45766 1774 45772 1806
rect 45696 1294 45772 1774
rect 45696 1230 45702 1294
rect 45766 1230 45772 1294
rect 45696 1224 45772 1230
rect 45832 0 45908 2590
rect 46920 2590 46926 2622
rect 46990 2622 46991 2654
rect 48013 2654 48079 2655
rect 48013 2622 48014 2654
rect 46990 2590 46996 2622
rect 46920 0 46996 2590
rect 48008 2590 48014 2622
rect 48078 2622 48079 2654
rect 49101 2654 49167 2655
rect 49101 2622 49102 2654
rect 48078 2590 48084 2622
rect 47469 1838 47535 1839
rect 47469 1806 47470 1838
rect 47464 1774 47470 1806
rect 47534 1806 47535 1838
rect 47534 1774 47540 1806
rect 47464 1294 47540 1774
rect 47464 1230 47470 1294
rect 47534 1230 47540 1294
rect 47464 1224 47540 1230
rect 48008 0 48084 2590
rect 49096 2590 49102 2622
rect 49166 2622 49167 2654
rect 49166 2590 49172 2622
rect 48965 1838 49031 1839
rect 48965 1806 48966 1838
rect 48960 1774 48966 1806
rect 49030 1806 49031 1838
rect 49030 1774 49036 1806
rect 48960 1294 49036 1774
rect 48960 1230 48966 1294
rect 49030 1230 49036 1294
rect 48960 1224 49036 1230
rect 49096 0 49172 2590
rect 49504 0 49580 17550
rect 49776 16526 49852 17958
rect 49912 17886 49988 19590
rect 50053 19590 50054 19622
rect 50118 19622 50124 19654
rect 50118 19590 50119 19622
rect 50053 19589 50119 19590
rect 54264 18974 54340 23534
rect 60792 23534 60798 23598
rect 60862 23534 60868 23598
rect 64605 23598 64671 23599
rect 64605 23566 64606 23598
rect 55080 22102 55156 22108
rect 55080 22038 55086 22102
rect 55150 22038 55156 22102
rect 59709 22102 59775 22103
rect 59709 22070 59710 22102
rect 54264 18910 54270 18974
rect 54334 18910 54340 18974
rect 54264 18904 54340 18910
rect 54944 19654 55020 19660
rect 54944 19590 54950 19654
rect 55014 19590 55020 19654
rect 55080 19654 55156 22038
rect 55080 19622 55086 19654
rect 54677 18838 54743 18839
rect 54677 18806 54678 18838
rect 54672 18774 54678 18806
rect 54742 18806 54743 18838
rect 54742 18774 54748 18806
rect 54672 18158 54748 18774
rect 54672 18094 54678 18158
rect 54742 18094 54748 18158
rect 54672 18088 54748 18094
rect 49912 17854 49918 17886
rect 49917 17822 49918 17854
rect 49982 17854 49988 17886
rect 54808 18022 54884 18028
rect 54808 17958 54814 18022
rect 54878 17958 54884 18022
rect 49982 17822 49983 17854
rect 49917 17821 49983 17822
rect 49912 17614 49988 17620
rect 49912 17550 49918 17614
rect 49982 17550 49988 17614
rect 54541 17614 54607 17615
rect 54541 17582 54542 17614
rect 49912 17206 49988 17550
rect 49912 17174 49918 17206
rect 49917 17142 49918 17174
rect 49982 17174 49988 17206
rect 54536 17550 54542 17582
rect 54606 17582 54607 17614
rect 54606 17550 54612 17582
rect 49982 17142 49983 17174
rect 49917 17141 49983 17142
rect 50053 17070 50119 17071
rect 50053 17038 50054 17070
rect 50048 17006 50054 17038
rect 50118 17038 50119 17070
rect 50118 17006 50124 17038
rect 49776 16494 49782 16526
rect 49781 16462 49782 16494
rect 49846 16494 49852 16526
rect 49912 16934 49988 16940
rect 49912 16870 49918 16934
rect 49982 16870 49988 16934
rect 49846 16462 49847 16494
rect 49781 16461 49847 16462
rect 49781 16390 49847 16391
rect 49781 16358 49782 16390
rect 49776 16326 49782 16358
rect 49846 16358 49847 16390
rect 49846 16326 49852 16358
rect 49776 15574 49852 16326
rect 49912 15982 49988 16870
rect 50048 16254 50124 17006
rect 50048 16190 50054 16254
rect 50118 16190 50124 16254
rect 50048 16184 50124 16190
rect 49912 15950 49918 15982
rect 49917 15918 49918 15950
rect 49982 15950 49988 15982
rect 49982 15918 49983 15950
rect 49917 15917 49983 15918
rect 49776 15510 49782 15574
rect 49846 15510 49852 15574
rect 49776 15504 49852 15510
rect 50325 2654 50391 2655
rect 50325 2622 50326 2654
rect 50320 2590 50326 2622
rect 50390 2622 50391 2654
rect 51549 2654 51615 2655
rect 51549 2622 51550 2654
rect 50390 2590 50396 2622
rect 50320 0 50396 2590
rect 51544 2590 51550 2622
rect 51614 2622 51615 2654
rect 52773 2654 52839 2655
rect 52773 2622 52774 2654
rect 51614 2590 51620 2622
rect 50733 1838 50799 1839
rect 50733 1806 50734 1838
rect 50728 1774 50734 1806
rect 50798 1806 50799 1838
rect 50798 1774 50804 1806
rect 50728 1294 50804 1774
rect 50728 1230 50734 1294
rect 50798 1230 50804 1294
rect 50728 1224 50804 1230
rect 51544 0 51620 2590
rect 52768 2590 52774 2622
rect 52838 2622 52839 2654
rect 53861 2654 53927 2655
rect 53861 2622 53862 2654
rect 52838 2590 52844 2622
rect 52365 1838 52431 1839
rect 52365 1806 52366 1838
rect 52360 1774 52366 1806
rect 52430 1806 52431 1838
rect 52430 1774 52436 1806
rect 52360 1294 52436 1774
rect 52360 1230 52366 1294
rect 52430 1230 52436 1294
rect 52360 1224 52436 1230
rect 52768 0 52844 2590
rect 53856 2590 53862 2622
rect 53926 2622 53927 2654
rect 53926 2590 53932 2622
rect 53856 0 53932 2590
rect 54133 1838 54199 1839
rect 54133 1806 54134 1838
rect 54128 1774 54134 1806
rect 54198 1806 54199 1838
rect 54198 1774 54204 1806
rect 54128 1294 54204 1774
rect 54128 1230 54134 1294
rect 54198 1230 54204 1294
rect 54128 1224 54204 1230
rect 54536 0 54612 17550
rect 54808 16526 54884 17958
rect 54944 17886 55020 19590
rect 55085 19590 55086 19622
rect 55150 19622 55156 19654
rect 59704 22038 59710 22070
rect 59774 22070 59775 22102
rect 59774 22038 59780 22070
rect 59704 19654 59780 22038
rect 55150 19590 55151 19622
rect 55085 19589 55151 19590
rect 59704 19590 59710 19654
rect 59774 19590 59780 19654
rect 59704 19584 59780 19590
rect 59976 19654 60052 19660
rect 59976 19590 59982 19654
rect 60046 19590 60052 19654
rect 59709 18838 59775 18839
rect 59709 18806 59710 18838
rect 59704 18774 59710 18806
rect 59774 18806 59775 18838
rect 59774 18774 59780 18806
rect 59704 18158 59780 18774
rect 59704 18094 59710 18158
rect 59774 18094 59780 18158
rect 59704 18088 59780 18094
rect 54944 17854 54950 17886
rect 54949 17822 54950 17854
rect 55014 17854 55020 17886
rect 59840 18022 59916 18028
rect 59840 17958 59846 18022
rect 59910 17958 59916 18022
rect 55014 17822 55015 17854
rect 54949 17821 55015 17822
rect 54944 17614 55020 17620
rect 54944 17550 54950 17614
rect 55014 17550 55020 17614
rect 59301 17614 59367 17615
rect 59301 17582 59302 17614
rect 54944 17070 55020 17550
rect 54944 17038 54950 17070
rect 54949 17006 54950 17038
rect 55014 17038 55020 17070
rect 59296 17550 59302 17582
rect 59366 17582 59367 17614
rect 59366 17550 59372 17582
rect 55014 17006 55015 17038
rect 54949 17005 55015 17006
rect 54949 16934 55015 16935
rect 54949 16902 54950 16934
rect 54808 16494 54814 16526
rect 54813 16462 54814 16494
rect 54878 16494 54884 16526
rect 54944 16870 54950 16902
rect 55014 16902 55015 16934
rect 55014 16870 55020 16902
rect 54878 16462 54879 16494
rect 54813 16461 54879 16462
rect 54813 16390 54879 16391
rect 54813 16358 54814 16390
rect 54808 16326 54814 16358
rect 54878 16358 54879 16390
rect 54878 16326 54884 16358
rect 54808 15574 54884 16326
rect 54944 16254 55020 16870
rect 54944 16190 54950 16254
rect 55014 16190 55020 16254
rect 54944 16184 55020 16190
rect 54808 15510 54814 15574
rect 54878 15510 54884 15574
rect 54808 15504 54884 15510
rect 54949 2654 55015 2655
rect 54949 2622 54950 2654
rect 54944 2590 54950 2622
rect 55014 2622 55015 2654
rect 56173 2654 56239 2655
rect 56173 2622 56174 2654
rect 55014 2590 55020 2622
rect 54944 0 55020 2590
rect 56168 2590 56174 2622
rect 56238 2622 56239 2654
rect 57397 2654 57463 2655
rect 57397 2622 57398 2654
rect 56238 2590 56244 2622
rect 55901 1838 55967 1839
rect 55901 1806 55902 1838
rect 55896 1774 55902 1806
rect 55966 1806 55967 1838
rect 55966 1774 55972 1806
rect 55896 1294 55972 1774
rect 55896 1230 55902 1294
rect 55966 1230 55972 1294
rect 55896 1224 55972 1230
rect 56168 0 56244 2590
rect 57392 2590 57398 2622
rect 57462 2622 57463 2654
rect 58621 2654 58687 2655
rect 58621 2622 58622 2654
rect 57462 2590 57468 2622
rect 57392 0 57468 2590
rect 58616 2590 58622 2622
rect 58686 2622 58687 2654
rect 58686 2590 58692 2622
rect 57669 1838 57735 1839
rect 57669 1806 57670 1838
rect 57664 1774 57670 1806
rect 57734 1806 57735 1838
rect 57734 1774 57740 1806
rect 57664 1294 57740 1774
rect 57664 1230 57670 1294
rect 57734 1230 57740 1294
rect 57664 1224 57740 1230
rect 58616 0 58692 2590
rect 59165 1838 59231 1839
rect 59165 1806 59166 1838
rect 59160 1774 59166 1806
rect 59230 1806 59231 1838
rect 59230 1774 59236 1806
rect 59160 1294 59236 1774
rect 59160 1230 59166 1294
rect 59230 1230 59236 1294
rect 59160 1224 59236 1230
rect 59296 0 59372 17550
rect 59704 17478 59780 17484
rect 59704 17414 59710 17478
rect 59774 17414 59780 17478
rect 59704 17070 59780 17414
rect 59704 17038 59710 17070
rect 59709 17006 59710 17038
rect 59774 17038 59780 17070
rect 59774 17006 59775 17038
rect 59709 17005 59775 17006
rect 59573 16934 59639 16935
rect 59573 16902 59574 16934
rect 59568 16870 59574 16902
rect 59638 16902 59639 16934
rect 59638 16870 59644 16902
rect 59568 16254 59644 16870
rect 59840 16526 59916 17958
rect 59976 17886 60052 19590
rect 60792 18974 60868 23534
rect 60792 18942 60798 18974
rect 60797 18910 60798 18942
rect 60862 18942 60868 18974
rect 64600 23534 64606 23566
rect 64670 23566 64671 23598
rect 70312 23598 70388 23604
rect 64670 23534 64676 23566
rect 64600 18974 64676 23534
rect 70312 23534 70318 23598
rect 70382 23534 70388 23598
rect 64872 22102 64948 22108
rect 64872 22038 64878 22102
rect 64942 22038 64948 22102
rect 64872 19654 64948 22038
rect 70040 22102 70116 22108
rect 70040 22038 70046 22102
rect 70110 22038 70116 22102
rect 64872 19622 64878 19654
rect 64877 19590 64878 19622
rect 64942 19622 64948 19654
rect 65008 19654 65084 19660
rect 64942 19590 64943 19622
rect 64877 19589 64943 19590
rect 65008 19590 65014 19654
rect 65078 19590 65084 19654
rect 60862 18910 60863 18942
rect 60797 18909 60863 18910
rect 64600 18910 64606 18974
rect 64670 18910 64676 18974
rect 64600 18904 64676 18910
rect 64877 18838 64943 18839
rect 64877 18806 64878 18838
rect 64872 18774 64878 18806
rect 64942 18806 64943 18838
rect 64942 18774 64948 18806
rect 64872 18158 64948 18774
rect 64872 18094 64878 18158
rect 64942 18094 64948 18158
rect 64872 18088 64948 18094
rect 59976 17854 59982 17886
rect 59981 17822 59982 17854
rect 60046 17854 60052 17886
rect 64736 18022 64812 18028
rect 64736 17958 64742 18022
rect 64806 17958 64812 18022
rect 60046 17822 60047 17854
rect 59981 17821 60047 17822
rect 64469 17614 64535 17615
rect 64469 17582 64470 17614
rect 59840 16494 59846 16526
rect 59845 16462 59846 16494
rect 59910 16494 59916 16526
rect 64464 17550 64470 17582
rect 64534 17582 64535 17614
rect 64534 17550 64540 17582
rect 59910 16462 59911 16494
rect 59845 16461 59911 16462
rect 59709 16390 59775 16391
rect 59709 16358 59710 16390
rect 59568 16190 59574 16254
rect 59638 16190 59644 16254
rect 59568 16184 59644 16190
rect 59704 16326 59710 16358
rect 59774 16358 59775 16390
rect 59774 16326 59780 16358
rect 59704 15574 59780 16326
rect 59704 15510 59710 15574
rect 59774 15510 59780 15574
rect 59704 15504 59780 15510
rect 59845 2654 59911 2655
rect 59845 2622 59846 2654
rect 59840 2590 59846 2622
rect 59910 2622 59911 2654
rect 60797 2654 60863 2655
rect 60797 2622 60798 2654
rect 59910 2590 59916 2622
rect 59840 0 59916 2590
rect 60792 2590 60798 2622
rect 60862 2622 60863 2654
rect 60862 2590 60868 2622
rect 60792 0 60868 2590
rect 61069 1838 61135 1839
rect 61069 1806 61070 1838
rect 61064 1774 61070 1806
rect 61134 1806 61135 1838
rect 62429 1838 62495 1839
rect 62429 1806 62430 1838
rect 61134 1774 61140 1806
rect 61064 1294 61140 1774
rect 61064 1230 61070 1294
rect 61134 1230 61140 1294
rect 61064 1224 61140 1230
rect 62424 1774 62430 1806
rect 62494 1806 62495 1838
rect 64061 1838 64127 1839
rect 64061 1806 64062 1838
rect 62494 1774 62500 1806
rect 62424 1294 62500 1774
rect 62424 1230 62430 1294
rect 62494 1230 62500 1294
rect 62424 1224 62500 1230
rect 64056 1774 64062 1806
rect 64126 1806 64127 1838
rect 64126 1774 64132 1806
rect 64056 1294 64132 1774
rect 64056 1230 64062 1294
rect 64126 1230 64132 1294
rect 64056 1224 64132 1230
rect 64464 0 64540 17550
rect 64736 16526 64812 17958
rect 65008 17886 65084 19590
rect 69904 19654 69980 19660
rect 69904 19590 69910 19654
rect 69974 19590 69980 19654
rect 70040 19654 70116 22038
rect 70040 19622 70046 19654
rect 69773 18838 69839 18839
rect 69773 18806 69774 18838
rect 69768 18774 69774 18806
rect 69838 18806 69839 18838
rect 69838 18774 69844 18806
rect 69768 18158 69844 18774
rect 69768 18094 69774 18158
rect 69838 18094 69844 18158
rect 69768 18088 69844 18094
rect 65008 17854 65014 17886
rect 65013 17822 65014 17854
rect 65078 17854 65084 17886
rect 69768 18022 69844 18028
rect 69768 17958 69774 18022
rect 69838 17958 69844 18022
rect 65078 17822 65079 17854
rect 65013 17821 65079 17822
rect 64872 17614 64948 17620
rect 64872 17550 64878 17614
rect 64942 17550 64948 17614
rect 69501 17614 69567 17615
rect 69501 17582 69502 17614
rect 64872 17070 64948 17550
rect 64872 17038 64878 17070
rect 64877 17006 64878 17038
rect 64942 17038 64948 17070
rect 69496 17550 69502 17582
rect 69566 17582 69567 17614
rect 69566 17550 69572 17582
rect 64942 17006 64943 17038
rect 64877 17005 64943 17006
rect 64877 16934 64943 16935
rect 64877 16902 64878 16934
rect 64736 16494 64742 16526
rect 64741 16462 64742 16494
rect 64806 16494 64812 16526
rect 64872 16870 64878 16902
rect 64942 16902 64943 16934
rect 64942 16870 64948 16902
rect 64806 16462 64807 16494
rect 64741 16461 64807 16462
rect 64741 16390 64807 16391
rect 64741 16358 64742 16390
rect 64736 16326 64742 16358
rect 64806 16358 64807 16390
rect 64806 16326 64812 16358
rect 64736 15574 64812 16326
rect 64872 16254 64948 16870
rect 64872 16190 64878 16254
rect 64942 16190 64948 16254
rect 64872 16184 64948 16190
rect 64736 15510 64742 15574
rect 64806 15510 64812 15574
rect 64736 15504 64812 15510
rect 65965 1838 66031 1839
rect 65965 1806 65966 1838
rect 65960 1774 65966 1806
rect 66030 1806 66031 1838
rect 67461 1838 67527 1839
rect 67461 1806 67462 1838
rect 66030 1774 66036 1806
rect 65960 1294 66036 1774
rect 65960 1230 65966 1294
rect 66030 1230 66036 1294
rect 65960 1224 66036 1230
rect 67456 1774 67462 1806
rect 67526 1806 67527 1838
rect 69229 1838 69295 1839
rect 69229 1806 69230 1838
rect 67526 1774 67532 1806
rect 67456 1294 67532 1774
rect 67456 1230 67462 1294
rect 67526 1230 67532 1294
rect 67456 1224 67532 1230
rect 69224 1774 69230 1806
rect 69294 1806 69295 1838
rect 69294 1774 69300 1806
rect 69224 1294 69300 1774
rect 69224 1230 69230 1294
rect 69294 1230 69300 1294
rect 69224 1224 69300 1230
rect 69496 0 69572 17550
rect 69768 16526 69844 17958
rect 69904 17886 69980 19590
rect 70045 19590 70046 19622
rect 70110 19622 70116 19654
rect 70110 19590 70111 19622
rect 70045 19589 70111 19590
rect 70312 18974 70388 23534
rect 75344 23598 75420 23604
rect 75344 23534 75350 23598
rect 75414 23534 75420 23598
rect 84189 23598 84255 23599
rect 84189 23566 84190 23598
rect 75072 22102 75148 22108
rect 75072 22038 75078 22102
rect 75142 22038 75148 22102
rect 70312 18942 70318 18974
rect 70317 18910 70318 18942
rect 70382 18942 70388 18974
rect 74936 19654 75012 19660
rect 74936 19590 74942 19654
rect 75006 19590 75012 19654
rect 75072 19654 75148 22038
rect 75072 19622 75078 19654
rect 70382 18910 70383 18942
rect 70317 18909 70383 18910
rect 74669 18838 74735 18839
rect 74669 18806 74670 18838
rect 74664 18774 74670 18806
rect 74734 18806 74735 18838
rect 74734 18774 74740 18806
rect 74664 18158 74740 18774
rect 74664 18094 74670 18158
rect 74734 18094 74740 18158
rect 74664 18088 74740 18094
rect 69904 17854 69910 17886
rect 69909 17822 69910 17854
rect 69974 17854 69980 17886
rect 74800 18022 74876 18028
rect 74800 17958 74806 18022
rect 74870 17958 74876 18022
rect 69974 17822 69975 17854
rect 69909 17821 69975 17822
rect 69904 17614 69980 17620
rect 69904 17550 69910 17614
rect 69974 17550 69980 17614
rect 74397 17614 74463 17615
rect 74397 17582 74398 17614
rect 69904 17070 69980 17550
rect 69904 17038 69910 17070
rect 69909 17006 69910 17038
rect 69974 17038 69980 17070
rect 74392 17550 74398 17582
rect 74462 17582 74463 17614
rect 74462 17550 74468 17582
rect 69974 17006 69975 17038
rect 69909 17005 69975 17006
rect 69909 16934 69975 16935
rect 69909 16902 69910 16934
rect 69768 16494 69774 16526
rect 69773 16462 69774 16494
rect 69838 16494 69844 16526
rect 69904 16870 69910 16902
rect 69974 16902 69975 16934
rect 69974 16870 69980 16902
rect 69838 16462 69839 16494
rect 69773 16461 69839 16462
rect 69773 16390 69839 16391
rect 69773 16358 69774 16390
rect 69768 16326 69774 16358
rect 69838 16358 69839 16390
rect 69838 16326 69844 16358
rect 69768 15574 69844 16326
rect 69904 16254 69980 16870
rect 69904 16190 69910 16254
rect 69974 16190 69980 16254
rect 69904 16184 69980 16190
rect 69768 15510 69774 15574
rect 69838 15510 69844 15574
rect 69768 15504 69844 15510
rect 70861 1838 70927 1839
rect 70861 1806 70862 1838
rect 70856 1774 70862 1806
rect 70926 1806 70927 1838
rect 72493 1838 72559 1839
rect 72493 1806 72494 1838
rect 70926 1774 70932 1806
rect 70856 1294 70932 1774
rect 70856 1230 70862 1294
rect 70926 1230 70932 1294
rect 70856 1224 70932 1230
rect 72488 1774 72494 1806
rect 72558 1806 72559 1838
rect 74261 1838 74327 1839
rect 74261 1806 74262 1838
rect 72558 1774 72564 1806
rect 72488 1294 72564 1774
rect 72488 1230 72494 1294
rect 72558 1230 72564 1294
rect 72488 1224 72564 1230
rect 74256 1774 74262 1806
rect 74326 1806 74327 1838
rect 74326 1774 74332 1806
rect 74256 1294 74332 1774
rect 74256 1230 74262 1294
rect 74326 1230 74332 1294
rect 74256 1224 74332 1230
rect 74392 0 74468 17550
rect 74664 17478 74740 17484
rect 74664 17414 74670 17478
rect 74734 17414 74740 17478
rect 74664 17070 74740 17414
rect 74664 17038 74670 17070
rect 74669 17006 74670 17038
rect 74734 17038 74740 17070
rect 74734 17006 74735 17038
rect 74669 17005 74735 17006
rect 74669 16934 74735 16935
rect 74669 16902 74670 16934
rect 74664 16870 74670 16902
rect 74734 16902 74735 16934
rect 74734 16870 74740 16902
rect 74533 16390 74599 16391
rect 74533 16358 74534 16390
rect 74528 16326 74534 16358
rect 74598 16358 74599 16390
rect 74598 16326 74604 16358
rect 74528 15574 74604 16326
rect 74664 16254 74740 16870
rect 74800 16526 74876 17958
rect 74936 17886 75012 19590
rect 75077 19590 75078 19622
rect 75142 19622 75148 19654
rect 75142 19590 75143 19622
rect 75077 19589 75143 19590
rect 75344 18974 75420 23534
rect 84184 23534 84190 23566
rect 84254 23566 84255 23598
rect 89629 23598 89695 23599
rect 89629 23566 89630 23598
rect 84254 23534 84260 23566
rect 79832 22102 79908 22108
rect 79832 22038 79838 22102
rect 79902 22038 79908 22102
rect 79832 19654 79908 22038
rect 79832 19622 79838 19654
rect 79837 19590 79838 19622
rect 79902 19622 79908 19654
rect 79968 19654 80044 19660
rect 79902 19590 79903 19622
rect 79837 19589 79903 19590
rect 79968 19590 79974 19654
rect 80038 19590 80044 19654
rect 75344 18942 75350 18974
rect 75349 18910 75350 18942
rect 75414 18942 75420 18974
rect 75414 18910 75415 18942
rect 75349 18909 75415 18910
rect 79701 18838 79767 18839
rect 79701 18806 79702 18838
rect 79696 18774 79702 18806
rect 79766 18806 79767 18838
rect 79766 18774 79772 18806
rect 79696 18158 79772 18774
rect 79696 18094 79702 18158
rect 79766 18094 79772 18158
rect 79696 18088 79772 18094
rect 74936 17854 74942 17886
rect 74941 17822 74942 17854
rect 75006 17854 75012 17886
rect 79832 18022 79908 18028
rect 79832 17958 79838 18022
rect 79902 17958 79908 18022
rect 75006 17822 75007 17854
rect 74941 17821 75007 17822
rect 79429 17614 79495 17615
rect 79429 17582 79430 17614
rect 79424 17550 79430 17582
rect 79494 17582 79495 17614
rect 79494 17550 79500 17582
rect 74800 16494 74806 16526
rect 74805 16462 74806 16494
rect 74870 16494 74876 16526
rect 79288 16934 79364 16940
rect 79288 16870 79294 16934
rect 79358 16870 79364 16934
rect 74870 16462 74871 16494
rect 74805 16461 74871 16462
rect 74664 16190 74670 16254
rect 74734 16190 74740 16254
rect 74664 16184 74740 16190
rect 79288 16118 79364 16870
rect 79288 16086 79294 16118
rect 79293 16054 79294 16086
rect 79358 16086 79364 16118
rect 79358 16054 79359 16086
rect 79293 16053 79359 16054
rect 74528 15510 74534 15574
rect 74598 15510 74604 15574
rect 74528 15504 74604 15510
rect 75893 1838 75959 1839
rect 75893 1806 75894 1838
rect 75888 1774 75894 1806
rect 75958 1806 75959 1838
rect 77661 1838 77727 1839
rect 77661 1806 77662 1838
rect 75958 1774 75964 1806
rect 75888 1294 75964 1774
rect 75888 1230 75894 1294
rect 75958 1230 75964 1294
rect 75888 1224 75964 1230
rect 77656 1774 77662 1806
rect 77726 1806 77727 1838
rect 79293 1838 79359 1839
rect 79293 1806 79294 1838
rect 77726 1774 77732 1806
rect 77656 1294 77732 1774
rect 77656 1230 77662 1294
rect 77726 1230 77732 1294
rect 77656 1224 77732 1230
rect 79288 1774 79294 1806
rect 79358 1806 79359 1838
rect 79358 1774 79364 1806
rect 79288 1294 79364 1774
rect 79288 1230 79294 1294
rect 79358 1230 79364 1294
rect 79288 1224 79364 1230
rect 79424 0 79500 17550
rect 79696 17478 79772 17484
rect 79696 17414 79702 17478
rect 79766 17414 79772 17478
rect 79696 17070 79772 17414
rect 79696 17038 79702 17070
rect 79701 17006 79702 17038
rect 79766 17038 79772 17070
rect 79766 17006 79767 17038
rect 79701 17005 79767 17006
rect 79832 16526 79908 17958
rect 79968 17886 80044 19590
rect 84184 18974 84260 23534
rect 89624 23534 89630 23566
rect 89694 23566 89695 23598
rect 95336 23598 95412 23604
rect 89694 23534 89700 23566
rect 85000 22102 85076 22108
rect 85000 22038 85006 22102
rect 85070 22038 85076 22102
rect 84184 18910 84190 18974
rect 84254 18910 84260 18974
rect 84184 18904 84260 18910
rect 84864 19654 84940 19660
rect 84864 19590 84870 19654
rect 84934 19590 84940 19654
rect 85000 19654 85076 22038
rect 85000 19622 85006 19654
rect 84733 18838 84799 18839
rect 84733 18806 84734 18838
rect 84728 18774 84734 18806
rect 84798 18806 84799 18838
rect 84798 18774 84804 18806
rect 84728 18158 84804 18774
rect 84728 18094 84734 18158
rect 84798 18094 84804 18158
rect 84728 18088 84804 18094
rect 79968 17854 79974 17886
rect 79973 17822 79974 17854
rect 80038 17854 80044 17886
rect 84728 18022 84804 18028
rect 84728 17958 84734 18022
rect 84798 17958 84804 18022
rect 80038 17822 80039 17854
rect 79973 17821 80039 17822
rect 84325 17614 84391 17615
rect 84325 17582 84326 17614
rect 84320 17550 84326 17582
rect 84390 17582 84391 17614
rect 84390 17550 84396 17582
rect 79973 16934 80039 16935
rect 79973 16902 79974 16934
rect 79832 16494 79838 16526
rect 79837 16462 79838 16494
rect 79902 16494 79908 16526
rect 79968 16870 79974 16902
rect 80038 16902 80039 16934
rect 80038 16870 80044 16902
rect 79902 16462 79903 16494
rect 79837 16461 79903 16462
rect 79701 16390 79767 16391
rect 79701 16358 79702 16390
rect 79696 16326 79702 16358
rect 79766 16358 79767 16390
rect 79766 16326 79772 16358
rect 79696 15574 79772 16326
rect 79968 16254 80044 16870
rect 79968 16190 79974 16254
rect 80038 16190 80044 16254
rect 79968 16184 80044 16190
rect 79696 15510 79702 15574
rect 79766 15510 79772 15574
rect 79696 15504 79772 15510
rect 80925 1838 80991 1839
rect 80925 1806 80926 1838
rect 80920 1774 80926 1806
rect 80990 1806 80991 1838
rect 82693 1838 82759 1839
rect 82693 1806 82694 1838
rect 80990 1774 80996 1806
rect 80920 1294 80996 1774
rect 80920 1230 80926 1294
rect 80990 1230 80996 1294
rect 80920 1224 80996 1230
rect 82688 1774 82694 1806
rect 82758 1806 82759 1838
rect 82758 1774 82764 1806
rect 82688 1294 82764 1774
rect 82688 1230 82694 1294
rect 82758 1230 82764 1294
rect 82688 1224 82764 1230
rect 84320 0 84396 17550
rect 84728 16526 84804 17958
rect 84864 17886 84940 19590
rect 85005 19590 85006 19622
rect 85070 19622 85076 19654
rect 85070 19590 85071 19622
rect 85005 19589 85071 19590
rect 89624 18974 89700 23534
rect 95336 23534 95342 23598
rect 95406 23534 95412 23598
rect 99557 23598 99623 23599
rect 99557 23566 99558 23598
rect 90032 22102 90108 22108
rect 90032 22038 90038 22102
rect 90102 22038 90108 22102
rect 89624 18910 89630 18974
rect 89694 18910 89700 18974
rect 89624 18904 89700 18910
rect 89896 19654 89972 19660
rect 89896 19590 89902 19654
rect 89966 19590 89972 19654
rect 90032 19654 90108 22038
rect 90032 19622 90038 19654
rect 89765 18838 89831 18839
rect 89765 18806 89766 18838
rect 89760 18774 89766 18806
rect 89830 18806 89831 18838
rect 89830 18774 89836 18806
rect 89760 18158 89836 18774
rect 89760 18094 89766 18158
rect 89830 18094 89836 18158
rect 89760 18088 89836 18094
rect 84864 17854 84870 17886
rect 84869 17822 84870 17854
rect 84934 17854 84940 17886
rect 89760 18022 89836 18028
rect 89760 17958 89766 18022
rect 89830 17958 89836 18022
rect 84934 17822 84935 17854
rect 84869 17821 84935 17822
rect 84864 17614 84940 17620
rect 84864 17550 84870 17614
rect 84934 17550 84940 17614
rect 89357 17614 89423 17615
rect 89357 17582 89358 17614
rect 84864 17070 84940 17550
rect 84864 17038 84870 17070
rect 84869 17006 84870 17038
rect 84934 17038 84940 17070
rect 89352 17550 89358 17582
rect 89422 17582 89423 17614
rect 89422 17550 89428 17582
rect 84934 17006 84935 17038
rect 84869 17005 84935 17006
rect 84869 16934 84935 16935
rect 84869 16902 84870 16934
rect 84728 16494 84734 16526
rect 84733 16462 84734 16494
rect 84798 16494 84804 16526
rect 84864 16870 84870 16902
rect 84934 16902 84935 16934
rect 84934 16870 84940 16902
rect 84798 16462 84799 16494
rect 84733 16461 84799 16462
rect 84597 16390 84663 16391
rect 84597 16358 84598 16390
rect 84592 16326 84598 16358
rect 84662 16358 84663 16390
rect 84662 16326 84668 16358
rect 84592 15574 84668 16326
rect 84864 16254 84940 16870
rect 84864 16190 84870 16254
rect 84934 16190 84940 16254
rect 84864 16184 84940 16190
rect 84592 15510 84598 15574
rect 84662 15510 84668 15574
rect 84592 15504 84668 15510
rect 84597 1838 84663 1839
rect 84597 1806 84598 1838
rect 84592 1774 84598 1806
rect 84662 1806 84663 1838
rect 85957 1838 86023 1839
rect 85957 1806 85958 1838
rect 84662 1774 84668 1806
rect 84592 1294 84668 1774
rect 84592 1230 84598 1294
rect 84662 1230 84668 1294
rect 84592 1224 84668 1230
rect 85952 1774 85958 1806
rect 86022 1806 86023 1838
rect 87725 1838 87791 1839
rect 87725 1806 87726 1838
rect 86022 1774 86028 1806
rect 85952 1294 86028 1774
rect 85952 1230 85958 1294
rect 86022 1230 86028 1294
rect 85952 1224 86028 1230
rect 87720 1774 87726 1806
rect 87790 1806 87791 1838
rect 87790 1774 87796 1806
rect 87720 1294 87796 1774
rect 87720 1230 87726 1294
rect 87790 1230 87796 1294
rect 87720 1224 87796 1230
rect 89352 0 89428 17550
rect 89624 17478 89700 17484
rect 89624 17414 89630 17478
rect 89694 17414 89700 17478
rect 89624 17070 89700 17414
rect 89624 17038 89630 17070
rect 89629 17006 89630 17038
rect 89694 17038 89700 17070
rect 89694 17006 89695 17038
rect 89629 17005 89695 17006
rect 89629 16934 89695 16935
rect 89629 16902 89630 16934
rect 89624 16870 89630 16902
rect 89694 16902 89695 16934
rect 89694 16870 89700 16902
rect 89493 16390 89559 16391
rect 89493 16358 89494 16390
rect 89488 16326 89494 16358
rect 89558 16358 89559 16390
rect 89558 16326 89564 16358
rect 89488 15574 89564 16326
rect 89624 16254 89700 16870
rect 89760 16526 89836 17958
rect 89896 17886 89972 19590
rect 90037 19590 90038 19622
rect 90102 19622 90108 19654
rect 94792 22102 94868 22108
rect 94792 22038 94798 22102
rect 94862 22038 94868 22102
rect 94792 19654 94868 22038
rect 94792 19622 94798 19654
rect 90102 19590 90103 19622
rect 90037 19589 90103 19590
rect 94797 19590 94798 19622
rect 94862 19622 94868 19654
rect 94928 19654 95004 19660
rect 94862 19590 94863 19622
rect 94797 19589 94863 19590
rect 94928 19590 94934 19654
rect 94998 19590 95004 19654
rect 94797 18838 94863 18839
rect 94797 18806 94798 18838
rect 94792 18774 94798 18806
rect 94862 18806 94863 18838
rect 94862 18774 94868 18806
rect 94792 18158 94868 18774
rect 94792 18094 94798 18158
rect 94862 18094 94868 18158
rect 94792 18088 94868 18094
rect 89896 17854 89902 17886
rect 89901 17822 89902 17854
rect 89966 17854 89972 17886
rect 94792 18022 94868 18028
rect 94792 17958 94798 18022
rect 94862 17958 94868 18022
rect 89966 17822 89967 17854
rect 89901 17821 89967 17822
rect 94389 17614 94455 17615
rect 94389 17582 94390 17614
rect 89760 16494 89766 16526
rect 89765 16462 89766 16494
rect 89830 16494 89836 16526
rect 94384 17550 94390 17582
rect 94454 17582 94455 17614
rect 94454 17550 94460 17582
rect 89830 16462 89831 16494
rect 89765 16461 89831 16462
rect 89624 16190 89630 16254
rect 89694 16190 89700 16254
rect 89624 16184 89700 16190
rect 89488 15510 89494 15574
rect 89558 15510 89564 15574
rect 89488 15504 89564 15510
rect 89493 1838 89559 1839
rect 89493 1806 89494 1838
rect 89488 1774 89494 1806
rect 89558 1806 89559 1838
rect 91125 1838 91191 1839
rect 91125 1806 91126 1838
rect 89558 1774 89564 1806
rect 89488 1294 89564 1774
rect 89488 1230 89494 1294
rect 89558 1230 89564 1294
rect 89488 1224 89564 1230
rect 91120 1774 91126 1806
rect 91190 1806 91191 1838
rect 92621 1838 92687 1839
rect 92621 1806 92622 1838
rect 91190 1774 91196 1806
rect 91120 1294 91196 1774
rect 91120 1230 91126 1294
rect 91190 1230 91196 1294
rect 91120 1224 91196 1230
rect 92616 1774 92622 1806
rect 92686 1806 92687 1838
rect 92686 1774 92692 1806
rect 92616 1294 92692 1774
rect 92616 1230 92622 1294
rect 92686 1230 92692 1294
rect 92616 1224 92692 1230
rect 94384 0 94460 17550
rect 94656 17478 94732 17484
rect 94656 17414 94662 17478
rect 94726 17414 94732 17478
rect 94656 17070 94732 17414
rect 94656 17038 94662 17070
rect 94661 17006 94662 17038
rect 94726 17038 94732 17070
rect 94726 17006 94727 17038
rect 94661 17005 94727 17006
rect 94792 16526 94868 17958
rect 94928 17886 95004 19590
rect 95336 18974 95412 23534
rect 95336 18942 95342 18974
rect 95341 18910 95342 18942
rect 95406 18942 95412 18974
rect 99552 23534 99558 23566
rect 99622 23566 99623 23598
rect 105264 23598 105340 23604
rect 99622 23534 99628 23566
rect 99552 18974 99628 23534
rect 105264 23534 105270 23598
rect 105334 23534 105340 23598
rect 99960 22102 100036 22108
rect 99960 22038 99966 22102
rect 100030 22038 100036 22102
rect 95406 18910 95407 18942
rect 95341 18909 95407 18910
rect 99552 18910 99558 18974
rect 99622 18910 99628 18974
rect 99552 18904 99628 18910
rect 99824 19654 99900 19660
rect 99824 19590 99830 19654
rect 99894 19590 99900 19654
rect 99960 19654 100036 22038
rect 104992 22102 105068 22108
rect 104992 22038 104998 22102
rect 105062 22038 105068 22102
rect 99960 19622 99966 19654
rect 99693 18838 99759 18839
rect 99693 18806 99694 18838
rect 99688 18774 99694 18806
rect 99758 18806 99759 18838
rect 99758 18774 99764 18806
rect 99688 18158 99764 18774
rect 99688 18094 99694 18158
rect 99758 18094 99764 18158
rect 99688 18088 99764 18094
rect 94928 17854 94934 17886
rect 94933 17822 94934 17854
rect 94998 17854 95004 17886
rect 99552 18022 99628 18028
rect 99552 17958 99558 18022
rect 99622 17958 99628 18022
rect 94998 17822 94999 17854
rect 94933 17821 94999 17822
rect 99421 17614 99487 17615
rect 99421 17582 99422 17614
rect 99416 17550 99422 17582
rect 99486 17582 99487 17614
rect 99486 17550 99492 17582
rect 94933 16934 94999 16935
rect 94933 16902 94934 16934
rect 94792 16494 94798 16526
rect 94797 16462 94798 16494
rect 94862 16494 94868 16526
rect 94928 16870 94934 16902
rect 94998 16902 94999 16934
rect 94998 16870 95004 16902
rect 94862 16462 94863 16494
rect 94797 16461 94863 16462
rect 94661 16390 94727 16391
rect 94661 16358 94662 16390
rect 94656 16326 94662 16358
rect 94726 16358 94727 16390
rect 94726 16326 94732 16358
rect 94656 15574 94732 16326
rect 94928 16254 95004 16870
rect 94928 16190 94934 16254
rect 94998 16190 95004 16254
rect 94928 16184 95004 16190
rect 94656 15510 94662 15574
rect 94726 15510 94732 15574
rect 94656 15504 94732 15510
rect 94661 1838 94727 1839
rect 94661 1806 94662 1838
rect 94656 1774 94662 1806
rect 94726 1806 94727 1838
rect 96157 1838 96223 1839
rect 96157 1806 96158 1838
rect 94726 1774 94732 1806
rect 94656 1294 94732 1774
rect 94656 1230 94662 1294
rect 94726 1230 94732 1294
rect 94656 1224 94732 1230
rect 96152 1774 96158 1806
rect 96222 1806 96223 1838
rect 97789 1838 97855 1839
rect 97789 1806 97790 1838
rect 96222 1774 96228 1806
rect 96152 1294 96228 1774
rect 96152 1230 96158 1294
rect 96222 1230 96228 1294
rect 96152 1224 96228 1230
rect 97784 1774 97790 1806
rect 97854 1806 97855 1838
rect 97854 1774 97860 1806
rect 97784 1294 97860 1774
rect 97784 1230 97790 1294
rect 97854 1230 97860 1294
rect 97784 1224 97860 1230
rect 99416 0 99492 17550
rect 99552 16526 99628 17958
rect 99824 17886 99900 19590
rect 99965 19590 99966 19622
rect 100030 19622 100036 19654
rect 104856 19654 104932 19660
rect 100030 19590 100031 19622
rect 99965 19589 100031 19590
rect 104856 19590 104862 19654
rect 104926 19590 104932 19654
rect 104992 19654 105068 22038
rect 104992 19622 104998 19654
rect 104589 18838 104655 18839
rect 104589 18806 104590 18838
rect 104584 18774 104590 18806
rect 104654 18806 104655 18838
rect 104654 18774 104660 18806
rect 104584 18158 104660 18774
rect 104584 18094 104590 18158
rect 104654 18094 104660 18158
rect 104584 18088 104660 18094
rect 99824 17854 99830 17886
rect 99829 17822 99830 17854
rect 99894 17854 99900 17886
rect 104720 18022 104796 18028
rect 104720 17958 104726 18022
rect 104790 17958 104796 18022
rect 99894 17822 99895 17854
rect 99829 17821 99895 17822
rect 99688 17614 99764 17620
rect 99688 17550 99694 17614
rect 99758 17550 99764 17614
rect 104317 17614 104383 17615
rect 104317 17582 104318 17614
rect 99688 17070 99764 17550
rect 99688 17038 99694 17070
rect 99693 17006 99694 17038
rect 99758 17038 99764 17070
rect 104312 17550 104318 17582
rect 104382 17582 104383 17614
rect 104382 17550 104388 17582
rect 99758 17006 99759 17038
rect 99693 17005 99759 17006
rect 99552 16494 99558 16526
rect 99557 16462 99558 16494
rect 99622 16494 99628 16526
rect 99688 16934 99764 16940
rect 99688 16870 99694 16934
rect 99758 16870 99764 16934
rect 99829 16934 99895 16935
rect 99829 16902 99830 16934
rect 99622 16462 99623 16494
rect 99557 16461 99623 16462
rect 99557 16390 99623 16391
rect 99557 16358 99558 16390
rect 99552 16326 99558 16358
rect 99622 16358 99623 16390
rect 99622 16326 99628 16358
rect 99552 15574 99628 16326
rect 99688 16118 99764 16870
rect 99824 16870 99830 16902
rect 99894 16902 99895 16934
rect 99894 16870 99900 16902
rect 99824 16254 99900 16870
rect 99824 16190 99830 16254
rect 99894 16190 99900 16254
rect 99824 16184 99900 16190
rect 99688 16086 99694 16118
rect 99693 16054 99694 16086
rect 99758 16086 99764 16118
rect 99758 16054 99759 16086
rect 99693 16053 99759 16054
rect 99552 15510 99558 15574
rect 99622 15510 99628 15574
rect 99552 15504 99628 15510
rect 99557 1838 99623 1839
rect 99557 1806 99558 1838
rect 99552 1774 99558 1806
rect 99622 1806 99623 1838
rect 101189 1838 101255 1839
rect 101189 1806 101190 1838
rect 99622 1774 99628 1806
rect 99552 1294 99628 1774
rect 99552 1230 99558 1294
rect 99622 1230 99628 1294
rect 99552 1224 99628 1230
rect 101184 1774 101190 1806
rect 101254 1806 101255 1838
rect 102957 1838 103023 1839
rect 102957 1806 102958 1838
rect 101254 1774 101260 1806
rect 101184 1294 101260 1774
rect 101184 1230 101190 1294
rect 101254 1230 101260 1294
rect 101184 1224 101260 1230
rect 102952 1774 102958 1806
rect 103022 1806 103023 1838
rect 103022 1774 103028 1806
rect 102952 1294 103028 1774
rect 102952 1230 102958 1294
rect 103022 1230 103028 1294
rect 102952 1224 103028 1230
rect 104312 0 104388 17550
rect 104584 17478 104660 17484
rect 104584 17414 104590 17478
rect 104654 17414 104660 17478
rect 104584 17070 104660 17414
rect 104584 17038 104590 17070
rect 104589 17006 104590 17038
rect 104654 17038 104660 17070
rect 104654 17006 104655 17038
rect 104589 17005 104655 17006
rect 104453 16934 104519 16935
rect 104453 16902 104454 16934
rect 104448 16870 104454 16902
rect 104518 16902 104519 16934
rect 104518 16870 104524 16902
rect 104448 16254 104524 16870
rect 104720 16526 104796 17958
rect 104856 17886 104932 19590
rect 104997 19590 104998 19622
rect 105062 19622 105068 19654
rect 105062 19590 105063 19622
rect 104997 19589 105063 19590
rect 105264 18974 105340 23534
rect 110296 23598 110372 23604
rect 110296 23534 110302 23598
rect 110366 23534 110372 23598
rect 114517 23598 114583 23599
rect 114517 23566 114518 23598
rect 110024 22102 110100 22108
rect 110024 22038 110030 22102
rect 110094 22038 110100 22102
rect 105264 18942 105270 18974
rect 105269 18910 105270 18942
rect 105334 18942 105340 18974
rect 109888 19654 109964 19660
rect 109888 19590 109894 19654
rect 109958 19590 109964 19654
rect 110024 19654 110100 22038
rect 110024 19622 110030 19654
rect 105334 18910 105335 18942
rect 105269 18909 105335 18910
rect 109757 18838 109823 18839
rect 109757 18806 109758 18838
rect 109752 18774 109758 18806
rect 109822 18806 109823 18838
rect 109822 18774 109828 18806
rect 109752 18158 109828 18774
rect 109752 18094 109758 18158
rect 109822 18094 109828 18158
rect 109752 18088 109828 18094
rect 104856 17854 104862 17886
rect 104861 17822 104862 17854
rect 104926 17854 104932 17886
rect 109752 18022 109828 18028
rect 109752 17958 109758 18022
rect 109822 17958 109828 18022
rect 104926 17822 104927 17854
rect 104861 17821 104927 17822
rect 109077 17614 109143 17615
rect 109077 17582 109078 17614
rect 104720 16494 104726 16526
rect 104725 16462 104726 16494
rect 104790 16494 104796 16526
rect 109072 17550 109078 17582
rect 109142 17582 109143 17614
rect 109142 17550 109148 17582
rect 104790 16462 104791 16494
rect 104725 16461 104791 16462
rect 104589 16390 104655 16391
rect 104589 16358 104590 16390
rect 104448 16190 104454 16254
rect 104518 16190 104524 16254
rect 104448 16184 104524 16190
rect 104584 16326 104590 16358
rect 104654 16358 104655 16390
rect 104654 16326 104660 16358
rect 104584 15574 104660 16326
rect 104584 15510 104590 15574
rect 104654 15510 104660 15574
rect 104584 15504 104660 15510
rect 104453 1838 104519 1839
rect 104453 1806 104454 1838
rect 104448 1774 104454 1806
rect 104518 1806 104519 1838
rect 106221 1838 106287 1839
rect 106221 1806 106222 1838
rect 104518 1774 104524 1806
rect 104448 1294 104524 1774
rect 104448 1230 104454 1294
rect 104518 1230 104524 1294
rect 104448 1224 104524 1230
rect 106216 1774 106222 1806
rect 106286 1806 106287 1838
rect 107853 1838 107919 1839
rect 107853 1806 107854 1838
rect 106286 1774 106292 1806
rect 106216 1294 106292 1774
rect 106216 1230 106222 1294
rect 106286 1230 106292 1294
rect 106216 1224 106292 1230
rect 107848 1774 107854 1806
rect 107918 1806 107919 1838
rect 107918 1774 107924 1806
rect 107848 1294 107924 1774
rect 107848 1230 107854 1294
rect 107918 1230 107924 1294
rect 107848 1224 107924 1230
rect 109072 0 109148 17550
rect 109616 17478 109692 17484
rect 109616 17414 109622 17478
rect 109686 17414 109692 17478
rect 109616 17070 109692 17414
rect 109616 17038 109622 17070
rect 109621 17006 109622 17038
rect 109686 17038 109692 17070
rect 109686 17006 109687 17038
rect 109621 17005 109687 17006
rect 109485 16934 109551 16935
rect 109485 16902 109486 16934
rect 109480 16870 109486 16902
rect 109550 16902 109551 16934
rect 109550 16870 109556 16902
rect 109480 16254 109556 16870
rect 109752 16526 109828 17958
rect 109888 17886 109964 19590
rect 110029 19590 110030 19622
rect 110094 19622 110100 19654
rect 110094 19590 110095 19622
rect 110029 19589 110095 19590
rect 110296 18974 110372 23534
rect 110296 18942 110302 18974
rect 110301 18910 110302 18942
rect 110366 18942 110372 18974
rect 114512 23534 114518 23566
rect 114582 23566 114583 23598
rect 119277 23598 119343 23599
rect 119277 23566 119278 23598
rect 114582 23534 114588 23566
rect 114512 18974 114588 23534
rect 119272 23534 119278 23566
rect 119342 23566 119343 23598
rect 124581 23598 124647 23599
rect 124581 23566 124582 23598
rect 119342 23534 119348 23566
rect 114784 22102 114860 22108
rect 114784 22038 114790 22102
rect 114854 22038 114860 22102
rect 114784 19654 114860 22038
rect 114784 19622 114790 19654
rect 114789 19590 114790 19622
rect 114854 19622 114860 19654
rect 114920 19654 114996 19660
rect 114854 19590 114855 19622
rect 114789 19589 114855 19590
rect 114920 19590 114926 19654
rect 114990 19590 114996 19654
rect 110366 18910 110367 18942
rect 110301 18909 110367 18910
rect 114512 18910 114518 18974
rect 114582 18910 114588 18974
rect 114512 18904 114588 18910
rect 114789 18838 114855 18839
rect 114789 18806 114790 18838
rect 114784 18774 114790 18806
rect 114854 18806 114855 18838
rect 114854 18774 114860 18806
rect 114784 18158 114860 18774
rect 114784 18094 114790 18158
rect 114854 18094 114860 18158
rect 114784 18088 114860 18094
rect 109888 17854 109894 17886
rect 109893 17822 109894 17854
rect 109958 17854 109964 17886
rect 114784 18022 114860 18028
rect 114784 17958 114790 18022
rect 114854 17958 114860 18022
rect 109958 17822 109959 17854
rect 109893 17821 109959 17822
rect 114381 17614 114447 17615
rect 114381 17582 114382 17614
rect 109752 16494 109758 16526
rect 109757 16462 109758 16494
rect 109822 16494 109828 16526
rect 114376 17550 114382 17582
rect 114446 17582 114447 17614
rect 114446 17550 114452 17582
rect 109822 16462 109823 16494
rect 109757 16461 109823 16462
rect 109621 16390 109687 16391
rect 109621 16358 109622 16390
rect 109480 16190 109486 16254
rect 109550 16190 109556 16254
rect 109480 16184 109556 16190
rect 109616 16326 109622 16358
rect 109686 16358 109687 16390
rect 109686 16326 109692 16358
rect 109616 15574 109692 16326
rect 109616 15510 109622 15574
rect 109686 15510 109692 15574
rect 109616 15504 109692 15510
rect 109485 1838 109551 1839
rect 109485 1806 109486 1838
rect 109480 1774 109486 1806
rect 109550 1806 109551 1838
rect 111117 1838 111183 1839
rect 111117 1806 111118 1838
rect 109550 1774 109556 1806
rect 109480 1294 109556 1774
rect 109480 1230 109486 1294
rect 109550 1230 109556 1294
rect 109480 1224 109556 1230
rect 111112 1774 111118 1806
rect 111182 1806 111183 1838
rect 112885 1838 112951 1839
rect 112885 1806 112886 1838
rect 111182 1774 111188 1806
rect 111112 1294 111188 1774
rect 111112 1230 111118 1294
rect 111182 1230 111188 1294
rect 111112 1224 111188 1230
rect 112880 1774 112886 1806
rect 112950 1806 112951 1838
rect 112950 1774 112956 1806
rect 112880 1294 112956 1774
rect 112880 1230 112886 1294
rect 112950 1230 112956 1294
rect 112880 1224 112956 1230
rect 114376 0 114452 17550
rect 114648 17478 114724 17484
rect 114648 17414 114654 17478
rect 114718 17414 114724 17478
rect 114648 17070 114724 17414
rect 114648 17038 114654 17070
rect 114653 17006 114654 17038
rect 114718 17038 114724 17070
rect 114718 17006 114719 17038
rect 114653 17005 114719 17006
rect 114653 16934 114719 16935
rect 114653 16902 114654 16934
rect 114648 16870 114654 16902
rect 114718 16902 114719 16934
rect 114718 16870 114724 16902
rect 114517 16390 114583 16391
rect 114517 16358 114518 16390
rect 114512 16326 114518 16358
rect 114582 16358 114583 16390
rect 114582 16326 114588 16358
rect 114512 15574 114588 16326
rect 114648 16254 114724 16870
rect 114784 16526 114860 17958
rect 114920 17886 114996 19590
rect 119272 18974 119348 23534
rect 124576 23534 124582 23566
rect 124646 23566 124647 23598
rect 130288 23598 130364 23604
rect 124646 23534 124652 23566
rect 119952 22102 120028 22108
rect 119952 22038 119958 22102
rect 120022 22038 120028 22102
rect 119272 18910 119278 18974
rect 119342 18910 119348 18974
rect 119272 18904 119348 18910
rect 119816 19654 119892 19660
rect 119816 19590 119822 19654
rect 119886 19590 119892 19654
rect 119952 19654 120028 22038
rect 119952 19622 119958 19654
rect 119549 18838 119615 18839
rect 119549 18806 119550 18838
rect 119544 18774 119550 18806
rect 119614 18806 119615 18838
rect 119614 18774 119620 18806
rect 119544 18158 119620 18774
rect 119544 18094 119550 18158
rect 119614 18094 119620 18158
rect 119544 18088 119620 18094
rect 114920 17854 114926 17886
rect 114925 17822 114926 17854
rect 114990 17854 114996 17886
rect 119680 18022 119756 18028
rect 119680 17958 119686 18022
rect 119750 17958 119756 18022
rect 114990 17822 114991 17854
rect 114925 17821 114991 17822
rect 119277 17614 119343 17615
rect 119277 17582 119278 17614
rect 114784 16494 114790 16526
rect 114789 16462 114790 16494
rect 114854 16494 114860 16526
rect 119272 17550 119278 17582
rect 119342 17582 119343 17614
rect 119342 17550 119348 17582
rect 114854 16462 114855 16494
rect 114789 16461 114855 16462
rect 114648 16190 114654 16254
rect 114718 16190 114724 16254
rect 114648 16184 114724 16190
rect 114512 15510 114518 15574
rect 114582 15510 114588 15574
rect 114512 15504 114588 15510
rect 114653 1838 114719 1839
rect 114653 1806 114654 1838
rect 114648 1774 114654 1806
rect 114718 1806 114719 1838
rect 116149 1838 116215 1839
rect 116149 1806 116150 1838
rect 114718 1774 114724 1806
rect 114648 1294 114724 1774
rect 114648 1230 114654 1294
rect 114718 1230 114724 1294
rect 114648 1224 114724 1230
rect 116144 1774 116150 1806
rect 116214 1806 116215 1838
rect 117917 1838 117983 1839
rect 117917 1806 117918 1838
rect 116214 1774 116220 1806
rect 116144 1294 116220 1774
rect 116144 1230 116150 1294
rect 116214 1230 116220 1294
rect 116144 1224 116220 1230
rect 117912 1774 117918 1806
rect 117982 1806 117983 1838
rect 117982 1774 117988 1806
rect 117912 1294 117988 1774
rect 117912 1230 117918 1294
rect 117982 1230 117988 1294
rect 117912 1224 117988 1230
rect 119272 0 119348 17550
rect 119544 16934 119620 16940
rect 119544 16870 119550 16934
rect 119614 16870 119620 16934
rect 119544 16118 119620 16870
rect 119680 16526 119756 17958
rect 119816 17886 119892 19590
rect 119957 19590 119958 19622
rect 120022 19622 120028 19654
rect 120022 19590 120023 19622
rect 119957 19589 120023 19590
rect 124576 18974 124652 23534
rect 130288 23534 130294 23598
rect 130358 23534 130364 23598
rect 134101 23598 134167 23599
rect 134101 23566 134102 23598
rect 124984 22102 125060 22108
rect 124984 22038 124990 22102
rect 125054 22038 125060 22102
rect 124576 18910 124582 18974
rect 124646 18910 124652 18974
rect 124576 18904 124652 18910
rect 124848 19654 124924 19660
rect 124848 19590 124854 19654
rect 124918 19590 124924 19654
rect 124984 19654 125060 22038
rect 124984 19622 124990 19654
rect 124581 18838 124647 18839
rect 124581 18806 124582 18838
rect 124576 18774 124582 18806
rect 124646 18806 124647 18838
rect 124646 18774 124652 18806
rect 124576 18158 124652 18774
rect 124576 18094 124582 18158
rect 124646 18094 124652 18158
rect 124576 18088 124652 18094
rect 119816 17854 119822 17886
rect 119821 17822 119822 17854
rect 119886 17854 119892 17886
rect 124712 18022 124788 18028
rect 124712 17958 124718 18022
rect 124782 17958 124788 18022
rect 119886 17822 119887 17854
rect 119821 17821 119887 17822
rect 119816 17614 119892 17620
rect 119816 17550 119822 17614
rect 119886 17550 119892 17614
rect 124309 17614 124375 17615
rect 124309 17582 124310 17614
rect 119816 17070 119892 17550
rect 119816 17038 119822 17070
rect 119821 17006 119822 17038
rect 119886 17038 119892 17070
rect 124304 17550 124310 17582
rect 124374 17582 124375 17614
rect 124374 17550 124380 17582
rect 119886 17006 119887 17038
rect 119821 17005 119887 17006
rect 119821 16934 119887 16935
rect 119821 16902 119822 16934
rect 119680 16494 119686 16526
rect 119685 16462 119686 16494
rect 119750 16494 119756 16526
rect 119816 16870 119822 16902
rect 119886 16902 119887 16934
rect 119886 16870 119892 16902
rect 119750 16462 119751 16494
rect 119685 16461 119751 16462
rect 119685 16390 119751 16391
rect 119685 16358 119686 16390
rect 119544 16086 119550 16118
rect 119549 16054 119550 16086
rect 119614 16086 119620 16118
rect 119680 16326 119686 16358
rect 119750 16358 119751 16390
rect 119750 16326 119756 16358
rect 119614 16054 119615 16086
rect 119549 16053 119615 16054
rect 119680 15574 119756 16326
rect 119816 16254 119892 16870
rect 119816 16190 119822 16254
rect 119886 16190 119892 16254
rect 119816 16184 119892 16190
rect 119680 15510 119686 15574
rect 119750 15510 119756 15574
rect 119680 15504 119756 15510
rect 119685 1838 119751 1839
rect 119685 1806 119686 1838
rect 119680 1774 119686 1806
rect 119750 1806 119751 1838
rect 121453 1838 121519 1839
rect 121453 1806 121454 1838
rect 119750 1774 119756 1806
rect 119680 1294 119756 1774
rect 119680 1230 119686 1294
rect 119750 1230 119756 1294
rect 119680 1224 119756 1230
rect 121448 1774 121454 1806
rect 121518 1806 121519 1838
rect 122949 1838 123015 1839
rect 122949 1806 122950 1838
rect 121518 1774 121524 1806
rect 121448 1294 121524 1774
rect 121448 1230 121454 1294
rect 121518 1230 121524 1294
rect 121448 1224 121524 1230
rect 122944 1774 122950 1806
rect 123014 1806 123015 1838
rect 123014 1774 123020 1806
rect 122944 1294 123020 1774
rect 122944 1230 122950 1294
rect 123014 1230 123020 1294
rect 122944 1224 123020 1230
rect 124304 0 124380 17550
rect 124576 17478 124652 17484
rect 124576 17414 124582 17478
rect 124646 17414 124652 17478
rect 124576 17070 124652 17414
rect 124576 17038 124582 17070
rect 124581 17006 124582 17038
rect 124646 17038 124652 17070
rect 124646 17006 124647 17038
rect 124581 17005 124647 17006
rect 124712 16526 124788 17958
rect 124848 17886 124924 19590
rect 124989 19590 124990 19622
rect 125054 19622 125060 19654
rect 129744 22102 129820 22108
rect 129744 22038 129750 22102
rect 129814 22038 129820 22102
rect 129744 19654 129820 22038
rect 129744 19622 129750 19654
rect 125054 19590 125055 19622
rect 124989 19589 125055 19590
rect 129749 19590 129750 19622
rect 129814 19622 129820 19654
rect 129880 19654 129956 19660
rect 129814 19590 129815 19622
rect 129749 19589 129815 19590
rect 129880 19590 129886 19654
rect 129950 19590 129956 19654
rect 129613 18838 129679 18839
rect 129613 18806 129614 18838
rect 129608 18774 129614 18806
rect 129678 18806 129679 18838
rect 129678 18774 129684 18806
rect 129608 18158 129684 18774
rect 129608 18094 129614 18158
rect 129678 18094 129684 18158
rect 129608 18088 129684 18094
rect 124848 17854 124854 17886
rect 124853 17822 124854 17854
rect 124918 17854 124924 17886
rect 129744 18022 129820 18028
rect 129744 17958 129750 18022
rect 129814 17958 129820 18022
rect 124918 17822 124919 17854
rect 124853 17821 124919 17822
rect 129341 17614 129407 17615
rect 129341 17582 129342 17614
rect 129336 17550 129342 17582
rect 129406 17582 129407 17614
rect 129406 17550 129412 17582
rect 124853 16934 124919 16935
rect 124853 16902 124854 16934
rect 124712 16494 124718 16526
rect 124717 16462 124718 16494
rect 124782 16494 124788 16526
rect 124848 16870 124854 16902
rect 124918 16902 124919 16934
rect 124918 16870 124924 16902
rect 124782 16462 124783 16494
rect 124717 16461 124783 16462
rect 124581 16390 124647 16391
rect 124581 16358 124582 16390
rect 124576 16326 124582 16358
rect 124646 16358 124647 16390
rect 124646 16326 124652 16358
rect 124576 15574 124652 16326
rect 124848 16254 124924 16870
rect 124848 16190 124854 16254
rect 124918 16190 124924 16254
rect 124848 16184 124924 16190
rect 124576 15510 124582 15574
rect 124646 15510 124652 15574
rect 124576 15504 124652 15510
rect 124717 1838 124783 1839
rect 124717 1806 124718 1838
rect 124712 1774 124718 1806
rect 124782 1806 124783 1838
rect 126213 1838 126279 1839
rect 126213 1806 126214 1838
rect 124782 1774 124788 1806
rect 124712 1294 124788 1774
rect 124712 1230 124718 1294
rect 124782 1230 124788 1294
rect 124712 1224 124788 1230
rect 126208 1774 126214 1806
rect 126278 1806 126279 1838
rect 127981 1838 128047 1839
rect 127981 1806 127982 1838
rect 126278 1774 126284 1806
rect 126208 1294 126284 1774
rect 126208 1230 126214 1294
rect 126278 1230 126284 1294
rect 126208 1224 126284 1230
rect 127976 1774 127982 1806
rect 128046 1806 128047 1838
rect 128046 1774 128052 1806
rect 127976 1294 128052 1774
rect 127976 1230 127982 1294
rect 128046 1230 128052 1294
rect 127976 1224 128052 1230
rect 129336 0 129412 17550
rect 129608 17478 129684 17484
rect 129608 17414 129614 17478
rect 129678 17414 129684 17478
rect 129608 17070 129684 17414
rect 129608 17038 129614 17070
rect 129613 17006 129614 17038
rect 129678 17038 129684 17070
rect 129678 17006 129679 17038
rect 129613 17005 129679 17006
rect 129744 16526 129820 17958
rect 129880 17886 129956 19590
rect 130288 18974 130364 23534
rect 130288 18942 130294 18974
rect 130293 18910 130294 18942
rect 130358 18942 130364 18974
rect 134096 23534 134102 23566
rect 134166 23566 134167 23598
rect 139133 23598 139199 23599
rect 139133 23566 139134 23598
rect 134166 23534 134172 23566
rect 134096 18974 134172 23534
rect 139128 23534 139134 23566
rect 139198 23566 139199 23598
rect 145656 23598 145732 23604
rect 139198 23534 139204 23566
rect 134912 22102 134988 22108
rect 134912 22038 134918 22102
rect 134982 22038 134988 22102
rect 130358 18910 130359 18942
rect 130293 18909 130359 18910
rect 134096 18910 134102 18974
rect 134166 18910 134172 18974
rect 134096 18904 134172 18910
rect 134776 19654 134852 19660
rect 134776 19590 134782 19654
rect 134846 19590 134852 19654
rect 134912 19654 134988 22038
rect 134912 19622 134918 19654
rect 134509 18838 134575 18839
rect 134509 18806 134510 18838
rect 134504 18774 134510 18806
rect 134574 18806 134575 18838
rect 134574 18774 134580 18806
rect 134504 18158 134580 18774
rect 134504 18094 134510 18158
rect 134574 18094 134580 18158
rect 134504 18088 134580 18094
rect 129880 17854 129886 17886
rect 129885 17822 129886 17854
rect 129950 17854 129956 17886
rect 134640 18022 134716 18028
rect 134640 17958 134646 18022
rect 134710 17958 134716 18022
rect 129950 17822 129951 17854
rect 129885 17821 129951 17822
rect 134373 17614 134439 17615
rect 134373 17582 134374 17614
rect 134368 17550 134374 17582
rect 134438 17582 134439 17614
rect 134438 17550 134444 17582
rect 129885 16934 129951 16935
rect 129885 16902 129886 16934
rect 129744 16494 129750 16526
rect 129749 16462 129750 16494
rect 129814 16494 129820 16526
rect 129880 16870 129886 16902
rect 129950 16902 129951 16934
rect 129950 16870 129956 16902
rect 129814 16462 129815 16494
rect 129749 16461 129815 16462
rect 129613 16390 129679 16391
rect 129613 16358 129614 16390
rect 129608 16326 129614 16358
rect 129678 16358 129679 16390
rect 129678 16326 129684 16358
rect 129608 15574 129684 16326
rect 129880 16254 129956 16870
rect 129880 16190 129886 16254
rect 129950 16190 129956 16254
rect 129880 16184 129956 16190
rect 129608 15510 129614 15574
rect 129678 15510 129684 15574
rect 129608 15504 129684 15510
rect 129613 1838 129679 1839
rect 129613 1806 129614 1838
rect 129608 1774 129614 1806
rect 129678 1806 129679 1838
rect 131381 1838 131447 1839
rect 131381 1806 131382 1838
rect 129678 1774 129684 1806
rect 129608 1294 129684 1774
rect 129608 1230 129614 1294
rect 129678 1230 129684 1294
rect 129608 1224 129684 1230
rect 131376 1774 131382 1806
rect 131446 1806 131447 1838
rect 133149 1838 133215 1839
rect 133149 1806 133150 1838
rect 131446 1774 131452 1806
rect 131376 1294 131452 1774
rect 131376 1230 131382 1294
rect 131446 1230 131452 1294
rect 131376 1224 131452 1230
rect 133144 1774 133150 1806
rect 133214 1806 133215 1838
rect 133214 1774 133220 1806
rect 133144 1294 133220 1774
rect 133144 1230 133150 1294
rect 133214 1230 133220 1294
rect 133144 1224 133220 1230
rect 134368 0 134444 17550
rect 134640 16526 134716 17958
rect 134776 17886 134852 19590
rect 134917 19590 134918 19622
rect 134982 19622 134988 19654
rect 134982 19590 134983 19622
rect 134917 19589 134983 19590
rect 139128 18974 139204 23534
rect 145656 23534 145662 23598
rect 145726 23534 145732 23598
rect 149469 23598 149535 23599
rect 149469 23566 149470 23598
rect 139944 22102 140020 22108
rect 139944 22038 139950 22102
rect 140014 22038 140020 22102
rect 139128 18910 139134 18974
rect 139198 18910 139204 18974
rect 139128 18904 139204 18910
rect 139808 19654 139884 19660
rect 139808 19590 139814 19654
rect 139878 19590 139884 19654
rect 139944 19654 140020 22038
rect 139944 19622 139950 19654
rect 139541 18838 139607 18839
rect 139541 18806 139542 18838
rect 139536 18774 139542 18806
rect 139606 18806 139607 18838
rect 139606 18774 139612 18806
rect 139536 18158 139612 18774
rect 139536 18094 139542 18158
rect 139606 18094 139612 18158
rect 139536 18088 139612 18094
rect 134776 17854 134782 17886
rect 134781 17822 134782 17854
rect 134846 17854 134852 17886
rect 139672 18022 139748 18028
rect 139672 17958 139678 18022
rect 139742 17958 139748 18022
rect 134846 17822 134847 17854
rect 134781 17821 134847 17822
rect 134776 17614 134852 17620
rect 134776 17550 134782 17614
rect 134846 17550 134852 17614
rect 139269 17614 139335 17615
rect 139269 17582 139270 17614
rect 134776 17206 134852 17550
rect 134776 17174 134782 17206
rect 134781 17142 134782 17174
rect 134846 17174 134852 17206
rect 139264 17550 139270 17582
rect 139334 17582 139335 17614
rect 139334 17550 139340 17582
rect 134846 17142 134847 17174
rect 134781 17141 134847 17142
rect 134917 17070 134983 17071
rect 134917 17038 134918 17070
rect 134912 17006 134918 17038
rect 134982 17038 134983 17070
rect 134982 17006 134988 17038
rect 134640 16494 134646 16526
rect 134645 16462 134646 16494
rect 134710 16494 134716 16526
rect 134776 16934 134852 16940
rect 134776 16870 134782 16934
rect 134846 16870 134852 16934
rect 134710 16462 134711 16494
rect 134645 16461 134711 16462
rect 134645 16390 134711 16391
rect 134645 16358 134646 16390
rect 134640 16326 134646 16358
rect 134710 16358 134711 16390
rect 134710 16326 134716 16358
rect 134640 15574 134716 16326
rect 134776 15982 134852 16870
rect 134912 16254 134988 17006
rect 134912 16190 134918 16254
rect 134982 16190 134988 16254
rect 134912 16184 134988 16190
rect 134776 15950 134782 15982
rect 134781 15918 134782 15950
rect 134846 15950 134852 15982
rect 134846 15918 134847 15950
rect 134781 15917 134847 15918
rect 134640 15510 134646 15574
rect 134710 15510 134716 15574
rect 134640 15504 134716 15510
rect 134645 1838 134711 1839
rect 134645 1806 134646 1838
rect 134640 1774 134646 1806
rect 134710 1806 134711 1838
rect 136413 1838 136479 1839
rect 136413 1806 136414 1838
rect 134710 1774 134716 1806
rect 134640 1294 134716 1774
rect 134640 1230 134646 1294
rect 134710 1230 134716 1294
rect 134640 1224 134716 1230
rect 136408 1774 136414 1806
rect 136478 1806 136479 1838
rect 138181 1838 138247 1839
rect 138181 1806 138182 1838
rect 136478 1774 136484 1806
rect 136408 1294 136484 1774
rect 136408 1230 136414 1294
rect 136478 1230 136484 1294
rect 136408 1224 136484 1230
rect 138176 1774 138182 1806
rect 138246 1806 138247 1838
rect 138246 1774 138252 1806
rect 138176 1294 138252 1774
rect 138176 1230 138182 1294
rect 138246 1230 138252 1294
rect 138176 1224 138252 1230
rect 139264 0 139340 17550
rect 139536 17478 139612 17484
rect 139536 17414 139542 17478
rect 139606 17414 139612 17478
rect 139536 17070 139612 17414
rect 139536 17038 139542 17070
rect 139541 17006 139542 17038
rect 139606 17038 139612 17070
rect 139606 17006 139607 17038
rect 139541 17005 139607 17006
rect 139672 16526 139748 17958
rect 139808 17886 139884 19590
rect 139949 19590 139950 19622
rect 140014 19622 140020 19654
rect 144704 22102 144916 22108
rect 144704 22038 144846 22102
rect 144910 22038 144916 22102
rect 144704 22032 144916 22038
rect 144704 19654 144780 22032
rect 144704 19622 144710 19654
rect 140014 19590 140015 19622
rect 139949 19589 140015 19590
rect 144709 19590 144710 19622
rect 144774 19622 144780 19654
rect 144840 19654 144916 19660
rect 144774 19590 144775 19622
rect 144709 19589 144775 19590
rect 144840 19590 144846 19654
rect 144910 19590 144916 19654
rect 144573 18838 144639 18839
rect 144573 18806 144574 18838
rect 144568 18774 144574 18806
rect 144638 18806 144639 18838
rect 144638 18774 144644 18806
rect 144568 18158 144644 18774
rect 144568 18094 144574 18158
rect 144638 18094 144644 18158
rect 144568 18088 144644 18094
rect 139808 17854 139814 17886
rect 139813 17822 139814 17854
rect 139878 17854 139884 17886
rect 144704 18022 144780 18028
rect 144704 17958 144710 18022
rect 144774 17958 144780 18022
rect 139878 17822 139879 17854
rect 139813 17821 139879 17822
rect 144301 17614 144367 17615
rect 144301 17582 144302 17614
rect 144296 17550 144302 17582
rect 144366 17582 144367 17614
rect 144366 17550 144372 17582
rect 139813 16934 139879 16935
rect 139813 16902 139814 16934
rect 139672 16494 139678 16526
rect 139677 16462 139678 16494
rect 139742 16494 139748 16526
rect 139808 16870 139814 16902
rect 139878 16902 139879 16934
rect 139878 16870 139884 16902
rect 139742 16462 139743 16494
rect 139677 16461 139743 16462
rect 139541 16390 139607 16391
rect 139541 16358 139542 16390
rect 139536 16326 139542 16358
rect 139606 16358 139607 16390
rect 139606 16326 139612 16358
rect 139536 15574 139612 16326
rect 139808 16254 139884 16870
rect 139808 16190 139814 16254
rect 139878 16190 139884 16254
rect 139808 16184 139884 16190
rect 139536 15510 139542 15574
rect 139606 15510 139612 15574
rect 139536 15504 139612 15510
rect 139677 1838 139743 1839
rect 139677 1806 139678 1838
rect 139672 1774 139678 1806
rect 139742 1806 139743 1838
rect 141445 1838 141511 1839
rect 141445 1806 141446 1838
rect 139742 1774 139748 1806
rect 139672 1294 139748 1774
rect 139672 1230 139678 1294
rect 139742 1230 139748 1294
rect 139672 1224 139748 1230
rect 141440 1774 141446 1806
rect 141510 1806 141511 1838
rect 143213 1838 143279 1839
rect 143213 1806 143214 1838
rect 141510 1774 141516 1806
rect 141440 1294 141516 1774
rect 141440 1230 141446 1294
rect 141510 1230 141516 1294
rect 141440 1224 141516 1230
rect 143208 1774 143214 1806
rect 143278 1806 143279 1838
rect 143278 1774 143284 1806
rect 143208 1294 143284 1774
rect 143208 1230 143214 1294
rect 143278 1230 143284 1294
rect 143208 1224 143284 1230
rect 144296 0 144372 17550
rect 144568 17478 144644 17484
rect 144568 17414 144574 17478
rect 144638 17414 144644 17478
rect 144568 17070 144644 17414
rect 144568 17038 144574 17070
rect 144573 17006 144574 17038
rect 144638 17038 144644 17070
rect 144638 17006 144639 17038
rect 144573 17005 144639 17006
rect 144704 16526 144780 17958
rect 144840 17886 144916 19590
rect 145656 18974 145732 23534
rect 145656 18942 145662 18974
rect 145661 18910 145662 18942
rect 145726 18942 145732 18974
rect 149464 23534 149470 23566
rect 149534 23566 149535 23598
rect 155176 23598 155252 23604
rect 149534 23534 149540 23566
rect 149464 18974 149540 23534
rect 155176 23534 155182 23598
rect 155246 23534 155252 23598
rect 149736 22102 149812 22108
rect 149736 22038 149742 22102
rect 149806 22038 149812 22102
rect 149736 19654 149812 22038
rect 154904 22102 154980 22108
rect 154904 22038 154910 22102
rect 154974 22038 154980 22102
rect 149736 19622 149742 19654
rect 149741 19590 149742 19622
rect 149806 19622 149812 19654
rect 149872 19654 149948 19660
rect 149806 19590 149807 19622
rect 149741 19589 149807 19590
rect 149872 19590 149878 19654
rect 149942 19590 149948 19654
rect 145726 18910 145727 18942
rect 145661 18909 145727 18910
rect 149464 18910 149470 18974
rect 149534 18910 149540 18974
rect 149464 18904 149540 18910
rect 149605 18838 149671 18839
rect 149605 18806 149606 18838
rect 149600 18774 149606 18806
rect 149670 18806 149671 18838
rect 149670 18774 149676 18806
rect 149600 18158 149676 18774
rect 149600 18094 149606 18158
rect 149670 18094 149676 18158
rect 149600 18088 149676 18094
rect 144840 17854 144846 17886
rect 144845 17822 144846 17854
rect 144910 17854 144916 17886
rect 149736 18022 149812 18028
rect 149736 17958 149742 18022
rect 149806 17958 149812 18022
rect 144910 17822 144911 17854
rect 144845 17821 144911 17822
rect 149061 17614 149127 17615
rect 149061 17582 149062 17614
rect 149056 17550 149062 17582
rect 149126 17582 149127 17614
rect 149126 17550 149132 17582
rect 144845 16934 144911 16935
rect 144845 16902 144846 16934
rect 144704 16494 144710 16526
rect 144709 16462 144710 16494
rect 144774 16494 144780 16526
rect 144840 16870 144846 16902
rect 144910 16902 144911 16934
rect 144910 16870 144916 16902
rect 144774 16462 144775 16494
rect 144709 16461 144775 16462
rect 144573 16390 144639 16391
rect 144573 16358 144574 16390
rect 144568 16326 144574 16358
rect 144638 16358 144639 16390
rect 144638 16326 144644 16358
rect 144568 15574 144644 16326
rect 144840 16254 144916 16870
rect 144840 16190 144846 16254
rect 144910 16190 144916 16254
rect 144840 16184 144916 16190
rect 144568 15510 144574 15574
rect 144638 15510 144644 15574
rect 144568 15504 144644 15510
rect 144709 1838 144775 1839
rect 144709 1806 144710 1838
rect 144704 1774 144710 1806
rect 144774 1806 144775 1838
rect 146477 1838 146543 1839
rect 146477 1806 146478 1838
rect 144774 1774 144780 1806
rect 144704 1294 144780 1774
rect 144704 1230 144710 1294
rect 144774 1230 144780 1294
rect 144704 1224 144780 1230
rect 146472 1774 146478 1806
rect 146542 1806 146543 1838
rect 148109 1838 148175 1839
rect 148109 1806 148110 1838
rect 146542 1774 146548 1806
rect 146472 1294 146548 1774
rect 146472 1230 146478 1294
rect 146542 1230 146548 1294
rect 146472 1224 146548 1230
rect 148104 1774 148110 1806
rect 148174 1806 148175 1838
rect 148174 1774 148180 1806
rect 148104 1294 148180 1774
rect 148104 1230 148110 1294
rect 148174 1230 148180 1294
rect 148104 1224 148180 1230
rect 149056 0 149132 17550
rect 149600 17478 149676 17484
rect 149600 17414 149606 17478
rect 149670 17414 149676 17478
rect 149600 17070 149676 17414
rect 149600 17038 149606 17070
rect 149605 17006 149606 17038
rect 149670 17038 149676 17070
rect 149670 17006 149671 17038
rect 149605 17005 149671 17006
rect 149469 16934 149535 16935
rect 149469 16902 149470 16934
rect 149464 16870 149470 16902
rect 149534 16902 149535 16934
rect 149534 16870 149540 16902
rect 149464 16254 149540 16870
rect 149736 16526 149812 17958
rect 149872 17886 149948 19590
rect 154768 19654 154844 19660
rect 154768 19590 154774 19654
rect 154838 19590 154844 19654
rect 154904 19654 154980 22038
rect 154904 19622 154910 19654
rect 154637 18838 154703 18839
rect 154637 18806 154638 18838
rect 154632 18774 154638 18806
rect 154702 18806 154703 18838
rect 154702 18774 154708 18806
rect 154632 18158 154708 18774
rect 154632 18094 154638 18158
rect 154702 18094 154708 18158
rect 154632 18088 154708 18094
rect 149872 17854 149878 17886
rect 149877 17822 149878 17854
rect 149942 17854 149948 17886
rect 154632 18022 154708 18028
rect 154632 17958 154638 18022
rect 154702 17958 154708 18022
rect 149942 17822 149943 17854
rect 149877 17821 149943 17822
rect 154229 17614 154295 17615
rect 154229 17582 154230 17614
rect 149736 16494 149742 16526
rect 149741 16462 149742 16494
rect 149806 16494 149812 16526
rect 154224 17550 154230 17582
rect 154294 17582 154295 17614
rect 154294 17550 154300 17582
rect 149806 16462 149807 16494
rect 149741 16461 149807 16462
rect 149605 16390 149671 16391
rect 149605 16358 149606 16390
rect 149464 16190 149470 16254
rect 149534 16190 149540 16254
rect 149464 16184 149540 16190
rect 149600 16326 149606 16358
rect 149670 16358 149671 16390
rect 149670 16326 149676 16358
rect 149600 15574 149676 16326
rect 149600 15510 149606 15574
rect 149670 15510 149676 15574
rect 149600 15504 149676 15510
rect 150013 1838 150079 1839
rect 150013 1806 150014 1838
rect 150008 1774 150014 1806
rect 150078 1806 150079 1838
rect 151645 1838 151711 1839
rect 151645 1806 151646 1838
rect 150078 1774 150084 1806
rect 150008 1294 150084 1774
rect 150008 1230 150014 1294
rect 150078 1230 150084 1294
rect 150008 1224 150084 1230
rect 151640 1774 151646 1806
rect 151710 1806 151711 1838
rect 153141 1838 153207 1839
rect 153141 1806 153142 1838
rect 151710 1774 151716 1806
rect 151640 1294 151716 1774
rect 151640 1230 151646 1294
rect 151710 1230 151716 1294
rect 151640 1224 151716 1230
rect 153136 1774 153142 1806
rect 153206 1806 153207 1838
rect 153206 1774 153212 1806
rect 153136 1294 153212 1774
rect 153136 1230 153142 1294
rect 153206 1230 153212 1294
rect 153136 1224 153212 1230
rect 154224 0 154300 17550
rect 154632 16526 154708 17958
rect 154768 17886 154844 19590
rect 154909 19590 154910 19622
rect 154974 19622 154980 19654
rect 154974 19590 154975 19622
rect 154909 19589 154975 19590
rect 155176 18974 155252 23534
rect 160208 23598 160284 23604
rect 160208 23534 160214 23598
rect 160278 23534 160284 23598
rect 164157 23598 164223 23599
rect 164157 23566 164158 23598
rect 159936 22102 160012 22108
rect 159936 22038 159942 22102
rect 160006 22038 160012 22102
rect 155176 18942 155182 18974
rect 155181 18910 155182 18942
rect 155246 18942 155252 18974
rect 159800 19654 159876 19660
rect 159800 19590 159806 19654
rect 159870 19590 159876 19654
rect 159936 19654 160012 22038
rect 159936 19622 159942 19654
rect 155246 18910 155247 18942
rect 155181 18909 155247 18910
rect 159533 18838 159599 18839
rect 159533 18806 159534 18838
rect 159528 18774 159534 18806
rect 159598 18806 159599 18838
rect 159598 18774 159604 18806
rect 159528 18158 159604 18774
rect 159528 18094 159534 18158
rect 159598 18094 159604 18158
rect 159528 18088 159604 18094
rect 154768 17854 154774 17886
rect 154773 17822 154774 17854
rect 154838 17854 154844 17886
rect 159664 18022 159740 18028
rect 159664 17958 159670 18022
rect 159734 17958 159740 18022
rect 154838 17822 154839 17854
rect 154773 17821 154839 17822
rect 154768 17614 154844 17620
rect 154768 17550 154774 17614
rect 154838 17550 154844 17614
rect 159261 17614 159327 17615
rect 159261 17582 159262 17614
rect 154768 17070 154844 17550
rect 154768 17038 154774 17070
rect 154773 17006 154774 17038
rect 154838 17038 154844 17070
rect 159256 17550 159262 17582
rect 159326 17582 159327 17614
rect 159326 17550 159332 17582
rect 154838 17006 154839 17038
rect 154773 17005 154839 17006
rect 154773 16934 154839 16935
rect 154773 16902 154774 16934
rect 154632 16494 154638 16526
rect 154637 16462 154638 16494
rect 154702 16494 154708 16526
rect 154768 16870 154774 16902
rect 154838 16902 154839 16934
rect 154838 16870 154844 16902
rect 154702 16462 154703 16494
rect 154637 16461 154703 16462
rect 154501 16390 154567 16391
rect 154501 16358 154502 16390
rect 154496 16326 154502 16358
rect 154566 16358 154567 16390
rect 154566 16326 154572 16358
rect 154496 15574 154572 16326
rect 154768 16254 154844 16870
rect 154768 16190 154774 16254
rect 154838 16190 154844 16254
rect 154768 16184 154844 16190
rect 154496 15510 154502 15574
rect 154566 15510 154572 15574
rect 154496 15504 154572 15510
rect 154909 1838 154975 1839
rect 154909 1806 154910 1838
rect 154904 1774 154910 1806
rect 154974 1806 154975 1838
rect 156677 1838 156743 1839
rect 156677 1806 156678 1838
rect 154974 1774 154980 1806
rect 154904 1294 154980 1774
rect 154904 1230 154910 1294
rect 154974 1230 154980 1294
rect 154904 1224 154980 1230
rect 156672 1774 156678 1806
rect 156742 1806 156743 1838
rect 158173 1838 158239 1839
rect 158173 1806 158174 1838
rect 156742 1774 156748 1806
rect 156672 1294 156748 1774
rect 156672 1230 156678 1294
rect 156742 1230 156748 1294
rect 156672 1224 156748 1230
rect 158168 1774 158174 1806
rect 158238 1806 158239 1838
rect 158238 1774 158244 1806
rect 158168 1294 158244 1774
rect 158168 1230 158174 1294
rect 158238 1230 158244 1294
rect 158168 1224 158244 1230
rect 159256 0 159332 17550
rect 159528 17478 159604 17484
rect 159528 17414 159534 17478
rect 159598 17414 159604 17478
rect 159528 17070 159604 17414
rect 159528 17038 159534 17070
rect 159533 17006 159534 17038
rect 159598 17038 159604 17070
rect 159598 17006 159599 17038
rect 159533 17005 159599 17006
rect 159533 16934 159599 16935
rect 159533 16902 159534 16934
rect 159528 16870 159534 16902
rect 159598 16902 159599 16934
rect 159598 16870 159604 16902
rect 159397 16390 159463 16391
rect 159397 16358 159398 16390
rect 159392 16326 159398 16358
rect 159462 16358 159463 16390
rect 159462 16326 159468 16358
rect 159392 15574 159468 16326
rect 159528 16254 159604 16870
rect 159664 16526 159740 17958
rect 159800 17886 159876 19590
rect 159941 19590 159942 19622
rect 160006 19622 160012 19654
rect 160006 19590 160007 19622
rect 159941 19589 160007 19590
rect 160208 18974 160284 23534
rect 160208 18942 160214 18974
rect 160213 18910 160214 18942
rect 160278 18942 160284 18974
rect 164152 23534 164158 23566
rect 164222 23566 164223 23598
rect 170136 23598 170212 23604
rect 164222 23534 164228 23566
rect 164152 18974 164228 23534
rect 170136 23534 170142 23598
rect 170206 23534 170212 23598
rect 174493 23598 174559 23599
rect 174493 23566 174494 23598
rect 164832 22102 164908 22108
rect 164832 22038 164838 22102
rect 164902 22038 164908 22102
rect 160278 18910 160279 18942
rect 160213 18909 160279 18910
rect 164152 18910 164158 18974
rect 164222 18910 164228 18974
rect 164152 18904 164228 18910
rect 164696 19654 164772 19660
rect 164696 19590 164702 19654
rect 164766 19590 164772 19654
rect 164832 19654 164908 22038
rect 169864 22102 169940 22108
rect 169864 22038 169870 22102
rect 169934 22038 169940 22102
rect 164832 19622 164838 19654
rect 164565 18838 164631 18839
rect 164565 18806 164566 18838
rect 164560 18774 164566 18806
rect 164630 18806 164631 18838
rect 164630 18774 164636 18806
rect 164560 18158 164636 18774
rect 164560 18094 164566 18158
rect 164630 18094 164636 18158
rect 164560 18088 164636 18094
rect 159800 17854 159806 17886
rect 159805 17822 159806 17854
rect 159870 17854 159876 17886
rect 164560 18022 164636 18028
rect 164560 17958 164566 18022
rect 164630 17958 164636 18022
rect 159870 17822 159871 17854
rect 159805 17821 159871 17822
rect 164293 17614 164359 17615
rect 164293 17582 164294 17614
rect 159664 16494 159670 16526
rect 159669 16462 159670 16494
rect 159734 16494 159740 16526
rect 164288 17550 164294 17582
rect 164358 17582 164359 17614
rect 164358 17550 164364 17582
rect 159734 16462 159735 16494
rect 159669 16461 159735 16462
rect 159528 16190 159534 16254
rect 159598 16190 159604 16254
rect 159528 16184 159604 16190
rect 159392 15510 159398 15574
rect 159462 15510 159468 15574
rect 159392 15504 159468 15510
rect 159941 1838 160007 1839
rect 159941 1806 159942 1838
rect 159936 1774 159942 1806
rect 160006 1806 160007 1838
rect 161709 1838 161775 1839
rect 161709 1806 161710 1838
rect 160006 1774 160012 1806
rect 159936 1294 160012 1774
rect 159936 1230 159942 1294
rect 160006 1230 160012 1294
rect 159936 1224 160012 1230
rect 161704 1774 161710 1806
rect 161774 1806 161775 1838
rect 163205 1838 163271 1839
rect 163205 1806 163206 1838
rect 161774 1774 161780 1806
rect 161704 1294 161780 1774
rect 161704 1230 161710 1294
rect 161774 1230 161780 1294
rect 161704 1224 161780 1230
rect 163200 1774 163206 1806
rect 163270 1806 163271 1838
rect 163270 1774 163276 1806
rect 163200 1294 163276 1774
rect 163200 1230 163206 1294
rect 163270 1230 163276 1294
rect 163200 1224 163276 1230
rect 164288 0 164364 17550
rect 164560 16526 164636 17958
rect 164696 17886 164772 19590
rect 164837 19590 164838 19622
rect 164902 19622 164908 19654
rect 169728 19654 169804 19660
rect 164902 19590 164903 19622
rect 164837 19589 164903 19590
rect 169728 19590 169734 19654
rect 169798 19590 169804 19654
rect 169864 19654 169940 22038
rect 169864 19622 169870 19654
rect 169597 18838 169663 18839
rect 169597 18806 169598 18838
rect 169592 18774 169598 18806
rect 169662 18806 169663 18838
rect 169662 18774 169668 18806
rect 169592 18158 169668 18774
rect 169592 18094 169598 18158
rect 169662 18094 169668 18158
rect 169592 18088 169668 18094
rect 164696 17854 164702 17886
rect 164701 17822 164702 17854
rect 164766 17854 164772 17886
rect 169592 18022 169668 18028
rect 169592 17958 169598 18022
rect 169662 17958 169668 18022
rect 164766 17822 164767 17854
rect 164701 17821 164767 17822
rect 164696 17614 164772 17620
rect 164696 17550 164702 17614
rect 164766 17550 164772 17614
rect 169189 17614 169255 17615
rect 169189 17582 169190 17614
rect 164696 17070 164772 17550
rect 164696 17038 164702 17070
rect 164701 17006 164702 17038
rect 164766 17038 164772 17070
rect 169184 17550 169190 17582
rect 169254 17582 169255 17614
rect 169254 17550 169260 17582
rect 164766 17006 164767 17038
rect 164701 17005 164767 17006
rect 164701 16934 164767 16935
rect 164701 16902 164702 16934
rect 164560 16494 164566 16526
rect 164565 16462 164566 16494
rect 164630 16494 164636 16526
rect 164696 16870 164702 16902
rect 164766 16902 164767 16934
rect 164766 16870 164772 16902
rect 164630 16462 164631 16494
rect 164565 16461 164631 16462
rect 164565 16390 164631 16391
rect 164565 16358 164566 16390
rect 164560 16326 164566 16358
rect 164630 16358 164631 16390
rect 164630 16326 164636 16358
rect 164560 15574 164636 16326
rect 164696 16254 164772 16870
rect 164696 16190 164702 16254
rect 164766 16190 164772 16254
rect 164696 16184 164772 16190
rect 164560 15510 164566 15574
rect 164630 15510 164636 15574
rect 164560 15504 164636 15510
rect 164973 1838 165039 1839
rect 164973 1806 164974 1838
rect 164968 1774 164974 1806
rect 165038 1806 165039 1838
rect 166605 1838 166671 1839
rect 166605 1806 166606 1838
rect 165038 1774 165044 1806
rect 164968 1294 165044 1774
rect 164968 1230 164974 1294
rect 165038 1230 165044 1294
rect 164968 1224 165044 1230
rect 166600 1774 166606 1806
rect 166670 1806 166671 1838
rect 168373 1838 168439 1839
rect 168373 1806 168374 1838
rect 166670 1774 166676 1806
rect 166600 1294 166676 1774
rect 166600 1230 166606 1294
rect 166670 1230 166676 1294
rect 166600 1224 166676 1230
rect 168368 1774 168374 1806
rect 168438 1806 168439 1838
rect 168438 1774 168444 1806
rect 168368 1294 168444 1774
rect 168368 1230 168374 1294
rect 168438 1230 168444 1294
rect 168368 1224 168444 1230
rect 169184 0 169260 17550
rect 169461 16934 169527 16935
rect 169461 16902 169462 16934
rect 169456 16870 169462 16902
rect 169526 16902 169527 16934
rect 169526 16870 169532 16902
rect 169456 16254 169532 16870
rect 169592 16526 169668 17958
rect 169728 17886 169804 19590
rect 169869 19590 169870 19622
rect 169934 19622 169940 19654
rect 169934 19590 169935 19622
rect 169869 19589 169935 19590
rect 170136 18974 170212 23534
rect 170136 18942 170142 18974
rect 170141 18910 170142 18942
rect 170206 18942 170212 18974
rect 174488 23534 174494 23566
rect 174558 23566 174559 23598
rect 180200 23598 180276 23604
rect 174558 23534 174564 23566
rect 174488 18974 174564 23534
rect 180200 23534 180206 23598
rect 180270 23534 180276 23598
rect 184421 23598 184487 23599
rect 184421 23566 184422 23598
rect 174896 22102 174972 22108
rect 174896 22038 174902 22102
rect 174966 22038 174972 22102
rect 170206 18910 170207 18942
rect 170141 18909 170207 18910
rect 174488 18910 174494 18974
rect 174558 18910 174564 18974
rect 174488 18904 174564 18910
rect 174760 19654 174836 19660
rect 174760 19590 174766 19654
rect 174830 19590 174836 19654
rect 174896 19654 174972 22038
rect 174896 19622 174902 19654
rect 174629 18838 174695 18839
rect 174629 18806 174630 18838
rect 174624 18774 174630 18806
rect 174694 18806 174695 18838
rect 174694 18774 174700 18806
rect 174624 18158 174700 18774
rect 174624 18094 174630 18158
rect 174694 18094 174700 18158
rect 174624 18088 174700 18094
rect 169728 17854 169734 17886
rect 169733 17822 169734 17854
rect 169798 17854 169804 17886
rect 174624 18022 174700 18028
rect 174624 17958 174630 18022
rect 174694 17958 174700 18022
rect 169798 17822 169799 17854
rect 169733 17821 169799 17822
rect 169728 17614 169804 17620
rect 169728 17550 169734 17614
rect 169798 17550 169804 17614
rect 174221 17614 174287 17615
rect 174221 17582 174222 17614
rect 169728 17070 169804 17550
rect 169728 17038 169734 17070
rect 169733 17006 169734 17038
rect 169798 17038 169804 17070
rect 174216 17550 174222 17582
rect 174286 17582 174287 17614
rect 174286 17550 174292 17582
rect 169798 17006 169799 17038
rect 169733 17005 169799 17006
rect 169592 16494 169598 16526
rect 169597 16462 169598 16494
rect 169662 16494 169668 16526
rect 169662 16462 169663 16494
rect 169597 16461 169663 16462
rect 169597 16390 169663 16391
rect 169597 16358 169598 16390
rect 169456 16190 169462 16254
rect 169526 16190 169532 16254
rect 169456 16184 169532 16190
rect 169592 16326 169598 16358
rect 169662 16358 169663 16390
rect 169662 16326 169668 16358
rect 169592 15574 169668 16326
rect 169592 15510 169598 15574
rect 169662 15510 169668 15574
rect 169592 15504 169668 15510
rect 170141 1838 170207 1839
rect 170141 1806 170142 1838
rect 170136 1774 170142 1806
rect 170206 1806 170207 1838
rect 171637 1838 171703 1839
rect 171637 1806 171638 1838
rect 170206 1774 170212 1806
rect 170136 1294 170212 1774
rect 170136 1230 170142 1294
rect 170206 1230 170212 1294
rect 170136 1224 170212 1230
rect 171632 1774 171638 1806
rect 171702 1806 171703 1838
rect 173405 1838 173471 1839
rect 173405 1806 173406 1838
rect 171702 1774 171708 1806
rect 171632 1294 171708 1774
rect 171632 1230 171638 1294
rect 171702 1230 171708 1294
rect 171632 1224 171708 1230
rect 173400 1774 173406 1806
rect 173470 1806 173471 1838
rect 173470 1774 173476 1806
rect 173400 1294 173476 1774
rect 173400 1230 173406 1294
rect 173470 1230 173476 1294
rect 173400 1224 173476 1230
rect 174216 0 174292 17550
rect 174488 17478 174564 17484
rect 174488 17414 174494 17478
rect 174558 17414 174564 17478
rect 174488 17070 174564 17414
rect 174488 17038 174494 17070
rect 174493 17006 174494 17038
rect 174558 17038 174564 17070
rect 174558 17006 174559 17038
rect 174493 17005 174559 17006
rect 174624 16526 174700 17958
rect 174760 17886 174836 19590
rect 174901 19590 174902 19622
rect 174966 19622 174972 19654
rect 179656 22102 179732 22108
rect 179656 22038 179662 22102
rect 179726 22038 179732 22102
rect 179656 19654 179732 22038
rect 179656 19622 179662 19654
rect 174966 19590 174967 19622
rect 174901 19589 174967 19590
rect 179661 19590 179662 19622
rect 179726 19622 179732 19654
rect 179792 19654 179868 19660
rect 179726 19590 179727 19622
rect 179661 19589 179727 19590
rect 179792 19590 179798 19654
rect 179862 19590 179868 19654
rect 179661 18838 179727 18839
rect 179661 18806 179662 18838
rect 179656 18774 179662 18806
rect 179726 18806 179727 18838
rect 179726 18774 179732 18806
rect 179656 18158 179732 18774
rect 179656 18094 179662 18158
rect 179726 18094 179732 18158
rect 179656 18088 179732 18094
rect 174760 17854 174766 17886
rect 174765 17822 174766 17854
rect 174830 17854 174836 17886
rect 179656 18022 179732 18028
rect 179656 17958 179662 18022
rect 179726 17958 179732 18022
rect 174830 17822 174831 17854
rect 174765 17821 174831 17822
rect 179253 17614 179319 17615
rect 179253 17582 179254 17614
rect 179248 17550 179254 17582
rect 179318 17582 179319 17614
rect 179318 17550 179324 17582
rect 174765 16934 174831 16935
rect 174765 16902 174766 16934
rect 174624 16494 174630 16526
rect 174629 16462 174630 16494
rect 174694 16494 174700 16526
rect 174760 16870 174766 16902
rect 174830 16902 174831 16934
rect 174830 16870 174836 16902
rect 174694 16462 174695 16494
rect 174629 16461 174695 16462
rect 174493 16390 174559 16391
rect 174493 16358 174494 16390
rect 174488 16326 174494 16358
rect 174558 16358 174559 16390
rect 174558 16326 174564 16358
rect 174488 15574 174564 16326
rect 174760 16254 174836 16870
rect 174760 16190 174766 16254
rect 174830 16190 174836 16254
rect 174760 16184 174836 16190
rect 174488 15510 174494 15574
rect 174558 15510 174564 15574
rect 174488 15504 174564 15510
rect 175173 1838 175239 1839
rect 175173 1806 175174 1838
rect 175168 1774 175174 1806
rect 175238 1806 175239 1838
rect 176669 1838 176735 1839
rect 176669 1806 176670 1838
rect 175238 1774 175244 1806
rect 175168 1294 175244 1774
rect 175168 1230 175174 1294
rect 175238 1230 175244 1294
rect 175168 1224 175244 1230
rect 176664 1774 176670 1806
rect 176734 1806 176735 1838
rect 178437 1838 178503 1839
rect 178437 1806 178438 1838
rect 176734 1774 176740 1806
rect 176664 1294 176740 1774
rect 176664 1230 176670 1294
rect 176734 1230 176740 1294
rect 176664 1224 176740 1230
rect 178432 1774 178438 1806
rect 178502 1806 178503 1838
rect 178502 1774 178508 1806
rect 178432 1294 178508 1774
rect 178432 1230 178438 1294
rect 178502 1230 178508 1294
rect 178432 1224 178508 1230
rect 179248 0 179324 17550
rect 179520 17478 179596 17484
rect 179520 17414 179526 17478
rect 179590 17414 179596 17478
rect 179520 17070 179596 17414
rect 179520 17038 179526 17070
rect 179525 17006 179526 17038
rect 179590 17038 179596 17070
rect 179590 17006 179591 17038
rect 179525 17005 179591 17006
rect 179656 16526 179732 17958
rect 179792 17886 179868 19590
rect 180200 18974 180276 23534
rect 180200 18942 180206 18974
rect 180205 18910 180206 18942
rect 180270 18942 180276 18974
rect 184416 23534 184422 23566
rect 184486 23566 184487 23598
rect 201144 23598 201220 25166
rect 204000 25166 204006 25198
rect 204070 25198 204071 25230
rect 204070 25166 204076 25198
rect 204000 24958 204076 25166
rect 204000 24894 204006 24958
rect 204070 24894 204076 24958
rect 204000 24888 204076 24894
rect 184486 23534 184492 23566
rect 184416 18974 184492 23534
rect 201144 23534 201150 23598
rect 201214 23534 201220 23598
rect 201144 23528 201220 23534
rect 204136 24822 204212 24828
rect 204136 24758 204142 24822
rect 204206 24758 204212 24822
rect 204005 23326 204071 23327
rect 204005 23294 204006 23326
rect 204000 23262 204006 23294
rect 204070 23294 204071 23326
rect 204070 23262 204076 23294
rect 184688 22102 184764 22108
rect 184688 22038 184694 22102
rect 184758 22038 184764 22102
rect 180270 18910 180271 18942
rect 180205 18909 180271 18910
rect 184416 18910 184422 18974
rect 184486 18910 184492 18974
rect 184416 18904 184492 18910
rect 184552 19654 184628 19660
rect 184552 19590 184558 19654
rect 184622 19590 184628 19654
rect 184688 19654 184764 22038
rect 204000 20742 204076 23262
rect 204136 22102 204212 24758
rect 204136 22070 204142 22102
rect 204141 22038 204142 22070
rect 204206 22070 204212 22102
rect 217464 24142 217812 25710
rect 217464 24078 217470 24142
rect 217534 24078 217812 24142
rect 217464 22374 217812 24078
rect 217464 22310 217470 22374
rect 217534 22310 217812 22374
rect 204206 22038 204207 22070
rect 204141 22037 204207 22038
rect 204000 20678 204006 20742
rect 204070 20678 204076 20742
rect 204000 20672 204076 20678
rect 204136 21966 204212 21972
rect 204136 21902 204142 21966
rect 204206 21902 204212 21966
rect 184688 19622 184694 19654
rect 184421 18838 184487 18839
rect 184421 18806 184422 18838
rect 184416 18774 184422 18806
rect 184486 18806 184487 18838
rect 184486 18774 184492 18806
rect 184416 18158 184492 18774
rect 184416 18094 184422 18158
rect 184486 18094 184492 18158
rect 184416 18088 184492 18094
rect 179792 17854 179798 17886
rect 179797 17822 179798 17854
rect 179862 17854 179868 17886
rect 184416 18022 184492 18028
rect 184416 17958 184422 18022
rect 184486 17958 184492 18022
rect 179862 17822 179863 17854
rect 179797 17821 179863 17822
rect 184285 17614 184351 17615
rect 184285 17582 184286 17614
rect 184280 17550 184286 17582
rect 184350 17582 184351 17614
rect 184350 17550 184356 17582
rect 179797 16934 179863 16935
rect 179797 16902 179798 16934
rect 179656 16494 179662 16526
rect 179661 16462 179662 16494
rect 179726 16494 179732 16526
rect 179792 16870 179798 16902
rect 179862 16902 179863 16934
rect 179862 16870 179868 16902
rect 179726 16462 179727 16494
rect 179661 16461 179727 16462
rect 179525 16390 179591 16391
rect 179525 16358 179526 16390
rect 179520 16326 179526 16358
rect 179590 16358 179591 16390
rect 179590 16326 179596 16358
rect 179520 15574 179596 16326
rect 179792 16254 179868 16870
rect 179792 16190 179798 16254
rect 179862 16190 179868 16254
rect 179792 16184 179868 16190
rect 179520 15510 179526 15574
rect 179590 15510 179596 15574
rect 179520 15504 179596 15510
rect 180205 1838 180271 1839
rect 180205 1806 180206 1838
rect 180200 1774 180206 1806
rect 180270 1806 180271 1838
rect 181701 1838 181767 1839
rect 181701 1806 181702 1838
rect 180270 1774 180276 1806
rect 180200 1294 180276 1774
rect 180200 1230 180206 1294
rect 180270 1230 180276 1294
rect 180200 1224 180276 1230
rect 181696 1774 181702 1806
rect 181766 1806 181767 1838
rect 183469 1838 183535 1839
rect 183469 1806 183470 1838
rect 181766 1774 181772 1806
rect 181696 1294 181772 1774
rect 181696 1230 181702 1294
rect 181766 1230 181772 1294
rect 181696 1224 181772 1230
rect 183464 1774 183470 1806
rect 183534 1806 183535 1838
rect 183534 1774 183540 1806
rect 183464 1294 183540 1774
rect 183464 1230 183470 1294
rect 183534 1230 183540 1294
rect 183464 1224 183540 1230
rect 184280 0 184356 17550
rect 184416 16526 184492 17958
rect 184552 17886 184628 19590
rect 184693 19590 184694 19622
rect 184758 19622 184764 19654
rect 204000 20606 204076 20612
rect 204000 20542 204006 20606
rect 204070 20542 204076 20606
rect 184758 19590 184759 19622
rect 184693 19589 184759 19590
rect 184552 17854 184558 17886
rect 184557 17822 184558 17854
rect 184622 17854 184628 17886
rect 204000 17886 204076 20542
rect 204136 19246 204212 21902
rect 204136 19214 204142 19246
rect 204141 19182 204142 19214
rect 204206 19214 204212 19246
rect 217464 20606 217812 22310
rect 217464 20542 217470 20606
rect 217534 20542 217812 20606
rect 204206 19182 204207 19214
rect 204141 19181 204207 19182
rect 204277 19110 204343 19111
rect 204277 19078 204278 19110
rect 204000 17854 204006 17886
rect 184622 17822 184623 17854
rect 184557 17821 184623 17822
rect 204005 17822 204006 17854
rect 204070 17854 204076 17886
rect 204272 19046 204278 19078
rect 204342 19078 204343 19110
rect 217464 19110 217812 20542
rect 204342 19046 204348 19078
rect 204070 17822 204071 17854
rect 204005 17821 204071 17822
rect 204136 17750 204212 17756
rect 204136 17686 204142 17750
rect 204206 17686 204212 17750
rect 184552 17614 184628 17620
rect 184552 17550 184558 17614
rect 184622 17550 184628 17614
rect 184552 17070 184628 17550
rect 184552 17038 184558 17070
rect 184557 17006 184558 17038
rect 184622 17038 184628 17070
rect 184622 17006 184623 17038
rect 184557 17005 184623 17006
rect 184416 16494 184422 16526
rect 184421 16462 184422 16494
rect 184486 16494 184492 16526
rect 184552 16934 184628 16940
rect 184552 16870 184558 16934
rect 184622 16870 184628 16934
rect 184693 16934 184759 16935
rect 184693 16902 184694 16934
rect 184486 16462 184487 16494
rect 184421 16461 184487 16462
rect 184421 16390 184487 16391
rect 184421 16358 184422 16390
rect 184416 16326 184422 16358
rect 184486 16358 184487 16390
rect 184486 16326 184492 16358
rect 184416 15574 184492 16326
rect 184552 16118 184628 16870
rect 184688 16870 184694 16902
rect 184758 16902 184759 16934
rect 184758 16870 184764 16902
rect 184688 16254 184764 16870
rect 184688 16190 184694 16254
rect 184758 16190 184764 16254
rect 184688 16184 184764 16190
rect 204000 16254 204076 16260
rect 204000 16190 204006 16254
rect 204070 16190 204076 16254
rect 184552 16086 184558 16118
rect 184557 16054 184558 16086
rect 184622 16086 184628 16118
rect 184622 16054 184623 16086
rect 184557 16053 184623 16054
rect 189181 15846 189247 15847
rect 189181 15814 189182 15846
rect 189176 15782 189182 15814
rect 189246 15814 189247 15846
rect 189246 15782 189252 15814
rect 184416 15510 184422 15574
rect 184486 15510 184492 15574
rect 189045 15574 189111 15575
rect 189045 15542 189046 15574
rect 184416 15504 184492 15510
rect 189040 15510 189046 15542
rect 189110 15542 189111 15574
rect 189110 15510 189116 15542
rect 189040 15166 189116 15510
rect 189040 15102 189046 15166
rect 189110 15102 189116 15166
rect 189040 15096 189116 15102
rect 189176 14078 189252 15782
rect 189176 14014 189182 14078
rect 189246 14014 189252 14078
rect 189176 14008 189252 14014
rect 204000 13670 204076 16190
rect 204136 15030 204212 17686
rect 204272 16526 204348 19046
rect 204272 16462 204278 16526
rect 204342 16462 204348 16526
rect 204272 16456 204348 16462
rect 217464 19046 217470 19110
rect 217534 19046 217812 19110
rect 217464 17206 217812 19046
rect 217464 17142 217470 17206
rect 217534 17142 217812 17206
rect 204136 14998 204142 15030
rect 204141 14966 204142 14998
rect 204206 14998 204212 15030
rect 217464 15710 217812 17142
rect 217464 15646 217470 15710
rect 217534 15646 217812 15710
rect 204206 14966 204207 14998
rect 204141 14965 204207 14966
rect 204000 13638 204006 13670
rect 204005 13606 204006 13638
rect 204070 13638 204076 13670
rect 217464 14078 217812 15646
rect 217464 14014 217470 14078
rect 217534 14014 217812 14078
rect 204070 13606 204071 13638
rect 204005 13605 204071 13606
rect 217464 12174 217812 14014
rect 217464 12110 217470 12174
rect 217534 12110 217812 12174
rect 217464 10542 217812 12110
rect 217464 10478 217470 10542
rect 217534 10478 217812 10542
rect 217464 8910 217812 10478
rect 217464 8846 217470 8910
rect 217534 8846 217812 8910
rect 217464 7278 217812 8846
rect 217464 7214 217470 7278
rect 217534 7214 217812 7278
rect 217464 5646 217812 7214
rect 217464 5582 217470 5646
rect 217534 5582 217812 5646
rect 217464 4014 217812 5582
rect 217464 3950 217470 4014
rect 217534 3950 217812 4014
rect 217464 2110 217812 3950
rect 217464 2046 217470 2110
rect 217534 2046 217812 2110
rect 185101 1838 185167 1839
rect 185101 1806 185102 1838
rect 185096 1774 185102 1806
rect 185166 1806 185167 1838
rect 186869 1838 186935 1839
rect 186869 1806 186870 1838
rect 185166 1774 185172 1806
rect 185096 1294 185172 1774
rect 185096 1230 185102 1294
rect 185166 1230 185172 1294
rect 185096 1224 185172 1230
rect 186864 1774 186870 1806
rect 186934 1806 186935 1838
rect 188637 1838 188703 1839
rect 188637 1806 188638 1838
rect 186934 1774 186940 1806
rect 186864 1294 186940 1774
rect 186864 1230 186870 1294
rect 186934 1230 186940 1294
rect 186864 1224 186940 1230
rect 188632 1774 188638 1806
rect 188702 1806 188703 1838
rect 190133 1838 190199 1839
rect 190133 1806 190134 1838
rect 188702 1774 188708 1806
rect 188632 1294 188708 1774
rect 188632 1230 188638 1294
rect 188702 1230 188708 1294
rect 188632 1224 188708 1230
rect 190128 1774 190134 1806
rect 190198 1806 190199 1838
rect 191901 1838 191967 1839
rect 191901 1806 191902 1838
rect 190198 1774 190204 1806
rect 190128 1294 190204 1774
rect 190128 1230 190134 1294
rect 190198 1230 190204 1294
rect 190128 1224 190204 1230
rect 191896 1774 191902 1806
rect 191966 1806 191967 1838
rect 193669 1838 193735 1839
rect 193669 1806 193670 1838
rect 191966 1774 191972 1806
rect 191896 1294 191972 1774
rect 191896 1230 191902 1294
rect 191966 1230 191972 1294
rect 191896 1224 191972 1230
rect 193664 1774 193670 1806
rect 193734 1806 193735 1838
rect 195165 1838 195231 1839
rect 195165 1806 195166 1838
rect 193734 1774 193740 1806
rect 193664 1294 193740 1774
rect 193664 1230 193670 1294
rect 193734 1230 193740 1294
rect 193664 1224 193740 1230
rect 195160 1774 195166 1806
rect 195230 1806 195231 1838
rect 196933 1838 196999 1839
rect 196933 1806 196934 1838
rect 195230 1774 195236 1806
rect 195160 1294 195236 1774
rect 195160 1230 195166 1294
rect 195230 1230 195236 1294
rect 195160 1224 195236 1230
rect 196928 1774 196934 1806
rect 196998 1806 196999 1838
rect 198701 1838 198767 1839
rect 198701 1806 198702 1838
rect 196998 1774 197004 1806
rect 196928 1294 197004 1774
rect 196928 1230 196934 1294
rect 196998 1230 197004 1294
rect 196928 1224 197004 1230
rect 198696 1774 198702 1806
rect 198766 1806 198767 1838
rect 200197 1838 200263 1839
rect 200197 1806 200198 1838
rect 198766 1774 198772 1806
rect 198696 1294 198772 1774
rect 198696 1230 198702 1294
rect 198766 1230 198772 1294
rect 198696 1224 198772 1230
rect 200192 1774 200198 1806
rect 200262 1806 200263 1838
rect 201965 1838 202031 1839
rect 201965 1806 201966 1838
rect 200262 1774 200268 1806
rect 200192 1294 200268 1774
rect 200192 1230 200198 1294
rect 200262 1230 200268 1294
rect 200192 1224 200268 1230
rect 201960 1774 201966 1806
rect 202030 1806 202031 1838
rect 203597 1838 203663 1839
rect 203597 1806 203598 1838
rect 202030 1774 202036 1806
rect 201960 1294 202036 1774
rect 201960 1230 201966 1294
rect 202030 1230 202036 1294
rect 201960 1224 202036 1230
rect 203592 1774 203598 1806
rect 203662 1806 203663 1838
rect 205229 1838 205295 1839
rect 205229 1806 205230 1838
rect 203662 1774 203668 1806
rect 203592 1294 203668 1774
rect 203592 1230 203598 1294
rect 203662 1230 203668 1294
rect 203592 1224 203668 1230
rect 205224 1774 205230 1806
rect 205294 1806 205295 1838
rect 207133 1838 207199 1839
rect 207133 1806 207134 1838
rect 205294 1774 205300 1806
rect 205224 1294 205300 1774
rect 205224 1230 205230 1294
rect 205294 1230 205300 1294
rect 205224 1224 205300 1230
rect 207128 1774 207134 1806
rect 207198 1806 207199 1838
rect 208629 1838 208695 1839
rect 208629 1806 208630 1838
rect 207198 1774 207204 1806
rect 207128 1294 207204 1774
rect 207128 1230 207134 1294
rect 207198 1230 207204 1294
rect 207128 1224 207204 1230
rect 208624 1774 208630 1806
rect 208694 1806 208695 1838
rect 210397 1838 210463 1839
rect 210397 1806 210398 1838
rect 208694 1774 208700 1806
rect 208624 1294 208700 1774
rect 208624 1230 208630 1294
rect 208694 1230 208700 1294
rect 208624 1224 208700 1230
rect 210392 1774 210398 1806
rect 210462 1806 210463 1838
rect 211893 1838 211959 1839
rect 211893 1806 211894 1838
rect 210462 1774 210468 1806
rect 210392 1294 210468 1774
rect 210392 1230 210398 1294
rect 210462 1230 210468 1294
rect 210392 1224 210468 1230
rect 211888 1774 211894 1806
rect 211958 1806 211959 1838
rect 213661 1838 213727 1839
rect 213661 1806 213662 1838
rect 211958 1774 211964 1806
rect 211888 1294 211964 1774
rect 211888 1230 211894 1294
rect 211958 1230 211964 1294
rect 211888 1224 211964 1230
rect 213656 1774 213662 1806
rect 213726 1806 213727 1838
rect 215429 1838 215495 1839
rect 215429 1806 215430 1838
rect 213726 1774 213732 1806
rect 213656 1294 213732 1774
rect 213656 1230 213662 1294
rect 213726 1230 213732 1294
rect 213656 1224 213732 1230
rect 215424 1774 215430 1806
rect 215494 1806 215495 1838
rect 215494 1774 215500 1806
rect 215424 1294 215500 1774
rect 215424 1230 215430 1294
rect 215494 1230 215500 1294
rect 215424 1224 215500 1230
rect 217464 1294 217812 2046
rect 217464 1230 217470 1294
rect 217534 1230 217606 1294
rect 217670 1230 217742 1294
rect 217806 1230 217812 1294
rect 217464 1158 217812 1230
rect 217464 1094 217470 1158
rect 217534 1094 217606 1158
rect 217670 1094 217742 1158
rect 217806 1094 217812 1158
rect 217464 1022 217812 1094
rect 217464 958 217470 1022
rect 217534 958 217606 1022
rect 217670 958 217742 1022
rect 217806 958 217812 1022
rect 217464 952 217812 958
rect 218144 133894 218492 143486
rect 218144 133830 218150 133894
rect 218214 133830 218492 133894
rect 218144 129678 218492 133830
rect 218144 129614 218150 129678
rect 218214 129614 218492 129678
rect 218144 126958 218492 129614
rect 218144 126894 218150 126958
rect 218214 126894 218492 126958
rect 218144 123966 218492 126894
rect 218144 123902 218150 123966
rect 218214 123902 218492 123966
rect 218144 121110 218492 123902
rect 218144 121046 218150 121110
rect 218214 121046 218492 121110
rect 218144 118526 218492 121046
rect 218144 118462 218150 118526
rect 218214 118462 218492 118526
rect 218144 614 218492 118462
rect 218144 550 218150 614
rect 218214 550 218286 614
rect 218350 550 218422 614
rect 218486 550 218492 614
rect 218144 478 218492 550
rect 218144 414 218150 478
rect 218214 414 218286 478
rect 218350 414 218422 478
rect 218486 414 218492 478
rect 218144 342 218492 414
rect 218144 278 218150 342
rect 218214 278 218286 342
rect 218350 278 218422 342
rect 218486 278 218492 342
rect 218144 272 218492 278
use cr_5  cr_5_0
timestamp 1624857261
transform 1 0 15406 0 1 10918
box 61024 65420 64083 68762
use cr_4  cr_4_0
timestamp 1624857261
transform 1 0 15406 0 1 10918
box 3208 -3962 52705 1462
use cr_3  cr_3_0
timestamp 1624857261
transform 1 0 15406 0 1 10918
box 2083 -3939 6102 5492
use data_dff  data_dff_0
timestamp 1624857261
transform 1 0 24582 0 1 2184
box -36 -49 37412 1467
use wmask_dff  wmask_dff_0
timestamp 1624857261
transform 1 0 19910 0 1 2184
box -36 -49 4708 1467
use col_addr_dff  col_addr_dff_1
timestamp 1624857261
transform 1 0 16406 0 1 2184
box -36 -49 1204 1467
use col_addr_dff  col_addr_dff_0
timestamp 1624857261
transform -1 0 201176 0 -1 142008
box -36 -49 1204 1467
use row_addr_dff  row_addr_dff_1
timestamp 1624857261
transform 1 0 14070 0 1 34317
box -36 -49 1204 9951
use row_addr_dff  row_addr_dff_0
timestamp 1624857261
transform -1 0 204680 0 -1 24837
box -36 -49 1204 9951
use control_logic_r  control_logic_r_0
timestamp 1624857261
transform -1 0 216482 0 -1 135355
box -75 -49 11458 18431
use control_logic_rw  control_logic_rw_0
timestamp 1624857261
transform 1 0 2184 0 1 12611
box -75 -49 11650 18431
use bank  bank_0
timestamp 1624857261
transform 1 0 15406 0 1 10918
box 0 0 67334 67312
use contact_13  contact_13_2111
timestamp 1624857261
transform 1 0 2041 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2110
timestamp 1624857261
transform 1 0 2377 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2109
timestamp 1624857261
transform 1 0 2713 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2108
timestamp 1624857261
transform 1 0 3049 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2107
timestamp 1624857261
transform 1 0 3385 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2106
timestamp 1624857261
transform 1 0 3721 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2105
timestamp 1624857261
transform 1 0 4057 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2104
timestamp 1624857261
transform 1 0 4393 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2103
timestamp 1624857261
transform 1 0 4729 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2102
timestamp 1624857261
transform 1 0 5065 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2101
timestamp 1624857261
transform 1 0 5401 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2100
timestamp 1624857261
transform 1 0 5737 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2099
timestamp 1624857261
transform 1 0 6073 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2098
timestamp 1624857261
transform 1 0 6409 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2097
timestamp 1624857261
transform 1 0 6745 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2096
timestamp 1624857261
transform 1 0 7081 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2095
timestamp 1624857261
transform 1 0 7417 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2094
timestamp 1624857261
transform 1 0 7753 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2093
timestamp 1624857261
transform 1 0 8089 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2092
timestamp 1624857261
transform 1 0 8425 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2091
timestamp 1624857261
transform 1 0 8761 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2090
timestamp 1624857261
transform 1 0 9097 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2089
timestamp 1624857261
transform 1 0 9433 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2088
timestamp 1624857261
transform 1 0 9769 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2087
timestamp 1624857261
transform 1 0 10105 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2086
timestamp 1624857261
transform 1 0 10441 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2085
timestamp 1624857261
transform 1 0 10777 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2084
timestamp 1624857261
transform 1 0 11113 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2083
timestamp 1624857261
transform 1 0 11449 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2082
timestamp 1624857261
transform 1 0 11785 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2081
timestamp 1624857261
transform 1 0 12121 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2080
timestamp 1624857261
transform 1 0 12457 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2079
timestamp 1624857261
transform 1 0 12793 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2078
timestamp 1624857261
transform 1 0 13129 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2077
timestamp 1624857261
transform 1 0 13465 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2076
timestamp 1624857261
transform 1 0 13801 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2075
timestamp 1624857261
transform 1 0 14137 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2074
timestamp 1624857261
transform 1 0 14473 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2073
timestamp 1624857261
transform 1 0 14809 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2072
timestamp 1624857261
transform 1 0 15145 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2071
timestamp 1624857261
transform 1 0 15481 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2070
timestamp 1624857261
transform 1 0 15817 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2069
timestamp 1624857261
transform 1 0 16153 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2068
timestamp 1624857261
transform 1 0 16489 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2067
timestamp 1624857261
transform 1 0 16825 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2066
timestamp 1624857261
transform 1 0 17161 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2065
timestamp 1624857261
transform 1 0 17497 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2064
timestamp 1624857261
transform 1 0 17833 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2063
timestamp 1624857261
transform 1 0 18169 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2062
timestamp 1624857261
transform 1 0 18505 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2061
timestamp 1624857261
transform 1 0 18841 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2060
timestamp 1624857261
transform 1 0 19177 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2059
timestamp 1624857261
transform 1 0 19513 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2058
timestamp 1624857261
transform 1 0 19849 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2057
timestamp 1624857261
transform 1 0 20185 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2056
timestamp 1624857261
transform 1 0 20521 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2055
timestamp 1624857261
transform 1 0 20857 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2054
timestamp 1624857261
transform 1 0 21193 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2053
timestamp 1624857261
transform 1 0 21529 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2052
timestamp 1624857261
transform 1 0 21865 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2051
timestamp 1624857261
transform 1 0 22201 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2050
timestamp 1624857261
transform 1 0 22537 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2049
timestamp 1624857261
transform 1 0 22873 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2048
timestamp 1624857261
transform 1 0 23209 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2047
timestamp 1624857261
transform 1 0 23545 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2046
timestamp 1624857261
transform 1 0 23881 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2045
timestamp 1624857261
transform 1 0 24217 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2044
timestamp 1624857261
transform 1 0 24553 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2043
timestamp 1624857261
transform 1 0 24889 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2042
timestamp 1624857261
transform 1 0 25225 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2041
timestamp 1624857261
transform 1 0 25561 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2040
timestamp 1624857261
transform 1 0 25897 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2039
timestamp 1624857261
transform 1 0 26233 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2038
timestamp 1624857261
transform 1 0 26569 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2037
timestamp 1624857261
transform 1 0 26905 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2036
timestamp 1624857261
transform 1 0 27241 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2035
timestamp 1624857261
transform 1 0 27577 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2034
timestamp 1624857261
transform 1 0 27913 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2033
timestamp 1624857261
transform 1 0 28249 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2032
timestamp 1624857261
transform 1 0 28585 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2031
timestamp 1624857261
transform 1 0 28921 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2030
timestamp 1624857261
transform 1 0 29257 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2029
timestamp 1624857261
transform 1 0 29593 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2028
timestamp 1624857261
transform 1 0 29929 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2027
timestamp 1624857261
transform 1 0 30265 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2026
timestamp 1624857261
transform 1 0 30601 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2025
timestamp 1624857261
transform 1 0 30937 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2024
timestamp 1624857261
transform 1 0 31273 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2023
timestamp 1624857261
transform 1 0 31609 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2022
timestamp 1624857261
transform 1 0 31945 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2021
timestamp 1624857261
transform 1 0 32281 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2020
timestamp 1624857261
transform 1 0 32617 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2019
timestamp 1624857261
transform 1 0 32953 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2018
timestamp 1624857261
transform 1 0 33289 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2017
timestamp 1624857261
transform 1 0 33625 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2016
timestamp 1624857261
transform 1 0 33961 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2015
timestamp 1624857261
transform 1 0 34297 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2014
timestamp 1624857261
transform 1 0 34633 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2013
timestamp 1624857261
transform 1 0 34969 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2012
timestamp 1624857261
transform 1 0 35305 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2011
timestamp 1624857261
transform 1 0 35641 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2010
timestamp 1624857261
transform 1 0 35977 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2009
timestamp 1624857261
transform 1 0 36313 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2008
timestamp 1624857261
transform 1 0 36649 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2007
timestamp 1624857261
transform 1 0 36985 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2006
timestamp 1624857261
transform 1 0 37321 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2005
timestamp 1624857261
transform 1 0 37657 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2004
timestamp 1624857261
transform 1 0 37993 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2003
timestamp 1624857261
transform 1 0 38329 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2002
timestamp 1624857261
transform 1 0 38665 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2001
timestamp 1624857261
transform 1 0 39001 0 1 1807
box 0 0 1 1
use contact_13  contact_13_2000
timestamp 1624857261
transform 1 0 39337 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1999
timestamp 1624857261
transform 1 0 39673 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1998
timestamp 1624857261
transform 1 0 40009 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1997
timestamp 1624857261
transform 1 0 40345 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1996
timestamp 1624857261
transform 1 0 40681 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1995
timestamp 1624857261
transform 1 0 41017 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1994
timestamp 1624857261
transform 1 0 41353 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1993
timestamp 1624857261
transform 1 0 41689 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1992
timestamp 1624857261
transform 1 0 42025 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1991
timestamp 1624857261
transform 1 0 42361 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1990
timestamp 1624857261
transform 1 0 42697 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1989
timestamp 1624857261
transform 1 0 43033 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1988
timestamp 1624857261
transform 1 0 43369 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1987
timestamp 1624857261
transform 1 0 43705 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1986
timestamp 1624857261
transform 1 0 44041 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1985
timestamp 1624857261
transform 1 0 44377 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1984
timestamp 1624857261
transform 1 0 44713 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1983
timestamp 1624857261
transform 1 0 45049 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1982
timestamp 1624857261
transform 1 0 45385 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1981
timestamp 1624857261
transform 1 0 45721 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1980
timestamp 1624857261
transform 1 0 46057 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1979
timestamp 1624857261
transform 1 0 46393 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1978
timestamp 1624857261
transform 1 0 46729 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1977
timestamp 1624857261
transform 1 0 47065 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1976
timestamp 1624857261
transform 1 0 47401 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1975
timestamp 1624857261
transform 1 0 47737 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1974
timestamp 1624857261
transform 1 0 48073 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1973
timestamp 1624857261
transform 1 0 48409 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1972
timestamp 1624857261
transform 1 0 48745 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1971
timestamp 1624857261
transform 1 0 49081 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1970
timestamp 1624857261
transform 1 0 49417 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1969
timestamp 1624857261
transform 1 0 49753 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1968
timestamp 1624857261
transform 1 0 50089 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1967
timestamp 1624857261
transform 1 0 50425 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1966
timestamp 1624857261
transform 1 0 50761 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1965
timestamp 1624857261
transform 1 0 51097 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1964
timestamp 1624857261
transform 1 0 51433 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1963
timestamp 1624857261
transform 1 0 51769 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1962
timestamp 1624857261
transform 1 0 52105 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1961
timestamp 1624857261
transform 1 0 52441 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1960
timestamp 1624857261
transform 1 0 52777 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1959
timestamp 1624857261
transform 1 0 53113 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1958
timestamp 1624857261
transform 1 0 53449 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1957
timestamp 1624857261
transform 1 0 53785 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1956
timestamp 1624857261
transform 1 0 54121 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1955
timestamp 1624857261
transform 1 0 54457 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1954
timestamp 1624857261
transform 1 0 54793 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1953
timestamp 1624857261
transform 1 0 55129 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1952
timestamp 1624857261
transform 1 0 55465 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1951
timestamp 1624857261
transform 1 0 55801 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1950
timestamp 1624857261
transform 1 0 56137 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1949
timestamp 1624857261
transform 1 0 56473 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1948
timestamp 1624857261
transform 1 0 56809 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1947
timestamp 1624857261
transform 1 0 57145 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1946
timestamp 1624857261
transform 1 0 57481 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1945
timestamp 1624857261
transform 1 0 57817 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1944
timestamp 1624857261
transform 1 0 58153 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1943
timestamp 1624857261
transform 1 0 58489 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1942
timestamp 1624857261
transform 1 0 58825 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1941
timestamp 1624857261
transform 1 0 59161 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1940
timestamp 1624857261
transform 1 0 59497 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1939
timestamp 1624857261
transform 1 0 59833 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1938
timestamp 1624857261
transform 1 0 60169 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1937
timestamp 1624857261
transform 1 0 60505 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1936
timestamp 1624857261
transform 1 0 60841 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1935
timestamp 1624857261
transform 1 0 61177 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1934
timestamp 1624857261
transform 1 0 61513 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1933
timestamp 1624857261
transform 1 0 61849 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1932
timestamp 1624857261
transform 1 0 62185 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1931
timestamp 1624857261
transform 1 0 62521 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1930
timestamp 1624857261
transform 1 0 62857 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1929
timestamp 1624857261
transform 1 0 63193 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1928
timestamp 1624857261
transform 1 0 63529 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1927
timestamp 1624857261
transform 1 0 63865 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1926
timestamp 1624857261
transform 1 0 64201 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1925
timestamp 1624857261
transform 1 0 64537 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1924
timestamp 1624857261
transform 1 0 64873 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1923
timestamp 1624857261
transform 1 0 65209 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1922
timestamp 1624857261
transform 1 0 65545 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1921
timestamp 1624857261
transform 1 0 65881 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1920
timestamp 1624857261
transform 1 0 66217 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1919
timestamp 1624857261
transform 1 0 66553 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1918
timestamp 1624857261
transform 1 0 66889 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1917
timestamp 1624857261
transform 1 0 67225 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1916
timestamp 1624857261
transform 1 0 67561 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1915
timestamp 1624857261
transform 1 0 67897 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1914
timestamp 1624857261
transform 1 0 68233 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1913
timestamp 1624857261
transform 1 0 68569 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1912
timestamp 1624857261
transform 1 0 68905 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1911
timestamp 1624857261
transform 1 0 69241 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1910
timestamp 1624857261
transform 1 0 69577 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1909
timestamp 1624857261
transform 1 0 69913 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1908
timestamp 1624857261
transform 1 0 70249 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1907
timestamp 1624857261
transform 1 0 70585 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1906
timestamp 1624857261
transform 1 0 70921 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1905
timestamp 1624857261
transform 1 0 71257 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1904
timestamp 1624857261
transform 1 0 71593 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1903
timestamp 1624857261
transform 1 0 71929 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1902
timestamp 1624857261
transform 1 0 72265 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1901
timestamp 1624857261
transform 1 0 72601 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1900
timestamp 1624857261
transform 1 0 72937 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1899
timestamp 1624857261
transform 1 0 73273 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1898
timestamp 1624857261
transform 1 0 73609 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1897
timestamp 1624857261
transform 1 0 73945 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1896
timestamp 1624857261
transform 1 0 74281 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1895
timestamp 1624857261
transform 1 0 74617 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1894
timestamp 1624857261
transform 1 0 74953 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1893
timestamp 1624857261
transform 1 0 75289 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1892
timestamp 1624857261
transform 1 0 75625 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1891
timestamp 1624857261
transform 1 0 75961 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1890
timestamp 1624857261
transform 1 0 76297 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1889
timestamp 1624857261
transform 1 0 76633 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1888
timestamp 1624857261
transform 1 0 76969 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1887
timestamp 1624857261
transform 1 0 77305 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1886
timestamp 1624857261
transform 1 0 77641 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1885
timestamp 1624857261
transform 1 0 77977 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1884
timestamp 1624857261
transform 1 0 78313 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1883
timestamp 1624857261
transform 1 0 78649 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1882
timestamp 1624857261
transform 1 0 78985 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1881
timestamp 1624857261
transform 1 0 79321 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1880
timestamp 1624857261
transform 1 0 79657 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1879
timestamp 1624857261
transform 1 0 79993 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1878
timestamp 1624857261
transform 1 0 80329 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1877
timestamp 1624857261
transform 1 0 80665 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1876
timestamp 1624857261
transform 1 0 81001 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1875
timestamp 1624857261
transform 1 0 81337 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1874
timestamp 1624857261
transform 1 0 81673 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1873
timestamp 1624857261
transform 1 0 82009 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1872
timestamp 1624857261
transform 1 0 82345 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1871
timestamp 1624857261
transform 1 0 82681 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1870
timestamp 1624857261
transform 1 0 83017 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1869
timestamp 1624857261
transform 1 0 83353 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1868
timestamp 1624857261
transform 1 0 83689 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1867
timestamp 1624857261
transform 1 0 84025 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1866
timestamp 1624857261
transform 1 0 84361 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1865
timestamp 1624857261
transform 1 0 84697 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1864
timestamp 1624857261
transform 1 0 85033 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1863
timestamp 1624857261
transform 1 0 85369 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1862
timestamp 1624857261
transform 1 0 85705 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1861
timestamp 1624857261
transform 1 0 86041 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1860
timestamp 1624857261
transform 1 0 86377 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1859
timestamp 1624857261
transform 1 0 86713 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1858
timestamp 1624857261
transform 1 0 87049 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1857
timestamp 1624857261
transform 1 0 87385 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1856
timestamp 1624857261
transform 1 0 87721 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1855
timestamp 1624857261
transform 1 0 88057 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1854
timestamp 1624857261
transform 1 0 88393 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1853
timestamp 1624857261
transform 1 0 88729 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1852
timestamp 1624857261
transform 1 0 89065 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1851
timestamp 1624857261
transform 1 0 89401 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1850
timestamp 1624857261
transform 1 0 89737 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1849
timestamp 1624857261
transform 1 0 90073 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1848
timestamp 1624857261
transform 1 0 90409 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1847
timestamp 1624857261
transform 1 0 90745 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1846
timestamp 1624857261
transform 1 0 91081 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1845
timestamp 1624857261
transform 1 0 91417 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1844
timestamp 1624857261
transform 1 0 91753 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1843
timestamp 1624857261
transform 1 0 92089 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1842
timestamp 1624857261
transform 1 0 92425 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1841
timestamp 1624857261
transform 1 0 92761 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1840
timestamp 1624857261
transform 1 0 93097 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1839
timestamp 1624857261
transform 1 0 93433 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1838
timestamp 1624857261
transform 1 0 93769 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1837
timestamp 1624857261
transform 1 0 94105 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1836
timestamp 1624857261
transform 1 0 94441 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1835
timestamp 1624857261
transform 1 0 94777 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1834
timestamp 1624857261
transform 1 0 95113 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1833
timestamp 1624857261
transform 1 0 95449 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1832
timestamp 1624857261
transform 1 0 95785 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1831
timestamp 1624857261
transform 1 0 96121 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1830
timestamp 1624857261
transform 1 0 96457 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1829
timestamp 1624857261
transform 1 0 96793 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1828
timestamp 1624857261
transform 1 0 97129 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1827
timestamp 1624857261
transform 1 0 97465 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1826
timestamp 1624857261
transform 1 0 97801 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1825
timestamp 1624857261
transform 1 0 98137 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1824
timestamp 1624857261
transform 1 0 98473 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1823
timestamp 1624857261
transform 1 0 98809 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1822
timestamp 1624857261
transform 1 0 99145 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1821
timestamp 1624857261
transform 1 0 99481 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1820
timestamp 1624857261
transform 1 0 99817 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1819
timestamp 1624857261
transform 1 0 100153 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1818
timestamp 1624857261
transform 1 0 100489 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1817
timestamp 1624857261
transform 1 0 100825 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1816
timestamp 1624857261
transform 1 0 101161 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1815
timestamp 1624857261
transform 1 0 101497 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1814
timestamp 1624857261
transform 1 0 101833 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1813
timestamp 1624857261
transform 1 0 102169 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1812
timestamp 1624857261
transform 1 0 102505 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1811
timestamp 1624857261
transform 1 0 102841 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1810
timestamp 1624857261
transform 1 0 103177 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1809
timestamp 1624857261
transform 1 0 103513 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1808
timestamp 1624857261
transform 1 0 103849 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1807
timestamp 1624857261
transform 1 0 104185 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1806
timestamp 1624857261
transform 1 0 104521 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1805
timestamp 1624857261
transform 1 0 104857 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1804
timestamp 1624857261
transform 1 0 105193 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1803
timestamp 1624857261
transform 1 0 105529 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1802
timestamp 1624857261
transform 1 0 105865 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1801
timestamp 1624857261
transform 1 0 106201 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1800
timestamp 1624857261
transform 1 0 106537 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1799
timestamp 1624857261
transform 1 0 106873 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1798
timestamp 1624857261
transform 1 0 107209 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1797
timestamp 1624857261
transform 1 0 107545 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1796
timestamp 1624857261
transform 1 0 107881 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1795
timestamp 1624857261
transform 1 0 108217 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1794
timestamp 1624857261
transform 1 0 108553 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1793
timestamp 1624857261
transform 1 0 108889 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1792
timestamp 1624857261
transform 1 0 109225 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1791
timestamp 1624857261
transform 1 0 109561 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1790
timestamp 1624857261
transform 1 0 109897 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1789
timestamp 1624857261
transform 1 0 110233 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1788
timestamp 1624857261
transform 1 0 110569 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1787
timestamp 1624857261
transform 1 0 110905 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1786
timestamp 1624857261
transform 1 0 111241 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1785
timestamp 1624857261
transform 1 0 111577 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1784
timestamp 1624857261
transform 1 0 111913 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1783
timestamp 1624857261
transform 1 0 112249 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1782
timestamp 1624857261
transform 1 0 112585 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1781
timestamp 1624857261
transform 1 0 112921 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1780
timestamp 1624857261
transform 1 0 113257 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1779
timestamp 1624857261
transform 1 0 113593 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1778
timestamp 1624857261
transform 1 0 113929 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1777
timestamp 1624857261
transform 1 0 114265 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1776
timestamp 1624857261
transform 1 0 114601 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1775
timestamp 1624857261
transform 1 0 114937 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1774
timestamp 1624857261
transform 1 0 115273 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1773
timestamp 1624857261
transform 1 0 115609 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1772
timestamp 1624857261
transform 1 0 115945 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1771
timestamp 1624857261
transform 1 0 116281 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1770
timestamp 1624857261
transform 1 0 116617 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1769
timestamp 1624857261
transform 1 0 116953 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1768
timestamp 1624857261
transform 1 0 117289 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1767
timestamp 1624857261
transform 1 0 117625 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1766
timestamp 1624857261
transform 1 0 117961 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1765
timestamp 1624857261
transform 1 0 118297 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1764
timestamp 1624857261
transform 1 0 118633 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1763
timestamp 1624857261
transform 1 0 118969 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1762
timestamp 1624857261
transform 1 0 119305 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1761
timestamp 1624857261
transform 1 0 119641 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1760
timestamp 1624857261
transform 1 0 119977 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1759
timestamp 1624857261
transform 1 0 120313 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1758
timestamp 1624857261
transform 1 0 120649 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1757
timestamp 1624857261
transform 1 0 120985 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1756
timestamp 1624857261
transform 1 0 121321 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1755
timestamp 1624857261
transform 1 0 121657 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1754
timestamp 1624857261
transform 1 0 121993 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1753
timestamp 1624857261
transform 1 0 122329 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1752
timestamp 1624857261
transform 1 0 122665 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1751
timestamp 1624857261
transform 1 0 123001 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1750
timestamp 1624857261
transform 1 0 123337 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1749
timestamp 1624857261
transform 1 0 123673 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1748
timestamp 1624857261
transform 1 0 124009 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1747
timestamp 1624857261
transform 1 0 124345 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1746
timestamp 1624857261
transform 1 0 124681 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1745
timestamp 1624857261
transform 1 0 125017 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1744
timestamp 1624857261
transform 1 0 125353 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1743
timestamp 1624857261
transform 1 0 125689 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1742
timestamp 1624857261
transform 1 0 126025 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1741
timestamp 1624857261
transform 1 0 126361 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1740
timestamp 1624857261
transform 1 0 126697 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1739
timestamp 1624857261
transform 1 0 127033 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1738
timestamp 1624857261
transform 1 0 127369 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1737
timestamp 1624857261
transform 1 0 127705 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1736
timestamp 1624857261
transform 1 0 128041 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1735
timestamp 1624857261
transform 1 0 128377 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1734
timestamp 1624857261
transform 1 0 128713 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1733
timestamp 1624857261
transform 1 0 129049 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1732
timestamp 1624857261
transform 1 0 129385 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1731
timestamp 1624857261
transform 1 0 129721 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1730
timestamp 1624857261
transform 1 0 130057 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1729
timestamp 1624857261
transform 1 0 130393 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1728
timestamp 1624857261
transform 1 0 130729 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1727
timestamp 1624857261
transform 1 0 131065 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1726
timestamp 1624857261
transform 1 0 131401 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1725
timestamp 1624857261
transform 1 0 131737 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1724
timestamp 1624857261
transform 1 0 132073 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1723
timestamp 1624857261
transform 1 0 132409 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1722
timestamp 1624857261
transform 1 0 132745 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1721
timestamp 1624857261
transform 1 0 133081 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1720
timestamp 1624857261
transform 1 0 133417 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1719
timestamp 1624857261
transform 1 0 133753 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1718
timestamp 1624857261
transform 1 0 134089 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1717
timestamp 1624857261
transform 1 0 134425 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1716
timestamp 1624857261
transform 1 0 134761 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1715
timestamp 1624857261
transform 1 0 135097 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1714
timestamp 1624857261
transform 1 0 135433 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1713
timestamp 1624857261
transform 1 0 135769 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1712
timestamp 1624857261
transform 1 0 136105 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1711
timestamp 1624857261
transform 1 0 136441 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1710
timestamp 1624857261
transform 1 0 136777 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1709
timestamp 1624857261
transform 1 0 137113 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1708
timestamp 1624857261
transform 1 0 137449 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1707
timestamp 1624857261
transform 1 0 137785 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1706
timestamp 1624857261
transform 1 0 138121 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1705
timestamp 1624857261
transform 1 0 138457 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1704
timestamp 1624857261
transform 1 0 138793 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1703
timestamp 1624857261
transform 1 0 139129 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1702
timestamp 1624857261
transform 1 0 139465 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1701
timestamp 1624857261
transform 1 0 139801 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1700
timestamp 1624857261
transform 1 0 140137 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1699
timestamp 1624857261
transform 1 0 140473 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1698
timestamp 1624857261
transform 1 0 140809 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1697
timestamp 1624857261
transform 1 0 141145 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1696
timestamp 1624857261
transform 1 0 141481 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1695
timestamp 1624857261
transform 1 0 141817 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1694
timestamp 1624857261
transform 1 0 142153 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1693
timestamp 1624857261
transform 1 0 142489 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1692
timestamp 1624857261
transform 1 0 142825 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1691
timestamp 1624857261
transform 1 0 143161 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1690
timestamp 1624857261
transform 1 0 143497 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1689
timestamp 1624857261
transform 1 0 143833 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1688
timestamp 1624857261
transform 1 0 144169 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1687
timestamp 1624857261
transform 1 0 144505 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1686
timestamp 1624857261
transform 1 0 144841 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1685
timestamp 1624857261
transform 1 0 145177 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1684
timestamp 1624857261
transform 1 0 145513 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1683
timestamp 1624857261
transform 1 0 145849 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1682
timestamp 1624857261
transform 1 0 146185 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1681
timestamp 1624857261
transform 1 0 146521 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1680
timestamp 1624857261
transform 1 0 146857 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1679
timestamp 1624857261
transform 1 0 147193 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1678
timestamp 1624857261
transform 1 0 147529 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1677
timestamp 1624857261
transform 1 0 147865 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1676
timestamp 1624857261
transform 1 0 148201 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1675
timestamp 1624857261
transform 1 0 148537 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1674
timestamp 1624857261
transform 1 0 148873 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1673
timestamp 1624857261
transform 1 0 149209 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1672
timestamp 1624857261
transform 1 0 149545 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1671
timestamp 1624857261
transform 1 0 149881 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1670
timestamp 1624857261
transform 1 0 150217 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1669
timestamp 1624857261
transform 1 0 150553 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1668
timestamp 1624857261
transform 1 0 150889 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1667
timestamp 1624857261
transform 1 0 151225 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1666
timestamp 1624857261
transform 1 0 151561 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1665
timestamp 1624857261
transform 1 0 151897 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1664
timestamp 1624857261
transform 1 0 152233 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1663
timestamp 1624857261
transform 1 0 152569 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1662
timestamp 1624857261
transform 1 0 152905 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1661
timestamp 1624857261
transform 1 0 153241 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1660
timestamp 1624857261
transform 1 0 153577 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1659
timestamp 1624857261
transform 1 0 153913 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1658
timestamp 1624857261
transform 1 0 154249 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1657
timestamp 1624857261
transform 1 0 154585 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1656
timestamp 1624857261
transform 1 0 154921 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1655
timestamp 1624857261
transform 1 0 155257 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1654
timestamp 1624857261
transform 1 0 155593 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1653
timestamp 1624857261
transform 1 0 155929 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1652
timestamp 1624857261
transform 1 0 156265 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1651
timestamp 1624857261
transform 1 0 156601 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1650
timestamp 1624857261
transform 1 0 156937 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1649
timestamp 1624857261
transform 1 0 157273 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1648
timestamp 1624857261
transform 1 0 157609 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1647
timestamp 1624857261
transform 1 0 157945 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1646
timestamp 1624857261
transform 1 0 158281 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1645
timestamp 1624857261
transform 1 0 158617 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1644
timestamp 1624857261
transform 1 0 158953 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1643
timestamp 1624857261
transform 1 0 159289 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1642
timestamp 1624857261
transform 1 0 159625 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1641
timestamp 1624857261
transform 1 0 159961 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1640
timestamp 1624857261
transform 1 0 160297 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1639
timestamp 1624857261
transform 1 0 160633 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1638
timestamp 1624857261
transform 1 0 160969 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1637
timestamp 1624857261
transform 1 0 161305 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1636
timestamp 1624857261
transform 1 0 161641 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1635
timestamp 1624857261
transform 1 0 161977 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1634
timestamp 1624857261
transform 1 0 162313 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1633
timestamp 1624857261
transform 1 0 162649 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1632
timestamp 1624857261
transform 1 0 162985 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1631
timestamp 1624857261
transform 1 0 163321 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1630
timestamp 1624857261
transform 1 0 163657 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1629
timestamp 1624857261
transform 1 0 163993 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1628
timestamp 1624857261
transform 1 0 164329 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1627
timestamp 1624857261
transform 1 0 164665 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1626
timestamp 1624857261
transform 1 0 165001 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1625
timestamp 1624857261
transform 1 0 165337 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1624
timestamp 1624857261
transform 1 0 165673 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1623
timestamp 1624857261
transform 1 0 166009 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1622
timestamp 1624857261
transform 1 0 166345 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1621
timestamp 1624857261
transform 1 0 166681 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1620
timestamp 1624857261
transform 1 0 167017 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1619
timestamp 1624857261
transform 1 0 167353 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1618
timestamp 1624857261
transform 1 0 167689 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1617
timestamp 1624857261
transform 1 0 168025 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1616
timestamp 1624857261
transform 1 0 168361 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1615
timestamp 1624857261
transform 1 0 168697 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1614
timestamp 1624857261
transform 1 0 169033 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1613
timestamp 1624857261
transform 1 0 169369 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1612
timestamp 1624857261
transform 1 0 169705 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1611
timestamp 1624857261
transform 1 0 170041 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1610
timestamp 1624857261
transform 1 0 170377 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1609
timestamp 1624857261
transform 1 0 170713 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1608
timestamp 1624857261
transform 1 0 171049 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1607
timestamp 1624857261
transform 1 0 171385 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1606
timestamp 1624857261
transform 1 0 171721 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1605
timestamp 1624857261
transform 1 0 172057 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1604
timestamp 1624857261
transform 1 0 172393 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1603
timestamp 1624857261
transform 1 0 172729 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1602
timestamp 1624857261
transform 1 0 173065 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1601
timestamp 1624857261
transform 1 0 173401 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1600
timestamp 1624857261
transform 1 0 173737 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1599
timestamp 1624857261
transform 1 0 174073 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1598
timestamp 1624857261
transform 1 0 174409 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1597
timestamp 1624857261
transform 1 0 174745 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1596
timestamp 1624857261
transform 1 0 175081 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1595
timestamp 1624857261
transform 1 0 175417 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1594
timestamp 1624857261
transform 1 0 175753 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1593
timestamp 1624857261
transform 1 0 176089 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1592
timestamp 1624857261
transform 1 0 176425 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1591
timestamp 1624857261
transform 1 0 176761 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1590
timestamp 1624857261
transform 1 0 177097 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1589
timestamp 1624857261
transform 1 0 177433 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1588
timestamp 1624857261
transform 1 0 177769 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1587
timestamp 1624857261
transform 1 0 178105 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1586
timestamp 1624857261
transform 1 0 178441 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1585
timestamp 1624857261
transform 1 0 178777 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1584
timestamp 1624857261
transform 1 0 179113 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1583
timestamp 1624857261
transform 1 0 179449 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1582
timestamp 1624857261
transform 1 0 179785 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1581
timestamp 1624857261
transform 1 0 180121 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1580
timestamp 1624857261
transform 1 0 180457 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1579
timestamp 1624857261
transform 1 0 180793 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1578
timestamp 1624857261
transform 1 0 181129 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1577
timestamp 1624857261
transform 1 0 181465 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1576
timestamp 1624857261
transform 1 0 181801 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1575
timestamp 1624857261
transform 1 0 182137 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1574
timestamp 1624857261
transform 1 0 182473 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1573
timestamp 1624857261
transform 1 0 182809 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1572
timestamp 1624857261
transform 1 0 183145 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1571
timestamp 1624857261
transform 1 0 183481 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1570
timestamp 1624857261
transform 1 0 183817 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1569
timestamp 1624857261
transform 1 0 184153 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1568
timestamp 1624857261
transform 1 0 184489 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1567
timestamp 1624857261
transform 1 0 184825 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1566
timestamp 1624857261
transform 1 0 185161 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1565
timestamp 1624857261
transform 1 0 185497 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1564
timestamp 1624857261
transform 1 0 185833 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1563
timestamp 1624857261
transform 1 0 186169 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1562
timestamp 1624857261
transform 1 0 186505 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1561
timestamp 1624857261
transform 1 0 186841 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1560
timestamp 1624857261
transform 1 0 187177 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1559
timestamp 1624857261
transform 1 0 187513 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1558
timestamp 1624857261
transform 1 0 187849 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1557
timestamp 1624857261
transform 1 0 188185 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1556
timestamp 1624857261
transform 1 0 188521 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1555
timestamp 1624857261
transform 1 0 188857 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1554
timestamp 1624857261
transform 1 0 189193 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1553
timestamp 1624857261
transform 1 0 189529 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1552
timestamp 1624857261
transform 1 0 189865 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1551
timestamp 1624857261
transform 1 0 190201 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1550
timestamp 1624857261
transform 1 0 190537 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1549
timestamp 1624857261
transform 1 0 190873 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1548
timestamp 1624857261
transform 1 0 191209 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1547
timestamp 1624857261
transform 1 0 191545 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1546
timestamp 1624857261
transform 1 0 191881 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1545
timestamp 1624857261
transform 1 0 192217 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1544
timestamp 1624857261
transform 1 0 192553 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1543
timestamp 1624857261
transform 1 0 192889 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1542
timestamp 1624857261
transform 1 0 193225 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1541
timestamp 1624857261
transform 1 0 193561 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1540
timestamp 1624857261
transform 1 0 193897 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1539
timestamp 1624857261
transform 1 0 194233 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1538
timestamp 1624857261
transform 1 0 194569 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1537
timestamp 1624857261
transform 1 0 194905 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1536
timestamp 1624857261
transform 1 0 195241 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1535
timestamp 1624857261
transform 1 0 195577 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1534
timestamp 1624857261
transform 1 0 195913 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1533
timestamp 1624857261
transform 1 0 196249 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1532
timestamp 1624857261
transform 1 0 196585 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1531
timestamp 1624857261
transform 1 0 196921 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1530
timestamp 1624857261
transform 1 0 197257 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1529
timestamp 1624857261
transform 1 0 197593 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1528
timestamp 1624857261
transform 1 0 197929 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1527
timestamp 1624857261
transform 1 0 198265 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1526
timestamp 1624857261
transform 1 0 198601 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1525
timestamp 1624857261
transform 1 0 198937 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1524
timestamp 1624857261
transform 1 0 199273 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1523
timestamp 1624857261
transform 1 0 199609 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1522
timestamp 1624857261
transform 1 0 199945 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1521
timestamp 1624857261
transform 1 0 200281 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1520
timestamp 1624857261
transform 1 0 200617 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1519
timestamp 1624857261
transform 1 0 200953 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1518
timestamp 1624857261
transform 1 0 201289 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1517
timestamp 1624857261
transform 1 0 201625 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1516
timestamp 1624857261
transform 1 0 201961 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1515
timestamp 1624857261
transform 1 0 202297 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1514
timestamp 1624857261
transform 1 0 202633 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1513
timestamp 1624857261
transform 1 0 202969 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1512
timestamp 1624857261
transform 1 0 203305 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1511
timestamp 1624857261
transform 1 0 203641 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1510
timestamp 1624857261
transform 1 0 203977 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1509
timestamp 1624857261
transform 1 0 204313 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1508
timestamp 1624857261
transform 1 0 204649 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1507
timestamp 1624857261
transform 1 0 204985 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1506
timestamp 1624857261
transform 1 0 205321 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1505
timestamp 1624857261
transform 1 0 205657 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1504
timestamp 1624857261
transform 1 0 205993 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1503
timestamp 1624857261
transform 1 0 206329 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1502
timestamp 1624857261
transform 1 0 206665 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1501
timestamp 1624857261
transform 1 0 207001 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1500
timestamp 1624857261
transform 1 0 207337 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1499
timestamp 1624857261
transform 1 0 207673 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1498
timestamp 1624857261
transform 1 0 208009 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1497
timestamp 1624857261
transform 1 0 208345 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1496
timestamp 1624857261
transform 1 0 208681 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1495
timestamp 1624857261
transform 1 0 209017 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1494
timestamp 1624857261
transform 1 0 209353 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1493
timestamp 1624857261
transform 1 0 209689 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1492
timestamp 1624857261
transform 1 0 210025 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1491
timestamp 1624857261
transform 1 0 210361 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1490
timestamp 1624857261
transform 1 0 210697 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1489
timestamp 1624857261
transform 1 0 211033 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1488
timestamp 1624857261
transform 1 0 211369 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1487
timestamp 1624857261
transform 1 0 211705 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1486
timestamp 1624857261
transform 1 0 212041 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1485
timestamp 1624857261
transform 1 0 212377 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1484
timestamp 1624857261
transform 1 0 212713 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1483
timestamp 1624857261
transform 1 0 213049 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1482
timestamp 1624857261
transform 1 0 213385 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1481
timestamp 1624857261
transform 1 0 213721 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1480
timestamp 1624857261
transform 1 0 214057 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1479
timestamp 1624857261
transform 1 0 214393 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1478
timestamp 1624857261
transform 1 0 214729 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1477
timestamp 1624857261
transform 1 0 215065 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1476
timestamp 1624857261
transform 1 0 215401 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1475
timestamp 1624857261
transform 1 0 215737 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1474
timestamp 1624857261
transform 1 0 216073 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1473
timestamp 1624857261
transform 1 0 216409 0 1 1807
box 0 0 1 1
use contact_13  contact_13_1472
timestamp 1624857261
transform 1 0 2041 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1471
timestamp 1624857261
transform 1 0 2377 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1470
timestamp 1624857261
transform 1 0 2713 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1469
timestamp 1624857261
transform 1 0 3049 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1468
timestamp 1624857261
transform 1 0 3385 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1467
timestamp 1624857261
transform 1 0 3721 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1466
timestamp 1624857261
transform 1 0 4057 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1465
timestamp 1624857261
transform 1 0 4393 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1464
timestamp 1624857261
transform 1 0 4729 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1463
timestamp 1624857261
transform 1 0 5065 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1462
timestamp 1624857261
transform 1 0 5401 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1461
timestamp 1624857261
transform 1 0 5737 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1460
timestamp 1624857261
transform 1 0 6073 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1459
timestamp 1624857261
transform 1 0 6409 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1458
timestamp 1624857261
transform 1 0 6745 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1457
timestamp 1624857261
transform 1 0 7081 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1456
timestamp 1624857261
transform 1 0 7417 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1455
timestamp 1624857261
transform 1 0 7753 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1454
timestamp 1624857261
transform 1 0 8089 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1453
timestamp 1624857261
transform 1 0 8425 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1452
timestamp 1624857261
transform 1 0 8761 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1451
timestamp 1624857261
transform 1 0 9097 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1450
timestamp 1624857261
transform 1 0 9433 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1449
timestamp 1624857261
transform 1 0 9769 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1448
timestamp 1624857261
transform 1 0 10105 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1447
timestamp 1624857261
transform 1 0 10441 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1446
timestamp 1624857261
transform 1 0 10777 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1445
timestamp 1624857261
transform 1 0 11113 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1444
timestamp 1624857261
transform 1 0 11449 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1443
timestamp 1624857261
transform 1 0 11785 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1442
timestamp 1624857261
transform 1 0 12121 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1441
timestamp 1624857261
transform 1 0 12457 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1440
timestamp 1624857261
transform 1 0 12793 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1439
timestamp 1624857261
transform 1 0 13129 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1438
timestamp 1624857261
transform 1 0 13465 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1437
timestamp 1624857261
transform 1 0 13801 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1436
timestamp 1624857261
transform 1 0 14137 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1435
timestamp 1624857261
transform 1 0 14473 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1434
timestamp 1624857261
transform 1 0 14809 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1433
timestamp 1624857261
transform 1 0 15145 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1432
timestamp 1624857261
transform 1 0 15481 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1431
timestamp 1624857261
transform 1 0 15817 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1430
timestamp 1624857261
transform 1 0 16153 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1429
timestamp 1624857261
transform 1 0 16489 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1428
timestamp 1624857261
transform 1 0 16825 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1427
timestamp 1624857261
transform 1 0 17161 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1426
timestamp 1624857261
transform 1 0 17497 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1425
timestamp 1624857261
transform 1 0 17833 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1424
timestamp 1624857261
transform 1 0 18169 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1423
timestamp 1624857261
transform 1 0 18505 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1422
timestamp 1624857261
transform 1 0 18841 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1421
timestamp 1624857261
transform 1 0 19177 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1420
timestamp 1624857261
transform 1 0 19513 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1419
timestamp 1624857261
transform 1 0 19849 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1418
timestamp 1624857261
transform 1 0 20185 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1417
timestamp 1624857261
transform 1 0 20521 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1416
timestamp 1624857261
transform 1 0 20857 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1415
timestamp 1624857261
transform 1 0 21193 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1414
timestamp 1624857261
transform 1 0 21529 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1413
timestamp 1624857261
transform 1 0 21865 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1412
timestamp 1624857261
transform 1 0 22201 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1411
timestamp 1624857261
transform 1 0 22537 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1410
timestamp 1624857261
transform 1 0 22873 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1409
timestamp 1624857261
transform 1 0 23209 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1408
timestamp 1624857261
transform 1 0 23545 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1407
timestamp 1624857261
transform 1 0 23881 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1406
timestamp 1624857261
transform 1 0 24217 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1405
timestamp 1624857261
transform 1 0 24553 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1404
timestamp 1624857261
transform 1 0 24889 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1403
timestamp 1624857261
transform 1 0 25225 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1402
timestamp 1624857261
transform 1 0 25561 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1401
timestamp 1624857261
transform 1 0 25897 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1400
timestamp 1624857261
transform 1 0 26233 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1399
timestamp 1624857261
transform 1 0 26569 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1398
timestamp 1624857261
transform 1 0 26905 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1397
timestamp 1624857261
transform 1 0 27241 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1396
timestamp 1624857261
transform 1 0 27577 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1395
timestamp 1624857261
transform 1 0 27913 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1394
timestamp 1624857261
transform 1 0 28249 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1393
timestamp 1624857261
transform 1 0 28585 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1392
timestamp 1624857261
transform 1 0 28921 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1391
timestamp 1624857261
transform 1 0 29257 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1390
timestamp 1624857261
transform 1 0 29593 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1389
timestamp 1624857261
transform 1 0 29929 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1388
timestamp 1624857261
transform 1 0 30265 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1387
timestamp 1624857261
transform 1 0 30601 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1386
timestamp 1624857261
transform 1 0 30937 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1385
timestamp 1624857261
transform 1 0 31273 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1384
timestamp 1624857261
transform 1 0 31609 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1383
timestamp 1624857261
transform 1 0 31945 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1382
timestamp 1624857261
transform 1 0 32281 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1381
timestamp 1624857261
transform 1 0 32617 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1380
timestamp 1624857261
transform 1 0 32953 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1379
timestamp 1624857261
transform 1 0 33289 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1378
timestamp 1624857261
transform 1 0 33625 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1377
timestamp 1624857261
transform 1 0 33961 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1376
timestamp 1624857261
transform 1 0 34297 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1375
timestamp 1624857261
transform 1 0 34633 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1374
timestamp 1624857261
transform 1 0 34969 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1373
timestamp 1624857261
transform 1 0 35305 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1372
timestamp 1624857261
transform 1 0 35641 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1371
timestamp 1624857261
transform 1 0 35977 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1370
timestamp 1624857261
transform 1 0 36313 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1369
timestamp 1624857261
transform 1 0 36649 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1368
timestamp 1624857261
transform 1 0 36985 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1367
timestamp 1624857261
transform 1 0 37321 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1366
timestamp 1624857261
transform 1 0 37657 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1365
timestamp 1624857261
transform 1 0 37993 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1364
timestamp 1624857261
transform 1 0 38329 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1363
timestamp 1624857261
transform 1 0 38665 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1362
timestamp 1624857261
transform 1 0 39001 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1361
timestamp 1624857261
transform 1 0 39337 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1360
timestamp 1624857261
transform 1 0 39673 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1359
timestamp 1624857261
transform 1 0 40009 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1358
timestamp 1624857261
transform 1 0 40345 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1357
timestamp 1624857261
transform 1 0 40681 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1356
timestamp 1624857261
transform 1 0 41017 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1355
timestamp 1624857261
transform 1 0 41353 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1354
timestamp 1624857261
transform 1 0 41689 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1353
timestamp 1624857261
transform 1 0 42025 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1352
timestamp 1624857261
transform 1 0 42361 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1351
timestamp 1624857261
transform 1 0 42697 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1350
timestamp 1624857261
transform 1 0 43033 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1349
timestamp 1624857261
transform 1 0 43369 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1348
timestamp 1624857261
transform 1 0 43705 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1347
timestamp 1624857261
transform 1 0 44041 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1346
timestamp 1624857261
transform 1 0 44377 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1345
timestamp 1624857261
transform 1 0 44713 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1344
timestamp 1624857261
transform 1 0 45049 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1343
timestamp 1624857261
transform 1 0 45385 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1342
timestamp 1624857261
transform 1 0 45721 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1341
timestamp 1624857261
transform 1 0 46057 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1340
timestamp 1624857261
transform 1 0 46393 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1339
timestamp 1624857261
transform 1 0 46729 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1338
timestamp 1624857261
transform 1 0 47065 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1337
timestamp 1624857261
transform 1 0 47401 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1336
timestamp 1624857261
transform 1 0 47737 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1335
timestamp 1624857261
transform 1 0 48073 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1334
timestamp 1624857261
transform 1 0 48409 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1333
timestamp 1624857261
transform 1 0 48745 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1332
timestamp 1624857261
transform 1 0 49081 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1331
timestamp 1624857261
transform 1 0 49417 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1330
timestamp 1624857261
transform 1 0 49753 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1329
timestamp 1624857261
transform 1 0 50089 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1328
timestamp 1624857261
transform 1 0 50425 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1327
timestamp 1624857261
transform 1 0 50761 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1326
timestamp 1624857261
transform 1 0 51097 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1325
timestamp 1624857261
transform 1 0 51433 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1324
timestamp 1624857261
transform 1 0 51769 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1323
timestamp 1624857261
transform 1 0 52105 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1322
timestamp 1624857261
transform 1 0 52441 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1321
timestamp 1624857261
transform 1 0 52777 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1320
timestamp 1624857261
transform 1 0 53113 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1319
timestamp 1624857261
transform 1 0 53449 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1318
timestamp 1624857261
transform 1 0 53785 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1317
timestamp 1624857261
transform 1 0 54121 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1316
timestamp 1624857261
transform 1 0 54457 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1315
timestamp 1624857261
transform 1 0 54793 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1314
timestamp 1624857261
transform 1 0 55129 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1313
timestamp 1624857261
transform 1 0 55465 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1312
timestamp 1624857261
transform 1 0 55801 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1311
timestamp 1624857261
transform 1 0 56137 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1310
timestamp 1624857261
transform 1 0 56473 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1309
timestamp 1624857261
transform 1 0 56809 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1308
timestamp 1624857261
transform 1 0 57145 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1307
timestamp 1624857261
transform 1 0 57481 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1306
timestamp 1624857261
transform 1 0 57817 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1305
timestamp 1624857261
transform 1 0 58153 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1304
timestamp 1624857261
transform 1 0 58489 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1303
timestamp 1624857261
transform 1 0 58825 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1302
timestamp 1624857261
transform 1 0 59161 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1301
timestamp 1624857261
transform 1 0 59497 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1300
timestamp 1624857261
transform 1 0 59833 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1299
timestamp 1624857261
transform 1 0 60169 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1298
timestamp 1624857261
transform 1 0 60505 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1297
timestamp 1624857261
transform 1 0 60841 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1296
timestamp 1624857261
transform 1 0 61177 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1295
timestamp 1624857261
transform 1 0 61513 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1294
timestamp 1624857261
transform 1 0 61849 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1293
timestamp 1624857261
transform 1 0 62185 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1292
timestamp 1624857261
transform 1 0 62521 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1291
timestamp 1624857261
transform 1 0 62857 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1290
timestamp 1624857261
transform 1 0 63193 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1289
timestamp 1624857261
transform 1 0 63529 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1288
timestamp 1624857261
transform 1 0 63865 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1287
timestamp 1624857261
transform 1 0 64201 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1286
timestamp 1624857261
transform 1 0 64537 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1285
timestamp 1624857261
transform 1 0 64873 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1284
timestamp 1624857261
transform 1 0 65209 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1283
timestamp 1624857261
transform 1 0 65545 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1282
timestamp 1624857261
transform 1 0 65881 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1281
timestamp 1624857261
transform 1 0 66217 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1280
timestamp 1624857261
transform 1 0 66553 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1279
timestamp 1624857261
transform 1 0 66889 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1278
timestamp 1624857261
transform 1 0 67225 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1277
timestamp 1624857261
transform 1 0 67561 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1276
timestamp 1624857261
transform 1 0 67897 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1275
timestamp 1624857261
transform 1 0 68233 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1274
timestamp 1624857261
transform 1 0 68569 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1273
timestamp 1624857261
transform 1 0 68905 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1272
timestamp 1624857261
transform 1 0 69241 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1271
timestamp 1624857261
transform 1 0 69577 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1270
timestamp 1624857261
transform 1 0 69913 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1269
timestamp 1624857261
transform 1 0 70249 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1268
timestamp 1624857261
transform 1 0 70585 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1267
timestamp 1624857261
transform 1 0 70921 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1266
timestamp 1624857261
transform 1 0 71257 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1265
timestamp 1624857261
transform 1 0 71593 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1264
timestamp 1624857261
transform 1 0 71929 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1263
timestamp 1624857261
transform 1 0 72265 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1262
timestamp 1624857261
transform 1 0 72601 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1261
timestamp 1624857261
transform 1 0 72937 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1260
timestamp 1624857261
transform 1 0 73273 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1259
timestamp 1624857261
transform 1 0 73609 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1258
timestamp 1624857261
transform 1 0 73945 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1257
timestamp 1624857261
transform 1 0 74281 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1256
timestamp 1624857261
transform 1 0 74617 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1255
timestamp 1624857261
transform 1 0 74953 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1254
timestamp 1624857261
transform 1 0 75289 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1253
timestamp 1624857261
transform 1 0 75625 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1252
timestamp 1624857261
transform 1 0 75961 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1251
timestamp 1624857261
transform 1 0 76297 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1250
timestamp 1624857261
transform 1 0 76633 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1249
timestamp 1624857261
transform 1 0 76969 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1248
timestamp 1624857261
transform 1 0 77305 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1247
timestamp 1624857261
transform 1 0 77641 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1246
timestamp 1624857261
transform 1 0 77977 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1245
timestamp 1624857261
transform 1 0 78313 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1244
timestamp 1624857261
transform 1 0 78649 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1243
timestamp 1624857261
transform 1 0 78985 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1242
timestamp 1624857261
transform 1 0 79321 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1241
timestamp 1624857261
transform 1 0 79657 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1240
timestamp 1624857261
transform 1 0 79993 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1239
timestamp 1624857261
transform 1 0 80329 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1238
timestamp 1624857261
transform 1 0 80665 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1237
timestamp 1624857261
transform 1 0 81001 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1236
timestamp 1624857261
transform 1 0 81337 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1235
timestamp 1624857261
transform 1 0 81673 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1234
timestamp 1624857261
transform 1 0 82009 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1233
timestamp 1624857261
transform 1 0 82345 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1232
timestamp 1624857261
transform 1 0 82681 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1231
timestamp 1624857261
transform 1 0 83017 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1230
timestamp 1624857261
transform 1 0 83353 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1229
timestamp 1624857261
transform 1 0 83689 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1228
timestamp 1624857261
transform 1 0 84025 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1227
timestamp 1624857261
transform 1 0 84361 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1226
timestamp 1624857261
transform 1 0 84697 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1225
timestamp 1624857261
transform 1 0 85033 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1224
timestamp 1624857261
transform 1 0 85369 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1223
timestamp 1624857261
transform 1 0 85705 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1222
timestamp 1624857261
transform 1 0 86041 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1221
timestamp 1624857261
transform 1 0 86377 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1220
timestamp 1624857261
transform 1 0 86713 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1219
timestamp 1624857261
transform 1 0 87049 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1218
timestamp 1624857261
transform 1 0 87385 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1217
timestamp 1624857261
transform 1 0 87721 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1216
timestamp 1624857261
transform 1 0 88057 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1215
timestamp 1624857261
transform 1 0 88393 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1214
timestamp 1624857261
transform 1 0 88729 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1213
timestamp 1624857261
transform 1 0 89065 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1212
timestamp 1624857261
transform 1 0 89401 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1211
timestamp 1624857261
transform 1 0 89737 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1210
timestamp 1624857261
transform 1 0 90073 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1209
timestamp 1624857261
transform 1 0 90409 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1208
timestamp 1624857261
transform 1 0 90745 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1207
timestamp 1624857261
transform 1 0 91081 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1206
timestamp 1624857261
transform 1 0 91417 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1205
timestamp 1624857261
transform 1 0 91753 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1204
timestamp 1624857261
transform 1 0 92089 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1203
timestamp 1624857261
transform 1 0 92425 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1202
timestamp 1624857261
transform 1 0 92761 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1201
timestamp 1624857261
transform 1 0 93097 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1200
timestamp 1624857261
transform 1 0 93433 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1199
timestamp 1624857261
transform 1 0 93769 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1198
timestamp 1624857261
transform 1 0 94105 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1197
timestamp 1624857261
transform 1 0 94441 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1196
timestamp 1624857261
transform 1 0 94777 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1195
timestamp 1624857261
transform 1 0 95113 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1194
timestamp 1624857261
transform 1 0 95449 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1193
timestamp 1624857261
transform 1 0 95785 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1192
timestamp 1624857261
transform 1 0 96121 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1191
timestamp 1624857261
transform 1 0 96457 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1190
timestamp 1624857261
transform 1 0 96793 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1189
timestamp 1624857261
transform 1 0 97129 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1188
timestamp 1624857261
transform 1 0 97465 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1187
timestamp 1624857261
transform 1 0 97801 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1186
timestamp 1624857261
transform 1 0 98137 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1185
timestamp 1624857261
transform 1 0 98473 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1184
timestamp 1624857261
transform 1 0 98809 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1183
timestamp 1624857261
transform 1 0 99145 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1182
timestamp 1624857261
transform 1 0 99481 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1181
timestamp 1624857261
transform 1 0 99817 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1180
timestamp 1624857261
transform 1 0 100153 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1179
timestamp 1624857261
transform 1 0 100489 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1178
timestamp 1624857261
transform 1 0 100825 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1177
timestamp 1624857261
transform 1 0 101161 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1176
timestamp 1624857261
transform 1 0 101497 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1175
timestamp 1624857261
transform 1 0 101833 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1174
timestamp 1624857261
transform 1 0 102169 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1173
timestamp 1624857261
transform 1 0 102505 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1172
timestamp 1624857261
transform 1 0 102841 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1171
timestamp 1624857261
transform 1 0 103177 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1170
timestamp 1624857261
transform 1 0 103513 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1169
timestamp 1624857261
transform 1 0 103849 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1168
timestamp 1624857261
transform 1 0 104185 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1167
timestamp 1624857261
transform 1 0 104521 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1166
timestamp 1624857261
transform 1 0 104857 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1165
timestamp 1624857261
transform 1 0 105193 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1164
timestamp 1624857261
transform 1 0 105529 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1163
timestamp 1624857261
transform 1 0 105865 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1162
timestamp 1624857261
transform 1 0 106201 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1161
timestamp 1624857261
transform 1 0 106537 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1160
timestamp 1624857261
transform 1 0 106873 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1159
timestamp 1624857261
transform 1 0 107209 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1158
timestamp 1624857261
transform 1 0 107545 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1157
timestamp 1624857261
transform 1 0 107881 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1156
timestamp 1624857261
transform 1 0 108217 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1155
timestamp 1624857261
transform 1 0 108553 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1154
timestamp 1624857261
transform 1 0 108889 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1153
timestamp 1624857261
transform 1 0 109225 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1152
timestamp 1624857261
transform 1 0 109561 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1151
timestamp 1624857261
transform 1 0 109897 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1150
timestamp 1624857261
transform 1 0 110233 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1149
timestamp 1624857261
transform 1 0 110569 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1148
timestamp 1624857261
transform 1 0 110905 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1147
timestamp 1624857261
transform 1 0 111241 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1146
timestamp 1624857261
transform 1 0 111577 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1145
timestamp 1624857261
transform 1 0 111913 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1144
timestamp 1624857261
transform 1 0 112249 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1143
timestamp 1624857261
transform 1 0 112585 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1142
timestamp 1624857261
transform 1 0 112921 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1141
timestamp 1624857261
transform 1 0 113257 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1140
timestamp 1624857261
transform 1 0 113593 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1139
timestamp 1624857261
transform 1 0 113929 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1138
timestamp 1624857261
transform 1 0 114265 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1137
timestamp 1624857261
transform 1 0 114601 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1136
timestamp 1624857261
transform 1 0 114937 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1135
timestamp 1624857261
transform 1 0 115273 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1134
timestamp 1624857261
transform 1 0 115609 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1133
timestamp 1624857261
transform 1 0 115945 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1132
timestamp 1624857261
transform 1 0 116281 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1131
timestamp 1624857261
transform 1 0 116617 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1130
timestamp 1624857261
transform 1 0 116953 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1129
timestamp 1624857261
transform 1 0 117289 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1128
timestamp 1624857261
transform 1 0 117625 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1127
timestamp 1624857261
transform 1 0 117961 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1126
timestamp 1624857261
transform 1 0 118297 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1125
timestamp 1624857261
transform 1 0 118633 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1124
timestamp 1624857261
transform 1 0 118969 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1123
timestamp 1624857261
transform 1 0 119305 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1122
timestamp 1624857261
transform 1 0 119641 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1121
timestamp 1624857261
transform 1 0 119977 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1120
timestamp 1624857261
transform 1 0 120313 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1119
timestamp 1624857261
transform 1 0 120649 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1118
timestamp 1624857261
transform 1 0 120985 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1117
timestamp 1624857261
transform 1 0 121321 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1116
timestamp 1624857261
transform 1 0 121657 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1115
timestamp 1624857261
transform 1 0 121993 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1114
timestamp 1624857261
transform 1 0 122329 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1113
timestamp 1624857261
transform 1 0 122665 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1112
timestamp 1624857261
transform 1 0 123001 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1111
timestamp 1624857261
transform 1 0 123337 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1110
timestamp 1624857261
transform 1 0 123673 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1109
timestamp 1624857261
transform 1 0 124009 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1108
timestamp 1624857261
transform 1 0 124345 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1107
timestamp 1624857261
transform 1 0 124681 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1106
timestamp 1624857261
transform 1 0 125017 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1105
timestamp 1624857261
transform 1 0 125353 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1104
timestamp 1624857261
transform 1 0 125689 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1103
timestamp 1624857261
transform 1 0 126025 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1102
timestamp 1624857261
transform 1 0 126361 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1101
timestamp 1624857261
transform 1 0 126697 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1100
timestamp 1624857261
transform 1 0 127033 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1099
timestamp 1624857261
transform 1 0 127369 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1098
timestamp 1624857261
transform 1 0 127705 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1097
timestamp 1624857261
transform 1 0 128041 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1096
timestamp 1624857261
transform 1 0 128377 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1095
timestamp 1624857261
transform 1 0 128713 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1094
timestamp 1624857261
transform 1 0 129049 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1093
timestamp 1624857261
transform 1 0 129385 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1092
timestamp 1624857261
transform 1 0 129721 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1091
timestamp 1624857261
transform 1 0 130057 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1090
timestamp 1624857261
transform 1 0 130393 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1089
timestamp 1624857261
transform 1 0 130729 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1088
timestamp 1624857261
transform 1 0 131065 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1087
timestamp 1624857261
transform 1 0 131401 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1086
timestamp 1624857261
transform 1 0 131737 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1085
timestamp 1624857261
transform 1 0 132073 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1084
timestamp 1624857261
transform 1 0 132409 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1083
timestamp 1624857261
transform 1 0 132745 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1082
timestamp 1624857261
transform 1 0 133081 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1081
timestamp 1624857261
transform 1 0 133417 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1080
timestamp 1624857261
transform 1 0 133753 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1079
timestamp 1624857261
transform 1 0 134089 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1078
timestamp 1624857261
transform 1 0 134425 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1077
timestamp 1624857261
transform 1 0 134761 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1076
timestamp 1624857261
transform 1 0 135097 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1075
timestamp 1624857261
transform 1 0 135433 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1074
timestamp 1624857261
transform 1 0 135769 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1073
timestamp 1624857261
transform 1 0 136105 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1072
timestamp 1624857261
transform 1 0 136441 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1071
timestamp 1624857261
transform 1 0 136777 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1070
timestamp 1624857261
transform 1 0 137113 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1069
timestamp 1624857261
transform 1 0 137449 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1068
timestamp 1624857261
transform 1 0 137785 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1067
timestamp 1624857261
transform 1 0 138121 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1066
timestamp 1624857261
transform 1 0 138457 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1065
timestamp 1624857261
transform 1 0 138793 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1064
timestamp 1624857261
transform 1 0 139129 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1063
timestamp 1624857261
transform 1 0 139465 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1062
timestamp 1624857261
transform 1 0 139801 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1061
timestamp 1624857261
transform 1 0 140137 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1060
timestamp 1624857261
transform 1 0 140473 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1059
timestamp 1624857261
transform 1 0 140809 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1058
timestamp 1624857261
transform 1 0 141145 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1057
timestamp 1624857261
transform 1 0 141481 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1056
timestamp 1624857261
transform 1 0 141817 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1055
timestamp 1624857261
transform 1 0 142153 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1054
timestamp 1624857261
transform 1 0 142489 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1053
timestamp 1624857261
transform 1 0 142825 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1052
timestamp 1624857261
transform 1 0 143161 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1051
timestamp 1624857261
transform 1 0 143497 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1050
timestamp 1624857261
transform 1 0 143833 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1049
timestamp 1624857261
transform 1 0 144169 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1048
timestamp 1624857261
transform 1 0 144505 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1047
timestamp 1624857261
transform 1 0 144841 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1046
timestamp 1624857261
transform 1 0 145177 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1045
timestamp 1624857261
transform 1 0 145513 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1044
timestamp 1624857261
transform 1 0 145849 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1043
timestamp 1624857261
transform 1 0 146185 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1042
timestamp 1624857261
transform 1 0 146521 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1041
timestamp 1624857261
transform 1 0 146857 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1040
timestamp 1624857261
transform 1 0 147193 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1039
timestamp 1624857261
transform 1 0 147529 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1038
timestamp 1624857261
transform 1 0 147865 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1037
timestamp 1624857261
transform 1 0 148201 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1036
timestamp 1624857261
transform 1 0 148537 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1035
timestamp 1624857261
transform 1 0 148873 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1034
timestamp 1624857261
transform 1 0 149209 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1033
timestamp 1624857261
transform 1 0 149545 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1032
timestamp 1624857261
transform 1 0 149881 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1031
timestamp 1624857261
transform 1 0 150217 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1030
timestamp 1624857261
transform 1 0 150553 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1029
timestamp 1624857261
transform 1 0 150889 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1028
timestamp 1624857261
transform 1 0 151225 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1027
timestamp 1624857261
transform 1 0 151561 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1026
timestamp 1624857261
transform 1 0 151897 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1025
timestamp 1624857261
transform 1 0 152233 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1024
timestamp 1624857261
transform 1 0 152569 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1023
timestamp 1624857261
transform 1 0 152905 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1022
timestamp 1624857261
transform 1 0 153241 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1021
timestamp 1624857261
transform 1 0 153577 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1020
timestamp 1624857261
transform 1 0 153913 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1019
timestamp 1624857261
transform 1 0 154249 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1018
timestamp 1624857261
transform 1 0 154585 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1017
timestamp 1624857261
transform 1 0 154921 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1016
timestamp 1624857261
transform 1 0 155257 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1015
timestamp 1624857261
transform 1 0 155593 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1014
timestamp 1624857261
transform 1 0 155929 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1013
timestamp 1624857261
transform 1 0 156265 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1012
timestamp 1624857261
transform 1 0 156601 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1011
timestamp 1624857261
transform 1 0 156937 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1010
timestamp 1624857261
transform 1 0 157273 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1009
timestamp 1624857261
transform 1 0 157609 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1008
timestamp 1624857261
transform 1 0 157945 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1007
timestamp 1624857261
transform 1 0 158281 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1006
timestamp 1624857261
transform 1 0 158617 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1005
timestamp 1624857261
transform 1 0 158953 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1004
timestamp 1624857261
transform 1 0 159289 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1003
timestamp 1624857261
transform 1 0 159625 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1002
timestamp 1624857261
transform 1 0 159961 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1001
timestamp 1624857261
transform 1 0 160297 0 1 142303
box 0 0 1 1
use contact_13  contact_13_1000
timestamp 1624857261
transform 1 0 160633 0 1 142303
box 0 0 1 1
use contact_13  contact_13_999
timestamp 1624857261
transform 1 0 160969 0 1 142303
box 0 0 1 1
use contact_13  contact_13_998
timestamp 1624857261
transform 1 0 161305 0 1 142303
box 0 0 1 1
use contact_13  contact_13_997
timestamp 1624857261
transform 1 0 161641 0 1 142303
box 0 0 1 1
use contact_13  contact_13_996
timestamp 1624857261
transform 1 0 161977 0 1 142303
box 0 0 1 1
use contact_13  contact_13_995
timestamp 1624857261
transform 1 0 162313 0 1 142303
box 0 0 1 1
use contact_13  contact_13_994
timestamp 1624857261
transform 1 0 162649 0 1 142303
box 0 0 1 1
use contact_13  contact_13_993
timestamp 1624857261
transform 1 0 162985 0 1 142303
box 0 0 1 1
use contact_13  contact_13_992
timestamp 1624857261
transform 1 0 163321 0 1 142303
box 0 0 1 1
use contact_13  contact_13_991
timestamp 1624857261
transform 1 0 163657 0 1 142303
box 0 0 1 1
use contact_13  contact_13_990
timestamp 1624857261
transform 1 0 163993 0 1 142303
box 0 0 1 1
use contact_13  contact_13_989
timestamp 1624857261
transform 1 0 164329 0 1 142303
box 0 0 1 1
use contact_13  contact_13_988
timestamp 1624857261
transform 1 0 164665 0 1 142303
box 0 0 1 1
use contact_13  contact_13_987
timestamp 1624857261
transform 1 0 165001 0 1 142303
box 0 0 1 1
use contact_13  contact_13_986
timestamp 1624857261
transform 1 0 165337 0 1 142303
box 0 0 1 1
use contact_13  contact_13_985
timestamp 1624857261
transform 1 0 165673 0 1 142303
box 0 0 1 1
use contact_13  contact_13_984
timestamp 1624857261
transform 1 0 166009 0 1 142303
box 0 0 1 1
use contact_13  contact_13_983
timestamp 1624857261
transform 1 0 166345 0 1 142303
box 0 0 1 1
use contact_13  contact_13_982
timestamp 1624857261
transform 1 0 166681 0 1 142303
box 0 0 1 1
use contact_13  contact_13_981
timestamp 1624857261
transform 1 0 167017 0 1 142303
box 0 0 1 1
use contact_13  contact_13_980
timestamp 1624857261
transform 1 0 167353 0 1 142303
box 0 0 1 1
use contact_13  contact_13_979
timestamp 1624857261
transform 1 0 167689 0 1 142303
box 0 0 1 1
use contact_13  contact_13_978
timestamp 1624857261
transform 1 0 168025 0 1 142303
box 0 0 1 1
use contact_13  contact_13_977
timestamp 1624857261
transform 1 0 168361 0 1 142303
box 0 0 1 1
use contact_13  contact_13_976
timestamp 1624857261
transform 1 0 168697 0 1 142303
box 0 0 1 1
use contact_13  contact_13_975
timestamp 1624857261
transform 1 0 169033 0 1 142303
box 0 0 1 1
use contact_13  contact_13_974
timestamp 1624857261
transform 1 0 169369 0 1 142303
box 0 0 1 1
use contact_13  contact_13_973
timestamp 1624857261
transform 1 0 169705 0 1 142303
box 0 0 1 1
use contact_13  contact_13_972
timestamp 1624857261
transform 1 0 170041 0 1 142303
box 0 0 1 1
use contact_13  contact_13_971
timestamp 1624857261
transform 1 0 170377 0 1 142303
box 0 0 1 1
use contact_13  contact_13_970
timestamp 1624857261
transform 1 0 170713 0 1 142303
box 0 0 1 1
use contact_13  contact_13_969
timestamp 1624857261
transform 1 0 171049 0 1 142303
box 0 0 1 1
use contact_13  contact_13_968
timestamp 1624857261
transform 1 0 171385 0 1 142303
box 0 0 1 1
use contact_13  contact_13_967
timestamp 1624857261
transform 1 0 171721 0 1 142303
box 0 0 1 1
use contact_13  contact_13_966
timestamp 1624857261
transform 1 0 172057 0 1 142303
box 0 0 1 1
use contact_13  contact_13_965
timestamp 1624857261
transform 1 0 172393 0 1 142303
box 0 0 1 1
use contact_13  contact_13_964
timestamp 1624857261
transform 1 0 172729 0 1 142303
box 0 0 1 1
use contact_13  contact_13_963
timestamp 1624857261
transform 1 0 173065 0 1 142303
box 0 0 1 1
use contact_13  contact_13_962
timestamp 1624857261
transform 1 0 173401 0 1 142303
box 0 0 1 1
use contact_13  contact_13_961
timestamp 1624857261
transform 1 0 173737 0 1 142303
box 0 0 1 1
use contact_13  contact_13_960
timestamp 1624857261
transform 1 0 174073 0 1 142303
box 0 0 1 1
use contact_13  contact_13_959
timestamp 1624857261
transform 1 0 174409 0 1 142303
box 0 0 1 1
use contact_13  contact_13_958
timestamp 1624857261
transform 1 0 174745 0 1 142303
box 0 0 1 1
use contact_13  contact_13_957
timestamp 1624857261
transform 1 0 175081 0 1 142303
box 0 0 1 1
use contact_13  contact_13_956
timestamp 1624857261
transform 1 0 175417 0 1 142303
box 0 0 1 1
use contact_13  contact_13_955
timestamp 1624857261
transform 1 0 175753 0 1 142303
box 0 0 1 1
use contact_13  contact_13_954
timestamp 1624857261
transform 1 0 176089 0 1 142303
box 0 0 1 1
use contact_13  contact_13_953
timestamp 1624857261
transform 1 0 176425 0 1 142303
box 0 0 1 1
use contact_13  contact_13_952
timestamp 1624857261
transform 1 0 176761 0 1 142303
box 0 0 1 1
use contact_13  contact_13_951
timestamp 1624857261
transform 1 0 177097 0 1 142303
box 0 0 1 1
use contact_13  contact_13_950
timestamp 1624857261
transform 1 0 177433 0 1 142303
box 0 0 1 1
use contact_13  contact_13_949
timestamp 1624857261
transform 1 0 177769 0 1 142303
box 0 0 1 1
use contact_13  contact_13_948
timestamp 1624857261
transform 1 0 178105 0 1 142303
box 0 0 1 1
use contact_13  contact_13_947
timestamp 1624857261
transform 1 0 178441 0 1 142303
box 0 0 1 1
use contact_13  contact_13_946
timestamp 1624857261
transform 1 0 178777 0 1 142303
box 0 0 1 1
use contact_13  contact_13_945
timestamp 1624857261
transform 1 0 179113 0 1 142303
box 0 0 1 1
use contact_13  contact_13_944
timestamp 1624857261
transform 1 0 179449 0 1 142303
box 0 0 1 1
use contact_13  contact_13_943
timestamp 1624857261
transform 1 0 179785 0 1 142303
box 0 0 1 1
use contact_13  contact_13_942
timestamp 1624857261
transform 1 0 180121 0 1 142303
box 0 0 1 1
use contact_13  contact_13_941
timestamp 1624857261
transform 1 0 180457 0 1 142303
box 0 0 1 1
use contact_13  contact_13_940
timestamp 1624857261
transform 1 0 180793 0 1 142303
box 0 0 1 1
use contact_13  contact_13_939
timestamp 1624857261
transform 1 0 181129 0 1 142303
box 0 0 1 1
use contact_13  contact_13_938
timestamp 1624857261
transform 1 0 181465 0 1 142303
box 0 0 1 1
use contact_13  contact_13_937
timestamp 1624857261
transform 1 0 181801 0 1 142303
box 0 0 1 1
use contact_13  contact_13_936
timestamp 1624857261
transform 1 0 182137 0 1 142303
box 0 0 1 1
use contact_13  contact_13_935
timestamp 1624857261
transform 1 0 182473 0 1 142303
box 0 0 1 1
use contact_13  contact_13_934
timestamp 1624857261
transform 1 0 182809 0 1 142303
box 0 0 1 1
use contact_13  contact_13_933
timestamp 1624857261
transform 1 0 183145 0 1 142303
box 0 0 1 1
use contact_13  contact_13_932
timestamp 1624857261
transform 1 0 183481 0 1 142303
box 0 0 1 1
use contact_13  contact_13_931
timestamp 1624857261
transform 1 0 183817 0 1 142303
box 0 0 1 1
use contact_13  contact_13_930
timestamp 1624857261
transform 1 0 184153 0 1 142303
box 0 0 1 1
use contact_13  contact_13_929
timestamp 1624857261
transform 1 0 184489 0 1 142303
box 0 0 1 1
use contact_13  contact_13_928
timestamp 1624857261
transform 1 0 184825 0 1 142303
box 0 0 1 1
use contact_13  contact_13_927
timestamp 1624857261
transform 1 0 185161 0 1 142303
box 0 0 1 1
use contact_13  contact_13_926
timestamp 1624857261
transform 1 0 185497 0 1 142303
box 0 0 1 1
use contact_13  contact_13_925
timestamp 1624857261
transform 1 0 185833 0 1 142303
box 0 0 1 1
use contact_13  contact_13_924
timestamp 1624857261
transform 1 0 186169 0 1 142303
box 0 0 1 1
use contact_13  contact_13_923
timestamp 1624857261
transform 1 0 186505 0 1 142303
box 0 0 1 1
use contact_13  contact_13_922
timestamp 1624857261
transform 1 0 186841 0 1 142303
box 0 0 1 1
use contact_13  contact_13_921
timestamp 1624857261
transform 1 0 187177 0 1 142303
box 0 0 1 1
use contact_13  contact_13_920
timestamp 1624857261
transform 1 0 187513 0 1 142303
box 0 0 1 1
use contact_13  contact_13_919
timestamp 1624857261
transform 1 0 187849 0 1 142303
box 0 0 1 1
use contact_13  contact_13_918
timestamp 1624857261
transform 1 0 188185 0 1 142303
box 0 0 1 1
use contact_13  contact_13_917
timestamp 1624857261
transform 1 0 188521 0 1 142303
box 0 0 1 1
use contact_13  contact_13_916
timestamp 1624857261
transform 1 0 188857 0 1 142303
box 0 0 1 1
use contact_13  contact_13_915
timestamp 1624857261
transform 1 0 189193 0 1 142303
box 0 0 1 1
use contact_13  contact_13_914
timestamp 1624857261
transform 1 0 189529 0 1 142303
box 0 0 1 1
use contact_13  contact_13_913
timestamp 1624857261
transform 1 0 189865 0 1 142303
box 0 0 1 1
use contact_13  contact_13_912
timestamp 1624857261
transform 1 0 190201 0 1 142303
box 0 0 1 1
use contact_13  contact_13_911
timestamp 1624857261
transform 1 0 190537 0 1 142303
box 0 0 1 1
use contact_13  contact_13_910
timestamp 1624857261
transform 1 0 190873 0 1 142303
box 0 0 1 1
use contact_13  contact_13_909
timestamp 1624857261
transform 1 0 191209 0 1 142303
box 0 0 1 1
use contact_13  contact_13_908
timestamp 1624857261
transform 1 0 191545 0 1 142303
box 0 0 1 1
use contact_13  contact_13_907
timestamp 1624857261
transform 1 0 191881 0 1 142303
box 0 0 1 1
use contact_13  contact_13_906
timestamp 1624857261
transform 1 0 192217 0 1 142303
box 0 0 1 1
use contact_13  contact_13_905
timestamp 1624857261
transform 1 0 192553 0 1 142303
box 0 0 1 1
use contact_13  contact_13_904
timestamp 1624857261
transform 1 0 192889 0 1 142303
box 0 0 1 1
use contact_13  contact_13_903
timestamp 1624857261
transform 1 0 193225 0 1 142303
box 0 0 1 1
use contact_13  contact_13_902
timestamp 1624857261
transform 1 0 193561 0 1 142303
box 0 0 1 1
use contact_13  contact_13_901
timestamp 1624857261
transform 1 0 193897 0 1 142303
box 0 0 1 1
use contact_13  contact_13_900
timestamp 1624857261
transform 1 0 194233 0 1 142303
box 0 0 1 1
use contact_13  contact_13_899
timestamp 1624857261
transform 1 0 194569 0 1 142303
box 0 0 1 1
use contact_13  contact_13_898
timestamp 1624857261
transform 1 0 194905 0 1 142303
box 0 0 1 1
use contact_13  contact_13_897
timestamp 1624857261
transform 1 0 195241 0 1 142303
box 0 0 1 1
use contact_13  contact_13_896
timestamp 1624857261
transform 1 0 195577 0 1 142303
box 0 0 1 1
use contact_13  contact_13_895
timestamp 1624857261
transform 1 0 195913 0 1 142303
box 0 0 1 1
use contact_13  contact_13_894
timestamp 1624857261
transform 1 0 196249 0 1 142303
box 0 0 1 1
use contact_13  contact_13_893
timestamp 1624857261
transform 1 0 196585 0 1 142303
box 0 0 1 1
use contact_13  contact_13_892
timestamp 1624857261
transform 1 0 196921 0 1 142303
box 0 0 1 1
use contact_13  contact_13_891
timestamp 1624857261
transform 1 0 197257 0 1 142303
box 0 0 1 1
use contact_13  contact_13_890
timestamp 1624857261
transform 1 0 197593 0 1 142303
box 0 0 1 1
use contact_13  contact_13_889
timestamp 1624857261
transform 1 0 197929 0 1 142303
box 0 0 1 1
use contact_13  contact_13_888
timestamp 1624857261
transform 1 0 198265 0 1 142303
box 0 0 1 1
use contact_13  contact_13_887
timestamp 1624857261
transform 1 0 198601 0 1 142303
box 0 0 1 1
use contact_13  contact_13_886
timestamp 1624857261
transform 1 0 198937 0 1 142303
box 0 0 1 1
use contact_13  contact_13_885
timestamp 1624857261
transform 1 0 199273 0 1 142303
box 0 0 1 1
use contact_13  contact_13_884
timestamp 1624857261
transform 1 0 199609 0 1 142303
box 0 0 1 1
use contact_13  contact_13_883
timestamp 1624857261
transform 1 0 199945 0 1 142303
box 0 0 1 1
use contact_13  contact_13_882
timestamp 1624857261
transform 1 0 200281 0 1 142303
box 0 0 1 1
use contact_13  contact_13_881
timestamp 1624857261
transform 1 0 200617 0 1 142303
box 0 0 1 1
use contact_13  contact_13_880
timestamp 1624857261
transform 1 0 200953 0 1 142303
box 0 0 1 1
use contact_13  contact_13_879
timestamp 1624857261
transform 1 0 201289 0 1 142303
box 0 0 1 1
use contact_13  contact_13_878
timestamp 1624857261
transform 1 0 201625 0 1 142303
box 0 0 1 1
use contact_13  contact_13_877
timestamp 1624857261
transform 1 0 201961 0 1 142303
box 0 0 1 1
use contact_13  contact_13_876
timestamp 1624857261
transform 1 0 202297 0 1 142303
box 0 0 1 1
use contact_13  contact_13_875
timestamp 1624857261
transform 1 0 202633 0 1 142303
box 0 0 1 1
use contact_13  contact_13_874
timestamp 1624857261
transform 1 0 202969 0 1 142303
box 0 0 1 1
use contact_13  contact_13_873
timestamp 1624857261
transform 1 0 203305 0 1 142303
box 0 0 1 1
use contact_13  contact_13_872
timestamp 1624857261
transform 1 0 203641 0 1 142303
box 0 0 1 1
use contact_13  contact_13_871
timestamp 1624857261
transform 1 0 203977 0 1 142303
box 0 0 1 1
use contact_13  contact_13_870
timestamp 1624857261
transform 1 0 204313 0 1 142303
box 0 0 1 1
use contact_13  contact_13_869
timestamp 1624857261
transform 1 0 204649 0 1 142303
box 0 0 1 1
use contact_13  contact_13_868
timestamp 1624857261
transform 1 0 204985 0 1 142303
box 0 0 1 1
use contact_13  contact_13_867
timestamp 1624857261
transform 1 0 205321 0 1 142303
box 0 0 1 1
use contact_13  contact_13_866
timestamp 1624857261
transform 1 0 205657 0 1 142303
box 0 0 1 1
use contact_13  contact_13_865
timestamp 1624857261
transform 1 0 205993 0 1 142303
box 0 0 1 1
use contact_13  contact_13_864
timestamp 1624857261
transform 1 0 206329 0 1 142303
box 0 0 1 1
use contact_13  contact_13_863
timestamp 1624857261
transform 1 0 206665 0 1 142303
box 0 0 1 1
use contact_13  contact_13_862
timestamp 1624857261
transform 1 0 207001 0 1 142303
box 0 0 1 1
use contact_13  contact_13_861
timestamp 1624857261
transform 1 0 207337 0 1 142303
box 0 0 1 1
use contact_13  contact_13_860
timestamp 1624857261
transform 1 0 207673 0 1 142303
box 0 0 1 1
use contact_13  contact_13_859
timestamp 1624857261
transform 1 0 208009 0 1 142303
box 0 0 1 1
use contact_13  contact_13_858
timestamp 1624857261
transform 1 0 208345 0 1 142303
box 0 0 1 1
use contact_13  contact_13_857
timestamp 1624857261
transform 1 0 208681 0 1 142303
box 0 0 1 1
use contact_13  contact_13_856
timestamp 1624857261
transform 1 0 209017 0 1 142303
box 0 0 1 1
use contact_13  contact_13_855
timestamp 1624857261
transform 1 0 209353 0 1 142303
box 0 0 1 1
use contact_13  contact_13_854
timestamp 1624857261
transform 1 0 209689 0 1 142303
box 0 0 1 1
use contact_13  contact_13_853
timestamp 1624857261
transform 1 0 210025 0 1 142303
box 0 0 1 1
use contact_13  contact_13_852
timestamp 1624857261
transform 1 0 210361 0 1 142303
box 0 0 1 1
use contact_13  contact_13_851
timestamp 1624857261
transform 1 0 210697 0 1 142303
box 0 0 1 1
use contact_13  contact_13_850
timestamp 1624857261
transform 1 0 211033 0 1 142303
box 0 0 1 1
use contact_13  contact_13_849
timestamp 1624857261
transform 1 0 211369 0 1 142303
box 0 0 1 1
use contact_13  contact_13_848
timestamp 1624857261
transform 1 0 211705 0 1 142303
box 0 0 1 1
use contact_13  contact_13_847
timestamp 1624857261
transform 1 0 212041 0 1 142303
box 0 0 1 1
use contact_13  contact_13_846
timestamp 1624857261
transform 1 0 212377 0 1 142303
box 0 0 1 1
use contact_13  contact_13_845
timestamp 1624857261
transform 1 0 212713 0 1 142303
box 0 0 1 1
use contact_13  contact_13_844
timestamp 1624857261
transform 1 0 213049 0 1 142303
box 0 0 1 1
use contact_13  contact_13_843
timestamp 1624857261
transform 1 0 213385 0 1 142303
box 0 0 1 1
use contact_13  contact_13_842
timestamp 1624857261
transform 1 0 213721 0 1 142303
box 0 0 1 1
use contact_13  contact_13_841
timestamp 1624857261
transform 1 0 214057 0 1 142303
box 0 0 1 1
use contact_13  contact_13_840
timestamp 1624857261
transform 1 0 214393 0 1 142303
box 0 0 1 1
use contact_13  contact_13_839
timestamp 1624857261
transform 1 0 214729 0 1 142303
box 0 0 1 1
use contact_13  contact_13_838
timestamp 1624857261
transform 1 0 215065 0 1 142303
box 0 0 1 1
use contact_13  contact_13_837
timestamp 1624857261
transform 1 0 215401 0 1 142303
box 0 0 1 1
use contact_13  contact_13_836
timestamp 1624857261
transform 1 0 215737 0 1 142303
box 0 0 1 1
use contact_13  contact_13_835
timestamp 1624857261
transform 1 0 216073 0 1 142303
box 0 0 1 1
use contact_13  contact_13_834
timestamp 1624857261
transform 1 0 216409 0 1 142303
box 0 0 1 1
use contact_13  contact_13_833
timestamp 1624857261
transform 1 0 1705 0 1 2143
box 0 0 1 1
use contact_13  contact_13_832
timestamp 1624857261
transform 1 0 1705 0 1 2479
box 0 0 1 1
use contact_13  contact_13_831
timestamp 1624857261
transform 1 0 1705 0 1 2815
box 0 0 1 1
use contact_13  contact_13_830
timestamp 1624857261
transform 1 0 1705 0 1 3151
box 0 0 1 1
use contact_13  contact_13_829
timestamp 1624857261
transform 1 0 1705 0 1 3487
box 0 0 1 1
use contact_13  contact_13_828
timestamp 1624857261
transform 1 0 1705 0 1 3823
box 0 0 1 1
use contact_13  contact_13_827
timestamp 1624857261
transform 1 0 1705 0 1 4159
box 0 0 1 1
use contact_13  contact_13_826
timestamp 1624857261
transform 1 0 1705 0 1 4495
box 0 0 1 1
use contact_13  contact_13_825
timestamp 1624857261
transform 1 0 1705 0 1 4831
box 0 0 1 1
use contact_13  contact_13_824
timestamp 1624857261
transform 1 0 1705 0 1 5167
box 0 0 1 1
use contact_13  contact_13_823
timestamp 1624857261
transform 1 0 1705 0 1 5503
box 0 0 1 1
use contact_13  contact_13_822
timestamp 1624857261
transform 1 0 1705 0 1 5839
box 0 0 1 1
use contact_13  contact_13_821
timestamp 1624857261
transform 1 0 1705 0 1 6175
box 0 0 1 1
use contact_13  contact_13_820
timestamp 1624857261
transform 1 0 1705 0 1 6511
box 0 0 1 1
use contact_13  contact_13_819
timestamp 1624857261
transform 1 0 1705 0 1 6847
box 0 0 1 1
use contact_13  contact_13_818
timestamp 1624857261
transform 1 0 1705 0 1 7183
box 0 0 1 1
use contact_13  contact_13_817
timestamp 1624857261
transform 1 0 1705 0 1 7519
box 0 0 1 1
use contact_13  contact_13_816
timestamp 1624857261
transform 1 0 1705 0 1 7855
box 0 0 1 1
use contact_13  contact_13_815
timestamp 1624857261
transform 1 0 1705 0 1 8191
box 0 0 1 1
use contact_13  contact_13_814
timestamp 1624857261
transform 1 0 1705 0 1 8527
box 0 0 1 1
use contact_13  contact_13_813
timestamp 1624857261
transform 1 0 1705 0 1 8863
box 0 0 1 1
use contact_13  contact_13_812
timestamp 1624857261
transform 1 0 1705 0 1 9199
box 0 0 1 1
use contact_13  contact_13_811
timestamp 1624857261
transform 1 0 1705 0 1 9535
box 0 0 1 1
use contact_13  contact_13_810
timestamp 1624857261
transform 1 0 1705 0 1 9871
box 0 0 1 1
use contact_13  contact_13_809
timestamp 1624857261
transform 1 0 1705 0 1 10207
box 0 0 1 1
use contact_13  contact_13_808
timestamp 1624857261
transform 1 0 1705 0 1 10543
box 0 0 1 1
use contact_13  contact_13_807
timestamp 1624857261
transform 1 0 1705 0 1 10879
box 0 0 1 1
use contact_13  contact_13_806
timestamp 1624857261
transform 1 0 1705 0 1 11215
box 0 0 1 1
use contact_13  contact_13_805
timestamp 1624857261
transform 1 0 1705 0 1 11551
box 0 0 1 1
use contact_13  contact_13_804
timestamp 1624857261
transform 1 0 1705 0 1 11887
box 0 0 1 1
use contact_13  contact_13_803
timestamp 1624857261
transform 1 0 1705 0 1 12223
box 0 0 1 1
use contact_13  contact_13_802
timestamp 1624857261
transform 1 0 1705 0 1 12559
box 0 0 1 1
use contact_13  contact_13_801
timestamp 1624857261
transform 1 0 1705 0 1 12895
box 0 0 1 1
use contact_13  contact_13_800
timestamp 1624857261
transform 1 0 1705 0 1 13231
box 0 0 1 1
use contact_13  contact_13_799
timestamp 1624857261
transform 1 0 1705 0 1 13567
box 0 0 1 1
use contact_13  contact_13_798
timestamp 1624857261
transform 1 0 1705 0 1 13903
box 0 0 1 1
use contact_13  contact_13_797
timestamp 1624857261
transform 1 0 1705 0 1 14239
box 0 0 1 1
use contact_13  contact_13_796
timestamp 1624857261
transform 1 0 1705 0 1 14575
box 0 0 1 1
use contact_13  contact_13_795
timestamp 1624857261
transform 1 0 1705 0 1 14911
box 0 0 1 1
use contact_13  contact_13_794
timestamp 1624857261
transform 1 0 1705 0 1 15247
box 0 0 1 1
use contact_13  contact_13_793
timestamp 1624857261
transform 1 0 1705 0 1 15583
box 0 0 1 1
use contact_13  contact_13_792
timestamp 1624857261
transform 1 0 1705 0 1 15919
box 0 0 1 1
use contact_13  contact_13_791
timestamp 1624857261
transform 1 0 1705 0 1 16255
box 0 0 1 1
use contact_13  contact_13_790
timestamp 1624857261
transform 1 0 1705 0 1 16591
box 0 0 1 1
use contact_13  contact_13_789
timestamp 1624857261
transform 1 0 1705 0 1 16927
box 0 0 1 1
use contact_13  contact_13_788
timestamp 1624857261
transform 1 0 1705 0 1 17263
box 0 0 1 1
use contact_13  contact_13_787
timestamp 1624857261
transform 1 0 1705 0 1 17599
box 0 0 1 1
use contact_13  contact_13_786
timestamp 1624857261
transform 1 0 1705 0 1 17935
box 0 0 1 1
use contact_13  contact_13_785
timestamp 1624857261
transform 1 0 1705 0 1 18271
box 0 0 1 1
use contact_13  contact_13_784
timestamp 1624857261
transform 1 0 1705 0 1 18607
box 0 0 1 1
use contact_13  contact_13_783
timestamp 1624857261
transform 1 0 1705 0 1 18943
box 0 0 1 1
use contact_13  contact_13_782
timestamp 1624857261
transform 1 0 1705 0 1 19279
box 0 0 1 1
use contact_13  contact_13_781
timestamp 1624857261
transform 1 0 1705 0 1 19615
box 0 0 1 1
use contact_13  contact_13_780
timestamp 1624857261
transform 1 0 1705 0 1 19951
box 0 0 1 1
use contact_13  contact_13_779
timestamp 1624857261
transform 1 0 1705 0 1 20287
box 0 0 1 1
use contact_13  contact_13_778
timestamp 1624857261
transform 1 0 1705 0 1 20623
box 0 0 1 1
use contact_13  contact_13_777
timestamp 1624857261
transform 1 0 1705 0 1 20959
box 0 0 1 1
use contact_13  contact_13_776
timestamp 1624857261
transform 1 0 1705 0 1 21295
box 0 0 1 1
use contact_13  contact_13_775
timestamp 1624857261
transform 1 0 1705 0 1 21631
box 0 0 1 1
use contact_13  contact_13_774
timestamp 1624857261
transform 1 0 1705 0 1 21967
box 0 0 1 1
use contact_13  contact_13_773
timestamp 1624857261
transform 1 0 1705 0 1 22303
box 0 0 1 1
use contact_13  contact_13_772
timestamp 1624857261
transform 1 0 1705 0 1 22639
box 0 0 1 1
use contact_13  contact_13_771
timestamp 1624857261
transform 1 0 1705 0 1 22975
box 0 0 1 1
use contact_13  contact_13_770
timestamp 1624857261
transform 1 0 1705 0 1 23311
box 0 0 1 1
use contact_13  contact_13_769
timestamp 1624857261
transform 1 0 1705 0 1 23647
box 0 0 1 1
use contact_13  contact_13_768
timestamp 1624857261
transform 1 0 1705 0 1 23983
box 0 0 1 1
use contact_13  contact_13_767
timestamp 1624857261
transform 1 0 1705 0 1 24319
box 0 0 1 1
use contact_13  contact_13_766
timestamp 1624857261
transform 1 0 1705 0 1 24655
box 0 0 1 1
use contact_13  contact_13_765
timestamp 1624857261
transform 1 0 1705 0 1 24991
box 0 0 1 1
use contact_13  contact_13_764
timestamp 1624857261
transform 1 0 1705 0 1 25327
box 0 0 1 1
use contact_13  contact_13_763
timestamp 1624857261
transform 1 0 1705 0 1 25663
box 0 0 1 1
use contact_13  contact_13_762
timestamp 1624857261
transform 1 0 1705 0 1 25999
box 0 0 1 1
use contact_13  contact_13_761
timestamp 1624857261
transform 1 0 1705 0 1 26335
box 0 0 1 1
use contact_13  contact_13_760
timestamp 1624857261
transform 1 0 1705 0 1 26671
box 0 0 1 1
use contact_13  contact_13_759
timestamp 1624857261
transform 1 0 1705 0 1 27007
box 0 0 1 1
use contact_13  contact_13_758
timestamp 1624857261
transform 1 0 1705 0 1 27343
box 0 0 1 1
use contact_13  contact_13_757
timestamp 1624857261
transform 1 0 1705 0 1 27679
box 0 0 1 1
use contact_13  contact_13_756
timestamp 1624857261
transform 1 0 1705 0 1 28015
box 0 0 1 1
use contact_13  contact_13_755
timestamp 1624857261
transform 1 0 1705 0 1 28351
box 0 0 1 1
use contact_13  contact_13_754
timestamp 1624857261
transform 1 0 1705 0 1 28687
box 0 0 1 1
use contact_13  contact_13_753
timestamp 1624857261
transform 1 0 1705 0 1 29023
box 0 0 1 1
use contact_13  contact_13_752
timestamp 1624857261
transform 1 0 1705 0 1 29359
box 0 0 1 1
use contact_13  contact_13_751
timestamp 1624857261
transform 1 0 1705 0 1 29695
box 0 0 1 1
use contact_13  contact_13_750
timestamp 1624857261
transform 1 0 1705 0 1 30031
box 0 0 1 1
use contact_13  contact_13_749
timestamp 1624857261
transform 1 0 1705 0 1 30367
box 0 0 1 1
use contact_13  contact_13_748
timestamp 1624857261
transform 1 0 1705 0 1 30703
box 0 0 1 1
use contact_13  contact_13_747
timestamp 1624857261
transform 1 0 1705 0 1 31039
box 0 0 1 1
use contact_13  contact_13_746
timestamp 1624857261
transform 1 0 1705 0 1 31375
box 0 0 1 1
use contact_13  contact_13_745
timestamp 1624857261
transform 1 0 1705 0 1 31711
box 0 0 1 1
use contact_13  contact_13_744
timestamp 1624857261
transform 1 0 1705 0 1 32047
box 0 0 1 1
use contact_13  contact_13_743
timestamp 1624857261
transform 1 0 1705 0 1 32383
box 0 0 1 1
use contact_13  contact_13_742
timestamp 1624857261
transform 1 0 1705 0 1 32719
box 0 0 1 1
use contact_13  contact_13_741
timestamp 1624857261
transform 1 0 1705 0 1 33055
box 0 0 1 1
use contact_13  contact_13_740
timestamp 1624857261
transform 1 0 1705 0 1 33391
box 0 0 1 1
use contact_13  contact_13_739
timestamp 1624857261
transform 1 0 1705 0 1 33727
box 0 0 1 1
use contact_13  contact_13_738
timestamp 1624857261
transform 1 0 1705 0 1 34063
box 0 0 1 1
use contact_13  contact_13_737
timestamp 1624857261
transform 1 0 1705 0 1 34399
box 0 0 1 1
use contact_13  contact_13_736
timestamp 1624857261
transform 1 0 1705 0 1 34735
box 0 0 1 1
use contact_13  contact_13_735
timestamp 1624857261
transform 1 0 1705 0 1 35071
box 0 0 1 1
use contact_13  contact_13_734
timestamp 1624857261
transform 1 0 1705 0 1 35407
box 0 0 1 1
use contact_13  contact_13_733
timestamp 1624857261
transform 1 0 1705 0 1 35743
box 0 0 1 1
use contact_13  contact_13_732
timestamp 1624857261
transform 1 0 1705 0 1 36079
box 0 0 1 1
use contact_13  contact_13_731
timestamp 1624857261
transform 1 0 1705 0 1 36415
box 0 0 1 1
use contact_13  contact_13_730
timestamp 1624857261
transform 1 0 1705 0 1 36751
box 0 0 1 1
use contact_13  contact_13_729
timestamp 1624857261
transform 1 0 1705 0 1 37087
box 0 0 1 1
use contact_13  contact_13_728
timestamp 1624857261
transform 1 0 1705 0 1 37423
box 0 0 1 1
use contact_13  contact_13_727
timestamp 1624857261
transform 1 0 1705 0 1 37759
box 0 0 1 1
use contact_13  contact_13_726
timestamp 1624857261
transform 1 0 1705 0 1 38095
box 0 0 1 1
use contact_13  contact_13_725
timestamp 1624857261
transform 1 0 1705 0 1 38431
box 0 0 1 1
use contact_13  contact_13_724
timestamp 1624857261
transform 1 0 1705 0 1 38767
box 0 0 1 1
use contact_13  contact_13_723
timestamp 1624857261
transform 1 0 1705 0 1 39103
box 0 0 1 1
use contact_13  contact_13_722
timestamp 1624857261
transform 1 0 1705 0 1 39439
box 0 0 1 1
use contact_13  contact_13_721
timestamp 1624857261
transform 1 0 1705 0 1 39775
box 0 0 1 1
use contact_13  contact_13_720
timestamp 1624857261
transform 1 0 1705 0 1 40111
box 0 0 1 1
use contact_13  contact_13_719
timestamp 1624857261
transform 1 0 1705 0 1 40447
box 0 0 1 1
use contact_13  contact_13_718
timestamp 1624857261
transform 1 0 1705 0 1 40783
box 0 0 1 1
use contact_13  contact_13_717
timestamp 1624857261
transform 1 0 1705 0 1 41119
box 0 0 1 1
use contact_13  contact_13_716
timestamp 1624857261
transform 1 0 1705 0 1 41455
box 0 0 1 1
use contact_13  contact_13_715
timestamp 1624857261
transform 1 0 1705 0 1 41791
box 0 0 1 1
use contact_13  contact_13_714
timestamp 1624857261
transform 1 0 1705 0 1 42127
box 0 0 1 1
use contact_13  contact_13_713
timestamp 1624857261
transform 1 0 1705 0 1 42463
box 0 0 1 1
use contact_13  contact_13_712
timestamp 1624857261
transform 1 0 1705 0 1 42799
box 0 0 1 1
use contact_13  contact_13_711
timestamp 1624857261
transform 1 0 1705 0 1 43135
box 0 0 1 1
use contact_13  contact_13_710
timestamp 1624857261
transform 1 0 1705 0 1 43471
box 0 0 1 1
use contact_13  contact_13_709
timestamp 1624857261
transform 1 0 1705 0 1 43807
box 0 0 1 1
use contact_13  contact_13_708
timestamp 1624857261
transform 1 0 1705 0 1 44143
box 0 0 1 1
use contact_13  contact_13_707
timestamp 1624857261
transform 1 0 1705 0 1 44479
box 0 0 1 1
use contact_13  contact_13_706
timestamp 1624857261
transform 1 0 1705 0 1 44815
box 0 0 1 1
use contact_13  contact_13_705
timestamp 1624857261
transform 1 0 1705 0 1 45151
box 0 0 1 1
use contact_13  contact_13_704
timestamp 1624857261
transform 1 0 1705 0 1 45487
box 0 0 1 1
use contact_13  contact_13_703
timestamp 1624857261
transform 1 0 1705 0 1 45823
box 0 0 1 1
use contact_13  contact_13_702
timestamp 1624857261
transform 1 0 1705 0 1 46159
box 0 0 1 1
use contact_13  contact_13_701
timestamp 1624857261
transform 1 0 1705 0 1 46495
box 0 0 1 1
use contact_13  contact_13_700
timestamp 1624857261
transform 1 0 1705 0 1 46831
box 0 0 1 1
use contact_13  contact_13_699
timestamp 1624857261
transform 1 0 1705 0 1 47167
box 0 0 1 1
use contact_13  contact_13_698
timestamp 1624857261
transform 1 0 1705 0 1 47503
box 0 0 1 1
use contact_13  contact_13_697
timestamp 1624857261
transform 1 0 1705 0 1 47839
box 0 0 1 1
use contact_13  contact_13_696
timestamp 1624857261
transform 1 0 1705 0 1 48175
box 0 0 1 1
use contact_13  contact_13_695
timestamp 1624857261
transform 1 0 1705 0 1 48511
box 0 0 1 1
use contact_13  contact_13_694
timestamp 1624857261
transform 1 0 1705 0 1 48847
box 0 0 1 1
use contact_13  contact_13_693
timestamp 1624857261
transform 1 0 1705 0 1 49183
box 0 0 1 1
use contact_13  contact_13_692
timestamp 1624857261
transform 1 0 1705 0 1 49519
box 0 0 1 1
use contact_13  contact_13_691
timestamp 1624857261
transform 1 0 1705 0 1 49855
box 0 0 1 1
use contact_13  contact_13_690
timestamp 1624857261
transform 1 0 1705 0 1 50191
box 0 0 1 1
use contact_13  contact_13_689
timestamp 1624857261
transform 1 0 1705 0 1 50527
box 0 0 1 1
use contact_13  contact_13_688
timestamp 1624857261
transform 1 0 1705 0 1 50863
box 0 0 1 1
use contact_13  contact_13_687
timestamp 1624857261
transform 1 0 1705 0 1 51199
box 0 0 1 1
use contact_13  contact_13_686
timestamp 1624857261
transform 1 0 1705 0 1 51535
box 0 0 1 1
use contact_13  contact_13_685
timestamp 1624857261
transform 1 0 1705 0 1 51871
box 0 0 1 1
use contact_13  contact_13_684
timestamp 1624857261
transform 1 0 1705 0 1 52207
box 0 0 1 1
use contact_13  contact_13_683
timestamp 1624857261
transform 1 0 1705 0 1 52543
box 0 0 1 1
use contact_13  contact_13_682
timestamp 1624857261
transform 1 0 1705 0 1 52879
box 0 0 1 1
use contact_13  contact_13_681
timestamp 1624857261
transform 1 0 1705 0 1 53215
box 0 0 1 1
use contact_13  contact_13_680
timestamp 1624857261
transform 1 0 1705 0 1 53551
box 0 0 1 1
use contact_13  contact_13_679
timestamp 1624857261
transform 1 0 1705 0 1 53887
box 0 0 1 1
use contact_13  contact_13_678
timestamp 1624857261
transform 1 0 1705 0 1 54223
box 0 0 1 1
use contact_13  contact_13_677
timestamp 1624857261
transform 1 0 1705 0 1 54559
box 0 0 1 1
use contact_13  contact_13_676
timestamp 1624857261
transform 1 0 1705 0 1 54895
box 0 0 1 1
use contact_13  contact_13_675
timestamp 1624857261
transform 1 0 1705 0 1 55231
box 0 0 1 1
use contact_13  contact_13_674
timestamp 1624857261
transform 1 0 1705 0 1 55567
box 0 0 1 1
use contact_13  contact_13_673
timestamp 1624857261
transform 1 0 1705 0 1 55903
box 0 0 1 1
use contact_13  contact_13_672
timestamp 1624857261
transform 1 0 1705 0 1 56239
box 0 0 1 1
use contact_13  contact_13_671
timestamp 1624857261
transform 1 0 1705 0 1 56575
box 0 0 1 1
use contact_13  contact_13_670
timestamp 1624857261
transform 1 0 1705 0 1 56911
box 0 0 1 1
use contact_13  contact_13_669
timestamp 1624857261
transform 1 0 1705 0 1 57247
box 0 0 1 1
use contact_13  contact_13_668
timestamp 1624857261
transform 1 0 1705 0 1 57583
box 0 0 1 1
use contact_13  contact_13_667
timestamp 1624857261
transform 1 0 1705 0 1 57919
box 0 0 1 1
use contact_13  contact_13_666
timestamp 1624857261
transform 1 0 1705 0 1 58255
box 0 0 1 1
use contact_13  contact_13_665
timestamp 1624857261
transform 1 0 1705 0 1 58591
box 0 0 1 1
use contact_13  contact_13_664
timestamp 1624857261
transform 1 0 1705 0 1 58927
box 0 0 1 1
use contact_13  contact_13_663
timestamp 1624857261
transform 1 0 1705 0 1 59263
box 0 0 1 1
use contact_13  contact_13_662
timestamp 1624857261
transform 1 0 1705 0 1 59599
box 0 0 1 1
use contact_13  contact_13_661
timestamp 1624857261
transform 1 0 1705 0 1 59935
box 0 0 1 1
use contact_13  contact_13_660
timestamp 1624857261
transform 1 0 1705 0 1 60271
box 0 0 1 1
use contact_13  contact_13_659
timestamp 1624857261
transform 1 0 1705 0 1 60607
box 0 0 1 1
use contact_13  contact_13_658
timestamp 1624857261
transform 1 0 1705 0 1 60943
box 0 0 1 1
use contact_13  contact_13_657
timestamp 1624857261
transform 1 0 1705 0 1 61279
box 0 0 1 1
use contact_13  contact_13_656
timestamp 1624857261
transform 1 0 1705 0 1 61615
box 0 0 1 1
use contact_13  contact_13_655
timestamp 1624857261
transform 1 0 1705 0 1 61951
box 0 0 1 1
use contact_13  contact_13_654
timestamp 1624857261
transform 1 0 1705 0 1 62287
box 0 0 1 1
use contact_13  contact_13_653
timestamp 1624857261
transform 1 0 1705 0 1 62623
box 0 0 1 1
use contact_13  contact_13_652
timestamp 1624857261
transform 1 0 1705 0 1 62959
box 0 0 1 1
use contact_13  contact_13_651
timestamp 1624857261
transform 1 0 1705 0 1 63295
box 0 0 1 1
use contact_13  contact_13_650
timestamp 1624857261
transform 1 0 1705 0 1 63631
box 0 0 1 1
use contact_13  contact_13_649
timestamp 1624857261
transform 1 0 1705 0 1 63967
box 0 0 1 1
use contact_13  contact_13_648
timestamp 1624857261
transform 1 0 1705 0 1 64303
box 0 0 1 1
use contact_13  contact_13_647
timestamp 1624857261
transform 1 0 1705 0 1 64639
box 0 0 1 1
use contact_13  contact_13_646
timestamp 1624857261
transform 1 0 1705 0 1 64975
box 0 0 1 1
use contact_13  contact_13_645
timestamp 1624857261
transform 1 0 1705 0 1 65311
box 0 0 1 1
use contact_13  contact_13_644
timestamp 1624857261
transform 1 0 1705 0 1 65647
box 0 0 1 1
use contact_13  contact_13_643
timestamp 1624857261
transform 1 0 1705 0 1 65983
box 0 0 1 1
use contact_13  contact_13_642
timestamp 1624857261
transform 1 0 1705 0 1 66319
box 0 0 1 1
use contact_13  contact_13_641
timestamp 1624857261
transform 1 0 1705 0 1 66655
box 0 0 1 1
use contact_13  contact_13_640
timestamp 1624857261
transform 1 0 1705 0 1 66991
box 0 0 1 1
use contact_13  contact_13_639
timestamp 1624857261
transform 1 0 1705 0 1 67327
box 0 0 1 1
use contact_13  contact_13_638
timestamp 1624857261
transform 1 0 1705 0 1 67663
box 0 0 1 1
use contact_13  contact_13_637
timestamp 1624857261
transform 1 0 1705 0 1 67999
box 0 0 1 1
use contact_13  contact_13_636
timestamp 1624857261
transform 1 0 1705 0 1 68335
box 0 0 1 1
use contact_13  contact_13_635
timestamp 1624857261
transform 1 0 1705 0 1 68671
box 0 0 1 1
use contact_13  contact_13_634
timestamp 1624857261
transform 1 0 1705 0 1 69007
box 0 0 1 1
use contact_13  contact_13_633
timestamp 1624857261
transform 1 0 1705 0 1 69343
box 0 0 1 1
use contact_13  contact_13_632
timestamp 1624857261
transform 1 0 1705 0 1 69679
box 0 0 1 1
use contact_13  contact_13_631
timestamp 1624857261
transform 1 0 1705 0 1 70015
box 0 0 1 1
use contact_13  contact_13_630
timestamp 1624857261
transform 1 0 1705 0 1 70351
box 0 0 1 1
use contact_13  contact_13_629
timestamp 1624857261
transform 1 0 1705 0 1 70687
box 0 0 1 1
use contact_13  contact_13_628
timestamp 1624857261
transform 1 0 1705 0 1 71023
box 0 0 1 1
use contact_13  contact_13_627
timestamp 1624857261
transform 1 0 1705 0 1 71359
box 0 0 1 1
use contact_13  contact_13_626
timestamp 1624857261
transform 1 0 1705 0 1 71695
box 0 0 1 1
use contact_13  contact_13_625
timestamp 1624857261
transform 1 0 1705 0 1 72031
box 0 0 1 1
use contact_13  contact_13_624
timestamp 1624857261
transform 1 0 1705 0 1 72367
box 0 0 1 1
use contact_13  contact_13_623
timestamp 1624857261
transform 1 0 1705 0 1 72703
box 0 0 1 1
use contact_13  contact_13_622
timestamp 1624857261
transform 1 0 1705 0 1 73039
box 0 0 1 1
use contact_13  contact_13_621
timestamp 1624857261
transform 1 0 1705 0 1 73375
box 0 0 1 1
use contact_13  contact_13_620
timestamp 1624857261
transform 1 0 1705 0 1 73711
box 0 0 1 1
use contact_13  contact_13_619
timestamp 1624857261
transform 1 0 1705 0 1 74047
box 0 0 1 1
use contact_13  contact_13_618
timestamp 1624857261
transform 1 0 1705 0 1 74383
box 0 0 1 1
use contact_13  contact_13_617
timestamp 1624857261
transform 1 0 1705 0 1 74719
box 0 0 1 1
use contact_13  contact_13_616
timestamp 1624857261
transform 1 0 1705 0 1 75055
box 0 0 1 1
use contact_13  contact_13_615
timestamp 1624857261
transform 1 0 1705 0 1 75391
box 0 0 1 1
use contact_13  contact_13_614
timestamp 1624857261
transform 1 0 1705 0 1 75727
box 0 0 1 1
use contact_13  contact_13_613
timestamp 1624857261
transform 1 0 1705 0 1 76063
box 0 0 1 1
use contact_13  contact_13_612
timestamp 1624857261
transform 1 0 1705 0 1 76399
box 0 0 1 1
use contact_13  contact_13_611
timestamp 1624857261
transform 1 0 1705 0 1 76735
box 0 0 1 1
use contact_13  contact_13_610
timestamp 1624857261
transform 1 0 1705 0 1 77071
box 0 0 1 1
use contact_13  contact_13_609
timestamp 1624857261
transform 1 0 1705 0 1 77407
box 0 0 1 1
use contact_13  contact_13_608
timestamp 1624857261
transform 1 0 1705 0 1 77743
box 0 0 1 1
use contact_13  contact_13_607
timestamp 1624857261
transform 1 0 1705 0 1 78079
box 0 0 1 1
use contact_13  contact_13_606
timestamp 1624857261
transform 1 0 1705 0 1 78415
box 0 0 1 1
use contact_13  contact_13_605
timestamp 1624857261
transform 1 0 1705 0 1 78751
box 0 0 1 1
use contact_13  contact_13_604
timestamp 1624857261
transform 1 0 1705 0 1 79087
box 0 0 1 1
use contact_13  contact_13_603
timestamp 1624857261
transform 1 0 1705 0 1 79423
box 0 0 1 1
use contact_13  contact_13_602
timestamp 1624857261
transform 1 0 1705 0 1 79759
box 0 0 1 1
use contact_13  contact_13_601
timestamp 1624857261
transform 1 0 1705 0 1 80095
box 0 0 1 1
use contact_13  contact_13_600
timestamp 1624857261
transform 1 0 1705 0 1 80431
box 0 0 1 1
use contact_13  contact_13_599
timestamp 1624857261
transform 1 0 1705 0 1 80767
box 0 0 1 1
use contact_13  contact_13_598
timestamp 1624857261
transform 1 0 1705 0 1 81103
box 0 0 1 1
use contact_13  contact_13_597
timestamp 1624857261
transform 1 0 1705 0 1 81439
box 0 0 1 1
use contact_13  contact_13_596
timestamp 1624857261
transform 1 0 1705 0 1 81775
box 0 0 1 1
use contact_13  contact_13_595
timestamp 1624857261
transform 1 0 1705 0 1 82111
box 0 0 1 1
use contact_13  contact_13_594
timestamp 1624857261
transform 1 0 1705 0 1 82447
box 0 0 1 1
use contact_13  contact_13_593
timestamp 1624857261
transform 1 0 1705 0 1 82783
box 0 0 1 1
use contact_13  contact_13_592
timestamp 1624857261
transform 1 0 1705 0 1 83119
box 0 0 1 1
use contact_13  contact_13_591
timestamp 1624857261
transform 1 0 1705 0 1 83455
box 0 0 1 1
use contact_13  contact_13_590
timestamp 1624857261
transform 1 0 1705 0 1 83791
box 0 0 1 1
use contact_13  contact_13_589
timestamp 1624857261
transform 1 0 1705 0 1 84127
box 0 0 1 1
use contact_13  contact_13_588
timestamp 1624857261
transform 1 0 1705 0 1 84463
box 0 0 1 1
use contact_13  contact_13_587
timestamp 1624857261
transform 1 0 1705 0 1 84799
box 0 0 1 1
use contact_13  contact_13_586
timestamp 1624857261
transform 1 0 1705 0 1 85135
box 0 0 1 1
use contact_13  contact_13_585
timestamp 1624857261
transform 1 0 1705 0 1 85471
box 0 0 1 1
use contact_13  contact_13_584
timestamp 1624857261
transform 1 0 1705 0 1 85807
box 0 0 1 1
use contact_13  contact_13_583
timestamp 1624857261
transform 1 0 1705 0 1 86143
box 0 0 1 1
use contact_13  contact_13_582
timestamp 1624857261
transform 1 0 1705 0 1 86479
box 0 0 1 1
use contact_13  contact_13_581
timestamp 1624857261
transform 1 0 1705 0 1 86815
box 0 0 1 1
use contact_13  contact_13_580
timestamp 1624857261
transform 1 0 1705 0 1 87151
box 0 0 1 1
use contact_13  contact_13_579
timestamp 1624857261
transform 1 0 1705 0 1 87487
box 0 0 1 1
use contact_13  contact_13_578
timestamp 1624857261
transform 1 0 1705 0 1 87823
box 0 0 1 1
use contact_13  contact_13_577
timestamp 1624857261
transform 1 0 1705 0 1 88159
box 0 0 1 1
use contact_13  contact_13_576
timestamp 1624857261
transform 1 0 1705 0 1 88495
box 0 0 1 1
use contact_13  contact_13_575
timestamp 1624857261
transform 1 0 1705 0 1 88831
box 0 0 1 1
use contact_13  contact_13_574
timestamp 1624857261
transform 1 0 1705 0 1 89167
box 0 0 1 1
use contact_13  contact_13_573
timestamp 1624857261
transform 1 0 1705 0 1 89503
box 0 0 1 1
use contact_13  contact_13_572
timestamp 1624857261
transform 1 0 1705 0 1 89839
box 0 0 1 1
use contact_13  contact_13_571
timestamp 1624857261
transform 1 0 1705 0 1 90175
box 0 0 1 1
use contact_13  contact_13_570
timestamp 1624857261
transform 1 0 1705 0 1 90511
box 0 0 1 1
use contact_13  contact_13_569
timestamp 1624857261
transform 1 0 1705 0 1 90847
box 0 0 1 1
use contact_13  contact_13_568
timestamp 1624857261
transform 1 0 1705 0 1 91183
box 0 0 1 1
use contact_13  contact_13_567
timestamp 1624857261
transform 1 0 1705 0 1 91519
box 0 0 1 1
use contact_13  contact_13_566
timestamp 1624857261
transform 1 0 1705 0 1 91855
box 0 0 1 1
use contact_13  contact_13_565
timestamp 1624857261
transform 1 0 1705 0 1 92191
box 0 0 1 1
use contact_13  contact_13_564
timestamp 1624857261
transform 1 0 1705 0 1 92527
box 0 0 1 1
use contact_13  contact_13_563
timestamp 1624857261
transform 1 0 1705 0 1 92863
box 0 0 1 1
use contact_13  contact_13_562
timestamp 1624857261
transform 1 0 1705 0 1 93199
box 0 0 1 1
use contact_13  contact_13_561
timestamp 1624857261
transform 1 0 1705 0 1 93535
box 0 0 1 1
use contact_13  contact_13_560
timestamp 1624857261
transform 1 0 1705 0 1 93871
box 0 0 1 1
use contact_13  contact_13_559
timestamp 1624857261
transform 1 0 1705 0 1 94207
box 0 0 1 1
use contact_13  contact_13_558
timestamp 1624857261
transform 1 0 1705 0 1 94543
box 0 0 1 1
use contact_13  contact_13_557
timestamp 1624857261
transform 1 0 1705 0 1 94879
box 0 0 1 1
use contact_13  contact_13_556
timestamp 1624857261
transform 1 0 1705 0 1 95215
box 0 0 1 1
use contact_13  contact_13_555
timestamp 1624857261
transform 1 0 1705 0 1 95551
box 0 0 1 1
use contact_13  contact_13_554
timestamp 1624857261
transform 1 0 1705 0 1 95887
box 0 0 1 1
use contact_13  contact_13_553
timestamp 1624857261
transform 1 0 1705 0 1 96223
box 0 0 1 1
use contact_13  contact_13_552
timestamp 1624857261
transform 1 0 1705 0 1 96559
box 0 0 1 1
use contact_13  contact_13_551
timestamp 1624857261
transform 1 0 1705 0 1 96895
box 0 0 1 1
use contact_13  contact_13_550
timestamp 1624857261
transform 1 0 1705 0 1 97231
box 0 0 1 1
use contact_13  contact_13_549
timestamp 1624857261
transform 1 0 1705 0 1 97567
box 0 0 1 1
use contact_13  contact_13_548
timestamp 1624857261
transform 1 0 1705 0 1 97903
box 0 0 1 1
use contact_13  contact_13_547
timestamp 1624857261
transform 1 0 1705 0 1 98239
box 0 0 1 1
use contact_13  contact_13_546
timestamp 1624857261
transform 1 0 1705 0 1 98575
box 0 0 1 1
use contact_13  contact_13_545
timestamp 1624857261
transform 1 0 1705 0 1 98911
box 0 0 1 1
use contact_13  contact_13_544
timestamp 1624857261
transform 1 0 1705 0 1 99247
box 0 0 1 1
use contact_13  contact_13_543
timestamp 1624857261
transform 1 0 1705 0 1 99583
box 0 0 1 1
use contact_13  contact_13_542
timestamp 1624857261
transform 1 0 1705 0 1 99919
box 0 0 1 1
use contact_13  contact_13_541
timestamp 1624857261
transform 1 0 1705 0 1 100255
box 0 0 1 1
use contact_13  contact_13_540
timestamp 1624857261
transform 1 0 1705 0 1 100591
box 0 0 1 1
use contact_13  contact_13_539
timestamp 1624857261
transform 1 0 1705 0 1 100927
box 0 0 1 1
use contact_13  contact_13_538
timestamp 1624857261
transform 1 0 1705 0 1 101263
box 0 0 1 1
use contact_13  contact_13_537
timestamp 1624857261
transform 1 0 1705 0 1 101599
box 0 0 1 1
use contact_13  contact_13_536
timestamp 1624857261
transform 1 0 1705 0 1 101935
box 0 0 1 1
use contact_13  contact_13_535
timestamp 1624857261
transform 1 0 1705 0 1 102271
box 0 0 1 1
use contact_13  contact_13_534
timestamp 1624857261
transform 1 0 1705 0 1 102607
box 0 0 1 1
use contact_13  contact_13_533
timestamp 1624857261
transform 1 0 1705 0 1 102943
box 0 0 1 1
use contact_13  contact_13_532
timestamp 1624857261
transform 1 0 1705 0 1 103279
box 0 0 1 1
use contact_13  contact_13_531
timestamp 1624857261
transform 1 0 1705 0 1 103615
box 0 0 1 1
use contact_13  contact_13_530
timestamp 1624857261
transform 1 0 1705 0 1 103951
box 0 0 1 1
use contact_13  contact_13_529
timestamp 1624857261
transform 1 0 1705 0 1 104287
box 0 0 1 1
use contact_13  contact_13_528
timestamp 1624857261
transform 1 0 1705 0 1 104623
box 0 0 1 1
use contact_13  contact_13_527
timestamp 1624857261
transform 1 0 1705 0 1 104959
box 0 0 1 1
use contact_13  contact_13_526
timestamp 1624857261
transform 1 0 1705 0 1 105295
box 0 0 1 1
use contact_13  contact_13_525
timestamp 1624857261
transform 1 0 1705 0 1 105631
box 0 0 1 1
use contact_13  contact_13_524
timestamp 1624857261
transform 1 0 1705 0 1 105967
box 0 0 1 1
use contact_13  contact_13_523
timestamp 1624857261
transform 1 0 1705 0 1 106303
box 0 0 1 1
use contact_13  contact_13_522
timestamp 1624857261
transform 1 0 1705 0 1 106639
box 0 0 1 1
use contact_13  contact_13_521
timestamp 1624857261
transform 1 0 1705 0 1 106975
box 0 0 1 1
use contact_13  contact_13_520
timestamp 1624857261
transform 1 0 1705 0 1 107311
box 0 0 1 1
use contact_13  contact_13_519
timestamp 1624857261
transform 1 0 1705 0 1 107647
box 0 0 1 1
use contact_13  contact_13_518
timestamp 1624857261
transform 1 0 1705 0 1 107983
box 0 0 1 1
use contact_13  contact_13_517
timestamp 1624857261
transform 1 0 1705 0 1 108319
box 0 0 1 1
use contact_13  contact_13_516
timestamp 1624857261
transform 1 0 1705 0 1 108655
box 0 0 1 1
use contact_13  contact_13_515
timestamp 1624857261
transform 1 0 1705 0 1 108991
box 0 0 1 1
use contact_13  contact_13_514
timestamp 1624857261
transform 1 0 1705 0 1 109327
box 0 0 1 1
use contact_13  contact_13_513
timestamp 1624857261
transform 1 0 1705 0 1 109663
box 0 0 1 1
use contact_13  contact_13_512
timestamp 1624857261
transform 1 0 1705 0 1 109999
box 0 0 1 1
use contact_13  contact_13_511
timestamp 1624857261
transform 1 0 1705 0 1 110335
box 0 0 1 1
use contact_13  contact_13_510
timestamp 1624857261
transform 1 0 1705 0 1 110671
box 0 0 1 1
use contact_13  contact_13_509
timestamp 1624857261
transform 1 0 1705 0 1 111007
box 0 0 1 1
use contact_13  contact_13_508
timestamp 1624857261
transform 1 0 1705 0 1 111343
box 0 0 1 1
use contact_13  contact_13_507
timestamp 1624857261
transform 1 0 1705 0 1 111679
box 0 0 1 1
use contact_13  contact_13_506
timestamp 1624857261
transform 1 0 1705 0 1 112015
box 0 0 1 1
use contact_13  contact_13_505
timestamp 1624857261
transform 1 0 1705 0 1 112351
box 0 0 1 1
use contact_13  contact_13_504
timestamp 1624857261
transform 1 0 1705 0 1 112687
box 0 0 1 1
use contact_13  contact_13_503
timestamp 1624857261
transform 1 0 1705 0 1 113023
box 0 0 1 1
use contact_13  contact_13_502
timestamp 1624857261
transform 1 0 1705 0 1 113359
box 0 0 1 1
use contact_13  contact_13_501
timestamp 1624857261
transform 1 0 1705 0 1 113695
box 0 0 1 1
use contact_13  contact_13_500
timestamp 1624857261
transform 1 0 1705 0 1 114031
box 0 0 1 1
use contact_13  contact_13_499
timestamp 1624857261
transform 1 0 1705 0 1 114367
box 0 0 1 1
use contact_13  contact_13_498
timestamp 1624857261
transform 1 0 1705 0 1 114703
box 0 0 1 1
use contact_13  contact_13_497
timestamp 1624857261
transform 1 0 1705 0 1 115039
box 0 0 1 1
use contact_13  contact_13_496
timestamp 1624857261
transform 1 0 1705 0 1 115375
box 0 0 1 1
use contact_13  contact_13_495
timestamp 1624857261
transform 1 0 1705 0 1 115711
box 0 0 1 1
use contact_13  contact_13_494
timestamp 1624857261
transform 1 0 1705 0 1 116047
box 0 0 1 1
use contact_13  contact_13_493
timestamp 1624857261
transform 1 0 1705 0 1 116383
box 0 0 1 1
use contact_13  contact_13_492
timestamp 1624857261
transform 1 0 1705 0 1 116719
box 0 0 1 1
use contact_13  contact_13_491
timestamp 1624857261
transform 1 0 1705 0 1 117055
box 0 0 1 1
use contact_13  contact_13_490
timestamp 1624857261
transform 1 0 1705 0 1 117391
box 0 0 1 1
use contact_13  contact_13_489
timestamp 1624857261
transform 1 0 1705 0 1 117727
box 0 0 1 1
use contact_13  contact_13_488
timestamp 1624857261
transform 1 0 1705 0 1 118063
box 0 0 1 1
use contact_13  contact_13_487
timestamp 1624857261
transform 1 0 1705 0 1 118399
box 0 0 1 1
use contact_13  contact_13_486
timestamp 1624857261
transform 1 0 1705 0 1 118735
box 0 0 1 1
use contact_13  contact_13_485
timestamp 1624857261
transform 1 0 1705 0 1 119071
box 0 0 1 1
use contact_13  contact_13_484
timestamp 1624857261
transform 1 0 1705 0 1 119407
box 0 0 1 1
use contact_13  contact_13_483
timestamp 1624857261
transform 1 0 1705 0 1 119743
box 0 0 1 1
use contact_13  contact_13_482
timestamp 1624857261
transform 1 0 1705 0 1 120079
box 0 0 1 1
use contact_13  contact_13_481
timestamp 1624857261
transform 1 0 1705 0 1 120415
box 0 0 1 1
use contact_13  contact_13_480
timestamp 1624857261
transform 1 0 1705 0 1 120751
box 0 0 1 1
use contact_13  contact_13_479
timestamp 1624857261
transform 1 0 1705 0 1 121087
box 0 0 1 1
use contact_13  contact_13_478
timestamp 1624857261
transform 1 0 1705 0 1 121423
box 0 0 1 1
use contact_13  contact_13_477
timestamp 1624857261
transform 1 0 1705 0 1 121759
box 0 0 1 1
use contact_13  contact_13_476
timestamp 1624857261
transform 1 0 1705 0 1 122095
box 0 0 1 1
use contact_13  contact_13_475
timestamp 1624857261
transform 1 0 1705 0 1 122431
box 0 0 1 1
use contact_13  contact_13_474
timestamp 1624857261
transform 1 0 1705 0 1 122767
box 0 0 1 1
use contact_13  contact_13_473
timestamp 1624857261
transform 1 0 1705 0 1 123103
box 0 0 1 1
use contact_13  contact_13_472
timestamp 1624857261
transform 1 0 1705 0 1 123439
box 0 0 1 1
use contact_13  contact_13_471
timestamp 1624857261
transform 1 0 1705 0 1 123775
box 0 0 1 1
use contact_13  contact_13_470
timestamp 1624857261
transform 1 0 1705 0 1 124111
box 0 0 1 1
use contact_13  contact_13_469
timestamp 1624857261
transform 1 0 1705 0 1 124447
box 0 0 1 1
use contact_13  contact_13_468
timestamp 1624857261
transform 1 0 1705 0 1 124783
box 0 0 1 1
use contact_13  contact_13_467
timestamp 1624857261
transform 1 0 1705 0 1 125119
box 0 0 1 1
use contact_13  contact_13_466
timestamp 1624857261
transform 1 0 1705 0 1 125455
box 0 0 1 1
use contact_13  contact_13_465
timestamp 1624857261
transform 1 0 1705 0 1 125791
box 0 0 1 1
use contact_13  contact_13_464
timestamp 1624857261
transform 1 0 1705 0 1 126127
box 0 0 1 1
use contact_13  contact_13_463
timestamp 1624857261
transform 1 0 1705 0 1 126463
box 0 0 1 1
use contact_13  contact_13_462
timestamp 1624857261
transform 1 0 1705 0 1 126799
box 0 0 1 1
use contact_13  contact_13_461
timestamp 1624857261
transform 1 0 1705 0 1 127135
box 0 0 1 1
use contact_13  contact_13_460
timestamp 1624857261
transform 1 0 1705 0 1 127471
box 0 0 1 1
use contact_13  contact_13_459
timestamp 1624857261
transform 1 0 1705 0 1 127807
box 0 0 1 1
use contact_13  contact_13_458
timestamp 1624857261
transform 1 0 1705 0 1 128143
box 0 0 1 1
use contact_13  contact_13_457
timestamp 1624857261
transform 1 0 1705 0 1 128479
box 0 0 1 1
use contact_13  contact_13_456
timestamp 1624857261
transform 1 0 1705 0 1 128815
box 0 0 1 1
use contact_13  contact_13_455
timestamp 1624857261
transform 1 0 1705 0 1 129151
box 0 0 1 1
use contact_13  contact_13_454
timestamp 1624857261
transform 1 0 1705 0 1 129487
box 0 0 1 1
use contact_13  contact_13_453
timestamp 1624857261
transform 1 0 1705 0 1 129823
box 0 0 1 1
use contact_13  contact_13_452
timestamp 1624857261
transform 1 0 1705 0 1 130159
box 0 0 1 1
use contact_13  contact_13_451
timestamp 1624857261
transform 1 0 1705 0 1 130495
box 0 0 1 1
use contact_13  contact_13_450
timestamp 1624857261
transform 1 0 1705 0 1 130831
box 0 0 1 1
use contact_13  contact_13_449
timestamp 1624857261
transform 1 0 1705 0 1 131167
box 0 0 1 1
use contact_13  contact_13_448
timestamp 1624857261
transform 1 0 1705 0 1 131503
box 0 0 1 1
use contact_13  contact_13_447
timestamp 1624857261
transform 1 0 1705 0 1 131839
box 0 0 1 1
use contact_13  contact_13_446
timestamp 1624857261
transform 1 0 1705 0 1 132175
box 0 0 1 1
use contact_13  contact_13_445
timestamp 1624857261
transform 1 0 1705 0 1 132511
box 0 0 1 1
use contact_13  contact_13_444
timestamp 1624857261
transform 1 0 1705 0 1 132847
box 0 0 1 1
use contact_13  contact_13_443
timestamp 1624857261
transform 1 0 1705 0 1 133183
box 0 0 1 1
use contact_13  contact_13_442
timestamp 1624857261
transform 1 0 1705 0 1 133519
box 0 0 1 1
use contact_13  contact_13_441
timestamp 1624857261
transform 1 0 1705 0 1 133855
box 0 0 1 1
use contact_13  contact_13_440
timestamp 1624857261
transform 1 0 1705 0 1 134191
box 0 0 1 1
use contact_13  contact_13_439
timestamp 1624857261
transform 1 0 1705 0 1 134527
box 0 0 1 1
use contact_13  contact_13_438
timestamp 1624857261
transform 1 0 1705 0 1 134863
box 0 0 1 1
use contact_13  contact_13_437
timestamp 1624857261
transform 1 0 1705 0 1 135199
box 0 0 1 1
use contact_13  contact_13_436
timestamp 1624857261
transform 1 0 1705 0 1 135535
box 0 0 1 1
use contact_13  contact_13_435
timestamp 1624857261
transform 1 0 1705 0 1 135871
box 0 0 1 1
use contact_13  contact_13_434
timestamp 1624857261
transform 1 0 1705 0 1 136207
box 0 0 1 1
use contact_13  contact_13_433
timestamp 1624857261
transform 1 0 1705 0 1 136543
box 0 0 1 1
use contact_13  contact_13_432
timestamp 1624857261
transform 1 0 1705 0 1 136879
box 0 0 1 1
use contact_13  contact_13_431
timestamp 1624857261
transform 1 0 1705 0 1 137215
box 0 0 1 1
use contact_13  contact_13_430
timestamp 1624857261
transform 1 0 1705 0 1 137551
box 0 0 1 1
use contact_13  contact_13_429
timestamp 1624857261
transform 1 0 1705 0 1 137887
box 0 0 1 1
use contact_13  contact_13_428
timestamp 1624857261
transform 1 0 1705 0 1 138223
box 0 0 1 1
use contact_13  contact_13_427
timestamp 1624857261
transform 1 0 1705 0 1 138559
box 0 0 1 1
use contact_13  contact_13_426
timestamp 1624857261
transform 1 0 1705 0 1 138895
box 0 0 1 1
use contact_13  contact_13_425
timestamp 1624857261
transform 1 0 1705 0 1 139231
box 0 0 1 1
use contact_13  contact_13_424
timestamp 1624857261
transform 1 0 1705 0 1 139567
box 0 0 1 1
use contact_13  contact_13_423
timestamp 1624857261
transform 1 0 1705 0 1 139903
box 0 0 1 1
use contact_13  contact_13_422
timestamp 1624857261
transform 1 0 1705 0 1 140239
box 0 0 1 1
use contact_13  contact_13_421
timestamp 1624857261
transform 1 0 1705 0 1 140575
box 0 0 1 1
use contact_13  contact_13_420
timestamp 1624857261
transform 1 0 1705 0 1 140911
box 0 0 1 1
use contact_13  contact_13_419
timestamp 1624857261
transform 1 0 1705 0 1 141247
box 0 0 1 1
use contact_13  contact_13_418
timestamp 1624857261
transform 1 0 1705 0 1 141583
box 0 0 1 1
use contact_13  contact_13_417
timestamp 1624857261
transform 1 0 1705 0 1 141919
box 0 0 1 1
use contact_13  contact_13_416
timestamp 1624857261
transform 1 0 216911 0 1 2143
box 0 0 1 1
use contact_13  contact_13_415
timestamp 1624857261
transform 1 0 216911 0 1 2479
box 0 0 1 1
use contact_13  contact_13_414
timestamp 1624857261
transform 1 0 216911 0 1 2815
box 0 0 1 1
use contact_13  contact_13_413
timestamp 1624857261
transform 1 0 216911 0 1 3151
box 0 0 1 1
use contact_13  contact_13_412
timestamp 1624857261
transform 1 0 216911 0 1 3487
box 0 0 1 1
use contact_13  contact_13_411
timestamp 1624857261
transform 1 0 216911 0 1 3823
box 0 0 1 1
use contact_13  contact_13_410
timestamp 1624857261
transform 1 0 216911 0 1 4159
box 0 0 1 1
use contact_13  contact_13_409
timestamp 1624857261
transform 1 0 216911 0 1 4495
box 0 0 1 1
use contact_13  contact_13_408
timestamp 1624857261
transform 1 0 216911 0 1 4831
box 0 0 1 1
use contact_13  contact_13_407
timestamp 1624857261
transform 1 0 216911 0 1 5167
box 0 0 1 1
use contact_13  contact_13_406
timestamp 1624857261
transform 1 0 216911 0 1 5503
box 0 0 1 1
use contact_13  contact_13_405
timestamp 1624857261
transform 1 0 216911 0 1 5839
box 0 0 1 1
use contact_13  contact_13_404
timestamp 1624857261
transform 1 0 216911 0 1 6175
box 0 0 1 1
use contact_13  contact_13_403
timestamp 1624857261
transform 1 0 216911 0 1 6511
box 0 0 1 1
use contact_13  contact_13_402
timestamp 1624857261
transform 1 0 216911 0 1 6847
box 0 0 1 1
use contact_13  contact_13_401
timestamp 1624857261
transform 1 0 216911 0 1 7183
box 0 0 1 1
use contact_13  contact_13_400
timestamp 1624857261
transform 1 0 216911 0 1 7519
box 0 0 1 1
use contact_13  contact_13_399
timestamp 1624857261
transform 1 0 216911 0 1 7855
box 0 0 1 1
use contact_13  contact_13_398
timestamp 1624857261
transform 1 0 216911 0 1 8191
box 0 0 1 1
use contact_13  contact_13_397
timestamp 1624857261
transform 1 0 216911 0 1 8527
box 0 0 1 1
use contact_13  contact_13_396
timestamp 1624857261
transform 1 0 216911 0 1 8863
box 0 0 1 1
use contact_13  contact_13_395
timestamp 1624857261
transform 1 0 216911 0 1 9199
box 0 0 1 1
use contact_13  contact_13_394
timestamp 1624857261
transform 1 0 216911 0 1 9535
box 0 0 1 1
use contact_13  contact_13_393
timestamp 1624857261
transform 1 0 216911 0 1 9871
box 0 0 1 1
use contact_13  contact_13_392
timestamp 1624857261
transform 1 0 216911 0 1 10207
box 0 0 1 1
use contact_13  contact_13_391
timestamp 1624857261
transform 1 0 216911 0 1 10543
box 0 0 1 1
use contact_13  contact_13_390
timestamp 1624857261
transform 1 0 216911 0 1 10879
box 0 0 1 1
use contact_13  contact_13_389
timestamp 1624857261
transform 1 0 216911 0 1 11215
box 0 0 1 1
use contact_13  contact_13_388
timestamp 1624857261
transform 1 0 216911 0 1 11551
box 0 0 1 1
use contact_13  contact_13_387
timestamp 1624857261
transform 1 0 216911 0 1 11887
box 0 0 1 1
use contact_13  contact_13_386
timestamp 1624857261
transform 1 0 216911 0 1 12223
box 0 0 1 1
use contact_13  contact_13_385
timestamp 1624857261
transform 1 0 216911 0 1 12559
box 0 0 1 1
use contact_13  contact_13_384
timestamp 1624857261
transform 1 0 216911 0 1 12895
box 0 0 1 1
use contact_13  contact_13_383
timestamp 1624857261
transform 1 0 216911 0 1 13231
box 0 0 1 1
use contact_13  contact_13_382
timestamp 1624857261
transform 1 0 216911 0 1 13567
box 0 0 1 1
use contact_13  contact_13_381
timestamp 1624857261
transform 1 0 216911 0 1 13903
box 0 0 1 1
use contact_13  contact_13_380
timestamp 1624857261
transform 1 0 216911 0 1 14239
box 0 0 1 1
use contact_13  contact_13_379
timestamp 1624857261
transform 1 0 216911 0 1 14575
box 0 0 1 1
use contact_13  contact_13_378
timestamp 1624857261
transform 1 0 216911 0 1 14911
box 0 0 1 1
use contact_13  contact_13_377
timestamp 1624857261
transform 1 0 216911 0 1 15247
box 0 0 1 1
use contact_13  contact_13_376
timestamp 1624857261
transform 1 0 216911 0 1 15583
box 0 0 1 1
use contact_13  contact_13_375
timestamp 1624857261
transform 1 0 216911 0 1 15919
box 0 0 1 1
use contact_13  contact_13_374
timestamp 1624857261
transform 1 0 216911 0 1 16255
box 0 0 1 1
use contact_13  contact_13_373
timestamp 1624857261
transform 1 0 216911 0 1 16591
box 0 0 1 1
use contact_13  contact_13_372
timestamp 1624857261
transform 1 0 216911 0 1 16927
box 0 0 1 1
use contact_13  contact_13_371
timestamp 1624857261
transform 1 0 216911 0 1 17263
box 0 0 1 1
use contact_13  contact_13_370
timestamp 1624857261
transform 1 0 216911 0 1 17599
box 0 0 1 1
use contact_13  contact_13_369
timestamp 1624857261
transform 1 0 216911 0 1 17935
box 0 0 1 1
use contact_13  contact_13_368
timestamp 1624857261
transform 1 0 216911 0 1 18271
box 0 0 1 1
use contact_13  contact_13_367
timestamp 1624857261
transform 1 0 216911 0 1 18607
box 0 0 1 1
use contact_13  contact_13_366
timestamp 1624857261
transform 1 0 216911 0 1 18943
box 0 0 1 1
use contact_13  contact_13_365
timestamp 1624857261
transform 1 0 216911 0 1 19279
box 0 0 1 1
use contact_13  contact_13_364
timestamp 1624857261
transform 1 0 216911 0 1 19615
box 0 0 1 1
use contact_13  contact_13_363
timestamp 1624857261
transform 1 0 216911 0 1 19951
box 0 0 1 1
use contact_13  contact_13_362
timestamp 1624857261
transform 1 0 216911 0 1 20287
box 0 0 1 1
use contact_13  contact_13_361
timestamp 1624857261
transform 1 0 216911 0 1 20623
box 0 0 1 1
use contact_13  contact_13_360
timestamp 1624857261
transform 1 0 216911 0 1 20959
box 0 0 1 1
use contact_13  contact_13_359
timestamp 1624857261
transform 1 0 216911 0 1 21295
box 0 0 1 1
use contact_13  contact_13_358
timestamp 1624857261
transform 1 0 216911 0 1 21631
box 0 0 1 1
use contact_13  contact_13_357
timestamp 1624857261
transform 1 0 216911 0 1 21967
box 0 0 1 1
use contact_13  contact_13_356
timestamp 1624857261
transform 1 0 216911 0 1 22303
box 0 0 1 1
use contact_13  contact_13_355
timestamp 1624857261
transform 1 0 216911 0 1 22639
box 0 0 1 1
use contact_13  contact_13_354
timestamp 1624857261
transform 1 0 216911 0 1 22975
box 0 0 1 1
use contact_13  contact_13_353
timestamp 1624857261
transform 1 0 216911 0 1 23311
box 0 0 1 1
use contact_13  contact_13_352
timestamp 1624857261
transform 1 0 216911 0 1 23647
box 0 0 1 1
use contact_13  contact_13_351
timestamp 1624857261
transform 1 0 216911 0 1 23983
box 0 0 1 1
use contact_13  contact_13_350
timestamp 1624857261
transform 1 0 216911 0 1 24319
box 0 0 1 1
use contact_13  contact_13_349
timestamp 1624857261
transform 1 0 216911 0 1 24655
box 0 0 1 1
use contact_13  contact_13_348
timestamp 1624857261
transform 1 0 216911 0 1 24991
box 0 0 1 1
use contact_13  contact_13_347
timestamp 1624857261
transform 1 0 216911 0 1 25327
box 0 0 1 1
use contact_13  contact_13_346
timestamp 1624857261
transform 1 0 216911 0 1 25663
box 0 0 1 1
use contact_13  contact_13_345
timestamp 1624857261
transform 1 0 216911 0 1 25999
box 0 0 1 1
use contact_13  contact_13_344
timestamp 1624857261
transform 1 0 216911 0 1 26335
box 0 0 1 1
use contact_13  contact_13_343
timestamp 1624857261
transform 1 0 216911 0 1 26671
box 0 0 1 1
use contact_13  contact_13_342
timestamp 1624857261
transform 1 0 216911 0 1 27007
box 0 0 1 1
use contact_13  contact_13_341
timestamp 1624857261
transform 1 0 216911 0 1 27343
box 0 0 1 1
use contact_13  contact_13_340
timestamp 1624857261
transform 1 0 216911 0 1 27679
box 0 0 1 1
use contact_13  contact_13_339
timestamp 1624857261
transform 1 0 216911 0 1 28015
box 0 0 1 1
use contact_13  contact_13_338
timestamp 1624857261
transform 1 0 216911 0 1 28351
box 0 0 1 1
use contact_13  contact_13_337
timestamp 1624857261
transform 1 0 216911 0 1 28687
box 0 0 1 1
use contact_13  contact_13_336
timestamp 1624857261
transform 1 0 216911 0 1 29023
box 0 0 1 1
use contact_13  contact_13_335
timestamp 1624857261
transform 1 0 216911 0 1 29359
box 0 0 1 1
use contact_13  contact_13_334
timestamp 1624857261
transform 1 0 216911 0 1 29695
box 0 0 1 1
use contact_13  contact_13_333
timestamp 1624857261
transform 1 0 216911 0 1 30031
box 0 0 1 1
use contact_13  contact_13_332
timestamp 1624857261
transform 1 0 216911 0 1 30367
box 0 0 1 1
use contact_13  contact_13_331
timestamp 1624857261
transform 1 0 216911 0 1 30703
box 0 0 1 1
use contact_13  contact_13_330
timestamp 1624857261
transform 1 0 216911 0 1 31039
box 0 0 1 1
use contact_13  contact_13_329
timestamp 1624857261
transform 1 0 216911 0 1 31375
box 0 0 1 1
use contact_13  contact_13_328
timestamp 1624857261
transform 1 0 216911 0 1 31711
box 0 0 1 1
use contact_13  contact_13_327
timestamp 1624857261
transform 1 0 216911 0 1 32047
box 0 0 1 1
use contact_13  contact_13_326
timestamp 1624857261
transform 1 0 216911 0 1 32383
box 0 0 1 1
use contact_13  contact_13_325
timestamp 1624857261
transform 1 0 216911 0 1 32719
box 0 0 1 1
use contact_13  contact_13_324
timestamp 1624857261
transform 1 0 216911 0 1 33055
box 0 0 1 1
use contact_13  contact_13_323
timestamp 1624857261
transform 1 0 216911 0 1 33391
box 0 0 1 1
use contact_13  contact_13_322
timestamp 1624857261
transform 1 0 216911 0 1 33727
box 0 0 1 1
use contact_13  contact_13_321
timestamp 1624857261
transform 1 0 216911 0 1 34063
box 0 0 1 1
use contact_13  contact_13_320
timestamp 1624857261
transform 1 0 216911 0 1 34399
box 0 0 1 1
use contact_13  contact_13_319
timestamp 1624857261
transform 1 0 216911 0 1 34735
box 0 0 1 1
use contact_13  contact_13_318
timestamp 1624857261
transform 1 0 216911 0 1 35071
box 0 0 1 1
use contact_13  contact_13_317
timestamp 1624857261
transform 1 0 216911 0 1 35407
box 0 0 1 1
use contact_13  contact_13_316
timestamp 1624857261
transform 1 0 216911 0 1 35743
box 0 0 1 1
use contact_13  contact_13_315
timestamp 1624857261
transform 1 0 216911 0 1 36079
box 0 0 1 1
use contact_13  contact_13_314
timestamp 1624857261
transform 1 0 216911 0 1 36415
box 0 0 1 1
use contact_13  contact_13_313
timestamp 1624857261
transform 1 0 216911 0 1 36751
box 0 0 1 1
use contact_13  contact_13_312
timestamp 1624857261
transform 1 0 216911 0 1 37087
box 0 0 1 1
use contact_13  contact_13_311
timestamp 1624857261
transform 1 0 216911 0 1 37423
box 0 0 1 1
use contact_13  contact_13_310
timestamp 1624857261
transform 1 0 216911 0 1 37759
box 0 0 1 1
use contact_13  contact_13_309
timestamp 1624857261
transform 1 0 216911 0 1 38095
box 0 0 1 1
use contact_13  contact_13_308
timestamp 1624857261
transform 1 0 216911 0 1 38431
box 0 0 1 1
use contact_13  contact_13_307
timestamp 1624857261
transform 1 0 216911 0 1 38767
box 0 0 1 1
use contact_13  contact_13_306
timestamp 1624857261
transform 1 0 216911 0 1 39103
box 0 0 1 1
use contact_13  contact_13_305
timestamp 1624857261
transform 1 0 216911 0 1 39439
box 0 0 1 1
use contact_13  contact_13_304
timestamp 1624857261
transform 1 0 216911 0 1 39775
box 0 0 1 1
use contact_13  contact_13_303
timestamp 1624857261
transform 1 0 216911 0 1 40111
box 0 0 1 1
use contact_13  contact_13_302
timestamp 1624857261
transform 1 0 216911 0 1 40447
box 0 0 1 1
use contact_13  contact_13_301
timestamp 1624857261
transform 1 0 216911 0 1 40783
box 0 0 1 1
use contact_13  contact_13_300
timestamp 1624857261
transform 1 0 216911 0 1 41119
box 0 0 1 1
use contact_13  contact_13_299
timestamp 1624857261
transform 1 0 216911 0 1 41455
box 0 0 1 1
use contact_13  contact_13_298
timestamp 1624857261
transform 1 0 216911 0 1 41791
box 0 0 1 1
use contact_13  contact_13_297
timestamp 1624857261
transform 1 0 216911 0 1 42127
box 0 0 1 1
use contact_13  contact_13_296
timestamp 1624857261
transform 1 0 216911 0 1 42463
box 0 0 1 1
use contact_13  contact_13_295
timestamp 1624857261
transform 1 0 216911 0 1 42799
box 0 0 1 1
use contact_13  contact_13_294
timestamp 1624857261
transform 1 0 216911 0 1 43135
box 0 0 1 1
use contact_13  contact_13_293
timestamp 1624857261
transform 1 0 216911 0 1 43471
box 0 0 1 1
use contact_13  contact_13_292
timestamp 1624857261
transform 1 0 216911 0 1 43807
box 0 0 1 1
use contact_13  contact_13_291
timestamp 1624857261
transform 1 0 216911 0 1 44143
box 0 0 1 1
use contact_13  contact_13_290
timestamp 1624857261
transform 1 0 216911 0 1 44479
box 0 0 1 1
use contact_13  contact_13_289
timestamp 1624857261
transform 1 0 216911 0 1 44815
box 0 0 1 1
use contact_13  contact_13_288
timestamp 1624857261
transform 1 0 216911 0 1 45151
box 0 0 1 1
use contact_13  contact_13_287
timestamp 1624857261
transform 1 0 216911 0 1 45487
box 0 0 1 1
use contact_13  contact_13_286
timestamp 1624857261
transform 1 0 216911 0 1 45823
box 0 0 1 1
use contact_13  contact_13_285
timestamp 1624857261
transform 1 0 216911 0 1 46159
box 0 0 1 1
use contact_13  contact_13_284
timestamp 1624857261
transform 1 0 216911 0 1 46495
box 0 0 1 1
use contact_13  contact_13_283
timestamp 1624857261
transform 1 0 216911 0 1 46831
box 0 0 1 1
use contact_13  contact_13_282
timestamp 1624857261
transform 1 0 216911 0 1 47167
box 0 0 1 1
use contact_13  contact_13_281
timestamp 1624857261
transform 1 0 216911 0 1 47503
box 0 0 1 1
use contact_13  contact_13_280
timestamp 1624857261
transform 1 0 216911 0 1 47839
box 0 0 1 1
use contact_13  contact_13_279
timestamp 1624857261
transform 1 0 216911 0 1 48175
box 0 0 1 1
use contact_13  contact_13_278
timestamp 1624857261
transform 1 0 216911 0 1 48511
box 0 0 1 1
use contact_13  contact_13_277
timestamp 1624857261
transform 1 0 216911 0 1 48847
box 0 0 1 1
use contact_13  contact_13_276
timestamp 1624857261
transform 1 0 216911 0 1 49183
box 0 0 1 1
use contact_13  contact_13_275
timestamp 1624857261
transform 1 0 216911 0 1 49519
box 0 0 1 1
use contact_13  contact_13_274
timestamp 1624857261
transform 1 0 216911 0 1 49855
box 0 0 1 1
use contact_13  contact_13_273
timestamp 1624857261
transform 1 0 216911 0 1 50191
box 0 0 1 1
use contact_13  contact_13_272
timestamp 1624857261
transform 1 0 216911 0 1 50527
box 0 0 1 1
use contact_13  contact_13_271
timestamp 1624857261
transform 1 0 216911 0 1 50863
box 0 0 1 1
use contact_13  contact_13_270
timestamp 1624857261
transform 1 0 216911 0 1 51199
box 0 0 1 1
use contact_13  contact_13_269
timestamp 1624857261
transform 1 0 216911 0 1 51535
box 0 0 1 1
use contact_13  contact_13_268
timestamp 1624857261
transform 1 0 216911 0 1 51871
box 0 0 1 1
use contact_13  contact_13_267
timestamp 1624857261
transform 1 0 216911 0 1 52207
box 0 0 1 1
use contact_13  contact_13_266
timestamp 1624857261
transform 1 0 216911 0 1 52543
box 0 0 1 1
use contact_13  contact_13_265
timestamp 1624857261
transform 1 0 216911 0 1 52879
box 0 0 1 1
use contact_13  contact_13_264
timestamp 1624857261
transform 1 0 216911 0 1 53215
box 0 0 1 1
use contact_13  contact_13_263
timestamp 1624857261
transform 1 0 216911 0 1 53551
box 0 0 1 1
use contact_13  contact_13_262
timestamp 1624857261
transform 1 0 216911 0 1 53887
box 0 0 1 1
use contact_13  contact_13_261
timestamp 1624857261
transform 1 0 216911 0 1 54223
box 0 0 1 1
use contact_13  contact_13_260
timestamp 1624857261
transform 1 0 216911 0 1 54559
box 0 0 1 1
use contact_13  contact_13_259
timestamp 1624857261
transform 1 0 216911 0 1 54895
box 0 0 1 1
use contact_13  contact_13_258
timestamp 1624857261
transform 1 0 216911 0 1 55231
box 0 0 1 1
use contact_13  contact_13_257
timestamp 1624857261
transform 1 0 216911 0 1 55567
box 0 0 1 1
use contact_13  contact_13_256
timestamp 1624857261
transform 1 0 216911 0 1 55903
box 0 0 1 1
use contact_13  contact_13_255
timestamp 1624857261
transform 1 0 216911 0 1 56239
box 0 0 1 1
use contact_13  contact_13_254
timestamp 1624857261
transform 1 0 216911 0 1 56575
box 0 0 1 1
use contact_13  contact_13_253
timestamp 1624857261
transform 1 0 216911 0 1 56911
box 0 0 1 1
use contact_13  contact_13_252
timestamp 1624857261
transform 1 0 216911 0 1 57247
box 0 0 1 1
use contact_13  contact_13_251
timestamp 1624857261
transform 1 0 216911 0 1 57583
box 0 0 1 1
use contact_13  contact_13_250
timestamp 1624857261
transform 1 0 216911 0 1 57919
box 0 0 1 1
use contact_13  contact_13_249
timestamp 1624857261
transform 1 0 216911 0 1 58255
box 0 0 1 1
use contact_13  contact_13_248
timestamp 1624857261
transform 1 0 216911 0 1 58591
box 0 0 1 1
use contact_13  contact_13_247
timestamp 1624857261
transform 1 0 216911 0 1 58927
box 0 0 1 1
use contact_13  contact_13_246
timestamp 1624857261
transform 1 0 216911 0 1 59263
box 0 0 1 1
use contact_13  contact_13_245
timestamp 1624857261
transform 1 0 216911 0 1 59599
box 0 0 1 1
use contact_13  contact_13_244
timestamp 1624857261
transform 1 0 216911 0 1 59935
box 0 0 1 1
use contact_13  contact_13_243
timestamp 1624857261
transform 1 0 216911 0 1 60271
box 0 0 1 1
use contact_13  contact_13_242
timestamp 1624857261
transform 1 0 216911 0 1 60607
box 0 0 1 1
use contact_13  contact_13_241
timestamp 1624857261
transform 1 0 216911 0 1 60943
box 0 0 1 1
use contact_13  contact_13_240
timestamp 1624857261
transform 1 0 216911 0 1 61279
box 0 0 1 1
use contact_13  contact_13_239
timestamp 1624857261
transform 1 0 216911 0 1 61615
box 0 0 1 1
use contact_13  contact_13_238
timestamp 1624857261
transform 1 0 216911 0 1 61951
box 0 0 1 1
use contact_13  contact_13_237
timestamp 1624857261
transform 1 0 216911 0 1 62287
box 0 0 1 1
use contact_13  contact_13_236
timestamp 1624857261
transform 1 0 216911 0 1 62623
box 0 0 1 1
use contact_13  contact_13_235
timestamp 1624857261
transform 1 0 216911 0 1 62959
box 0 0 1 1
use contact_13  contact_13_234
timestamp 1624857261
transform 1 0 216911 0 1 63295
box 0 0 1 1
use contact_13  contact_13_233
timestamp 1624857261
transform 1 0 216911 0 1 63631
box 0 0 1 1
use contact_13  contact_13_232
timestamp 1624857261
transform 1 0 216911 0 1 63967
box 0 0 1 1
use contact_13  contact_13_231
timestamp 1624857261
transform 1 0 216911 0 1 64303
box 0 0 1 1
use contact_13  contact_13_230
timestamp 1624857261
transform 1 0 216911 0 1 64639
box 0 0 1 1
use contact_13  contact_13_229
timestamp 1624857261
transform 1 0 216911 0 1 64975
box 0 0 1 1
use contact_13  contact_13_228
timestamp 1624857261
transform 1 0 216911 0 1 65311
box 0 0 1 1
use contact_13  contact_13_227
timestamp 1624857261
transform 1 0 216911 0 1 65647
box 0 0 1 1
use contact_13  contact_13_226
timestamp 1624857261
transform 1 0 216911 0 1 65983
box 0 0 1 1
use contact_13  contact_13_225
timestamp 1624857261
transform 1 0 216911 0 1 66319
box 0 0 1 1
use contact_13  contact_13_224
timestamp 1624857261
transform 1 0 216911 0 1 66655
box 0 0 1 1
use contact_13  contact_13_223
timestamp 1624857261
transform 1 0 216911 0 1 66991
box 0 0 1 1
use contact_13  contact_13_222
timestamp 1624857261
transform 1 0 216911 0 1 67327
box 0 0 1 1
use contact_13  contact_13_221
timestamp 1624857261
transform 1 0 216911 0 1 67663
box 0 0 1 1
use contact_13  contact_13_220
timestamp 1624857261
transform 1 0 216911 0 1 67999
box 0 0 1 1
use contact_13  contact_13_219
timestamp 1624857261
transform 1 0 216911 0 1 68335
box 0 0 1 1
use contact_13  contact_13_218
timestamp 1624857261
transform 1 0 216911 0 1 68671
box 0 0 1 1
use contact_13  contact_13_217
timestamp 1624857261
transform 1 0 216911 0 1 69007
box 0 0 1 1
use contact_13  contact_13_216
timestamp 1624857261
transform 1 0 216911 0 1 69343
box 0 0 1 1
use contact_13  contact_13_215
timestamp 1624857261
transform 1 0 216911 0 1 69679
box 0 0 1 1
use contact_13  contact_13_214
timestamp 1624857261
transform 1 0 216911 0 1 70015
box 0 0 1 1
use contact_13  contact_13_213
timestamp 1624857261
transform 1 0 216911 0 1 70351
box 0 0 1 1
use contact_13  contact_13_212
timestamp 1624857261
transform 1 0 216911 0 1 70687
box 0 0 1 1
use contact_13  contact_13_211
timestamp 1624857261
transform 1 0 216911 0 1 71023
box 0 0 1 1
use contact_13  contact_13_210
timestamp 1624857261
transform 1 0 216911 0 1 71359
box 0 0 1 1
use contact_13  contact_13_209
timestamp 1624857261
transform 1 0 216911 0 1 71695
box 0 0 1 1
use contact_13  contact_13_208
timestamp 1624857261
transform 1 0 216911 0 1 72031
box 0 0 1 1
use contact_13  contact_13_207
timestamp 1624857261
transform 1 0 216911 0 1 72367
box 0 0 1 1
use contact_13  contact_13_206
timestamp 1624857261
transform 1 0 216911 0 1 72703
box 0 0 1 1
use contact_13  contact_13_205
timestamp 1624857261
transform 1 0 216911 0 1 73039
box 0 0 1 1
use contact_13  contact_13_204
timestamp 1624857261
transform 1 0 216911 0 1 73375
box 0 0 1 1
use contact_13  contact_13_203
timestamp 1624857261
transform 1 0 216911 0 1 73711
box 0 0 1 1
use contact_13  contact_13_202
timestamp 1624857261
transform 1 0 216911 0 1 74047
box 0 0 1 1
use contact_13  contact_13_201
timestamp 1624857261
transform 1 0 216911 0 1 74383
box 0 0 1 1
use contact_13  contact_13_200
timestamp 1624857261
transform 1 0 216911 0 1 74719
box 0 0 1 1
use contact_13  contact_13_199
timestamp 1624857261
transform 1 0 216911 0 1 75055
box 0 0 1 1
use contact_13  contact_13_198
timestamp 1624857261
transform 1 0 216911 0 1 75391
box 0 0 1 1
use contact_13  contact_13_197
timestamp 1624857261
transform 1 0 216911 0 1 75727
box 0 0 1 1
use contact_13  contact_13_196
timestamp 1624857261
transform 1 0 216911 0 1 76063
box 0 0 1 1
use contact_13  contact_13_195
timestamp 1624857261
transform 1 0 216911 0 1 76399
box 0 0 1 1
use contact_13  contact_13_194
timestamp 1624857261
transform 1 0 216911 0 1 76735
box 0 0 1 1
use contact_13  contact_13_193
timestamp 1624857261
transform 1 0 216911 0 1 77071
box 0 0 1 1
use contact_13  contact_13_192
timestamp 1624857261
transform 1 0 216911 0 1 77407
box 0 0 1 1
use contact_13  contact_13_191
timestamp 1624857261
transform 1 0 216911 0 1 77743
box 0 0 1 1
use contact_13  contact_13_190
timestamp 1624857261
transform 1 0 216911 0 1 78079
box 0 0 1 1
use contact_13  contact_13_189
timestamp 1624857261
transform 1 0 216911 0 1 78415
box 0 0 1 1
use contact_13  contact_13_188
timestamp 1624857261
transform 1 0 216911 0 1 78751
box 0 0 1 1
use contact_13  contact_13_187
timestamp 1624857261
transform 1 0 216911 0 1 79087
box 0 0 1 1
use contact_13  contact_13_186
timestamp 1624857261
transform 1 0 216911 0 1 79423
box 0 0 1 1
use contact_13  contact_13_185
timestamp 1624857261
transform 1 0 216911 0 1 79759
box 0 0 1 1
use contact_13  contact_13_184
timestamp 1624857261
transform 1 0 216911 0 1 80095
box 0 0 1 1
use contact_13  contact_13_183
timestamp 1624857261
transform 1 0 216911 0 1 80431
box 0 0 1 1
use contact_13  contact_13_182
timestamp 1624857261
transform 1 0 216911 0 1 80767
box 0 0 1 1
use contact_13  contact_13_181
timestamp 1624857261
transform 1 0 216911 0 1 81103
box 0 0 1 1
use contact_13  contact_13_180
timestamp 1624857261
transform 1 0 216911 0 1 81439
box 0 0 1 1
use contact_13  contact_13_179
timestamp 1624857261
transform 1 0 216911 0 1 81775
box 0 0 1 1
use contact_13  contact_13_178
timestamp 1624857261
transform 1 0 216911 0 1 82111
box 0 0 1 1
use contact_13  contact_13_177
timestamp 1624857261
transform 1 0 216911 0 1 82447
box 0 0 1 1
use contact_13  contact_13_176
timestamp 1624857261
transform 1 0 216911 0 1 82783
box 0 0 1 1
use contact_13  contact_13_175
timestamp 1624857261
transform 1 0 216911 0 1 83119
box 0 0 1 1
use contact_13  contact_13_174
timestamp 1624857261
transform 1 0 216911 0 1 83455
box 0 0 1 1
use contact_13  contact_13_173
timestamp 1624857261
transform 1 0 216911 0 1 83791
box 0 0 1 1
use contact_13  contact_13_172
timestamp 1624857261
transform 1 0 216911 0 1 84127
box 0 0 1 1
use contact_13  contact_13_171
timestamp 1624857261
transform 1 0 216911 0 1 84463
box 0 0 1 1
use contact_13  contact_13_170
timestamp 1624857261
transform 1 0 216911 0 1 84799
box 0 0 1 1
use contact_13  contact_13_169
timestamp 1624857261
transform 1 0 216911 0 1 85135
box 0 0 1 1
use contact_13  contact_13_168
timestamp 1624857261
transform 1 0 216911 0 1 85471
box 0 0 1 1
use contact_13  contact_13_167
timestamp 1624857261
transform 1 0 216911 0 1 85807
box 0 0 1 1
use contact_13  contact_13_166
timestamp 1624857261
transform 1 0 216911 0 1 86143
box 0 0 1 1
use contact_13  contact_13_165
timestamp 1624857261
transform 1 0 216911 0 1 86479
box 0 0 1 1
use contact_13  contact_13_164
timestamp 1624857261
transform 1 0 216911 0 1 86815
box 0 0 1 1
use contact_13  contact_13_163
timestamp 1624857261
transform 1 0 216911 0 1 87151
box 0 0 1 1
use contact_13  contact_13_162
timestamp 1624857261
transform 1 0 216911 0 1 87487
box 0 0 1 1
use contact_13  contact_13_161
timestamp 1624857261
transform 1 0 216911 0 1 87823
box 0 0 1 1
use contact_13  contact_13_160
timestamp 1624857261
transform 1 0 216911 0 1 88159
box 0 0 1 1
use contact_13  contact_13_159
timestamp 1624857261
transform 1 0 216911 0 1 88495
box 0 0 1 1
use contact_13  contact_13_158
timestamp 1624857261
transform 1 0 216911 0 1 88831
box 0 0 1 1
use contact_13  contact_13_157
timestamp 1624857261
transform 1 0 216911 0 1 89167
box 0 0 1 1
use contact_13  contact_13_156
timestamp 1624857261
transform 1 0 216911 0 1 89503
box 0 0 1 1
use contact_13  contact_13_155
timestamp 1624857261
transform 1 0 216911 0 1 89839
box 0 0 1 1
use contact_13  contact_13_154
timestamp 1624857261
transform 1 0 216911 0 1 90175
box 0 0 1 1
use contact_13  contact_13_153
timestamp 1624857261
transform 1 0 216911 0 1 90511
box 0 0 1 1
use contact_13  contact_13_152
timestamp 1624857261
transform 1 0 216911 0 1 90847
box 0 0 1 1
use contact_13  contact_13_151
timestamp 1624857261
transform 1 0 216911 0 1 91183
box 0 0 1 1
use contact_13  contact_13_150
timestamp 1624857261
transform 1 0 216911 0 1 91519
box 0 0 1 1
use contact_13  contact_13_149
timestamp 1624857261
transform 1 0 216911 0 1 91855
box 0 0 1 1
use contact_13  contact_13_148
timestamp 1624857261
transform 1 0 216911 0 1 92191
box 0 0 1 1
use contact_13  contact_13_147
timestamp 1624857261
transform 1 0 216911 0 1 92527
box 0 0 1 1
use contact_13  contact_13_146
timestamp 1624857261
transform 1 0 216911 0 1 92863
box 0 0 1 1
use contact_13  contact_13_145
timestamp 1624857261
transform 1 0 216911 0 1 93199
box 0 0 1 1
use contact_13  contact_13_144
timestamp 1624857261
transform 1 0 216911 0 1 93535
box 0 0 1 1
use contact_13  contact_13_143
timestamp 1624857261
transform 1 0 216911 0 1 93871
box 0 0 1 1
use contact_13  contact_13_142
timestamp 1624857261
transform 1 0 216911 0 1 94207
box 0 0 1 1
use contact_13  contact_13_141
timestamp 1624857261
transform 1 0 216911 0 1 94543
box 0 0 1 1
use contact_13  contact_13_140
timestamp 1624857261
transform 1 0 216911 0 1 94879
box 0 0 1 1
use contact_13  contact_13_139
timestamp 1624857261
transform 1 0 216911 0 1 95215
box 0 0 1 1
use contact_13  contact_13_138
timestamp 1624857261
transform 1 0 216911 0 1 95551
box 0 0 1 1
use contact_13  contact_13_137
timestamp 1624857261
transform 1 0 216911 0 1 95887
box 0 0 1 1
use contact_13  contact_13_136
timestamp 1624857261
transform 1 0 216911 0 1 96223
box 0 0 1 1
use contact_13  contact_13_135
timestamp 1624857261
transform 1 0 216911 0 1 96559
box 0 0 1 1
use contact_13  contact_13_134
timestamp 1624857261
transform 1 0 216911 0 1 96895
box 0 0 1 1
use contact_13  contact_13_133
timestamp 1624857261
transform 1 0 216911 0 1 97231
box 0 0 1 1
use contact_13  contact_13_132
timestamp 1624857261
transform 1 0 216911 0 1 97567
box 0 0 1 1
use contact_13  contact_13_131
timestamp 1624857261
transform 1 0 216911 0 1 97903
box 0 0 1 1
use contact_13  contact_13_130
timestamp 1624857261
transform 1 0 216911 0 1 98239
box 0 0 1 1
use contact_13  contact_13_129
timestamp 1624857261
transform 1 0 216911 0 1 98575
box 0 0 1 1
use contact_13  contact_13_128
timestamp 1624857261
transform 1 0 216911 0 1 98911
box 0 0 1 1
use contact_13  contact_13_127
timestamp 1624857261
transform 1 0 216911 0 1 99247
box 0 0 1 1
use contact_13  contact_13_126
timestamp 1624857261
transform 1 0 216911 0 1 99583
box 0 0 1 1
use contact_13  contact_13_125
timestamp 1624857261
transform 1 0 216911 0 1 99919
box 0 0 1 1
use contact_13  contact_13_124
timestamp 1624857261
transform 1 0 216911 0 1 100255
box 0 0 1 1
use contact_13  contact_13_123
timestamp 1624857261
transform 1 0 216911 0 1 100591
box 0 0 1 1
use contact_13  contact_13_122
timestamp 1624857261
transform 1 0 216911 0 1 100927
box 0 0 1 1
use contact_13  contact_13_121
timestamp 1624857261
transform 1 0 216911 0 1 101263
box 0 0 1 1
use contact_13  contact_13_120
timestamp 1624857261
transform 1 0 216911 0 1 101599
box 0 0 1 1
use contact_13  contact_13_119
timestamp 1624857261
transform 1 0 216911 0 1 101935
box 0 0 1 1
use contact_13  contact_13_118
timestamp 1624857261
transform 1 0 216911 0 1 102271
box 0 0 1 1
use contact_13  contact_13_117
timestamp 1624857261
transform 1 0 216911 0 1 102607
box 0 0 1 1
use contact_13  contact_13_116
timestamp 1624857261
transform 1 0 216911 0 1 102943
box 0 0 1 1
use contact_13  contact_13_115
timestamp 1624857261
transform 1 0 216911 0 1 103279
box 0 0 1 1
use contact_13  contact_13_114
timestamp 1624857261
transform 1 0 216911 0 1 103615
box 0 0 1 1
use contact_13  contact_13_113
timestamp 1624857261
transform 1 0 216911 0 1 103951
box 0 0 1 1
use contact_13  contact_13_112
timestamp 1624857261
transform 1 0 216911 0 1 104287
box 0 0 1 1
use contact_13  contact_13_111
timestamp 1624857261
transform 1 0 216911 0 1 104623
box 0 0 1 1
use contact_13  contact_13_110
timestamp 1624857261
transform 1 0 216911 0 1 104959
box 0 0 1 1
use contact_13  contact_13_109
timestamp 1624857261
transform 1 0 216911 0 1 105295
box 0 0 1 1
use contact_13  contact_13_108
timestamp 1624857261
transform 1 0 216911 0 1 105631
box 0 0 1 1
use contact_13  contact_13_107
timestamp 1624857261
transform 1 0 216911 0 1 105967
box 0 0 1 1
use contact_13  contact_13_106
timestamp 1624857261
transform 1 0 216911 0 1 106303
box 0 0 1 1
use contact_13  contact_13_105
timestamp 1624857261
transform 1 0 216911 0 1 106639
box 0 0 1 1
use contact_13  contact_13_104
timestamp 1624857261
transform 1 0 216911 0 1 106975
box 0 0 1 1
use contact_13  contact_13_103
timestamp 1624857261
transform 1 0 216911 0 1 107311
box 0 0 1 1
use contact_13  contact_13_102
timestamp 1624857261
transform 1 0 216911 0 1 107647
box 0 0 1 1
use contact_13  contact_13_101
timestamp 1624857261
transform 1 0 216911 0 1 107983
box 0 0 1 1
use contact_13  contact_13_100
timestamp 1624857261
transform 1 0 216911 0 1 108319
box 0 0 1 1
use contact_13  contact_13_99
timestamp 1624857261
transform 1 0 216911 0 1 108655
box 0 0 1 1
use contact_13  contact_13_98
timestamp 1624857261
transform 1 0 216911 0 1 108991
box 0 0 1 1
use contact_13  contact_13_97
timestamp 1624857261
transform 1 0 216911 0 1 109327
box 0 0 1 1
use contact_13  contact_13_96
timestamp 1624857261
transform 1 0 216911 0 1 109663
box 0 0 1 1
use contact_13  contact_13_95
timestamp 1624857261
transform 1 0 216911 0 1 109999
box 0 0 1 1
use contact_13  contact_13_94
timestamp 1624857261
transform 1 0 216911 0 1 110335
box 0 0 1 1
use contact_13  contact_13_93
timestamp 1624857261
transform 1 0 216911 0 1 110671
box 0 0 1 1
use contact_13  contact_13_92
timestamp 1624857261
transform 1 0 216911 0 1 111007
box 0 0 1 1
use contact_13  contact_13_91
timestamp 1624857261
transform 1 0 216911 0 1 111343
box 0 0 1 1
use contact_13  contact_13_90
timestamp 1624857261
transform 1 0 216911 0 1 111679
box 0 0 1 1
use contact_13  contact_13_89
timestamp 1624857261
transform 1 0 216911 0 1 112015
box 0 0 1 1
use contact_13  contact_13_88
timestamp 1624857261
transform 1 0 216911 0 1 112351
box 0 0 1 1
use contact_13  contact_13_87
timestamp 1624857261
transform 1 0 216911 0 1 112687
box 0 0 1 1
use contact_13  contact_13_86
timestamp 1624857261
transform 1 0 216911 0 1 113023
box 0 0 1 1
use contact_13  contact_13_85
timestamp 1624857261
transform 1 0 216911 0 1 113359
box 0 0 1 1
use contact_13  contact_13_84
timestamp 1624857261
transform 1 0 216911 0 1 113695
box 0 0 1 1
use contact_13  contact_13_83
timestamp 1624857261
transform 1 0 216911 0 1 114031
box 0 0 1 1
use contact_13  contact_13_82
timestamp 1624857261
transform 1 0 216911 0 1 114367
box 0 0 1 1
use contact_13  contact_13_81
timestamp 1624857261
transform 1 0 216911 0 1 114703
box 0 0 1 1
use contact_13  contact_13_80
timestamp 1624857261
transform 1 0 216911 0 1 115039
box 0 0 1 1
use contact_13  contact_13_79
timestamp 1624857261
transform 1 0 216911 0 1 115375
box 0 0 1 1
use contact_13  contact_13_78
timestamp 1624857261
transform 1 0 216911 0 1 115711
box 0 0 1 1
use contact_13  contact_13_77
timestamp 1624857261
transform 1 0 216911 0 1 116047
box 0 0 1 1
use contact_13  contact_13_76
timestamp 1624857261
transform 1 0 216911 0 1 116383
box 0 0 1 1
use contact_13  contact_13_75
timestamp 1624857261
transform 1 0 216911 0 1 116719
box 0 0 1 1
use contact_13  contact_13_74
timestamp 1624857261
transform 1 0 216911 0 1 117055
box 0 0 1 1
use contact_13  contact_13_73
timestamp 1624857261
transform 1 0 216911 0 1 117391
box 0 0 1 1
use contact_13  contact_13_72
timestamp 1624857261
transform 1 0 216911 0 1 117727
box 0 0 1 1
use contact_13  contact_13_71
timestamp 1624857261
transform 1 0 216911 0 1 118063
box 0 0 1 1
use contact_13  contact_13_70
timestamp 1624857261
transform 1 0 216911 0 1 118399
box 0 0 1 1
use contact_13  contact_13_69
timestamp 1624857261
transform 1 0 216911 0 1 118735
box 0 0 1 1
use contact_13  contact_13_68
timestamp 1624857261
transform 1 0 216911 0 1 119071
box 0 0 1 1
use contact_13  contact_13_67
timestamp 1624857261
transform 1 0 216911 0 1 119407
box 0 0 1 1
use contact_13  contact_13_66
timestamp 1624857261
transform 1 0 216911 0 1 119743
box 0 0 1 1
use contact_13  contact_13_65
timestamp 1624857261
transform 1 0 216911 0 1 120079
box 0 0 1 1
use contact_13  contact_13_64
timestamp 1624857261
transform 1 0 216911 0 1 120415
box 0 0 1 1
use contact_13  contact_13_63
timestamp 1624857261
transform 1 0 216911 0 1 120751
box 0 0 1 1
use contact_13  contact_13_62
timestamp 1624857261
transform 1 0 216911 0 1 121087
box 0 0 1 1
use contact_13  contact_13_61
timestamp 1624857261
transform 1 0 216911 0 1 121423
box 0 0 1 1
use contact_13  contact_13_60
timestamp 1624857261
transform 1 0 216911 0 1 121759
box 0 0 1 1
use contact_13  contact_13_59
timestamp 1624857261
transform 1 0 216911 0 1 122095
box 0 0 1 1
use contact_13  contact_13_58
timestamp 1624857261
transform 1 0 216911 0 1 122431
box 0 0 1 1
use contact_13  contact_13_57
timestamp 1624857261
transform 1 0 216911 0 1 122767
box 0 0 1 1
use contact_13  contact_13_56
timestamp 1624857261
transform 1 0 216911 0 1 123103
box 0 0 1 1
use contact_13  contact_13_55
timestamp 1624857261
transform 1 0 216911 0 1 123439
box 0 0 1 1
use contact_13  contact_13_54
timestamp 1624857261
transform 1 0 216911 0 1 123775
box 0 0 1 1
use contact_13  contact_13_53
timestamp 1624857261
transform 1 0 216911 0 1 124111
box 0 0 1 1
use contact_13  contact_13_52
timestamp 1624857261
transform 1 0 216911 0 1 124447
box 0 0 1 1
use contact_13  contact_13_51
timestamp 1624857261
transform 1 0 216911 0 1 124783
box 0 0 1 1
use contact_13  contact_13_50
timestamp 1624857261
transform 1 0 216911 0 1 125119
box 0 0 1 1
use contact_13  contact_13_49
timestamp 1624857261
transform 1 0 216911 0 1 125455
box 0 0 1 1
use contact_13  contact_13_48
timestamp 1624857261
transform 1 0 216911 0 1 125791
box 0 0 1 1
use contact_13  contact_13_47
timestamp 1624857261
transform 1 0 216911 0 1 126127
box 0 0 1 1
use contact_13  contact_13_46
timestamp 1624857261
transform 1 0 216911 0 1 126463
box 0 0 1 1
use contact_13  contact_13_45
timestamp 1624857261
transform 1 0 216911 0 1 126799
box 0 0 1 1
use contact_13  contact_13_44
timestamp 1624857261
transform 1 0 216911 0 1 127135
box 0 0 1 1
use contact_13  contact_13_43
timestamp 1624857261
transform 1 0 216911 0 1 127471
box 0 0 1 1
use contact_13  contact_13_42
timestamp 1624857261
transform 1 0 216911 0 1 127807
box 0 0 1 1
use contact_13  contact_13_41
timestamp 1624857261
transform 1 0 216911 0 1 128143
box 0 0 1 1
use contact_13  contact_13_40
timestamp 1624857261
transform 1 0 216911 0 1 128479
box 0 0 1 1
use contact_13  contact_13_39
timestamp 1624857261
transform 1 0 216911 0 1 128815
box 0 0 1 1
use contact_13  contact_13_38
timestamp 1624857261
transform 1 0 216911 0 1 129151
box 0 0 1 1
use contact_13  contact_13_37
timestamp 1624857261
transform 1 0 216911 0 1 129487
box 0 0 1 1
use contact_13  contact_13_36
timestamp 1624857261
transform 1 0 216911 0 1 129823
box 0 0 1 1
use contact_13  contact_13_35
timestamp 1624857261
transform 1 0 216911 0 1 130159
box 0 0 1 1
use contact_13  contact_13_34
timestamp 1624857261
transform 1 0 216911 0 1 130495
box 0 0 1 1
use contact_13  contact_13_33
timestamp 1624857261
transform 1 0 216911 0 1 130831
box 0 0 1 1
use contact_13  contact_13_32
timestamp 1624857261
transform 1 0 216911 0 1 131167
box 0 0 1 1
use contact_13  contact_13_31
timestamp 1624857261
transform 1 0 216911 0 1 131503
box 0 0 1 1
use contact_13  contact_13_30
timestamp 1624857261
transform 1 0 216911 0 1 131839
box 0 0 1 1
use contact_13  contact_13_29
timestamp 1624857261
transform 1 0 216911 0 1 132175
box 0 0 1 1
use contact_13  contact_13_28
timestamp 1624857261
transform 1 0 216911 0 1 132511
box 0 0 1 1
use contact_13  contact_13_27
timestamp 1624857261
transform 1 0 216911 0 1 132847
box 0 0 1 1
use contact_13  contact_13_26
timestamp 1624857261
transform 1 0 216911 0 1 133183
box 0 0 1 1
use contact_13  contact_13_25
timestamp 1624857261
transform 1 0 216911 0 1 133519
box 0 0 1 1
use contact_13  contact_13_24
timestamp 1624857261
transform 1 0 216911 0 1 133855
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1624857261
transform 1 0 216911 0 1 134191
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1624857261
transform 1 0 216911 0 1 134527
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1624857261
transform 1 0 216911 0 1 134863
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1624857261
transform 1 0 216911 0 1 135199
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1624857261
transform 1 0 216911 0 1 135535
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1624857261
transform 1 0 216911 0 1 135871
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1624857261
transform 1 0 216911 0 1 136207
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1624857261
transform 1 0 216911 0 1 136543
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1624857261
transform 1 0 216911 0 1 136879
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1624857261
transform 1 0 216911 0 1 137215
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1624857261
transform 1 0 216911 0 1 137551
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1624857261
transform 1 0 216911 0 1 137887
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1624857261
transform 1 0 216911 0 1 138223
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1624857261
transform 1 0 216911 0 1 138559
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1624857261
transform 1 0 216911 0 1 138895
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1624857261
transform 1 0 216911 0 1 139231
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1624857261
transform 1 0 216911 0 1 139567
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1624857261
transform 1 0 216911 0 1 139903
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1624857261
transform 1 0 216911 0 1 140239
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1624857261
transform 1 0 216911 0 1 140575
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1624857261
transform 1 0 216911 0 1 140911
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1624857261
transform 1 0 216911 0 1 141247
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1624857261
transform 1 0 216911 0 1 141583
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1624857261
transform 1 0 216911 0 1 141919
box 0 0 1 1
use contact_9  contact_9_598
timestamp 1624857261
transform 1 0 15205 0 1 17523
box 0 0 1 1
use contact_9  contact_9_597
timestamp 1624857261
transform 1 0 27572 0 1 17523
box 0 0 1 1
use contact_9  contact_9_596
timestamp 1624857261
transform 1 0 15205 0 1 18937
box 0 0 1 1
use contact_9  contact_9_595
timestamp 1624857261
transform 1 0 27696 0 1 18937
box 0 0 1 1
use contact_9  contact_9_594
timestamp 1624857261
transform 1 0 15205 0 1 20351
box 0 0 1 1
use contact_9  contact_9_593
timestamp 1624857261
transform 1 0 27448 0 1 20351
box 0 0 1 1
use contact_9  contact_9_592
timestamp 1624857261
transform 1 0 15205 0 1 23179
box 0 0 1 1
use contact_9  contact_9_591
timestamp 1624857261
transform 1 0 23747 0 1 23179
box 0 0 1 1
use contact_9  contact_9_590
timestamp 1624857261
transform 1 0 203479 0 1 130369
box 0 0 1 1
use contact_9  contact_9_589
timestamp 1624857261
transform 1 0 190870 0 1 130369
box 0 0 1 1
use contact_9  contact_9_588
timestamp 1624857261
transform 1 0 203479 0 1 128955
box 0 0 1 1
use contact_9  contact_9_587
timestamp 1624857261
transform 1 0 190994 0 1 128955
box 0 0 1 1
use contact_9  contact_9_586
timestamp 1624857261
transform 1 0 203479 0 1 127541
box 0 0 1 1
use contact_9  contact_9_585
timestamp 1624857261
transform 1 0 194853 0 1 127541
box 0 0 1 1
use contact_9  contact_9_584
timestamp 1624857261
transform 1 0 2108 0 1 30287
box 0 0 1 1
use contact_9  contact_9_583
timestamp 1624857261
transform 1 0 216492 0 1 117605
box 0 0 1 1
use contact_9  contact_9_582
timestamp 1624857261
transform 1 0 15152 0 1 34915
box 0 0 1 1
use contact_9  contact_9_581
timestamp 1624857261
transform 1 0 15406 0 1 34915
box 0 0 1 1
use contact_9  contact_9_580
timestamp 1624857261
transform 1 0 15152 0 1 36473
box 0 0 1 1
use contact_9  contact_9_579
timestamp 1624857261
transform 1 0 15486 0 1 36473
box 0 0 1 1
use contact_9  contact_9_578
timestamp 1624857261
transform 1 0 15152 0 1 37743
box 0 0 1 1
use contact_9  contact_9_577
timestamp 1624857261
transform 1 0 15566 0 1 37743
box 0 0 1 1
use contact_9  contact_9_576
timestamp 1624857261
transform 1 0 15152 0 1 39301
box 0 0 1 1
use contact_9  contact_9_575
timestamp 1624857261
transform 1 0 15646 0 1 39301
box 0 0 1 1
use contact_9  contact_9_574
timestamp 1624857261
transform 1 0 15152 0 1 40571
box 0 0 1 1
use contact_9  contact_9_573
timestamp 1624857261
transform 1 0 15726 0 1 40571
box 0 0 1 1
use contact_9  contact_9_572
timestamp 1624857261
transform 1 0 15152 0 1 42129
box 0 0 1 1
use contact_9  contact_9_571
timestamp 1624857261
transform 1 0 15806 0 1 42129
box 0 0 1 1
use contact_9  contact_9_570
timestamp 1624857261
transform 1 0 15152 0 1 43399
box 0 0 1 1
use contact_9  contact_9_569
timestamp 1624857261
transform 1 0 15886 0 1 43399
box 0 0 1 1
use contact_9  contact_9_568
timestamp 1624857261
transform 1 0 15152 0 1 44957
box 0 0 1 1
use contact_9  contact_9_567
timestamp 1624857261
transform 1 0 15966 0 1 44957
box 0 0 1 1
use contact_9  contact_9_566
timestamp 1624857261
transform 1 0 203532 0 1 24165
box 0 0 1 1
use contact_9  contact_9_565
timestamp 1624857261
transform 1 0 203194 0 1 24165
box 0 0 1 1
use contact_9  contact_9_564
timestamp 1624857261
transform 1 0 203532 0 1 22607
box 0 0 1 1
use contact_9  contact_9_563
timestamp 1624857261
transform 1 0 203114 0 1 22607
box 0 0 1 1
use contact_9  contact_9_562
timestamp 1624857261
transform 1 0 203532 0 1 21337
box 0 0 1 1
use contact_9  contact_9_561
timestamp 1624857261
transform 1 0 203034 0 1 21337
box 0 0 1 1
use contact_9  contact_9_560
timestamp 1624857261
transform 1 0 203532 0 1 19779
box 0 0 1 1
use contact_9  contact_9_559
timestamp 1624857261
transform 1 0 202954 0 1 19779
box 0 0 1 1
use contact_9  contact_9_558
timestamp 1624857261
transform 1 0 203532 0 1 18509
box 0 0 1 1
use contact_9  contact_9_557
timestamp 1624857261
transform 1 0 202874 0 1 18509
box 0 0 1 1
use contact_9  contact_9_556
timestamp 1624857261
transform 1 0 203532 0 1 16951
box 0 0 1 1
use contact_9  contact_9_555
timestamp 1624857261
transform 1 0 202794 0 1 16951
box 0 0 1 1
use contact_9  contact_9_554
timestamp 1624857261
transform 1 0 203532 0 1 15681
box 0 0 1 1
use contact_9  contact_9_553
timestamp 1624857261
transform 1 0 202714 0 1 15681
box 0 0 1 1
use contact_9  contact_9_552
timestamp 1624857261
transform 1 0 203532 0 1 14123
box 0 0 1 1
use contact_9  contact_9_551
timestamp 1624857261
transform 1 0 202634 0 1 14123
box 0 0 1 1
use contact_9  contact_9_550
timestamp 1624857261
transform 1 0 2321 0 1 13138
box 0 0 1 1
use contact_9  contact_9_549
timestamp 1624857261
transform 1 0 2321 0 1 14838
box 0 0 1 1
use contact_9  contact_9_548
timestamp 1624857261
transform 1 0 5506 0 1 13243
box 0 0 1 1
use contact_9  contact_9_547
timestamp 1624857261
transform 1 0 24719 0 1 2711
box 0 0 1 1
use contact_9  contact_9_546
timestamp 1624857261
transform 1 0 25887 0 1 2711
box 0 0 1 1
use contact_9  contact_9_545
timestamp 1624857261
transform 1 0 27055 0 1 2711
box 0 0 1 1
use contact_9  contact_9_544
timestamp 1624857261
transform 1 0 28223 0 1 2711
box 0 0 1 1
use contact_9  contact_9_543
timestamp 1624857261
transform 1 0 29391 0 1 2711
box 0 0 1 1
use contact_9  contact_9_542
timestamp 1624857261
transform 1 0 30559 0 1 2711
box 0 0 1 1
use contact_9  contact_9_541
timestamp 1624857261
transform 1 0 31727 0 1 2711
box 0 0 1 1
use contact_9  contact_9_540
timestamp 1624857261
transform 1 0 32895 0 1 2711
box 0 0 1 1
use contact_9  contact_9_539
timestamp 1624857261
transform 1 0 34063 0 1 2711
box 0 0 1 1
use contact_9  contact_9_538
timestamp 1624857261
transform 1 0 35231 0 1 2711
box 0 0 1 1
use contact_9  contact_9_537
timestamp 1624857261
transform 1 0 36399 0 1 2711
box 0 0 1 1
use contact_9  contact_9_536
timestamp 1624857261
transform 1 0 37567 0 1 2711
box 0 0 1 1
use contact_9  contact_9_535
timestamp 1624857261
transform 1 0 38735 0 1 2711
box 0 0 1 1
use contact_9  contact_9_534
timestamp 1624857261
transform 1 0 39903 0 1 2711
box 0 0 1 1
use contact_9  contact_9_533
timestamp 1624857261
transform 1 0 41071 0 1 2711
box 0 0 1 1
use contact_9  contact_9_532
timestamp 1624857261
transform 1 0 42239 0 1 2711
box 0 0 1 1
use contact_9  contact_9_531
timestamp 1624857261
transform 1 0 43407 0 1 2711
box 0 0 1 1
use contact_9  contact_9_530
timestamp 1624857261
transform 1 0 44575 0 1 2711
box 0 0 1 1
use contact_9  contact_9_529
timestamp 1624857261
transform 1 0 45743 0 1 2711
box 0 0 1 1
use contact_9  contact_9_528
timestamp 1624857261
transform 1 0 46911 0 1 2711
box 0 0 1 1
use contact_9  contact_9_527
timestamp 1624857261
transform 1 0 48079 0 1 2711
box 0 0 1 1
use contact_9  contact_9_526
timestamp 1624857261
transform 1 0 49247 0 1 2711
box 0 0 1 1
use contact_9  contact_9_525
timestamp 1624857261
transform 1 0 50415 0 1 2711
box 0 0 1 1
use contact_9  contact_9_524
timestamp 1624857261
transform 1 0 51583 0 1 2711
box 0 0 1 1
use contact_9  contact_9_523
timestamp 1624857261
transform 1 0 52751 0 1 2711
box 0 0 1 1
use contact_9  contact_9_522
timestamp 1624857261
transform 1 0 53919 0 1 2711
box 0 0 1 1
use contact_9  contact_9_521
timestamp 1624857261
transform 1 0 55087 0 1 2711
box 0 0 1 1
use contact_9  contact_9_520
timestamp 1624857261
transform 1 0 56255 0 1 2711
box 0 0 1 1
use contact_9  contact_9_519
timestamp 1624857261
transform 1 0 57423 0 1 2711
box 0 0 1 1
use contact_9  contact_9_518
timestamp 1624857261
transform 1 0 58591 0 1 2711
box 0 0 1 1
use contact_9  contact_9_517
timestamp 1624857261
transform 1 0 59759 0 1 2711
box 0 0 1 1
use contact_9  contact_9_516
timestamp 1624857261
transform 1 0 60927 0 1 2711
box 0 0 1 1
use contact_9  contact_9_515
timestamp 1624857261
transform 1 0 29555 0 1 17691
box 0 0 1 1
use contact_9  contact_9_514
timestamp 1624857261
transform 1 0 34547 0 1 17691
box 0 0 1 1
use contact_9  contact_9_513
timestamp 1624857261
transform 1 0 39539 0 1 17691
box 0 0 1 1
use contact_9  contact_9_512
timestamp 1624857261
transform 1 0 44531 0 1 17691
box 0 0 1 1
use contact_9  contact_9_511
timestamp 1624857261
transform 1 0 49523 0 1 17691
box 0 0 1 1
use contact_9  contact_9_510
timestamp 1624857261
transform 1 0 54515 0 1 17691
box 0 0 1 1
use contact_9  contact_9_509
timestamp 1624857261
transform 1 0 59507 0 1 17691
box 0 0 1 1
use contact_9  contact_9_508
timestamp 1624857261
transform 1 0 64499 0 1 17691
box 0 0 1 1
use contact_9  contact_9_507
timestamp 1624857261
transform 1 0 69491 0 1 17691
box 0 0 1 1
use contact_9  contact_9_506
timestamp 1624857261
transform 1 0 74483 0 1 17691
box 0 0 1 1
use contact_9  contact_9_505
timestamp 1624857261
transform 1 0 79475 0 1 17691
box 0 0 1 1
use contact_9  contact_9_504
timestamp 1624857261
transform 1 0 84467 0 1 17691
box 0 0 1 1
use contact_9  contact_9_503
timestamp 1624857261
transform 1 0 89459 0 1 17691
box 0 0 1 1
use contact_9  contact_9_502
timestamp 1624857261
transform 1 0 94451 0 1 17691
box 0 0 1 1
use contact_9  contact_9_501
timestamp 1624857261
transform 1 0 99443 0 1 17691
box 0 0 1 1
use contact_9  contact_9_500
timestamp 1624857261
transform 1 0 104435 0 1 17691
box 0 0 1 1
use contact_9  contact_9_499
timestamp 1624857261
transform 1 0 109427 0 1 17691
box 0 0 1 1
use contact_9  contact_9_498
timestamp 1624857261
transform 1 0 114419 0 1 17691
box 0 0 1 1
use contact_9  contact_9_497
timestamp 1624857261
transform 1 0 119411 0 1 17691
box 0 0 1 1
use contact_9  contact_9_496
timestamp 1624857261
transform 1 0 124403 0 1 17691
box 0 0 1 1
use contact_9  contact_9_495
timestamp 1624857261
transform 1 0 129395 0 1 17691
box 0 0 1 1
use contact_9  contact_9_494
timestamp 1624857261
transform 1 0 134387 0 1 17691
box 0 0 1 1
use contact_9  contact_9_493
timestamp 1624857261
transform 1 0 139379 0 1 17691
box 0 0 1 1
use contact_9  contact_9_492
timestamp 1624857261
transform 1 0 144371 0 1 17691
box 0 0 1 1
use contact_9  contact_9_491
timestamp 1624857261
transform 1 0 149363 0 1 17691
box 0 0 1 1
use contact_9  contact_9_490
timestamp 1624857261
transform 1 0 154355 0 1 17691
box 0 0 1 1
use contact_9  contact_9_489
timestamp 1624857261
transform 1 0 159347 0 1 17691
box 0 0 1 1
use contact_9  contact_9_488
timestamp 1624857261
transform 1 0 164339 0 1 17691
box 0 0 1 1
use contact_9  contact_9_487
timestamp 1624857261
transform 1 0 169331 0 1 17691
box 0 0 1 1
use contact_9  contact_9_486
timestamp 1624857261
transform 1 0 174323 0 1 17691
box 0 0 1 1
use contact_9  contact_9_485
timestamp 1624857261
transform 1 0 179315 0 1 17691
box 0 0 1 1
use contact_9  contact_9_484
timestamp 1624857261
transform 1 0 184307 0 1 17691
box 0 0 1 1
use contact_9  contact_9_483
timestamp 1624857261
transform 1 0 16543 0 1 2711
box 0 0 1 1
use contact_9  contact_9_482
timestamp 1624857261
transform 1 0 17711 0 1 2711
box 0 0 1 1
use contact_9  contact_9_481
timestamp 1624857261
transform 1 0 18879 0 1 2711
box 0 0 1 1
use contact_9  contact_9_480
timestamp 1624857261
transform 1 0 14207 0 1 34844
box 0 0 1 1
use contact_9  contact_9_479
timestamp 1624857261
transform 1 0 14207 0 1 36544
box 0 0 1 1
use contact_9  contact_9_478
timestamp 1624857261
transform 1 0 14207 0 1 37672
box 0 0 1 1
use contact_9  contact_9_477
timestamp 1624857261
transform 1 0 14207 0 1 39372
box 0 0 1 1
use contact_9  contact_9_476
timestamp 1624857261
transform 1 0 14207 0 1 40500
box 0 0 1 1
use contact_9  contact_9_475
timestamp 1624857261
transform 1 0 14207 0 1 42200
box 0 0 1 1
use contact_9  contact_9_474
timestamp 1624857261
transform 1 0 14207 0 1 43328
box 0 0 1 1
use contact_9  contact_9_473
timestamp 1624857261
transform 1 0 14207 0 1 45028
box 0 0 1 1
use contact_9  contact_9_472
timestamp 1624857261
transform 1 0 20047 0 1 2711
box 0 0 1 1
use contact_9  contact_9_471
timestamp 1624857261
transform 1 0 21215 0 1 2711
box 0 0 1 1
use contact_9  contact_9_470
timestamp 1624857261
transform 1 0 22383 0 1 2711
box 0 0 1 1
use contact_9  contact_9_469
timestamp 1624857261
transform 1 0 23551 0 1 2711
box 0 0 1 1
use contact_9  contact_9_468
timestamp 1624857261
transform 1 0 216279 0 1 134754
box 0 0 1 1
use contact_9  contact_9_467
timestamp 1624857261
transform 1 0 213178 0 1 134649
box 0 0 1 1
use contact_9  contact_9_466
timestamp 1624857261
transform 1 0 29555 0 1 133029
box 0 0 1 1
use contact_9  contact_9_465
timestamp 1624857261
transform 1 0 34547 0 1 133029
box 0 0 1 1
use contact_9  contact_9_464
timestamp 1624857261
transform 1 0 39539 0 1 133029
box 0 0 1 1
use contact_9  contact_9_463
timestamp 1624857261
transform 1 0 44531 0 1 133029
box 0 0 1 1
use contact_9  contact_9_462
timestamp 1624857261
transform 1 0 49523 0 1 133029
box 0 0 1 1
use contact_9  contact_9_461
timestamp 1624857261
transform 1 0 54515 0 1 133029
box 0 0 1 1
use contact_9  contact_9_460
timestamp 1624857261
transform 1 0 59507 0 1 133029
box 0 0 1 1
use contact_9  contact_9_459
timestamp 1624857261
transform 1 0 64499 0 1 133029
box 0 0 1 1
use contact_9  contact_9_458
timestamp 1624857261
transform 1 0 69491 0 1 133029
box 0 0 1 1
use contact_9  contact_9_457
timestamp 1624857261
transform 1 0 74483 0 1 133029
box 0 0 1 1
use contact_9  contact_9_456
timestamp 1624857261
transform 1 0 79475 0 1 133029
box 0 0 1 1
use contact_9  contact_9_455
timestamp 1624857261
transform 1 0 84467 0 1 133029
box 0 0 1 1
use contact_9  contact_9_454
timestamp 1624857261
transform 1 0 89459 0 1 133029
box 0 0 1 1
use contact_9  contact_9_453
timestamp 1624857261
transform 1 0 94451 0 1 133029
box 0 0 1 1
use contact_9  contact_9_452
timestamp 1624857261
transform 1 0 99443 0 1 133029
box 0 0 1 1
use contact_9  contact_9_451
timestamp 1624857261
transform 1 0 104435 0 1 133029
box 0 0 1 1
use contact_9  contact_9_450
timestamp 1624857261
transform 1 0 109427 0 1 133029
box 0 0 1 1
use contact_9  contact_9_449
timestamp 1624857261
transform 1 0 114419 0 1 133029
box 0 0 1 1
use contact_9  contact_9_448
timestamp 1624857261
transform 1 0 119411 0 1 133029
box 0 0 1 1
use contact_9  contact_9_447
timestamp 1624857261
transform 1 0 124403 0 1 133029
box 0 0 1 1
use contact_9  contact_9_446
timestamp 1624857261
transform 1 0 129395 0 1 133029
box 0 0 1 1
use contact_9  contact_9_445
timestamp 1624857261
transform 1 0 134387 0 1 133029
box 0 0 1 1
use contact_9  contact_9_444
timestamp 1624857261
transform 1 0 139379 0 1 133029
box 0 0 1 1
use contact_9  contact_9_443
timestamp 1624857261
transform 1 0 144371 0 1 133029
box 0 0 1 1
use contact_9  contact_9_442
timestamp 1624857261
transform 1 0 149363 0 1 133029
box 0 0 1 1
use contact_9  contact_9_441
timestamp 1624857261
transform 1 0 154355 0 1 133029
box 0 0 1 1
use contact_9  contact_9_440
timestamp 1624857261
transform 1 0 159347 0 1 133029
box 0 0 1 1
use contact_9  contact_9_439
timestamp 1624857261
transform 1 0 164339 0 1 133029
box 0 0 1 1
use contact_9  contact_9_438
timestamp 1624857261
transform 1 0 169331 0 1 133029
box 0 0 1 1
use contact_9  contact_9_437
timestamp 1624857261
transform 1 0 174323 0 1 133029
box 0 0 1 1
use contact_9  contact_9_436
timestamp 1624857261
transform 1 0 179315 0 1 133029
box 0 0 1 1
use contact_9  contact_9_435
timestamp 1624857261
transform 1 0 184307 0 1 133029
box 0 0 1 1
use contact_9  contact_9_434
timestamp 1624857261
transform 1 0 200973 0 1 141407
box 0 0 1 1
use contact_9  contact_9_433
timestamp 1624857261
transform 1 0 199805 0 1 141407
box 0 0 1 1
use contact_9  contact_9_432
timestamp 1624857261
transform 1 0 198637 0 1 141407
box 0 0 1 1
use contact_9  contact_9_431
timestamp 1624857261
transform 1 0 204477 0 1 24236
box 0 0 1 1
use contact_9  contact_9_430
timestamp 1624857261
transform 1 0 204477 0 1 22536
box 0 0 1 1
use contact_9  contact_9_429
timestamp 1624857261
transform 1 0 204477 0 1 21408
box 0 0 1 1
use contact_9  contact_9_428
timestamp 1624857261
transform 1 0 204477 0 1 19708
box 0 0 1 1
use contact_9  contact_9_427
timestamp 1624857261
transform 1 0 204477 0 1 18580
box 0 0 1 1
use contact_9  contact_9_426
timestamp 1624857261
transform 1 0 204477 0 1 16880
box 0 0 1 1
use contact_9  contact_9_425
timestamp 1624857261
transform 1 0 204477 0 1 15752
box 0 0 1 1
use contact_9  contact_9_424
timestamp 1624857261
transform 1 0 204477 0 1 14052
box 0 0 1 1
use contact_9  contact_9_423
timestamp 1624857261
transform 1 0 2033 0 1 1811
box 0 0 1 1
use contact_9  contact_9_422
timestamp 1624857261
transform 1 0 3713 0 1 1811
box 0 0 1 1
use contact_9  contact_9_421
timestamp 1624857261
transform 1 0 5393 0 1 1811
box 0 0 1 1
use contact_9  contact_9_420
timestamp 1624857261
transform 1 0 7073 0 1 1811
box 0 0 1 1
use contact_9  contact_9_419
timestamp 1624857261
transform 1 0 8753 0 1 1811
box 0 0 1 1
use contact_9  contact_9_418
timestamp 1624857261
transform 1 0 10433 0 1 1811
box 0 0 1 1
use contact_9  contact_9_417
timestamp 1624857261
transform 1 0 12113 0 1 1811
box 0 0 1 1
use contact_9  contact_9_416
timestamp 1624857261
transform 1 0 13793 0 1 1811
box 0 0 1 1
use contact_9  contact_9_415
timestamp 1624857261
transform 1 0 15473 0 1 1811
box 0 0 1 1
use contact_9  contact_9_414
timestamp 1624857261
transform 1 0 17153 0 1 1811
box 0 0 1 1
use contact_9  contact_9_413
timestamp 1624857261
transform 1 0 18833 0 1 1811
box 0 0 1 1
use contact_9  contact_9_412
timestamp 1624857261
transform 1 0 20513 0 1 1811
box 0 0 1 1
use contact_9  contact_9_411
timestamp 1624857261
transform 1 0 22193 0 1 1811
box 0 0 1 1
use contact_9  contact_9_410
timestamp 1624857261
transform 1 0 23873 0 1 1811
box 0 0 1 1
use contact_9  contact_9_409
timestamp 1624857261
transform 1 0 25553 0 1 1811
box 0 0 1 1
use contact_9  contact_9_408
timestamp 1624857261
transform 1 0 27233 0 1 1811
box 0 0 1 1
use contact_9  contact_9_407
timestamp 1624857261
transform 1 0 28913 0 1 1811
box 0 0 1 1
use contact_9  contact_9_406
timestamp 1624857261
transform 1 0 30593 0 1 1811
box 0 0 1 1
use contact_9  contact_9_405
timestamp 1624857261
transform 1 0 32273 0 1 1811
box 0 0 1 1
use contact_9  contact_9_404
timestamp 1624857261
transform 1 0 33953 0 1 1811
box 0 0 1 1
use contact_9  contact_9_403
timestamp 1624857261
transform 1 0 35633 0 1 1811
box 0 0 1 1
use contact_9  contact_9_402
timestamp 1624857261
transform 1 0 37313 0 1 1811
box 0 0 1 1
use contact_9  contact_9_401
timestamp 1624857261
transform 1 0 38993 0 1 1811
box 0 0 1 1
use contact_9  contact_9_400
timestamp 1624857261
transform 1 0 40673 0 1 1811
box 0 0 1 1
use contact_9  contact_9_399
timestamp 1624857261
transform 1 0 42353 0 1 1811
box 0 0 1 1
use contact_9  contact_9_398
timestamp 1624857261
transform 1 0 44033 0 1 1811
box 0 0 1 1
use contact_9  contact_9_397
timestamp 1624857261
transform 1 0 45713 0 1 1811
box 0 0 1 1
use contact_9  contact_9_396
timestamp 1624857261
transform 1 0 47393 0 1 1811
box 0 0 1 1
use contact_9  contact_9_395
timestamp 1624857261
transform 1 0 49073 0 1 1811
box 0 0 1 1
use contact_9  contact_9_394
timestamp 1624857261
transform 1 0 50753 0 1 1811
box 0 0 1 1
use contact_9  contact_9_393
timestamp 1624857261
transform 1 0 52433 0 1 1811
box 0 0 1 1
use contact_9  contact_9_392
timestamp 1624857261
transform 1 0 54113 0 1 1811
box 0 0 1 1
use contact_9  contact_9_391
timestamp 1624857261
transform 1 0 55793 0 1 1811
box 0 0 1 1
use contact_9  contact_9_390
timestamp 1624857261
transform 1 0 57473 0 1 1811
box 0 0 1 1
use contact_9  contact_9_389
timestamp 1624857261
transform 1 0 59153 0 1 1811
box 0 0 1 1
use contact_9  contact_9_388
timestamp 1624857261
transform 1 0 60833 0 1 1811
box 0 0 1 1
use contact_9  contact_9_387
timestamp 1624857261
transform 1 0 62513 0 1 1811
box 0 0 1 1
use contact_9  contact_9_386
timestamp 1624857261
transform 1 0 64193 0 1 1811
box 0 0 1 1
use contact_9  contact_9_385
timestamp 1624857261
transform 1 0 65873 0 1 1811
box 0 0 1 1
use contact_9  contact_9_384
timestamp 1624857261
transform 1 0 67553 0 1 1811
box 0 0 1 1
use contact_9  contact_9_383
timestamp 1624857261
transform 1 0 69233 0 1 1811
box 0 0 1 1
use contact_9  contact_9_382
timestamp 1624857261
transform 1 0 70913 0 1 1811
box 0 0 1 1
use contact_9  contact_9_381
timestamp 1624857261
transform 1 0 72593 0 1 1811
box 0 0 1 1
use contact_9  contact_9_380
timestamp 1624857261
transform 1 0 74273 0 1 1811
box 0 0 1 1
use contact_9  contact_9_379
timestamp 1624857261
transform 1 0 75953 0 1 1811
box 0 0 1 1
use contact_9  contact_9_378
timestamp 1624857261
transform 1 0 77633 0 1 1811
box 0 0 1 1
use contact_9  contact_9_377
timestamp 1624857261
transform 1 0 79313 0 1 1811
box 0 0 1 1
use contact_9  contact_9_376
timestamp 1624857261
transform 1 0 80993 0 1 1811
box 0 0 1 1
use contact_9  contact_9_375
timestamp 1624857261
transform 1 0 82673 0 1 1811
box 0 0 1 1
use contact_9  contact_9_374
timestamp 1624857261
transform 1 0 84353 0 1 1811
box 0 0 1 1
use contact_9  contact_9_373
timestamp 1624857261
transform 1 0 86033 0 1 1811
box 0 0 1 1
use contact_9  contact_9_372
timestamp 1624857261
transform 1 0 87713 0 1 1811
box 0 0 1 1
use contact_9  contact_9_371
timestamp 1624857261
transform 1 0 89393 0 1 1811
box 0 0 1 1
use contact_9  contact_9_370
timestamp 1624857261
transform 1 0 91073 0 1 1811
box 0 0 1 1
use contact_9  contact_9_369
timestamp 1624857261
transform 1 0 92753 0 1 1811
box 0 0 1 1
use contact_9  contact_9_368
timestamp 1624857261
transform 1 0 94433 0 1 1811
box 0 0 1 1
use contact_9  contact_9_367
timestamp 1624857261
transform 1 0 96113 0 1 1811
box 0 0 1 1
use contact_9  contact_9_366
timestamp 1624857261
transform 1 0 97793 0 1 1811
box 0 0 1 1
use contact_9  contact_9_365
timestamp 1624857261
transform 1 0 99473 0 1 1811
box 0 0 1 1
use contact_9  contact_9_364
timestamp 1624857261
transform 1 0 101153 0 1 1811
box 0 0 1 1
use contact_9  contact_9_363
timestamp 1624857261
transform 1 0 102833 0 1 1811
box 0 0 1 1
use contact_9  contact_9_362
timestamp 1624857261
transform 1 0 104513 0 1 1811
box 0 0 1 1
use contact_9  contact_9_361
timestamp 1624857261
transform 1 0 106193 0 1 1811
box 0 0 1 1
use contact_9  contact_9_360
timestamp 1624857261
transform 1 0 107873 0 1 1811
box 0 0 1 1
use contact_9  contact_9_359
timestamp 1624857261
transform 1 0 109553 0 1 1811
box 0 0 1 1
use contact_9  contact_9_358
timestamp 1624857261
transform 1 0 111233 0 1 1811
box 0 0 1 1
use contact_9  contact_9_357
timestamp 1624857261
transform 1 0 112913 0 1 1811
box 0 0 1 1
use contact_9  contact_9_356
timestamp 1624857261
transform 1 0 114593 0 1 1811
box 0 0 1 1
use contact_9  contact_9_355
timestamp 1624857261
transform 1 0 116273 0 1 1811
box 0 0 1 1
use contact_9  contact_9_354
timestamp 1624857261
transform 1 0 117953 0 1 1811
box 0 0 1 1
use contact_9  contact_9_353
timestamp 1624857261
transform 1 0 119633 0 1 1811
box 0 0 1 1
use contact_9  contact_9_352
timestamp 1624857261
transform 1 0 121313 0 1 1811
box 0 0 1 1
use contact_9  contact_9_351
timestamp 1624857261
transform 1 0 122993 0 1 1811
box 0 0 1 1
use contact_9  contact_9_350
timestamp 1624857261
transform 1 0 124673 0 1 1811
box 0 0 1 1
use contact_9  contact_9_349
timestamp 1624857261
transform 1 0 126353 0 1 1811
box 0 0 1 1
use contact_9  contact_9_348
timestamp 1624857261
transform 1 0 128033 0 1 1811
box 0 0 1 1
use contact_9  contact_9_347
timestamp 1624857261
transform 1 0 129713 0 1 1811
box 0 0 1 1
use contact_9  contact_9_346
timestamp 1624857261
transform 1 0 131393 0 1 1811
box 0 0 1 1
use contact_9  contact_9_345
timestamp 1624857261
transform 1 0 133073 0 1 1811
box 0 0 1 1
use contact_9  contact_9_344
timestamp 1624857261
transform 1 0 134753 0 1 1811
box 0 0 1 1
use contact_9  contact_9_343
timestamp 1624857261
transform 1 0 136433 0 1 1811
box 0 0 1 1
use contact_9  contact_9_342
timestamp 1624857261
transform 1 0 138113 0 1 1811
box 0 0 1 1
use contact_9  contact_9_341
timestamp 1624857261
transform 1 0 139793 0 1 1811
box 0 0 1 1
use contact_9  contact_9_340
timestamp 1624857261
transform 1 0 141473 0 1 1811
box 0 0 1 1
use contact_9  contact_9_339
timestamp 1624857261
transform 1 0 143153 0 1 1811
box 0 0 1 1
use contact_9  contact_9_338
timestamp 1624857261
transform 1 0 144833 0 1 1811
box 0 0 1 1
use contact_9  contact_9_337
timestamp 1624857261
transform 1 0 146513 0 1 1811
box 0 0 1 1
use contact_9  contact_9_336
timestamp 1624857261
transform 1 0 148193 0 1 1811
box 0 0 1 1
use contact_9  contact_9_335
timestamp 1624857261
transform 1 0 149873 0 1 1811
box 0 0 1 1
use contact_9  contact_9_334
timestamp 1624857261
transform 1 0 151553 0 1 1811
box 0 0 1 1
use contact_9  contact_9_333
timestamp 1624857261
transform 1 0 153233 0 1 1811
box 0 0 1 1
use contact_9  contact_9_332
timestamp 1624857261
transform 1 0 154913 0 1 1811
box 0 0 1 1
use contact_9  contact_9_331
timestamp 1624857261
transform 1 0 156593 0 1 1811
box 0 0 1 1
use contact_9  contact_9_330
timestamp 1624857261
transform 1 0 158273 0 1 1811
box 0 0 1 1
use contact_9  contact_9_329
timestamp 1624857261
transform 1 0 159953 0 1 1811
box 0 0 1 1
use contact_9  contact_9_328
timestamp 1624857261
transform 1 0 161633 0 1 1811
box 0 0 1 1
use contact_9  contact_9_327
timestamp 1624857261
transform 1 0 163313 0 1 1811
box 0 0 1 1
use contact_9  contact_9_326
timestamp 1624857261
transform 1 0 164993 0 1 1811
box 0 0 1 1
use contact_9  contact_9_325
timestamp 1624857261
transform 1 0 166673 0 1 1811
box 0 0 1 1
use contact_9  contact_9_324
timestamp 1624857261
transform 1 0 168353 0 1 1811
box 0 0 1 1
use contact_9  contact_9_323
timestamp 1624857261
transform 1 0 170033 0 1 1811
box 0 0 1 1
use contact_9  contact_9_322
timestamp 1624857261
transform 1 0 171713 0 1 1811
box 0 0 1 1
use contact_9  contact_9_321
timestamp 1624857261
transform 1 0 173393 0 1 1811
box 0 0 1 1
use contact_9  contact_9_320
timestamp 1624857261
transform 1 0 175073 0 1 1811
box 0 0 1 1
use contact_9  contact_9_319
timestamp 1624857261
transform 1 0 176753 0 1 1811
box 0 0 1 1
use contact_9  contact_9_318
timestamp 1624857261
transform 1 0 178433 0 1 1811
box 0 0 1 1
use contact_9  contact_9_317
timestamp 1624857261
transform 1 0 180113 0 1 1811
box 0 0 1 1
use contact_9  contact_9_316
timestamp 1624857261
transform 1 0 181793 0 1 1811
box 0 0 1 1
use contact_9  contact_9_315
timestamp 1624857261
transform 1 0 183473 0 1 1811
box 0 0 1 1
use contact_9  contact_9_314
timestamp 1624857261
transform 1 0 185153 0 1 1811
box 0 0 1 1
use contact_9  contact_9_313
timestamp 1624857261
transform 1 0 186833 0 1 1811
box 0 0 1 1
use contact_9  contact_9_312
timestamp 1624857261
transform 1 0 188513 0 1 1811
box 0 0 1 1
use contact_9  contact_9_311
timestamp 1624857261
transform 1 0 190193 0 1 1811
box 0 0 1 1
use contact_9  contact_9_310
timestamp 1624857261
transform 1 0 191873 0 1 1811
box 0 0 1 1
use contact_9  contact_9_309
timestamp 1624857261
transform 1 0 193553 0 1 1811
box 0 0 1 1
use contact_9  contact_9_308
timestamp 1624857261
transform 1 0 195233 0 1 1811
box 0 0 1 1
use contact_9  contact_9_307
timestamp 1624857261
transform 1 0 196913 0 1 1811
box 0 0 1 1
use contact_9  contact_9_306
timestamp 1624857261
transform 1 0 198593 0 1 1811
box 0 0 1 1
use contact_9  contact_9_305
timestamp 1624857261
transform 1 0 200273 0 1 1811
box 0 0 1 1
use contact_9  contact_9_304
timestamp 1624857261
transform 1 0 201953 0 1 1811
box 0 0 1 1
use contact_9  contact_9_303
timestamp 1624857261
transform 1 0 203633 0 1 1811
box 0 0 1 1
use contact_9  contact_9_302
timestamp 1624857261
transform 1 0 205313 0 1 1811
box 0 0 1 1
use contact_9  contact_9_301
timestamp 1624857261
transform 1 0 206993 0 1 1811
box 0 0 1 1
use contact_9  contact_9_300
timestamp 1624857261
transform 1 0 208673 0 1 1811
box 0 0 1 1
use contact_9  contact_9_299
timestamp 1624857261
transform 1 0 210353 0 1 1811
box 0 0 1 1
use contact_9  contact_9_298
timestamp 1624857261
transform 1 0 212033 0 1 1811
box 0 0 1 1
use contact_9  contact_9_297
timestamp 1624857261
transform 1 0 213713 0 1 1811
box 0 0 1 1
use contact_9  contact_9_296
timestamp 1624857261
transform 1 0 215393 0 1 1811
box 0 0 1 1
use contact_9  contact_9_295
timestamp 1624857261
transform 1 0 2033 0 1 142307
box 0 0 1 1
use contact_9  contact_9_294
timestamp 1624857261
transform 1 0 3713 0 1 142307
box 0 0 1 1
use contact_9  contact_9_293
timestamp 1624857261
transform 1 0 5393 0 1 142307
box 0 0 1 1
use contact_9  contact_9_292
timestamp 1624857261
transform 1 0 7073 0 1 142307
box 0 0 1 1
use contact_9  contact_9_291
timestamp 1624857261
transform 1 0 8753 0 1 142307
box 0 0 1 1
use contact_9  contact_9_290
timestamp 1624857261
transform 1 0 10433 0 1 142307
box 0 0 1 1
use contact_9  contact_9_289
timestamp 1624857261
transform 1 0 12113 0 1 142307
box 0 0 1 1
use contact_9  contact_9_288
timestamp 1624857261
transform 1 0 13793 0 1 142307
box 0 0 1 1
use contact_9  contact_9_287
timestamp 1624857261
transform 1 0 15473 0 1 142307
box 0 0 1 1
use contact_9  contact_9_286
timestamp 1624857261
transform 1 0 17153 0 1 142307
box 0 0 1 1
use contact_9  contact_9_285
timestamp 1624857261
transform 1 0 18833 0 1 142307
box 0 0 1 1
use contact_9  contact_9_284
timestamp 1624857261
transform 1 0 20513 0 1 142307
box 0 0 1 1
use contact_9  contact_9_283
timestamp 1624857261
transform 1 0 22193 0 1 142307
box 0 0 1 1
use contact_9  contact_9_282
timestamp 1624857261
transform 1 0 23873 0 1 142307
box 0 0 1 1
use contact_9  contact_9_281
timestamp 1624857261
transform 1 0 25553 0 1 142307
box 0 0 1 1
use contact_9  contact_9_280
timestamp 1624857261
transform 1 0 27233 0 1 142307
box 0 0 1 1
use contact_9  contact_9_279
timestamp 1624857261
transform 1 0 28913 0 1 142307
box 0 0 1 1
use contact_9  contact_9_278
timestamp 1624857261
transform 1 0 30593 0 1 142307
box 0 0 1 1
use contact_9  contact_9_277
timestamp 1624857261
transform 1 0 32273 0 1 142307
box 0 0 1 1
use contact_9  contact_9_276
timestamp 1624857261
transform 1 0 33953 0 1 142307
box 0 0 1 1
use contact_9  contact_9_275
timestamp 1624857261
transform 1 0 35633 0 1 142307
box 0 0 1 1
use contact_9  contact_9_274
timestamp 1624857261
transform 1 0 37313 0 1 142307
box 0 0 1 1
use contact_9  contact_9_273
timestamp 1624857261
transform 1 0 38993 0 1 142307
box 0 0 1 1
use contact_9  contact_9_272
timestamp 1624857261
transform 1 0 40673 0 1 142307
box 0 0 1 1
use contact_9  contact_9_271
timestamp 1624857261
transform 1 0 42353 0 1 142307
box 0 0 1 1
use contact_9  contact_9_270
timestamp 1624857261
transform 1 0 44033 0 1 142307
box 0 0 1 1
use contact_9  contact_9_269
timestamp 1624857261
transform 1 0 45713 0 1 142307
box 0 0 1 1
use contact_9  contact_9_268
timestamp 1624857261
transform 1 0 47393 0 1 142307
box 0 0 1 1
use contact_9  contact_9_267
timestamp 1624857261
transform 1 0 49073 0 1 142307
box 0 0 1 1
use contact_9  contact_9_266
timestamp 1624857261
transform 1 0 50753 0 1 142307
box 0 0 1 1
use contact_9  contact_9_265
timestamp 1624857261
transform 1 0 52433 0 1 142307
box 0 0 1 1
use contact_9  contact_9_264
timestamp 1624857261
transform 1 0 54113 0 1 142307
box 0 0 1 1
use contact_9  contact_9_263
timestamp 1624857261
transform 1 0 55793 0 1 142307
box 0 0 1 1
use contact_9  contact_9_262
timestamp 1624857261
transform 1 0 57473 0 1 142307
box 0 0 1 1
use contact_9  contact_9_261
timestamp 1624857261
transform 1 0 59153 0 1 142307
box 0 0 1 1
use contact_9  contact_9_260
timestamp 1624857261
transform 1 0 60833 0 1 142307
box 0 0 1 1
use contact_9  contact_9_259
timestamp 1624857261
transform 1 0 62513 0 1 142307
box 0 0 1 1
use contact_9  contact_9_258
timestamp 1624857261
transform 1 0 64193 0 1 142307
box 0 0 1 1
use contact_9  contact_9_257
timestamp 1624857261
transform 1 0 65873 0 1 142307
box 0 0 1 1
use contact_9  contact_9_256
timestamp 1624857261
transform 1 0 67553 0 1 142307
box 0 0 1 1
use contact_9  contact_9_255
timestamp 1624857261
transform 1 0 69233 0 1 142307
box 0 0 1 1
use contact_9  contact_9_254
timestamp 1624857261
transform 1 0 70913 0 1 142307
box 0 0 1 1
use contact_9  contact_9_253
timestamp 1624857261
transform 1 0 72593 0 1 142307
box 0 0 1 1
use contact_9  contact_9_252
timestamp 1624857261
transform 1 0 74273 0 1 142307
box 0 0 1 1
use contact_9  contact_9_251
timestamp 1624857261
transform 1 0 75953 0 1 142307
box 0 0 1 1
use contact_9  contact_9_250
timestamp 1624857261
transform 1 0 77633 0 1 142307
box 0 0 1 1
use contact_9  contact_9_249
timestamp 1624857261
transform 1 0 79313 0 1 142307
box 0 0 1 1
use contact_9  contact_9_248
timestamp 1624857261
transform 1 0 80993 0 1 142307
box 0 0 1 1
use contact_9  contact_9_247
timestamp 1624857261
transform 1 0 82673 0 1 142307
box 0 0 1 1
use contact_9  contact_9_246
timestamp 1624857261
transform 1 0 84353 0 1 142307
box 0 0 1 1
use contact_9  contact_9_245
timestamp 1624857261
transform 1 0 86033 0 1 142307
box 0 0 1 1
use contact_9  contact_9_244
timestamp 1624857261
transform 1 0 87713 0 1 142307
box 0 0 1 1
use contact_9  contact_9_243
timestamp 1624857261
transform 1 0 89393 0 1 142307
box 0 0 1 1
use contact_9  contact_9_242
timestamp 1624857261
transform 1 0 91073 0 1 142307
box 0 0 1 1
use contact_9  contact_9_241
timestamp 1624857261
transform 1 0 92753 0 1 142307
box 0 0 1 1
use contact_9  contact_9_240
timestamp 1624857261
transform 1 0 94433 0 1 142307
box 0 0 1 1
use contact_9  contact_9_239
timestamp 1624857261
transform 1 0 96113 0 1 142307
box 0 0 1 1
use contact_9  contact_9_238
timestamp 1624857261
transform 1 0 97793 0 1 142307
box 0 0 1 1
use contact_9  contact_9_237
timestamp 1624857261
transform 1 0 99473 0 1 142307
box 0 0 1 1
use contact_9  contact_9_236
timestamp 1624857261
transform 1 0 101153 0 1 142307
box 0 0 1 1
use contact_9  contact_9_235
timestamp 1624857261
transform 1 0 102833 0 1 142307
box 0 0 1 1
use contact_9  contact_9_234
timestamp 1624857261
transform 1 0 104513 0 1 142307
box 0 0 1 1
use contact_9  contact_9_233
timestamp 1624857261
transform 1 0 106193 0 1 142307
box 0 0 1 1
use contact_9  contact_9_232
timestamp 1624857261
transform 1 0 107873 0 1 142307
box 0 0 1 1
use contact_9  contact_9_231
timestamp 1624857261
transform 1 0 109553 0 1 142307
box 0 0 1 1
use contact_9  contact_9_230
timestamp 1624857261
transform 1 0 111233 0 1 142307
box 0 0 1 1
use contact_9  contact_9_229
timestamp 1624857261
transform 1 0 112913 0 1 142307
box 0 0 1 1
use contact_9  contact_9_228
timestamp 1624857261
transform 1 0 114593 0 1 142307
box 0 0 1 1
use contact_9  contact_9_227
timestamp 1624857261
transform 1 0 116273 0 1 142307
box 0 0 1 1
use contact_9  contact_9_226
timestamp 1624857261
transform 1 0 117953 0 1 142307
box 0 0 1 1
use contact_9  contact_9_225
timestamp 1624857261
transform 1 0 119633 0 1 142307
box 0 0 1 1
use contact_9  contact_9_224
timestamp 1624857261
transform 1 0 121313 0 1 142307
box 0 0 1 1
use contact_9  contact_9_223
timestamp 1624857261
transform 1 0 122993 0 1 142307
box 0 0 1 1
use contact_9  contact_9_222
timestamp 1624857261
transform 1 0 124673 0 1 142307
box 0 0 1 1
use contact_9  contact_9_221
timestamp 1624857261
transform 1 0 126353 0 1 142307
box 0 0 1 1
use contact_9  contact_9_220
timestamp 1624857261
transform 1 0 128033 0 1 142307
box 0 0 1 1
use contact_9  contact_9_219
timestamp 1624857261
transform 1 0 129713 0 1 142307
box 0 0 1 1
use contact_9  contact_9_218
timestamp 1624857261
transform 1 0 131393 0 1 142307
box 0 0 1 1
use contact_9  contact_9_217
timestamp 1624857261
transform 1 0 133073 0 1 142307
box 0 0 1 1
use contact_9  contact_9_216
timestamp 1624857261
transform 1 0 134753 0 1 142307
box 0 0 1 1
use contact_9  contact_9_215
timestamp 1624857261
transform 1 0 136433 0 1 142307
box 0 0 1 1
use contact_9  contact_9_214
timestamp 1624857261
transform 1 0 138113 0 1 142307
box 0 0 1 1
use contact_9  contact_9_213
timestamp 1624857261
transform 1 0 139793 0 1 142307
box 0 0 1 1
use contact_9  contact_9_212
timestamp 1624857261
transform 1 0 141473 0 1 142307
box 0 0 1 1
use contact_9  contact_9_211
timestamp 1624857261
transform 1 0 143153 0 1 142307
box 0 0 1 1
use contact_9  contact_9_210
timestamp 1624857261
transform 1 0 144833 0 1 142307
box 0 0 1 1
use contact_9  contact_9_209
timestamp 1624857261
transform 1 0 146513 0 1 142307
box 0 0 1 1
use contact_9  contact_9_208
timestamp 1624857261
transform 1 0 148193 0 1 142307
box 0 0 1 1
use contact_9  contact_9_207
timestamp 1624857261
transform 1 0 149873 0 1 142307
box 0 0 1 1
use contact_9  contact_9_206
timestamp 1624857261
transform 1 0 151553 0 1 142307
box 0 0 1 1
use contact_9  contact_9_205
timestamp 1624857261
transform 1 0 153233 0 1 142307
box 0 0 1 1
use contact_9  contact_9_204
timestamp 1624857261
transform 1 0 154913 0 1 142307
box 0 0 1 1
use contact_9  contact_9_203
timestamp 1624857261
transform 1 0 156593 0 1 142307
box 0 0 1 1
use contact_9  contact_9_202
timestamp 1624857261
transform 1 0 158273 0 1 142307
box 0 0 1 1
use contact_9  contact_9_201
timestamp 1624857261
transform 1 0 159953 0 1 142307
box 0 0 1 1
use contact_9  contact_9_200
timestamp 1624857261
transform 1 0 161633 0 1 142307
box 0 0 1 1
use contact_9  contact_9_199
timestamp 1624857261
transform 1 0 163313 0 1 142307
box 0 0 1 1
use contact_9  contact_9_198
timestamp 1624857261
transform 1 0 164993 0 1 142307
box 0 0 1 1
use contact_9  contact_9_197
timestamp 1624857261
transform 1 0 166673 0 1 142307
box 0 0 1 1
use contact_9  contact_9_196
timestamp 1624857261
transform 1 0 168353 0 1 142307
box 0 0 1 1
use contact_9  contact_9_195
timestamp 1624857261
transform 1 0 170033 0 1 142307
box 0 0 1 1
use contact_9  contact_9_194
timestamp 1624857261
transform 1 0 171713 0 1 142307
box 0 0 1 1
use contact_9  contact_9_193
timestamp 1624857261
transform 1 0 173393 0 1 142307
box 0 0 1 1
use contact_9  contact_9_192
timestamp 1624857261
transform 1 0 175073 0 1 142307
box 0 0 1 1
use contact_9  contact_9_191
timestamp 1624857261
transform 1 0 176753 0 1 142307
box 0 0 1 1
use contact_9  contact_9_190
timestamp 1624857261
transform 1 0 178433 0 1 142307
box 0 0 1 1
use contact_9  contact_9_189
timestamp 1624857261
transform 1 0 180113 0 1 142307
box 0 0 1 1
use contact_9  contact_9_188
timestamp 1624857261
transform 1 0 181793 0 1 142307
box 0 0 1 1
use contact_9  contact_9_187
timestamp 1624857261
transform 1 0 183473 0 1 142307
box 0 0 1 1
use contact_9  contact_9_186
timestamp 1624857261
transform 1 0 185153 0 1 142307
box 0 0 1 1
use contact_9  contact_9_185
timestamp 1624857261
transform 1 0 186833 0 1 142307
box 0 0 1 1
use contact_9  contact_9_184
timestamp 1624857261
transform 1 0 188513 0 1 142307
box 0 0 1 1
use contact_9  contact_9_183
timestamp 1624857261
transform 1 0 190193 0 1 142307
box 0 0 1 1
use contact_9  contact_9_182
timestamp 1624857261
transform 1 0 191873 0 1 142307
box 0 0 1 1
use contact_9  contact_9_181
timestamp 1624857261
transform 1 0 193553 0 1 142307
box 0 0 1 1
use contact_9  contact_9_180
timestamp 1624857261
transform 1 0 195233 0 1 142307
box 0 0 1 1
use contact_9  contact_9_179
timestamp 1624857261
transform 1 0 196913 0 1 142307
box 0 0 1 1
use contact_9  contact_9_178
timestamp 1624857261
transform 1 0 198593 0 1 142307
box 0 0 1 1
use contact_9  contact_9_177
timestamp 1624857261
transform 1 0 200273 0 1 142307
box 0 0 1 1
use contact_9  contact_9_176
timestamp 1624857261
transform 1 0 201953 0 1 142307
box 0 0 1 1
use contact_9  contact_9_175
timestamp 1624857261
transform 1 0 203633 0 1 142307
box 0 0 1 1
use contact_9  contact_9_174
timestamp 1624857261
transform 1 0 205313 0 1 142307
box 0 0 1 1
use contact_9  contact_9_173
timestamp 1624857261
transform 1 0 206993 0 1 142307
box 0 0 1 1
use contact_9  contact_9_172
timestamp 1624857261
transform 1 0 208673 0 1 142307
box 0 0 1 1
use contact_9  contact_9_171
timestamp 1624857261
transform 1 0 210353 0 1 142307
box 0 0 1 1
use contact_9  contact_9_170
timestamp 1624857261
transform 1 0 212033 0 1 142307
box 0 0 1 1
use contact_9  contact_9_169
timestamp 1624857261
transform 1 0 213713 0 1 142307
box 0 0 1 1
use contact_9  contact_9_168
timestamp 1624857261
transform 1 0 215393 0 1 142307
box 0 0 1 1
use contact_9  contact_9_167
timestamp 1624857261
transform 1 0 1697 0 1 2147
box 0 0 1 1
use contact_9  contact_9_166
timestamp 1624857261
transform 1 0 1697 0 1 3827
box 0 0 1 1
use contact_9  contact_9_165
timestamp 1624857261
transform 1 0 1697 0 1 5507
box 0 0 1 1
use contact_9  contact_9_164
timestamp 1624857261
transform 1 0 1697 0 1 7187
box 0 0 1 1
use contact_9  contact_9_163
timestamp 1624857261
transform 1 0 1697 0 1 8867
box 0 0 1 1
use contact_9  contact_9_162
timestamp 1624857261
transform 1 0 1697 0 1 10547
box 0 0 1 1
use contact_9  contact_9_161
timestamp 1624857261
transform 1 0 1697 0 1 12227
box 0 0 1 1
use contact_9  contact_9_160
timestamp 1624857261
transform 1 0 1697 0 1 13907
box 0 0 1 1
use contact_9  contact_9_159
timestamp 1624857261
transform 1 0 1697 0 1 15587
box 0 0 1 1
use contact_9  contact_9_158
timestamp 1624857261
transform 1 0 1697 0 1 17267
box 0 0 1 1
use contact_9  contact_9_157
timestamp 1624857261
transform 1 0 1697 0 1 18947
box 0 0 1 1
use contact_9  contact_9_156
timestamp 1624857261
transform 1 0 1697 0 1 20627
box 0 0 1 1
use contact_9  contact_9_155
timestamp 1624857261
transform 1 0 1697 0 1 22307
box 0 0 1 1
use contact_9  contact_9_154
timestamp 1624857261
transform 1 0 1697 0 1 23987
box 0 0 1 1
use contact_9  contact_9_153
timestamp 1624857261
transform 1 0 1697 0 1 25667
box 0 0 1 1
use contact_9  contact_9_152
timestamp 1624857261
transform 1 0 1697 0 1 27347
box 0 0 1 1
use contact_9  contact_9_151
timestamp 1624857261
transform 1 0 1697 0 1 29027
box 0 0 1 1
use contact_9  contact_9_150
timestamp 1624857261
transform 1 0 1697 0 1 30707
box 0 0 1 1
use contact_9  contact_9_149
timestamp 1624857261
transform 1 0 1697 0 1 32387
box 0 0 1 1
use contact_9  contact_9_148
timestamp 1624857261
transform 1 0 1697 0 1 34067
box 0 0 1 1
use contact_9  contact_9_147
timestamp 1624857261
transform 1 0 1697 0 1 35747
box 0 0 1 1
use contact_9  contact_9_146
timestamp 1624857261
transform 1 0 1697 0 1 37427
box 0 0 1 1
use contact_9  contact_9_145
timestamp 1624857261
transform 1 0 1697 0 1 39107
box 0 0 1 1
use contact_9  contact_9_144
timestamp 1624857261
transform 1 0 1697 0 1 40787
box 0 0 1 1
use contact_9  contact_9_143
timestamp 1624857261
transform 1 0 1697 0 1 42467
box 0 0 1 1
use contact_9  contact_9_142
timestamp 1624857261
transform 1 0 1697 0 1 44147
box 0 0 1 1
use contact_9  contact_9_141
timestamp 1624857261
transform 1 0 1697 0 1 45827
box 0 0 1 1
use contact_9  contact_9_140
timestamp 1624857261
transform 1 0 1697 0 1 47507
box 0 0 1 1
use contact_9  contact_9_139
timestamp 1624857261
transform 1 0 1697 0 1 49187
box 0 0 1 1
use contact_9  contact_9_138
timestamp 1624857261
transform 1 0 1697 0 1 50867
box 0 0 1 1
use contact_9  contact_9_137
timestamp 1624857261
transform 1 0 1697 0 1 52547
box 0 0 1 1
use contact_9  contact_9_136
timestamp 1624857261
transform 1 0 1697 0 1 54227
box 0 0 1 1
use contact_9  contact_9_135
timestamp 1624857261
transform 1 0 1697 0 1 55907
box 0 0 1 1
use contact_9  contact_9_134
timestamp 1624857261
transform 1 0 1697 0 1 57587
box 0 0 1 1
use contact_9  contact_9_133
timestamp 1624857261
transform 1 0 1697 0 1 59267
box 0 0 1 1
use contact_9  contact_9_132
timestamp 1624857261
transform 1 0 1697 0 1 60947
box 0 0 1 1
use contact_9  contact_9_131
timestamp 1624857261
transform 1 0 1697 0 1 62627
box 0 0 1 1
use contact_9  contact_9_130
timestamp 1624857261
transform 1 0 1697 0 1 64307
box 0 0 1 1
use contact_9  contact_9_129
timestamp 1624857261
transform 1 0 1697 0 1 65987
box 0 0 1 1
use contact_9  contact_9_128
timestamp 1624857261
transform 1 0 1697 0 1 67667
box 0 0 1 1
use contact_9  contact_9_127
timestamp 1624857261
transform 1 0 1697 0 1 69347
box 0 0 1 1
use contact_9  contact_9_126
timestamp 1624857261
transform 1 0 1697 0 1 71027
box 0 0 1 1
use contact_9  contact_9_125
timestamp 1624857261
transform 1 0 1697 0 1 72707
box 0 0 1 1
use contact_9  contact_9_124
timestamp 1624857261
transform 1 0 1697 0 1 74387
box 0 0 1 1
use contact_9  contact_9_123
timestamp 1624857261
transform 1 0 1697 0 1 76067
box 0 0 1 1
use contact_9  contact_9_122
timestamp 1624857261
transform 1 0 1697 0 1 77747
box 0 0 1 1
use contact_9  contact_9_121
timestamp 1624857261
transform 1 0 1697 0 1 79427
box 0 0 1 1
use contact_9  contact_9_120
timestamp 1624857261
transform 1 0 1697 0 1 81107
box 0 0 1 1
use contact_9  contact_9_119
timestamp 1624857261
transform 1 0 1697 0 1 82787
box 0 0 1 1
use contact_9  contact_9_118
timestamp 1624857261
transform 1 0 1697 0 1 84467
box 0 0 1 1
use contact_9  contact_9_117
timestamp 1624857261
transform 1 0 1697 0 1 86147
box 0 0 1 1
use contact_9  contact_9_116
timestamp 1624857261
transform 1 0 1697 0 1 87827
box 0 0 1 1
use contact_9  contact_9_115
timestamp 1624857261
transform 1 0 1697 0 1 89507
box 0 0 1 1
use contact_9  contact_9_114
timestamp 1624857261
transform 1 0 1697 0 1 91187
box 0 0 1 1
use contact_9  contact_9_113
timestamp 1624857261
transform 1 0 1697 0 1 92867
box 0 0 1 1
use contact_9  contact_9_112
timestamp 1624857261
transform 1 0 1697 0 1 94547
box 0 0 1 1
use contact_9  contact_9_111
timestamp 1624857261
transform 1 0 1697 0 1 96227
box 0 0 1 1
use contact_9  contact_9_110
timestamp 1624857261
transform 1 0 1697 0 1 97907
box 0 0 1 1
use contact_9  contact_9_109
timestamp 1624857261
transform 1 0 1697 0 1 99587
box 0 0 1 1
use contact_9  contact_9_108
timestamp 1624857261
transform 1 0 1697 0 1 101267
box 0 0 1 1
use contact_9  contact_9_107
timestamp 1624857261
transform 1 0 1697 0 1 102947
box 0 0 1 1
use contact_9  contact_9_106
timestamp 1624857261
transform 1 0 1697 0 1 104627
box 0 0 1 1
use contact_9  contact_9_105
timestamp 1624857261
transform 1 0 1697 0 1 106307
box 0 0 1 1
use contact_9  contact_9_104
timestamp 1624857261
transform 1 0 1697 0 1 107987
box 0 0 1 1
use contact_9  contact_9_103
timestamp 1624857261
transform 1 0 1697 0 1 109667
box 0 0 1 1
use contact_9  contact_9_102
timestamp 1624857261
transform 1 0 1697 0 1 111347
box 0 0 1 1
use contact_9  contact_9_101
timestamp 1624857261
transform 1 0 1697 0 1 113027
box 0 0 1 1
use contact_9  contact_9_100
timestamp 1624857261
transform 1 0 1697 0 1 114707
box 0 0 1 1
use contact_9  contact_9_99
timestamp 1624857261
transform 1 0 1697 0 1 116387
box 0 0 1 1
use contact_9  contact_9_98
timestamp 1624857261
transform 1 0 1697 0 1 118067
box 0 0 1 1
use contact_9  contact_9_97
timestamp 1624857261
transform 1 0 1697 0 1 119747
box 0 0 1 1
use contact_9  contact_9_96
timestamp 1624857261
transform 1 0 1697 0 1 121427
box 0 0 1 1
use contact_9  contact_9_95
timestamp 1624857261
transform 1 0 1697 0 1 123107
box 0 0 1 1
use contact_9  contact_9_94
timestamp 1624857261
transform 1 0 1697 0 1 124787
box 0 0 1 1
use contact_9  contact_9_93
timestamp 1624857261
transform 1 0 1697 0 1 126467
box 0 0 1 1
use contact_9  contact_9_92
timestamp 1624857261
transform 1 0 1697 0 1 128147
box 0 0 1 1
use contact_9  contact_9_91
timestamp 1624857261
transform 1 0 1697 0 1 129827
box 0 0 1 1
use contact_9  contact_9_90
timestamp 1624857261
transform 1 0 1697 0 1 131507
box 0 0 1 1
use contact_9  contact_9_89
timestamp 1624857261
transform 1 0 1697 0 1 133187
box 0 0 1 1
use contact_9  contact_9_88
timestamp 1624857261
transform 1 0 1697 0 1 134867
box 0 0 1 1
use contact_9  contact_9_87
timestamp 1624857261
transform 1 0 1697 0 1 136547
box 0 0 1 1
use contact_9  contact_9_86
timestamp 1624857261
transform 1 0 1697 0 1 138227
box 0 0 1 1
use contact_9  contact_9_85
timestamp 1624857261
transform 1 0 1697 0 1 139907
box 0 0 1 1
use contact_9  contact_9_84
timestamp 1624857261
transform 1 0 1697 0 1 141587
box 0 0 1 1
use contact_9  contact_9_83
timestamp 1624857261
transform 1 0 216903 0 1 2147
box 0 0 1 1
use contact_9  contact_9_82
timestamp 1624857261
transform 1 0 216903 0 1 3827
box 0 0 1 1
use contact_9  contact_9_81
timestamp 1624857261
transform 1 0 216903 0 1 5507
box 0 0 1 1
use contact_9  contact_9_80
timestamp 1624857261
transform 1 0 216903 0 1 7187
box 0 0 1 1
use contact_9  contact_9_79
timestamp 1624857261
transform 1 0 216903 0 1 8867
box 0 0 1 1
use contact_9  contact_9_78
timestamp 1624857261
transform 1 0 216903 0 1 10547
box 0 0 1 1
use contact_9  contact_9_77
timestamp 1624857261
transform 1 0 216903 0 1 12227
box 0 0 1 1
use contact_9  contact_9_76
timestamp 1624857261
transform 1 0 216903 0 1 13907
box 0 0 1 1
use contact_9  contact_9_75
timestamp 1624857261
transform 1 0 216903 0 1 15587
box 0 0 1 1
use contact_9  contact_9_74
timestamp 1624857261
transform 1 0 216903 0 1 17267
box 0 0 1 1
use contact_9  contact_9_73
timestamp 1624857261
transform 1 0 216903 0 1 18947
box 0 0 1 1
use contact_9  contact_9_72
timestamp 1624857261
transform 1 0 216903 0 1 20627
box 0 0 1 1
use contact_9  contact_9_71
timestamp 1624857261
transform 1 0 216903 0 1 22307
box 0 0 1 1
use contact_9  contact_9_70
timestamp 1624857261
transform 1 0 216903 0 1 23987
box 0 0 1 1
use contact_9  contact_9_69
timestamp 1624857261
transform 1 0 216903 0 1 25667
box 0 0 1 1
use contact_9  contact_9_68
timestamp 1624857261
transform 1 0 216903 0 1 27347
box 0 0 1 1
use contact_9  contact_9_67
timestamp 1624857261
transform 1 0 216903 0 1 29027
box 0 0 1 1
use contact_9  contact_9_66
timestamp 1624857261
transform 1 0 216903 0 1 30707
box 0 0 1 1
use contact_9  contact_9_65
timestamp 1624857261
transform 1 0 216903 0 1 32387
box 0 0 1 1
use contact_9  contact_9_64
timestamp 1624857261
transform 1 0 216903 0 1 34067
box 0 0 1 1
use contact_9  contact_9_63
timestamp 1624857261
transform 1 0 216903 0 1 35747
box 0 0 1 1
use contact_9  contact_9_62
timestamp 1624857261
transform 1 0 216903 0 1 37427
box 0 0 1 1
use contact_9  contact_9_61
timestamp 1624857261
transform 1 0 216903 0 1 39107
box 0 0 1 1
use contact_9  contact_9_60
timestamp 1624857261
transform 1 0 216903 0 1 40787
box 0 0 1 1
use contact_9  contact_9_59
timestamp 1624857261
transform 1 0 216903 0 1 42467
box 0 0 1 1
use contact_9  contact_9_58
timestamp 1624857261
transform 1 0 216903 0 1 44147
box 0 0 1 1
use contact_9  contact_9_57
timestamp 1624857261
transform 1 0 216903 0 1 45827
box 0 0 1 1
use contact_9  contact_9_56
timestamp 1624857261
transform 1 0 216903 0 1 47507
box 0 0 1 1
use contact_9  contact_9_55
timestamp 1624857261
transform 1 0 216903 0 1 49187
box 0 0 1 1
use contact_9  contact_9_54
timestamp 1624857261
transform 1 0 216903 0 1 50867
box 0 0 1 1
use contact_9  contact_9_53
timestamp 1624857261
transform 1 0 216903 0 1 52547
box 0 0 1 1
use contact_9  contact_9_52
timestamp 1624857261
transform 1 0 216903 0 1 54227
box 0 0 1 1
use contact_9  contact_9_51
timestamp 1624857261
transform 1 0 216903 0 1 55907
box 0 0 1 1
use contact_9  contact_9_50
timestamp 1624857261
transform 1 0 216903 0 1 57587
box 0 0 1 1
use contact_9  contact_9_49
timestamp 1624857261
transform 1 0 216903 0 1 59267
box 0 0 1 1
use contact_9  contact_9_48
timestamp 1624857261
transform 1 0 216903 0 1 60947
box 0 0 1 1
use contact_9  contact_9_47
timestamp 1624857261
transform 1 0 216903 0 1 62627
box 0 0 1 1
use contact_9  contact_9_46
timestamp 1624857261
transform 1 0 216903 0 1 64307
box 0 0 1 1
use contact_9  contact_9_45
timestamp 1624857261
transform 1 0 216903 0 1 65987
box 0 0 1 1
use contact_9  contact_9_44
timestamp 1624857261
transform 1 0 216903 0 1 67667
box 0 0 1 1
use contact_9  contact_9_43
timestamp 1624857261
transform 1 0 216903 0 1 69347
box 0 0 1 1
use contact_9  contact_9_42
timestamp 1624857261
transform 1 0 216903 0 1 71027
box 0 0 1 1
use contact_9  contact_9_41
timestamp 1624857261
transform 1 0 216903 0 1 72707
box 0 0 1 1
use contact_9  contact_9_40
timestamp 1624857261
transform 1 0 216903 0 1 74387
box 0 0 1 1
use contact_9  contact_9_39
timestamp 1624857261
transform 1 0 216903 0 1 76067
box 0 0 1 1
use contact_9  contact_9_38
timestamp 1624857261
transform 1 0 216903 0 1 77747
box 0 0 1 1
use contact_9  contact_9_37
timestamp 1624857261
transform 1 0 216903 0 1 79427
box 0 0 1 1
use contact_9  contact_9_36
timestamp 1624857261
transform 1 0 216903 0 1 81107
box 0 0 1 1
use contact_9  contact_9_35
timestamp 1624857261
transform 1 0 216903 0 1 82787
box 0 0 1 1
use contact_9  contact_9_34
timestamp 1624857261
transform 1 0 216903 0 1 84467
box 0 0 1 1
use contact_9  contact_9_33
timestamp 1624857261
transform 1 0 216903 0 1 86147
box 0 0 1 1
use contact_9  contact_9_32
timestamp 1624857261
transform 1 0 216903 0 1 87827
box 0 0 1 1
use contact_9  contact_9_31
timestamp 1624857261
transform 1 0 216903 0 1 89507
box 0 0 1 1
use contact_9  contact_9_30
timestamp 1624857261
transform 1 0 216903 0 1 91187
box 0 0 1 1
use contact_9  contact_9_29
timestamp 1624857261
transform 1 0 216903 0 1 92867
box 0 0 1 1
use contact_9  contact_9_28
timestamp 1624857261
transform 1 0 216903 0 1 94547
box 0 0 1 1
use contact_9  contact_9_27
timestamp 1624857261
transform 1 0 216903 0 1 96227
box 0 0 1 1
use contact_9  contact_9_26
timestamp 1624857261
transform 1 0 216903 0 1 97907
box 0 0 1 1
use contact_9  contact_9_25
timestamp 1624857261
transform 1 0 216903 0 1 99587
box 0 0 1 1
use contact_9  contact_9_24
timestamp 1624857261
transform 1 0 216903 0 1 101267
box 0 0 1 1
use contact_9  contact_9_23
timestamp 1624857261
transform 1 0 216903 0 1 102947
box 0 0 1 1
use contact_9  contact_9_22
timestamp 1624857261
transform 1 0 216903 0 1 104627
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1624857261
transform 1 0 216903 0 1 106307
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1624857261
transform 1 0 216903 0 1 107987
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1624857261
transform 1 0 216903 0 1 109667
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1624857261
transform 1 0 216903 0 1 111347
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1624857261
transform 1 0 216903 0 1 113027
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1624857261
transform 1 0 216903 0 1 114707
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1624857261
transform 1 0 216903 0 1 116387
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1624857261
transform 1 0 216903 0 1 118067
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1624857261
transform 1 0 216903 0 1 119747
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1624857261
transform 1 0 216903 0 1 121427
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1624857261
transform 1 0 216903 0 1 123107
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1624857261
transform 1 0 216903 0 1 124787
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1624857261
transform 1 0 216903 0 1 126467
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1624857261
transform 1 0 216903 0 1 128147
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1624857261
transform 1 0 216903 0 1 129827
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1624857261
transform 1 0 216903 0 1 131507
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1624857261
transform 1 0 216903 0 1 133187
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1624857261
transform 1 0 216903 0 1 134867
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1624857261
transform 1 0 216903 0 1 136547
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1624857261
transform 1 0 216903 0 1 138227
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1624857261
transform 1 0 216903 0 1 139907
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1624857261
transform 1 0 216903 0 1 141587
box 0 0 1 1
use contact_8  contact_8_1169
timestamp 1624857261
transform 1 0 15407 0 1 34920
box 0 0 1 1
use contact_8  contact_8_1168
timestamp 1624857261
transform 1 0 15487 0 1 36478
box 0 0 1 1
use contact_8  contact_8_1167
timestamp 1624857261
transform 1 0 15567 0 1 37748
box 0 0 1 1
use contact_8  contact_8_1166
timestamp 1624857261
transform 1 0 15647 0 1 39306
box 0 0 1 1
use contact_8  contact_8_1165
timestamp 1624857261
transform 1 0 15727 0 1 40576
box 0 0 1 1
use contact_8  contact_8_1164
timestamp 1624857261
transform 1 0 15807 0 1 42134
box 0 0 1 1
use contact_8  contact_8_1163
timestamp 1624857261
transform 1 0 15887 0 1 43404
box 0 0 1 1
use contact_8  contact_8_1162
timestamp 1624857261
transform 1 0 15967 0 1 44962
box 0 0 1 1
use contact_8  contact_8_1161
timestamp 1624857261
transform 1 0 203195 0 1 24170
box 0 0 1 1
use contact_8  contact_8_1160
timestamp 1624857261
transform 1 0 203115 0 1 22612
box 0 0 1 1
use contact_8  contact_8_1159
timestamp 1624857261
transform 1 0 203035 0 1 21342
box 0 0 1 1
use contact_8  contact_8_1158
timestamp 1624857261
transform 1 0 202955 0 1 19784
box 0 0 1 1
use contact_8  contact_8_1157
timestamp 1624857261
transform 1 0 202875 0 1 18514
box 0 0 1 1
use contact_8  contact_8_1156
timestamp 1624857261
transform 1 0 202795 0 1 16956
box 0 0 1 1
use contact_8  contact_8_1155
timestamp 1624857261
transform 1 0 202715 0 1 15686
box 0 0 1 1
use contact_8  contact_8_1154
timestamp 1624857261
transform 1 0 202635 0 1 14128
box 0 0 1 1
use contact_8  contact_8_1153
timestamp 1624857261
transform 1 0 29556 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1152
timestamp 1624857261
transform 1 0 34548 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1151
timestamp 1624857261
transform 1 0 39540 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1150
timestamp 1624857261
transform 1 0 44532 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1149
timestamp 1624857261
transform 1 0 49524 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1148
timestamp 1624857261
transform 1 0 54516 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1147
timestamp 1624857261
transform 1 0 59508 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1146
timestamp 1624857261
transform 1 0 64500 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1145
timestamp 1624857261
transform 1 0 69492 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1144
timestamp 1624857261
transform 1 0 74484 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1143
timestamp 1624857261
transform 1 0 79476 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1142
timestamp 1624857261
transform 1 0 84468 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1141
timestamp 1624857261
transform 1 0 89460 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1140
timestamp 1624857261
transform 1 0 94452 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1139
timestamp 1624857261
transform 1 0 99444 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1138
timestamp 1624857261
transform 1 0 104436 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1137
timestamp 1624857261
transform 1 0 109428 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1136
timestamp 1624857261
transform 1 0 114420 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1135
timestamp 1624857261
transform 1 0 119412 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1134
timestamp 1624857261
transform 1 0 124404 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1133
timestamp 1624857261
transform 1 0 129396 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1132
timestamp 1624857261
transform 1 0 134388 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1131
timestamp 1624857261
transform 1 0 139380 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1130
timestamp 1624857261
transform 1 0 144372 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1129
timestamp 1624857261
transform 1 0 149364 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1128
timestamp 1624857261
transform 1 0 154356 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1127
timestamp 1624857261
transform 1 0 159348 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1126
timestamp 1624857261
transform 1 0 164340 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1125
timestamp 1624857261
transform 1 0 169332 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1124
timestamp 1624857261
transform 1 0 174324 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1123
timestamp 1624857261
transform 1 0 179316 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1122
timestamp 1624857261
transform 1 0 184308 0 1 17696
box 0 0 1 1
use contact_8  contact_8_1121
timestamp 1624857261
transform 1 0 29556 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1120
timestamp 1624857261
transform 1 0 34548 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1119
timestamp 1624857261
transform 1 0 39540 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1118
timestamp 1624857261
transform 1 0 44532 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1117
timestamp 1624857261
transform 1 0 49524 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1116
timestamp 1624857261
transform 1 0 54516 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1115
timestamp 1624857261
transform 1 0 59508 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1114
timestamp 1624857261
transform 1 0 64500 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1113
timestamp 1624857261
transform 1 0 69492 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1112
timestamp 1624857261
transform 1 0 74484 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1111
timestamp 1624857261
transform 1 0 79476 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1110
timestamp 1624857261
transform 1 0 84468 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1109
timestamp 1624857261
transform 1 0 89460 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1108
timestamp 1624857261
transform 1 0 94452 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1107
timestamp 1624857261
transform 1 0 99444 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1106
timestamp 1624857261
transform 1 0 104436 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1105
timestamp 1624857261
transform 1 0 109428 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1104
timestamp 1624857261
transform 1 0 114420 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1103
timestamp 1624857261
transform 1 0 119412 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1102
timestamp 1624857261
transform 1 0 124404 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1101
timestamp 1624857261
transform 1 0 129396 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1100
timestamp 1624857261
transform 1 0 134388 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1099
timestamp 1624857261
transform 1 0 139380 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1098
timestamp 1624857261
transform 1 0 144372 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1097
timestamp 1624857261
transform 1 0 149364 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1096
timestamp 1624857261
transform 1 0 154356 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1095
timestamp 1624857261
transform 1 0 159348 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1094
timestamp 1624857261
transform 1 0 164340 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1093
timestamp 1624857261
transform 1 0 169332 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1092
timestamp 1624857261
transform 1 0 174324 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1091
timestamp 1624857261
transform 1 0 179316 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1090
timestamp 1624857261
transform 1 0 184308 0 1 133034
box 0 0 1 1
use contact_8  contact_8_1089
timestamp 1624857261
transform 1 0 2034 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1088
timestamp 1624857261
transform 1 0 3714 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1087
timestamp 1624857261
transform 1 0 5394 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1086
timestamp 1624857261
transform 1 0 7074 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1085
timestamp 1624857261
transform 1 0 8754 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1084
timestamp 1624857261
transform 1 0 10434 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1083
timestamp 1624857261
transform 1 0 12114 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1082
timestamp 1624857261
transform 1 0 13794 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1081
timestamp 1624857261
transform 1 0 15474 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1080
timestamp 1624857261
transform 1 0 17154 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1079
timestamp 1624857261
transform 1 0 18834 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1078
timestamp 1624857261
transform 1 0 20514 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1077
timestamp 1624857261
transform 1 0 22194 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1076
timestamp 1624857261
transform 1 0 23874 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1075
timestamp 1624857261
transform 1 0 25554 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1074
timestamp 1624857261
transform 1 0 27234 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1073
timestamp 1624857261
transform 1 0 28914 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1072
timestamp 1624857261
transform 1 0 30594 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1071
timestamp 1624857261
transform 1 0 32274 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1070
timestamp 1624857261
transform 1 0 33954 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1069
timestamp 1624857261
transform 1 0 35634 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1068
timestamp 1624857261
transform 1 0 37314 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1067
timestamp 1624857261
transform 1 0 38994 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1066
timestamp 1624857261
transform 1 0 40674 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1065
timestamp 1624857261
transform 1 0 42354 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1064
timestamp 1624857261
transform 1 0 44034 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1063
timestamp 1624857261
transform 1 0 45714 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1062
timestamp 1624857261
transform 1 0 47394 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1061
timestamp 1624857261
transform 1 0 49074 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1060
timestamp 1624857261
transform 1 0 50754 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1059
timestamp 1624857261
transform 1 0 52434 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1058
timestamp 1624857261
transform 1 0 54114 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1057
timestamp 1624857261
transform 1 0 55794 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1056
timestamp 1624857261
transform 1 0 57474 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1055
timestamp 1624857261
transform 1 0 59154 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1054
timestamp 1624857261
transform 1 0 60834 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1053
timestamp 1624857261
transform 1 0 62514 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1052
timestamp 1624857261
transform 1 0 64194 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1051
timestamp 1624857261
transform 1 0 65874 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1050
timestamp 1624857261
transform 1 0 67554 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1049
timestamp 1624857261
transform 1 0 69234 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1048
timestamp 1624857261
transform 1 0 70914 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1047
timestamp 1624857261
transform 1 0 72594 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1046
timestamp 1624857261
transform 1 0 74274 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1045
timestamp 1624857261
transform 1 0 75954 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1044
timestamp 1624857261
transform 1 0 77634 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1043
timestamp 1624857261
transform 1 0 79314 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1042
timestamp 1624857261
transform 1 0 80994 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1041
timestamp 1624857261
transform 1 0 82674 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1040
timestamp 1624857261
transform 1 0 84354 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1039
timestamp 1624857261
transform 1 0 86034 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1038
timestamp 1624857261
transform 1 0 87714 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1037
timestamp 1624857261
transform 1 0 89394 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1036
timestamp 1624857261
transform 1 0 91074 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1035
timestamp 1624857261
transform 1 0 92754 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1034
timestamp 1624857261
transform 1 0 94434 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1033
timestamp 1624857261
transform 1 0 96114 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1032
timestamp 1624857261
transform 1 0 97794 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1031
timestamp 1624857261
transform 1 0 99474 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1030
timestamp 1624857261
transform 1 0 101154 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1029
timestamp 1624857261
transform 1 0 102834 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1028
timestamp 1624857261
transform 1 0 104514 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1027
timestamp 1624857261
transform 1 0 106194 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1026
timestamp 1624857261
transform 1 0 107874 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1025
timestamp 1624857261
transform 1 0 109554 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1024
timestamp 1624857261
transform 1 0 111234 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1023
timestamp 1624857261
transform 1 0 112914 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1022
timestamp 1624857261
transform 1 0 114594 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1021
timestamp 1624857261
transform 1 0 116274 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1020
timestamp 1624857261
transform 1 0 117954 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1019
timestamp 1624857261
transform 1 0 119634 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1018
timestamp 1624857261
transform 1 0 121314 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1017
timestamp 1624857261
transform 1 0 122994 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1016
timestamp 1624857261
transform 1 0 124674 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1015
timestamp 1624857261
transform 1 0 126354 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1014
timestamp 1624857261
transform 1 0 128034 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1013
timestamp 1624857261
transform 1 0 129714 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1012
timestamp 1624857261
transform 1 0 131394 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1011
timestamp 1624857261
transform 1 0 133074 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1010
timestamp 1624857261
transform 1 0 134754 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1009
timestamp 1624857261
transform 1 0 136434 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1008
timestamp 1624857261
transform 1 0 138114 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1007
timestamp 1624857261
transform 1 0 139794 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1006
timestamp 1624857261
transform 1 0 141474 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1005
timestamp 1624857261
transform 1 0 143154 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1004
timestamp 1624857261
transform 1 0 144834 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1003
timestamp 1624857261
transform 1 0 146514 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1002
timestamp 1624857261
transform 1 0 148194 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1001
timestamp 1624857261
transform 1 0 149874 0 1 1816
box 0 0 1 1
use contact_8  contact_8_1000
timestamp 1624857261
transform 1 0 151554 0 1 1816
box 0 0 1 1
use contact_8  contact_8_999
timestamp 1624857261
transform 1 0 153234 0 1 1816
box 0 0 1 1
use contact_8  contact_8_998
timestamp 1624857261
transform 1 0 154914 0 1 1816
box 0 0 1 1
use contact_8  contact_8_997
timestamp 1624857261
transform 1 0 156594 0 1 1816
box 0 0 1 1
use contact_8  contact_8_996
timestamp 1624857261
transform 1 0 158274 0 1 1816
box 0 0 1 1
use contact_8  contact_8_995
timestamp 1624857261
transform 1 0 159954 0 1 1816
box 0 0 1 1
use contact_8  contact_8_994
timestamp 1624857261
transform 1 0 161634 0 1 1816
box 0 0 1 1
use contact_8  contact_8_993
timestamp 1624857261
transform 1 0 163314 0 1 1816
box 0 0 1 1
use contact_8  contact_8_992
timestamp 1624857261
transform 1 0 164994 0 1 1816
box 0 0 1 1
use contact_8  contact_8_991
timestamp 1624857261
transform 1 0 166674 0 1 1816
box 0 0 1 1
use contact_8  contact_8_990
timestamp 1624857261
transform 1 0 168354 0 1 1816
box 0 0 1 1
use contact_8  contact_8_989
timestamp 1624857261
transform 1 0 170034 0 1 1816
box 0 0 1 1
use contact_8  contact_8_988
timestamp 1624857261
transform 1 0 171714 0 1 1816
box 0 0 1 1
use contact_8  contact_8_987
timestamp 1624857261
transform 1 0 173394 0 1 1816
box 0 0 1 1
use contact_8  contact_8_986
timestamp 1624857261
transform 1 0 175074 0 1 1816
box 0 0 1 1
use contact_8  contact_8_985
timestamp 1624857261
transform 1 0 176754 0 1 1816
box 0 0 1 1
use contact_8  contact_8_984
timestamp 1624857261
transform 1 0 178434 0 1 1816
box 0 0 1 1
use contact_8  contact_8_983
timestamp 1624857261
transform 1 0 180114 0 1 1816
box 0 0 1 1
use contact_8  contact_8_982
timestamp 1624857261
transform 1 0 181794 0 1 1816
box 0 0 1 1
use contact_8  contact_8_981
timestamp 1624857261
transform 1 0 183474 0 1 1816
box 0 0 1 1
use contact_8  contact_8_980
timestamp 1624857261
transform 1 0 185154 0 1 1816
box 0 0 1 1
use contact_8  contact_8_979
timestamp 1624857261
transform 1 0 186834 0 1 1816
box 0 0 1 1
use contact_8  contact_8_978
timestamp 1624857261
transform 1 0 188514 0 1 1816
box 0 0 1 1
use contact_8  contact_8_977
timestamp 1624857261
transform 1 0 190194 0 1 1816
box 0 0 1 1
use contact_8  contact_8_976
timestamp 1624857261
transform 1 0 191874 0 1 1816
box 0 0 1 1
use contact_8  contact_8_975
timestamp 1624857261
transform 1 0 193554 0 1 1816
box 0 0 1 1
use contact_8  contact_8_974
timestamp 1624857261
transform 1 0 195234 0 1 1816
box 0 0 1 1
use contact_8  contact_8_973
timestamp 1624857261
transform 1 0 196914 0 1 1816
box 0 0 1 1
use contact_8  contact_8_972
timestamp 1624857261
transform 1 0 198594 0 1 1816
box 0 0 1 1
use contact_8  contact_8_971
timestamp 1624857261
transform 1 0 200274 0 1 1816
box 0 0 1 1
use contact_8  contact_8_970
timestamp 1624857261
transform 1 0 201954 0 1 1816
box 0 0 1 1
use contact_8  contact_8_969
timestamp 1624857261
transform 1 0 203634 0 1 1816
box 0 0 1 1
use contact_8  contact_8_968
timestamp 1624857261
transform 1 0 205314 0 1 1816
box 0 0 1 1
use contact_8  contact_8_967
timestamp 1624857261
transform 1 0 206994 0 1 1816
box 0 0 1 1
use contact_8  contact_8_966
timestamp 1624857261
transform 1 0 208674 0 1 1816
box 0 0 1 1
use contact_8  contact_8_965
timestamp 1624857261
transform 1 0 210354 0 1 1816
box 0 0 1 1
use contact_8  contact_8_964
timestamp 1624857261
transform 1 0 212034 0 1 1816
box 0 0 1 1
use contact_8  contact_8_963
timestamp 1624857261
transform 1 0 213714 0 1 1816
box 0 0 1 1
use contact_8  contact_8_962
timestamp 1624857261
transform 1 0 215394 0 1 1816
box 0 0 1 1
use contact_8  contact_8_961
timestamp 1624857261
transform 1 0 2034 0 1 142312
box 0 0 1 1
use contact_8  contact_8_960
timestamp 1624857261
transform 1 0 3714 0 1 142312
box 0 0 1 1
use contact_8  contact_8_959
timestamp 1624857261
transform 1 0 5394 0 1 142312
box 0 0 1 1
use contact_8  contact_8_958
timestamp 1624857261
transform 1 0 7074 0 1 142312
box 0 0 1 1
use contact_8  contact_8_957
timestamp 1624857261
transform 1 0 8754 0 1 142312
box 0 0 1 1
use contact_8  contact_8_956
timestamp 1624857261
transform 1 0 10434 0 1 142312
box 0 0 1 1
use contact_8  contact_8_955
timestamp 1624857261
transform 1 0 12114 0 1 142312
box 0 0 1 1
use contact_8  contact_8_954
timestamp 1624857261
transform 1 0 13794 0 1 142312
box 0 0 1 1
use contact_8  contact_8_953
timestamp 1624857261
transform 1 0 15474 0 1 142312
box 0 0 1 1
use contact_8  contact_8_952
timestamp 1624857261
transform 1 0 17154 0 1 142312
box 0 0 1 1
use contact_8  contact_8_951
timestamp 1624857261
transform 1 0 18834 0 1 142312
box 0 0 1 1
use contact_8  contact_8_950
timestamp 1624857261
transform 1 0 20514 0 1 142312
box 0 0 1 1
use contact_8  contact_8_949
timestamp 1624857261
transform 1 0 22194 0 1 142312
box 0 0 1 1
use contact_8  contact_8_948
timestamp 1624857261
transform 1 0 23874 0 1 142312
box 0 0 1 1
use contact_8  contact_8_947
timestamp 1624857261
transform 1 0 25554 0 1 142312
box 0 0 1 1
use contact_8  contact_8_946
timestamp 1624857261
transform 1 0 27234 0 1 142312
box 0 0 1 1
use contact_8  contact_8_945
timestamp 1624857261
transform 1 0 28914 0 1 142312
box 0 0 1 1
use contact_8  contact_8_944
timestamp 1624857261
transform 1 0 30594 0 1 142312
box 0 0 1 1
use contact_8  contact_8_943
timestamp 1624857261
transform 1 0 32274 0 1 142312
box 0 0 1 1
use contact_8  contact_8_942
timestamp 1624857261
transform 1 0 33954 0 1 142312
box 0 0 1 1
use contact_8  contact_8_941
timestamp 1624857261
transform 1 0 35634 0 1 142312
box 0 0 1 1
use contact_8  contact_8_940
timestamp 1624857261
transform 1 0 37314 0 1 142312
box 0 0 1 1
use contact_8  contact_8_939
timestamp 1624857261
transform 1 0 38994 0 1 142312
box 0 0 1 1
use contact_8  contact_8_938
timestamp 1624857261
transform 1 0 40674 0 1 142312
box 0 0 1 1
use contact_8  contact_8_937
timestamp 1624857261
transform 1 0 42354 0 1 142312
box 0 0 1 1
use contact_8  contact_8_936
timestamp 1624857261
transform 1 0 44034 0 1 142312
box 0 0 1 1
use contact_8  contact_8_935
timestamp 1624857261
transform 1 0 45714 0 1 142312
box 0 0 1 1
use contact_8  contact_8_934
timestamp 1624857261
transform 1 0 47394 0 1 142312
box 0 0 1 1
use contact_8  contact_8_933
timestamp 1624857261
transform 1 0 49074 0 1 142312
box 0 0 1 1
use contact_8  contact_8_932
timestamp 1624857261
transform 1 0 50754 0 1 142312
box 0 0 1 1
use contact_8  contact_8_931
timestamp 1624857261
transform 1 0 52434 0 1 142312
box 0 0 1 1
use contact_8  contact_8_930
timestamp 1624857261
transform 1 0 54114 0 1 142312
box 0 0 1 1
use contact_8  contact_8_929
timestamp 1624857261
transform 1 0 55794 0 1 142312
box 0 0 1 1
use contact_8  contact_8_928
timestamp 1624857261
transform 1 0 57474 0 1 142312
box 0 0 1 1
use contact_8  contact_8_927
timestamp 1624857261
transform 1 0 59154 0 1 142312
box 0 0 1 1
use contact_8  contact_8_926
timestamp 1624857261
transform 1 0 60834 0 1 142312
box 0 0 1 1
use contact_8  contact_8_925
timestamp 1624857261
transform 1 0 62514 0 1 142312
box 0 0 1 1
use contact_8  contact_8_924
timestamp 1624857261
transform 1 0 64194 0 1 142312
box 0 0 1 1
use contact_8  contact_8_923
timestamp 1624857261
transform 1 0 65874 0 1 142312
box 0 0 1 1
use contact_8  contact_8_922
timestamp 1624857261
transform 1 0 67554 0 1 142312
box 0 0 1 1
use contact_8  contact_8_921
timestamp 1624857261
transform 1 0 69234 0 1 142312
box 0 0 1 1
use contact_8  contact_8_920
timestamp 1624857261
transform 1 0 70914 0 1 142312
box 0 0 1 1
use contact_8  contact_8_919
timestamp 1624857261
transform 1 0 72594 0 1 142312
box 0 0 1 1
use contact_8  contact_8_918
timestamp 1624857261
transform 1 0 74274 0 1 142312
box 0 0 1 1
use contact_8  contact_8_917
timestamp 1624857261
transform 1 0 75954 0 1 142312
box 0 0 1 1
use contact_8  contact_8_916
timestamp 1624857261
transform 1 0 77634 0 1 142312
box 0 0 1 1
use contact_8  contact_8_915
timestamp 1624857261
transform 1 0 79314 0 1 142312
box 0 0 1 1
use contact_8  contact_8_914
timestamp 1624857261
transform 1 0 80994 0 1 142312
box 0 0 1 1
use contact_8  contact_8_913
timestamp 1624857261
transform 1 0 82674 0 1 142312
box 0 0 1 1
use contact_8  contact_8_912
timestamp 1624857261
transform 1 0 84354 0 1 142312
box 0 0 1 1
use contact_8  contact_8_911
timestamp 1624857261
transform 1 0 86034 0 1 142312
box 0 0 1 1
use contact_8  contact_8_910
timestamp 1624857261
transform 1 0 87714 0 1 142312
box 0 0 1 1
use contact_8  contact_8_909
timestamp 1624857261
transform 1 0 89394 0 1 142312
box 0 0 1 1
use contact_8  contact_8_908
timestamp 1624857261
transform 1 0 91074 0 1 142312
box 0 0 1 1
use contact_8  contact_8_907
timestamp 1624857261
transform 1 0 92754 0 1 142312
box 0 0 1 1
use contact_8  contact_8_906
timestamp 1624857261
transform 1 0 94434 0 1 142312
box 0 0 1 1
use contact_8  contact_8_905
timestamp 1624857261
transform 1 0 96114 0 1 142312
box 0 0 1 1
use contact_8  contact_8_904
timestamp 1624857261
transform 1 0 97794 0 1 142312
box 0 0 1 1
use contact_8  contact_8_903
timestamp 1624857261
transform 1 0 99474 0 1 142312
box 0 0 1 1
use contact_8  contact_8_902
timestamp 1624857261
transform 1 0 101154 0 1 142312
box 0 0 1 1
use contact_8  contact_8_901
timestamp 1624857261
transform 1 0 102834 0 1 142312
box 0 0 1 1
use contact_8  contact_8_900
timestamp 1624857261
transform 1 0 104514 0 1 142312
box 0 0 1 1
use contact_8  contact_8_899
timestamp 1624857261
transform 1 0 106194 0 1 142312
box 0 0 1 1
use contact_8  contact_8_898
timestamp 1624857261
transform 1 0 107874 0 1 142312
box 0 0 1 1
use contact_8  contact_8_897
timestamp 1624857261
transform 1 0 109554 0 1 142312
box 0 0 1 1
use contact_8  contact_8_896
timestamp 1624857261
transform 1 0 111234 0 1 142312
box 0 0 1 1
use contact_8  contact_8_895
timestamp 1624857261
transform 1 0 112914 0 1 142312
box 0 0 1 1
use contact_8  contact_8_894
timestamp 1624857261
transform 1 0 114594 0 1 142312
box 0 0 1 1
use contact_8  contact_8_893
timestamp 1624857261
transform 1 0 116274 0 1 142312
box 0 0 1 1
use contact_8  contact_8_892
timestamp 1624857261
transform 1 0 117954 0 1 142312
box 0 0 1 1
use contact_8  contact_8_891
timestamp 1624857261
transform 1 0 119634 0 1 142312
box 0 0 1 1
use contact_8  contact_8_890
timestamp 1624857261
transform 1 0 121314 0 1 142312
box 0 0 1 1
use contact_8  contact_8_889
timestamp 1624857261
transform 1 0 122994 0 1 142312
box 0 0 1 1
use contact_8  contact_8_888
timestamp 1624857261
transform 1 0 124674 0 1 142312
box 0 0 1 1
use contact_8  contact_8_887
timestamp 1624857261
transform 1 0 126354 0 1 142312
box 0 0 1 1
use contact_8  contact_8_886
timestamp 1624857261
transform 1 0 128034 0 1 142312
box 0 0 1 1
use contact_8  contact_8_885
timestamp 1624857261
transform 1 0 129714 0 1 142312
box 0 0 1 1
use contact_8  contact_8_884
timestamp 1624857261
transform 1 0 131394 0 1 142312
box 0 0 1 1
use contact_8  contact_8_883
timestamp 1624857261
transform 1 0 133074 0 1 142312
box 0 0 1 1
use contact_8  contact_8_882
timestamp 1624857261
transform 1 0 134754 0 1 142312
box 0 0 1 1
use contact_8  contact_8_881
timestamp 1624857261
transform 1 0 136434 0 1 142312
box 0 0 1 1
use contact_8  contact_8_880
timestamp 1624857261
transform 1 0 138114 0 1 142312
box 0 0 1 1
use contact_8  contact_8_879
timestamp 1624857261
transform 1 0 139794 0 1 142312
box 0 0 1 1
use contact_8  contact_8_878
timestamp 1624857261
transform 1 0 141474 0 1 142312
box 0 0 1 1
use contact_8  contact_8_877
timestamp 1624857261
transform 1 0 143154 0 1 142312
box 0 0 1 1
use contact_8  contact_8_876
timestamp 1624857261
transform 1 0 144834 0 1 142312
box 0 0 1 1
use contact_8  contact_8_875
timestamp 1624857261
transform 1 0 146514 0 1 142312
box 0 0 1 1
use contact_8  contact_8_874
timestamp 1624857261
transform 1 0 148194 0 1 142312
box 0 0 1 1
use contact_8  contact_8_873
timestamp 1624857261
transform 1 0 149874 0 1 142312
box 0 0 1 1
use contact_8  contact_8_872
timestamp 1624857261
transform 1 0 151554 0 1 142312
box 0 0 1 1
use contact_8  contact_8_871
timestamp 1624857261
transform 1 0 153234 0 1 142312
box 0 0 1 1
use contact_8  contact_8_870
timestamp 1624857261
transform 1 0 154914 0 1 142312
box 0 0 1 1
use contact_8  contact_8_869
timestamp 1624857261
transform 1 0 156594 0 1 142312
box 0 0 1 1
use contact_8  contact_8_868
timestamp 1624857261
transform 1 0 158274 0 1 142312
box 0 0 1 1
use contact_8  contact_8_867
timestamp 1624857261
transform 1 0 159954 0 1 142312
box 0 0 1 1
use contact_8  contact_8_866
timestamp 1624857261
transform 1 0 161634 0 1 142312
box 0 0 1 1
use contact_8  contact_8_865
timestamp 1624857261
transform 1 0 163314 0 1 142312
box 0 0 1 1
use contact_8  contact_8_864
timestamp 1624857261
transform 1 0 164994 0 1 142312
box 0 0 1 1
use contact_8  contact_8_863
timestamp 1624857261
transform 1 0 166674 0 1 142312
box 0 0 1 1
use contact_8  contact_8_862
timestamp 1624857261
transform 1 0 168354 0 1 142312
box 0 0 1 1
use contact_8  contact_8_861
timestamp 1624857261
transform 1 0 170034 0 1 142312
box 0 0 1 1
use contact_8  contact_8_860
timestamp 1624857261
transform 1 0 171714 0 1 142312
box 0 0 1 1
use contact_8  contact_8_859
timestamp 1624857261
transform 1 0 173394 0 1 142312
box 0 0 1 1
use contact_8  contact_8_858
timestamp 1624857261
transform 1 0 175074 0 1 142312
box 0 0 1 1
use contact_8  contact_8_857
timestamp 1624857261
transform 1 0 176754 0 1 142312
box 0 0 1 1
use contact_8  contact_8_856
timestamp 1624857261
transform 1 0 178434 0 1 142312
box 0 0 1 1
use contact_8  contact_8_855
timestamp 1624857261
transform 1 0 180114 0 1 142312
box 0 0 1 1
use contact_8  contact_8_854
timestamp 1624857261
transform 1 0 181794 0 1 142312
box 0 0 1 1
use contact_8  contact_8_853
timestamp 1624857261
transform 1 0 183474 0 1 142312
box 0 0 1 1
use contact_8  contact_8_852
timestamp 1624857261
transform 1 0 185154 0 1 142312
box 0 0 1 1
use contact_8  contact_8_851
timestamp 1624857261
transform 1 0 186834 0 1 142312
box 0 0 1 1
use contact_8  contact_8_850
timestamp 1624857261
transform 1 0 188514 0 1 142312
box 0 0 1 1
use contact_8  contact_8_849
timestamp 1624857261
transform 1 0 190194 0 1 142312
box 0 0 1 1
use contact_8  contact_8_848
timestamp 1624857261
transform 1 0 191874 0 1 142312
box 0 0 1 1
use contact_8  contact_8_847
timestamp 1624857261
transform 1 0 193554 0 1 142312
box 0 0 1 1
use contact_8  contact_8_846
timestamp 1624857261
transform 1 0 195234 0 1 142312
box 0 0 1 1
use contact_8  contact_8_845
timestamp 1624857261
transform 1 0 196914 0 1 142312
box 0 0 1 1
use contact_8  contact_8_844
timestamp 1624857261
transform 1 0 198594 0 1 142312
box 0 0 1 1
use contact_8  contact_8_843
timestamp 1624857261
transform 1 0 200274 0 1 142312
box 0 0 1 1
use contact_8  contact_8_842
timestamp 1624857261
transform 1 0 201954 0 1 142312
box 0 0 1 1
use contact_8  contact_8_841
timestamp 1624857261
transform 1 0 203634 0 1 142312
box 0 0 1 1
use contact_8  contact_8_840
timestamp 1624857261
transform 1 0 205314 0 1 142312
box 0 0 1 1
use contact_8  contact_8_839
timestamp 1624857261
transform 1 0 206994 0 1 142312
box 0 0 1 1
use contact_8  contact_8_838
timestamp 1624857261
transform 1 0 208674 0 1 142312
box 0 0 1 1
use contact_8  contact_8_837
timestamp 1624857261
transform 1 0 210354 0 1 142312
box 0 0 1 1
use contact_8  contact_8_836
timestamp 1624857261
transform 1 0 212034 0 1 142312
box 0 0 1 1
use contact_8  contact_8_835
timestamp 1624857261
transform 1 0 213714 0 1 142312
box 0 0 1 1
use contact_8  contact_8_834
timestamp 1624857261
transform 1 0 215394 0 1 142312
box 0 0 1 1
use contact_8  contact_8_833
timestamp 1624857261
transform 1 0 1698 0 1 2152
box 0 0 1 1
use contact_8  contact_8_832
timestamp 1624857261
transform 1 0 1698 0 1 2488
box 0 0 1 1
use contact_8  contact_8_831
timestamp 1624857261
transform 1 0 1698 0 1 2824
box 0 0 1 1
use contact_8  contact_8_830
timestamp 1624857261
transform 1 0 1698 0 1 3160
box 0 0 1 1
use contact_8  contact_8_829
timestamp 1624857261
transform 1 0 1698 0 1 3496
box 0 0 1 1
use contact_8  contact_8_828
timestamp 1624857261
transform 1 0 1698 0 1 3832
box 0 0 1 1
use contact_8  contact_8_827
timestamp 1624857261
transform 1 0 1698 0 1 4168
box 0 0 1 1
use contact_8  contact_8_826
timestamp 1624857261
transform 1 0 1698 0 1 4504
box 0 0 1 1
use contact_8  contact_8_825
timestamp 1624857261
transform 1 0 1698 0 1 4840
box 0 0 1 1
use contact_8  contact_8_824
timestamp 1624857261
transform 1 0 1698 0 1 5176
box 0 0 1 1
use contact_8  contact_8_823
timestamp 1624857261
transform 1 0 1698 0 1 5512
box 0 0 1 1
use contact_8  contact_8_822
timestamp 1624857261
transform 1 0 1698 0 1 5848
box 0 0 1 1
use contact_8  contact_8_821
timestamp 1624857261
transform 1 0 1698 0 1 6184
box 0 0 1 1
use contact_8  contact_8_820
timestamp 1624857261
transform 1 0 1698 0 1 6520
box 0 0 1 1
use contact_8  contact_8_819
timestamp 1624857261
transform 1 0 1698 0 1 6856
box 0 0 1 1
use contact_8  contact_8_818
timestamp 1624857261
transform 1 0 1698 0 1 7192
box 0 0 1 1
use contact_8  contact_8_817
timestamp 1624857261
transform 1 0 1698 0 1 7528
box 0 0 1 1
use contact_8  contact_8_816
timestamp 1624857261
transform 1 0 1698 0 1 7864
box 0 0 1 1
use contact_8  contact_8_815
timestamp 1624857261
transform 1 0 1698 0 1 8200
box 0 0 1 1
use contact_8  contact_8_814
timestamp 1624857261
transform 1 0 1698 0 1 8536
box 0 0 1 1
use contact_8  contact_8_813
timestamp 1624857261
transform 1 0 1698 0 1 8872
box 0 0 1 1
use contact_8  contact_8_812
timestamp 1624857261
transform 1 0 1698 0 1 9208
box 0 0 1 1
use contact_8  contact_8_811
timestamp 1624857261
transform 1 0 1698 0 1 9544
box 0 0 1 1
use contact_8  contact_8_810
timestamp 1624857261
transform 1 0 1698 0 1 9880
box 0 0 1 1
use contact_8  contact_8_809
timestamp 1624857261
transform 1 0 1698 0 1 10216
box 0 0 1 1
use contact_8  contact_8_808
timestamp 1624857261
transform 1 0 1698 0 1 10552
box 0 0 1 1
use contact_8  contact_8_807
timestamp 1624857261
transform 1 0 1698 0 1 10888
box 0 0 1 1
use contact_8  contact_8_806
timestamp 1624857261
transform 1 0 1698 0 1 11224
box 0 0 1 1
use contact_8  contact_8_805
timestamp 1624857261
transform 1 0 1698 0 1 11560
box 0 0 1 1
use contact_8  contact_8_804
timestamp 1624857261
transform 1 0 1698 0 1 11896
box 0 0 1 1
use contact_8  contact_8_803
timestamp 1624857261
transform 1 0 1698 0 1 12232
box 0 0 1 1
use contact_8  contact_8_802
timestamp 1624857261
transform 1 0 1698 0 1 12568
box 0 0 1 1
use contact_8  contact_8_801
timestamp 1624857261
transform 1 0 1698 0 1 12904
box 0 0 1 1
use contact_8  contact_8_800
timestamp 1624857261
transform 1 0 1698 0 1 13240
box 0 0 1 1
use contact_8  contact_8_799
timestamp 1624857261
transform 1 0 1698 0 1 13576
box 0 0 1 1
use contact_8  contact_8_798
timestamp 1624857261
transform 1 0 1698 0 1 13912
box 0 0 1 1
use contact_8  contact_8_797
timestamp 1624857261
transform 1 0 1698 0 1 14248
box 0 0 1 1
use contact_8  contact_8_796
timestamp 1624857261
transform 1 0 1698 0 1 14584
box 0 0 1 1
use contact_8  contact_8_795
timestamp 1624857261
transform 1 0 1698 0 1 14920
box 0 0 1 1
use contact_8  contact_8_794
timestamp 1624857261
transform 1 0 1698 0 1 15256
box 0 0 1 1
use contact_8  contact_8_793
timestamp 1624857261
transform 1 0 1698 0 1 15592
box 0 0 1 1
use contact_8  contact_8_792
timestamp 1624857261
transform 1 0 1698 0 1 15928
box 0 0 1 1
use contact_8  contact_8_791
timestamp 1624857261
transform 1 0 1698 0 1 16264
box 0 0 1 1
use contact_8  contact_8_790
timestamp 1624857261
transform 1 0 1698 0 1 16600
box 0 0 1 1
use contact_8  contact_8_789
timestamp 1624857261
transform 1 0 1698 0 1 16936
box 0 0 1 1
use contact_8  contact_8_788
timestamp 1624857261
transform 1 0 1698 0 1 17272
box 0 0 1 1
use contact_8  contact_8_787
timestamp 1624857261
transform 1 0 1698 0 1 17608
box 0 0 1 1
use contact_8  contact_8_786
timestamp 1624857261
transform 1 0 1698 0 1 17944
box 0 0 1 1
use contact_8  contact_8_785
timestamp 1624857261
transform 1 0 1698 0 1 18280
box 0 0 1 1
use contact_8  contact_8_784
timestamp 1624857261
transform 1 0 1698 0 1 18616
box 0 0 1 1
use contact_8  contact_8_783
timestamp 1624857261
transform 1 0 1698 0 1 18952
box 0 0 1 1
use contact_8  contact_8_782
timestamp 1624857261
transform 1 0 1698 0 1 19288
box 0 0 1 1
use contact_8  contact_8_781
timestamp 1624857261
transform 1 0 1698 0 1 19624
box 0 0 1 1
use contact_8  contact_8_780
timestamp 1624857261
transform 1 0 1698 0 1 19960
box 0 0 1 1
use contact_8  contact_8_779
timestamp 1624857261
transform 1 0 1698 0 1 20296
box 0 0 1 1
use contact_8  contact_8_778
timestamp 1624857261
transform 1 0 1698 0 1 20632
box 0 0 1 1
use contact_8  contact_8_777
timestamp 1624857261
transform 1 0 1698 0 1 20968
box 0 0 1 1
use contact_8  contact_8_776
timestamp 1624857261
transform 1 0 1698 0 1 21304
box 0 0 1 1
use contact_8  contact_8_775
timestamp 1624857261
transform 1 0 1698 0 1 21640
box 0 0 1 1
use contact_8  contact_8_774
timestamp 1624857261
transform 1 0 1698 0 1 21976
box 0 0 1 1
use contact_8  contact_8_773
timestamp 1624857261
transform 1 0 1698 0 1 22312
box 0 0 1 1
use contact_8  contact_8_772
timestamp 1624857261
transform 1 0 1698 0 1 22648
box 0 0 1 1
use contact_8  contact_8_771
timestamp 1624857261
transform 1 0 1698 0 1 22984
box 0 0 1 1
use contact_8  contact_8_770
timestamp 1624857261
transform 1 0 1698 0 1 23320
box 0 0 1 1
use contact_8  contact_8_769
timestamp 1624857261
transform 1 0 1698 0 1 23656
box 0 0 1 1
use contact_8  contact_8_768
timestamp 1624857261
transform 1 0 1698 0 1 23992
box 0 0 1 1
use contact_8  contact_8_767
timestamp 1624857261
transform 1 0 1698 0 1 24328
box 0 0 1 1
use contact_8  contact_8_766
timestamp 1624857261
transform 1 0 1698 0 1 24664
box 0 0 1 1
use contact_8  contact_8_765
timestamp 1624857261
transform 1 0 1698 0 1 25000
box 0 0 1 1
use contact_8  contact_8_764
timestamp 1624857261
transform 1 0 1698 0 1 25336
box 0 0 1 1
use contact_8  contact_8_763
timestamp 1624857261
transform 1 0 1698 0 1 25672
box 0 0 1 1
use contact_8  contact_8_762
timestamp 1624857261
transform 1 0 1698 0 1 26008
box 0 0 1 1
use contact_8  contact_8_761
timestamp 1624857261
transform 1 0 1698 0 1 26344
box 0 0 1 1
use contact_8  contact_8_760
timestamp 1624857261
transform 1 0 1698 0 1 26680
box 0 0 1 1
use contact_8  contact_8_759
timestamp 1624857261
transform 1 0 1698 0 1 27016
box 0 0 1 1
use contact_8  contact_8_758
timestamp 1624857261
transform 1 0 1698 0 1 27352
box 0 0 1 1
use contact_8  contact_8_757
timestamp 1624857261
transform 1 0 1698 0 1 27688
box 0 0 1 1
use contact_8  contact_8_756
timestamp 1624857261
transform 1 0 1698 0 1 28024
box 0 0 1 1
use contact_8  contact_8_755
timestamp 1624857261
transform 1 0 1698 0 1 28360
box 0 0 1 1
use contact_8  contact_8_754
timestamp 1624857261
transform 1 0 1698 0 1 28696
box 0 0 1 1
use contact_8  contact_8_753
timestamp 1624857261
transform 1 0 1698 0 1 29032
box 0 0 1 1
use contact_8  contact_8_752
timestamp 1624857261
transform 1 0 1698 0 1 29368
box 0 0 1 1
use contact_8  contact_8_751
timestamp 1624857261
transform 1 0 1698 0 1 29704
box 0 0 1 1
use contact_8  contact_8_750
timestamp 1624857261
transform 1 0 1698 0 1 30040
box 0 0 1 1
use contact_8  contact_8_749
timestamp 1624857261
transform 1 0 1698 0 1 30376
box 0 0 1 1
use contact_8  contact_8_748
timestamp 1624857261
transform 1 0 1698 0 1 30712
box 0 0 1 1
use contact_8  contact_8_747
timestamp 1624857261
transform 1 0 1698 0 1 31048
box 0 0 1 1
use contact_8  contact_8_746
timestamp 1624857261
transform 1 0 1698 0 1 31384
box 0 0 1 1
use contact_8  contact_8_745
timestamp 1624857261
transform 1 0 1698 0 1 31720
box 0 0 1 1
use contact_8  contact_8_744
timestamp 1624857261
transform 1 0 1698 0 1 32056
box 0 0 1 1
use contact_8  contact_8_743
timestamp 1624857261
transform 1 0 1698 0 1 32392
box 0 0 1 1
use contact_8  contact_8_742
timestamp 1624857261
transform 1 0 1698 0 1 32728
box 0 0 1 1
use contact_8  contact_8_741
timestamp 1624857261
transform 1 0 1698 0 1 33064
box 0 0 1 1
use contact_8  contact_8_740
timestamp 1624857261
transform 1 0 1698 0 1 33400
box 0 0 1 1
use contact_8  contact_8_739
timestamp 1624857261
transform 1 0 1698 0 1 33736
box 0 0 1 1
use contact_8  contact_8_738
timestamp 1624857261
transform 1 0 1698 0 1 34072
box 0 0 1 1
use contact_8  contact_8_737
timestamp 1624857261
transform 1 0 1698 0 1 34408
box 0 0 1 1
use contact_8  contact_8_736
timestamp 1624857261
transform 1 0 1698 0 1 34744
box 0 0 1 1
use contact_8  contact_8_735
timestamp 1624857261
transform 1 0 1698 0 1 35080
box 0 0 1 1
use contact_8  contact_8_734
timestamp 1624857261
transform 1 0 1698 0 1 35416
box 0 0 1 1
use contact_8  contact_8_733
timestamp 1624857261
transform 1 0 1698 0 1 35752
box 0 0 1 1
use contact_8  contact_8_732
timestamp 1624857261
transform 1 0 1698 0 1 36088
box 0 0 1 1
use contact_8  contact_8_731
timestamp 1624857261
transform 1 0 1698 0 1 36424
box 0 0 1 1
use contact_8  contact_8_730
timestamp 1624857261
transform 1 0 1698 0 1 36760
box 0 0 1 1
use contact_8  contact_8_729
timestamp 1624857261
transform 1 0 1698 0 1 37096
box 0 0 1 1
use contact_8  contact_8_728
timestamp 1624857261
transform 1 0 1698 0 1 37432
box 0 0 1 1
use contact_8  contact_8_727
timestamp 1624857261
transform 1 0 1698 0 1 37768
box 0 0 1 1
use contact_8  contact_8_726
timestamp 1624857261
transform 1 0 1698 0 1 38104
box 0 0 1 1
use contact_8  contact_8_725
timestamp 1624857261
transform 1 0 1698 0 1 38440
box 0 0 1 1
use contact_8  contact_8_724
timestamp 1624857261
transform 1 0 1698 0 1 38776
box 0 0 1 1
use contact_8  contact_8_723
timestamp 1624857261
transform 1 0 1698 0 1 39112
box 0 0 1 1
use contact_8  contact_8_722
timestamp 1624857261
transform 1 0 1698 0 1 39448
box 0 0 1 1
use contact_8  contact_8_721
timestamp 1624857261
transform 1 0 1698 0 1 39784
box 0 0 1 1
use contact_8  contact_8_720
timestamp 1624857261
transform 1 0 1698 0 1 40120
box 0 0 1 1
use contact_8  contact_8_719
timestamp 1624857261
transform 1 0 1698 0 1 40456
box 0 0 1 1
use contact_8  contact_8_718
timestamp 1624857261
transform 1 0 1698 0 1 40792
box 0 0 1 1
use contact_8  contact_8_717
timestamp 1624857261
transform 1 0 1698 0 1 41128
box 0 0 1 1
use contact_8  contact_8_716
timestamp 1624857261
transform 1 0 1698 0 1 41464
box 0 0 1 1
use contact_8  contact_8_715
timestamp 1624857261
transform 1 0 1698 0 1 41800
box 0 0 1 1
use contact_8  contact_8_714
timestamp 1624857261
transform 1 0 1698 0 1 42136
box 0 0 1 1
use contact_8  contact_8_713
timestamp 1624857261
transform 1 0 1698 0 1 42472
box 0 0 1 1
use contact_8  contact_8_712
timestamp 1624857261
transform 1 0 1698 0 1 42808
box 0 0 1 1
use contact_8  contact_8_711
timestamp 1624857261
transform 1 0 1698 0 1 43144
box 0 0 1 1
use contact_8  contact_8_710
timestamp 1624857261
transform 1 0 1698 0 1 43480
box 0 0 1 1
use contact_8  contact_8_709
timestamp 1624857261
transform 1 0 1698 0 1 43816
box 0 0 1 1
use contact_8  contact_8_708
timestamp 1624857261
transform 1 0 1698 0 1 44152
box 0 0 1 1
use contact_8  contact_8_707
timestamp 1624857261
transform 1 0 1698 0 1 44488
box 0 0 1 1
use contact_8  contact_8_706
timestamp 1624857261
transform 1 0 1698 0 1 44824
box 0 0 1 1
use contact_8  contact_8_705
timestamp 1624857261
transform 1 0 1698 0 1 45160
box 0 0 1 1
use contact_8  contact_8_704
timestamp 1624857261
transform 1 0 1698 0 1 45496
box 0 0 1 1
use contact_8  contact_8_703
timestamp 1624857261
transform 1 0 1698 0 1 45832
box 0 0 1 1
use contact_8  contact_8_702
timestamp 1624857261
transform 1 0 1698 0 1 46168
box 0 0 1 1
use contact_8  contact_8_701
timestamp 1624857261
transform 1 0 1698 0 1 46504
box 0 0 1 1
use contact_8  contact_8_700
timestamp 1624857261
transform 1 0 1698 0 1 46840
box 0 0 1 1
use contact_8  contact_8_699
timestamp 1624857261
transform 1 0 1698 0 1 47176
box 0 0 1 1
use contact_8  contact_8_698
timestamp 1624857261
transform 1 0 1698 0 1 47512
box 0 0 1 1
use contact_8  contact_8_697
timestamp 1624857261
transform 1 0 1698 0 1 47848
box 0 0 1 1
use contact_8  contact_8_696
timestamp 1624857261
transform 1 0 1698 0 1 48184
box 0 0 1 1
use contact_8  contact_8_695
timestamp 1624857261
transform 1 0 1698 0 1 48520
box 0 0 1 1
use contact_8  contact_8_694
timestamp 1624857261
transform 1 0 1698 0 1 48856
box 0 0 1 1
use contact_8  contact_8_693
timestamp 1624857261
transform 1 0 1698 0 1 49192
box 0 0 1 1
use contact_8  contact_8_692
timestamp 1624857261
transform 1 0 1698 0 1 49528
box 0 0 1 1
use contact_8  contact_8_691
timestamp 1624857261
transform 1 0 1698 0 1 49864
box 0 0 1 1
use contact_8  contact_8_690
timestamp 1624857261
transform 1 0 1698 0 1 50200
box 0 0 1 1
use contact_8  contact_8_689
timestamp 1624857261
transform 1 0 1698 0 1 50536
box 0 0 1 1
use contact_8  contact_8_688
timestamp 1624857261
transform 1 0 1698 0 1 50872
box 0 0 1 1
use contact_8  contact_8_687
timestamp 1624857261
transform 1 0 1698 0 1 51208
box 0 0 1 1
use contact_8  contact_8_686
timestamp 1624857261
transform 1 0 1698 0 1 51544
box 0 0 1 1
use contact_8  contact_8_685
timestamp 1624857261
transform 1 0 1698 0 1 51880
box 0 0 1 1
use contact_8  contact_8_684
timestamp 1624857261
transform 1 0 1698 0 1 52216
box 0 0 1 1
use contact_8  contact_8_683
timestamp 1624857261
transform 1 0 1698 0 1 52552
box 0 0 1 1
use contact_8  contact_8_682
timestamp 1624857261
transform 1 0 1698 0 1 52888
box 0 0 1 1
use contact_8  contact_8_681
timestamp 1624857261
transform 1 0 1698 0 1 53224
box 0 0 1 1
use contact_8  contact_8_680
timestamp 1624857261
transform 1 0 1698 0 1 53560
box 0 0 1 1
use contact_8  contact_8_679
timestamp 1624857261
transform 1 0 1698 0 1 53896
box 0 0 1 1
use contact_8  contact_8_678
timestamp 1624857261
transform 1 0 1698 0 1 54232
box 0 0 1 1
use contact_8  contact_8_677
timestamp 1624857261
transform 1 0 1698 0 1 54568
box 0 0 1 1
use contact_8  contact_8_676
timestamp 1624857261
transform 1 0 1698 0 1 54904
box 0 0 1 1
use contact_8  contact_8_675
timestamp 1624857261
transform 1 0 1698 0 1 55240
box 0 0 1 1
use contact_8  contact_8_674
timestamp 1624857261
transform 1 0 1698 0 1 55576
box 0 0 1 1
use contact_8  contact_8_673
timestamp 1624857261
transform 1 0 1698 0 1 55912
box 0 0 1 1
use contact_8  contact_8_672
timestamp 1624857261
transform 1 0 1698 0 1 56248
box 0 0 1 1
use contact_8  contact_8_671
timestamp 1624857261
transform 1 0 1698 0 1 56584
box 0 0 1 1
use contact_8  contact_8_670
timestamp 1624857261
transform 1 0 1698 0 1 56920
box 0 0 1 1
use contact_8  contact_8_669
timestamp 1624857261
transform 1 0 1698 0 1 57256
box 0 0 1 1
use contact_8  contact_8_668
timestamp 1624857261
transform 1 0 1698 0 1 57592
box 0 0 1 1
use contact_8  contact_8_667
timestamp 1624857261
transform 1 0 1698 0 1 57928
box 0 0 1 1
use contact_8  contact_8_666
timestamp 1624857261
transform 1 0 1698 0 1 58264
box 0 0 1 1
use contact_8  contact_8_665
timestamp 1624857261
transform 1 0 1698 0 1 58600
box 0 0 1 1
use contact_8  contact_8_664
timestamp 1624857261
transform 1 0 1698 0 1 58936
box 0 0 1 1
use contact_8  contact_8_663
timestamp 1624857261
transform 1 0 1698 0 1 59272
box 0 0 1 1
use contact_8  contact_8_662
timestamp 1624857261
transform 1 0 1698 0 1 59608
box 0 0 1 1
use contact_8  contact_8_661
timestamp 1624857261
transform 1 0 1698 0 1 59944
box 0 0 1 1
use contact_8  contact_8_660
timestamp 1624857261
transform 1 0 1698 0 1 60280
box 0 0 1 1
use contact_8  contact_8_659
timestamp 1624857261
transform 1 0 1698 0 1 60616
box 0 0 1 1
use contact_8  contact_8_658
timestamp 1624857261
transform 1 0 1698 0 1 60952
box 0 0 1 1
use contact_8  contact_8_657
timestamp 1624857261
transform 1 0 1698 0 1 61288
box 0 0 1 1
use contact_8  contact_8_656
timestamp 1624857261
transform 1 0 1698 0 1 61624
box 0 0 1 1
use contact_8  contact_8_655
timestamp 1624857261
transform 1 0 1698 0 1 61960
box 0 0 1 1
use contact_8  contact_8_654
timestamp 1624857261
transform 1 0 1698 0 1 62296
box 0 0 1 1
use contact_8  contact_8_653
timestamp 1624857261
transform 1 0 1698 0 1 62632
box 0 0 1 1
use contact_8  contact_8_652
timestamp 1624857261
transform 1 0 1698 0 1 62968
box 0 0 1 1
use contact_8  contact_8_651
timestamp 1624857261
transform 1 0 1698 0 1 63304
box 0 0 1 1
use contact_8  contact_8_650
timestamp 1624857261
transform 1 0 1698 0 1 63640
box 0 0 1 1
use contact_8  contact_8_649
timestamp 1624857261
transform 1 0 1698 0 1 63976
box 0 0 1 1
use contact_8  contact_8_648
timestamp 1624857261
transform 1 0 1698 0 1 64312
box 0 0 1 1
use contact_8  contact_8_647
timestamp 1624857261
transform 1 0 1698 0 1 64648
box 0 0 1 1
use contact_8  contact_8_646
timestamp 1624857261
transform 1 0 1698 0 1 64984
box 0 0 1 1
use contact_8  contact_8_645
timestamp 1624857261
transform 1 0 1698 0 1 65320
box 0 0 1 1
use contact_8  contact_8_644
timestamp 1624857261
transform 1 0 1698 0 1 65656
box 0 0 1 1
use contact_8  contact_8_643
timestamp 1624857261
transform 1 0 1698 0 1 65992
box 0 0 1 1
use contact_8  contact_8_642
timestamp 1624857261
transform 1 0 1698 0 1 66328
box 0 0 1 1
use contact_8  contact_8_641
timestamp 1624857261
transform 1 0 1698 0 1 66664
box 0 0 1 1
use contact_8  contact_8_640
timestamp 1624857261
transform 1 0 1698 0 1 67000
box 0 0 1 1
use contact_8  contact_8_639
timestamp 1624857261
transform 1 0 1698 0 1 67336
box 0 0 1 1
use contact_8  contact_8_638
timestamp 1624857261
transform 1 0 1698 0 1 67672
box 0 0 1 1
use contact_8  contact_8_637
timestamp 1624857261
transform 1 0 1698 0 1 68008
box 0 0 1 1
use contact_8  contact_8_636
timestamp 1624857261
transform 1 0 1698 0 1 68344
box 0 0 1 1
use contact_8  contact_8_635
timestamp 1624857261
transform 1 0 1698 0 1 68680
box 0 0 1 1
use contact_8  contact_8_634
timestamp 1624857261
transform 1 0 1698 0 1 69016
box 0 0 1 1
use contact_8  contact_8_633
timestamp 1624857261
transform 1 0 1698 0 1 69352
box 0 0 1 1
use contact_8  contact_8_632
timestamp 1624857261
transform 1 0 1698 0 1 69688
box 0 0 1 1
use contact_8  contact_8_631
timestamp 1624857261
transform 1 0 1698 0 1 70024
box 0 0 1 1
use contact_8  contact_8_630
timestamp 1624857261
transform 1 0 1698 0 1 70360
box 0 0 1 1
use contact_8  contact_8_629
timestamp 1624857261
transform 1 0 1698 0 1 70696
box 0 0 1 1
use contact_8  contact_8_628
timestamp 1624857261
transform 1 0 1698 0 1 71032
box 0 0 1 1
use contact_8  contact_8_627
timestamp 1624857261
transform 1 0 1698 0 1 71368
box 0 0 1 1
use contact_8  contact_8_626
timestamp 1624857261
transform 1 0 1698 0 1 71704
box 0 0 1 1
use contact_8  contact_8_625
timestamp 1624857261
transform 1 0 1698 0 1 72040
box 0 0 1 1
use contact_8  contact_8_624
timestamp 1624857261
transform 1 0 1698 0 1 72376
box 0 0 1 1
use contact_8  contact_8_623
timestamp 1624857261
transform 1 0 1698 0 1 72712
box 0 0 1 1
use contact_8  contact_8_622
timestamp 1624857261
transform 1 0 1698 0 1 73048
box 0 0 1 1
use contact_8  contact_8_621
timestamp 1624857261
transform 1 0 1698 0 1 73384
box 0 0 1 1
use contact_8  contact_8_620
timestamp 1624857261
transform 1 0 1698 0 1 73720
box 0 0 1 1
use contact_8  contact_8_619
timestamp 1624857261
transform 1 0 1698 0 1 74056
box 0 0 1 1
use contact_8  contact_8_618
timestamp 1624857261
transform 1 0 1698 0 1 74392
box 0 0 1 1
use contact_8  contact_8_617
timestamp 1624857261
transform 1 0 1698 0 1 74728
box 0 0 1 1
use contact_8  contact_8_616
timestamp 1624857261
transform 1 0 1698 0 1 75064
box 0 0 1 1
use contact_8  contact_8_615
timestamp 1624857261
transform 1 0 1698 0 1 75400
box 0 0 1 1
use contact_8  contact_8_614
timestamp 1624857261
transform 1 0 1698 0 1 75736
box 0 0 1 1
use contact_8  contact_8_613
timestamp 1624857261
transform 1 0 1698 0 1 76072
box 0 0 1 1
use contact_8  contact_8_612
timestamp 1624857261
transform 1 0 1698 0 1 76408
box 0 0 1 1
use contact_8  contact_8_611
timestamp 1624857261
transform 1 0 1698 0 1 76744
box 0 0 1 1
use contact_8  contact_8_610
timestamp 1624857261
transform 1 0 1698 0 1 77080
box 0 0 1 1
use contact_8  contact_8_609
timestamp 1624857261
transform 1 0 1698 0 1 77416
box 0 0 1 1
use contact_8  contact_8_608
timestamp 1624857261
transform 1 0 1698 0 1 77752
box 0 0 1 1
use contact_8  contact_8_607
timestamp 1624857261
transform 1 0 1698 0 1 78088
box 0 0 1 1
use contact_8  contact_8_606
timestamp 1624857261
transform 1 0 1698 0 1 78424
box 0 0 1 1
use contact_8  contact_8_605
timestamp 1624857261
transform 1 0 1698 0 1 78760
box 0 0 1 1
use contact_8  contact_8_604
timestamp 1624857261
transform 1 0 1698 0 1 79096
box 0 0 1 1
use contact_8  contact_8_603
timestamp 1624857261
transform 1 0 1698 0 1 79432
box 0 0 1 1
use contact_8  contact_8_602
timestamp 1624857261
transform 1 0 1698 0 1 79768
box 0 0 1 1
use contact_8  contact_8_601
timestamp 1624857261
transform 1 0 1698 0 1 80104
box 0 0 1 1
use contact_8  contact_8_600
timestamp 1624857261
transform 1 0 1698 0 1 80440
box 0 0 1 1
use contact_8  contact_8_599
timestamp 1624857261
transform 1 0 1698 0 1 80776
box 0 0 1 1
use contact_8  contact_8_598
timestamp 1624857261
transform 1 0 1698 0 1 81112
box 0 0 1 1
use contact_8  contact_8_597
timestamp 1624857261
transform 1 0 1698 0 1 81448
box 0 0 1 1
use contact_8  contact_8_596
timestamp 1624857261
transform 1 0 1698 0 1 81784
box 0 0 1 1
use contact_8  contact_8_595
timestamp 1624857261
transform 1 0 1698 0 1 82120
box 0 0 1 1
use contact_8  contact_8_594
timestamp 1624857261
transform 1 0 1698 0 1 82456
box 0 0 1 1
use contact_8  contact_8_593
timestamp 1624857261
transform 1 0 1698 0 1 82792
box 0 0 1 1
use contact_8  contact_8_592
timestamp 1624857261
transform 1 0 1698 0 1 83128
box 0 0 1 1
use contact_8  contact_8_591
timestamp 1624857261
transform 1 0 1698 0 1 83464
box 0 0 1 1
use contact_8  contact_8_590
timestamp 1624857261
transform 1 0 1698 0 1 83800
box 0 0 1 1
use contact_8  contact_8_589
timestamp 1624857261
transform 1 0 1698 0 1 84136
box 0 0 1 1
use contact_8  contact_8_588
timestamp 1624857261
transform 1 0 1698 0 1 84472
box 0 0 1 1
use contact_8  contact_8_587
timestamp 1624857261
transform 1 0 1698 0 1 84808
box 0 0 1 1
use contact_8  contact_8_586
timestamp 1624857261
transform 1 0 1698 0 1 85144
box 0 0 1 1
use contact_8  contact_8_585
timestamp 1624857261
transform 1 0 1698 0 1 85480
box 0 0 1 1
use contact_8  contact_8_584
timestamp 1624857261
transform 1 0 1698 0 1 85816
box 0 0 1 1
use contact_8  contact_8_583
timestamp 1624857261
transform 1 0 1698 0 1 86152
box 0 0 1 1
use contact_8  contact_8_582
timestamp 1624857261
transform 1 0 1698 0 1 86488
box 0 0 1 1
use contact_8  contact_8_581
timestamp 1624857261
transform 1 0 1698 0 1 86824
box 0 0 1 1
use contact_8  contact_8_580
timestamp 1624857261
transform 1 0 1698 0 1 87160
box 0 0 1 1
use contact_8  contact_8_579
timestamp 1624857261
transform 1 0 1698 0 1 87496
box 0 0 1 1
use contact_8  contact_8_578
timestamp 1624857261
transform 1 0 1698 0 1 87832
box 0 0 1 1
use contact_8  contact_8_577
timestamp 1624857261
transform 1 0 1698 0 1 88168
box 0 0 1 1
use contact_8  contact_8_576
timestamp 1624857261
transform 1 0 1698 0 1 88504
box 0 0 1 1
use contact_8  contact_8_575
timestamp 1624857261
transform 1 0 1698 0 1 88840
box 0 0 1 1
use contact_8  contact_8_574
timestamp 1624857261
transform 1 0 1698 0 1 89176
box 0 0 1 1
use contact_8  contact_8_573
timestamp 1624857261
transform 1 0 1698 0 1 89512
box 0 0 1 1
use contact_8  contact_8_572
timestamp 1624857261
transform 1 0 1698 0 1 89848
box 0 0 1 1
use contact_8  contact_8_571
timestamp 1624857261
transform 1 0 1698 0 1 90184
box 0 0 1 1
use contact_8  contact_8_570
timestamp 1624857261
transform 1 0 1698 0 1 90520
box 0 0 1 1
use contact_8  contact_8_569
timestamp 1624857261
transform 1 0 1698 0 1 90856
box 0 0 1 1
use contact_8  contact_8_568
timestamp 1624857261
transform 1 0 1698 0 1 91192
box 0 0 1 1
use contact_8  contact_8_567
timestamp 1624857261
transform 1 0 1698 0 1 91528
box 0 0 1 1
use contact_8  contact_8_566
timestamp 1624857261
transform 1 0 1698 0 1 91864
box 0 0 1 1
use contact_8  contact_8_565
timestamp 1624857261
transform 1 0 1698 0 1 92200
box 0 0 1 1
use contact_8  contact_8_564
timestamp 1624857261
transform 1 0 1698 0 1 92536
box 0 0 1 1
use contact_8  contact_8_563
timestamp 1624857261
transform 1 0 1698 0 1 92872
box 0 0 1 1
use contact_8  contact_8_562
timestamp 1624857261
transform 1 0 1698 0 1 93208
box 0 0 1 1
use contact_8  contact_8_561
timestamp 1624857261
transform 1 0 1698 0 1 93544
box 0 0 1 1
use contact_8  contact_8_560
timestamp 1624857261
transform 1 0 1698 0 1 93880
box 0 0 1 1
use contact_8  contact_8_559
timestamp 1624857261
transform 1 0 1698 0 1 94216
box 0 0 1 1
use contact_8  contact_8_558
timestamp 1624857261
transform 1 0 1698 0 1 94552
box 0 0 1 1
use contact_8  contact_8_557
timestamp 1624857261
transform 1 0 1698 0 1 94888
box 0 0 1 1
use contact_8  contact_8_556
timestamp 1624857261
transform 1 0 1698 0 1 95224
box 0 0 1 1
use contact_8  contact_8_555
timestamp 1624857261
transform 1 0 1698 0 1 95560
box 0 0 1 1
use contact_8  contact_8_554
timestamp 1624857261
transform 1 0 1698 0 1 95896
box 0 0 1 1
use contact_8  contact_8_553
timestamp 1624857261
transform 1 0 1698 0 1 96232
box 0 0 1 1
use contact_8  contact_8_552
timestamp 1624857261
transform 1 0 1698 0 1 96568
box 0 0 1 1
use contact_8  contact_8_551
timestamp 1624857261
transform 1 0 1698 0 1 96904
box 0 0 1 1
use contact_8  contact_8_550
timestamp 1624857261
transform 1 0 1698 0 1 97240
box 0 0 1 1
use contact_8  contact_8_549
timestamp 1624857261
transform 1 0 1698 0 1 97576
box 0 0 1 1
use contact_8  contact_8_548
timestamp 1624857261
transform 1 0 1698 0 1 97912
box 0 0 1 1
use contact_8  contact_8_547
timestamp 1624857261
transform 1 0 1698 0 1 98248
box 0 0 1 1
use contact_8  contact_8_546
timestamp 1624857261
transform 1 0 1698 0 1 98584
box 0 0 1 1
use contact_8  contact_8_545
timestamp 1624857261
transform 1 0 1698 0 1 98920
box 0 0 1 1
use contact_8  contact_8_544
timestamp 1624857261
transform 1 0 1698 0 1 99256
box 0 0 1 1
use contact_8  contact_8_543
timestamp 1624857261
transform 1 0 1698 0 1 99592
box 0 0 1 1
use contact_8  contact_8_542
timestamp 1624857261
transform 1 0 1698 0 1 99928
box 0 0 1 1
use contact_8  contact_8_541
timestamp 1624857261
transform 1 0 1698 0 1 100264
box 0 0 1 1
use contact_8  contact_8_540
timestamp 1624857261
transform 1 0 1698 0 1 100600
box 0 0 1 1
use contact_8  contact_8_539
timestamp 1624857261
transform 1 0 1698 0 1 100936
box 0 0 1 1
use contact_8  contact_8_538
timestamp 1624857261
transform 1 0 1698 0 1 101272
box 0 0 1 1
use contact_8  contact_8_537
timestamp 1624857261
transform 1 0 1698 0 1 101608
box 0 0 1 1
use contact_8  contact_8_536
timestamp 1624857261
transform 1 0 1698 0 1 101944
box 0 0 1 1
use contact_8  contact_8_535
timestamp 1624857261
transform 1 0 1698 0 1 102280
box 0 0 1 1
use contact_8  contact_8_534
timestamp 1624857261
transform 1 0 1698 0 1 102616
box 0 0 1 1
use contact_8  contact_8_533
timestamp 1624857261
transform 1 0 1698 0 1 102952
box 0 0 1 1
use contact_8  contact_8_532
timestamp 1624857261
transform 1 0 1698 0 1 103288
box 0 0 1 1
use contact_8  contact_8_531
timestamp 1624857261
transform 1 0 1698 0 1 103624
box 0 0 1 1
use contact_8  contact_8_530
timestamp 1624857261
transform 1 0 1698 0 1 103960
box 0 0 1 1
use contact_8  contact_8_529
timestamp 1624857261
transform 1 0 1698 0 1 104296
box 0 0 1 1
use contact_8  contact_8_528
timestamp 1624857261
transform 1 0 1698 0 1 104632
box 0 0 1 1
use contact_8  contact_8_527
timestamp 1624857261
transform 1 0 1698 0 1 104968
box 0 0 1 1
use contact_8  contact_8_526
timestamp 1624857261
transform 1 0 1698 0 1 105304
box 0 0 1 1
use contact_8  contact_8_525
timestamp 1624857261
transform 1 0 1698 0 1 105640
box 0 0 1 1
use contact_8  contact_8_524
timestamp 1624857261
transform 1 0 1698 0 1 105976
box 0 0 1 1
use contact_8  contact_8_523
timestamp 1624857261
transform 1 0 1698 0 1 106312
box 0 0 1 1
use contact_8  contact_8_522
timestamp 1624857261
transform 1 0 1698 0 1 106648
box 0 0 1 1
use contact_8  contact_8_521
timestamp 1624857261
transform 1 0 1698 0 1 106984
box 0 0 1 1
use contact_8  contact_8_520
timestamp 1624857261
transform 1 0 1698 0 1 107320
box 0 0 1 1
use contact_8  contact_8_519
timestamp 1624857261
transform 1 0 1698 0 1 107656
box 0 0 1 1
use contact_8  contact_8_518
timestamp 1624857261
transform 1 0 1698 0 1 107992
box 0 0 1 1
use contact_8  contact_8_517
timestamp 1624857261
transform 1 0 1698 0 1 108328
box 0 0 1 1
use contact_8  contact_8_516
timestamp 1624857261
transform 1 0 1698 0 1 108664
box 0 0 1 1
use contact_8  contact_8_515
timestamp 1624857261
transform 1 0 1698 0 1 109000
box 0 0 1 1
use contact_8  contact_8_514
timestamp 1624857261
transform 1 0 1698 0 1 109336
box 0 0 1 1
use contact_8  contact_8_513
timestamp 1624857261
transform 1 0 1698 0 1 109672
box 0 0 1 1
use contact_8  contact_8_512
timestamp 1624857261
transform 1 0 1698 0 1 110008
box 0 0 1 1
use contact_8  contact_8_511
timestamp 1624857261
transform 1 0 1698 0 1 110344
box 0 0 1 1
use contact_8  contact_8_510
timestamp 1624857261
transform 1 0 1698 0 1 110680
box 0 0 1 1
use contact_8  contact_8_509
timestamp 1624857261
transform 1 0 1698 0 1 111016
box 0 0 1 1
use contact_8  contact_8_508
timestamp 1624857261
transform 1 0 1698 0 1 111352
box 0 0 1 1
use contact_8  contact_8_507
timestamp 1624857261
transform 1 0 1698 0 1 111688
box 0 0 1 1
use contact_8  contact_8_506
timestamp 1624857261
transform 1 0 1698 0 1 112024
box 0 0 1 1
use contact_8  contact_8_505
timestamp 1624857261
transform 1 0 1698 0 1 112360
box 0 0 1 1
use contact_8  contact_8_504
timestamp 1624857261
transform 1 0 1698 0 1 112696
box 0 0 1 1
use contact_8  contact_8_503
timestamp 1624857261
transform 1 0 1698 0 1 113032
box 0 0 1 1
use contact_8  contact_8_502
timestamp 1624857261
transform 1 0 1698 0 1 113368
box 0 0 1 1
use contact_8  contact_8_501
timestamp 1624857261
transform 1 0 1698 0 1 113704
box 0 0 1 1
use contact_8  contact_8_500
timestamp 1624857261
transform 1 0 1698 0 1 114040
box 0 0 1 1
use contact_8  contact_8_499
timestamp 1624857261
transform 1 0 1698 0 1 114376
box 0 0 1 1
use contact_8  contact_8_498
timestamp 1624857261
transform 1 0 1698 0 1 114712
box 0 0 1 1
use contact_8  contact_8_497
timestamp 1624857261
transform 1 0 1698 0 1 115048
box 0 0 1 1
use contact_8  contact_8_496
timestamp 1624857261
transform 1 0 1698 0 1 115384
box 0 0 1 1
use contact_8  contact_8_495
timestamp 1624857261
transform 1 0 1698 0 1 115720
box 0 0 1 1
use contact_8  contact_8_494
timestamp 1624857261
transform 1 0 1698 0 1 116056
box 0 0 1 1
use contact_8  contact_8_493
timestamp 1624857261
transform 1 0 1698 0 1 116392
box 0 0 1 1
use contact_8  contact_8_492
timestamp 1624857261
transform 1 0 1698 0 1 116728
box 0 0 1 1
use contact_8  contact_8_491
timestamp 1624857261
transform 1 0 1698 0 1 117064
box 0 0 1 1
use contact_8  contact_8_490
timestamp 1624857261
transform 1 0 1698 0 1 117400
box 0 0 1 1
use contact_8  contact_8_489
timestamp 1624857261
transform 1 0 1698 0 1 117736
box 0 0 1 1
use contact_8  contact_8_488
timestamp 1624857261
transform 1 0 1698 0 1 118072
box 0 0 1 1
use contact_8  contact_8_487
timestamp 1624857261
transform 1 0 1698 0 1 118408
box 0 0 1 1
use contact_8  contact_8_486
timestamp 1624857261
transform 1 0 1698 0 1 118744
box 0 0 1 1
use contact_8  contact_8_485
timestamp 1624857261
transform 1 0 1698 0 1 119080
box 0 0 1 1
use contact_8  contact_8_484
timestamp 1624857261
transform 1 0 1698 0 1 119416
box 0 0 1 1
use contact_8  contact_8_483
timestamp 1624857261
transform 1 0 1698 0 1 119752
box 0 0 1 1
use contact_8  contact_8_482
timestamp 1624857261
transform 1 0 1698 0 1 120088
box 0 0 1 1
use contact_8  contact_8_481
timestamp 1624857261
transform 1 0 1698 0 1 120424
box 0 0 1 1
use contact_8  contact_8_480
timestamp 1624857261
transform 1 0 1698 0 1 120760
box 0 0 1 1
use contact_8  contact_8_479
timestamp 1624857261
transform 1 0 1698 0 1 121096
box 0 0 1 1
use contact_8  contact_8_478
timestamp 1624857261
transform 1 0 1698 0 1 121432
box 0 0 1 1
use contact_8  contact_8_477
timestamp 1624857261
transform 1 0 1698 0 1 121768
box 0 0 1 1
use contact_8  contact_8_476
timestamp 1624857261
transform 1 0 1698 0 1 122104
box 0 0 1 1
use contact_8  contact_8_475
timestamp 1624857261
transform 1 0 1698 0 1 122440
box 0 0 1 1
use contact_8  contact_8_474
timestamp 1624857261
transform 1 0 1698 0 1 122776
box 0 0 1 1
use contact_8  contact_8_473
timestamp 1624857261
transform 1 0 1698 0 1 123112
box 0 0 1 1
use contact_8  contact_8_472
timestamp 1624857261
transform 1 0 1698 0 1 123448
box 0 0 1 1
use contact_8  contact_8_471
timestamp 1624857261
transform 1 0 1698 0 1 123784
box 0 0 1 1
use contact_8  contact_8_470
timestamp 1624857261
transform 1 0 1698 0 1 124120
box 0 0 1 1
use contact_8  contact_8_469
timestamp 1624857261
transform 1 0 1698 0 1 124456
box 0 0 1 1
use contact_8  contact_8_468
timestamp 1624857261
transform 1 0 1698 0 1 124792
box 0 0 1 1
use contact_8  contact_8_467
timestamp 1624857261
transform 1 0 1698 0 1 125128
box 0 0 1 1
use contact_8  contact_8_466
timestamp 1624857261
transform 1 0 1698 0 1 125464
box 0 0 1 1
use contact_8  contact_8_465
timestamp 1624857261
transform 1 0 1698 0 1 125800
box 0 0 1 1
use contact_8  contact_8_464
timestamp 1624857261
transform 1 0 1698 0 1 126136
box 0 0 1 1
use contact_8  contact_8_463
timestamp 1624857261
transform 1 0 1698 0 1 126472
box 0 0 1 1
use contact_8  contact_8_462
timestamp 1624857261
transform 1 0 1698 0 1 126808
box 0 0 1 1
use contact_8  contact_8_461
timestamp 1624857261
transform 1 0 1698 0 1 127144
box 0 0 1 1
use contact_8  contact_8_460
timestamp 1624857261
transform 1 0 1698 0 1 127480
box 0 0 1 1
use contact_8  contact_8_459
timestamp 1624857261
transform 1 0 1698 0 1 127816
box 0 0 1 1
use contact_8  contact_8_458
timestamp 1624857261
transform 1 0 1698 0 1 128152
box 0 0 1 1
use contact_8  contact_8_457
timestamp 1624857261
transform 1 0 1698 0 1 128488
box 0 0 1 1
use contact_8  contact_8_456
timestamp 1624857261
transform 1 0 1698 0 1 128824
box 0 0 1 1
use contact_8  contact_8_455
timestamp 1624857261
transform 1 0 1698 0 1 129160
box 0 0 1 1
use contact_8  contact_8_454
timestamp 1624857261
transform 1 0 1698 0 1 129496
box 0 0 1 1
use contact_8  contact_8_453
timestamp 1624857261
transform 1 0 1698 0 1 129832
box 0 0 1 1
use contact_8  contact_8_452
timestamp 1624857261
transform 1 0 1698 0 1 130168
box 0 0 1 1
use contact_8  contact_8_451
timestamp 1624857261
transform 1 0 1698 0 1 130504
box 0 0 1 1
use contact_8  contact_8_450
timestamp 1624857261
transform 1 0 1698 0 1 130840
box 0 0 1 1
use contact_8  contact_8_449
timestamp 1624857261
transform 1 0 1698 0 1 131176
box 0 0 1 1
use contact_8  contact_8_448
timestamp 1624857261
transform 1 0 1698 0 1 131512
box 0 0 1 1
use contact_8  contact_8_447
timestamp 1624857261
transform 1 0 1698 0 1 131848
box 0 0 1 1
use contact_8  contact_8_446
timestamp 1624857261
transform 1 0 1698 0 1 132184
box 0 0 1 1
use contact_8  contact_8_445
timestamp 1624857261
transform 1 0 1698 0 1 132520
box 0 0 1 1
use contact_8  contact_8_444
timestamp 1624857261
transform 1 0 1698 0 1 132856
box 0 0 1 1
use contact_8  contact_8_443
timestamp 1624857261
transform 1 0 1698 0 1 133192
box 0 0 1 1
use contact_8  contact_8_442
timestamp 1624857261
transform 1 0 1698 0 1 133528
box 0 0 1 1
use contact_8  contact_8_441
timestamp 1624857261
transform 1 0 1698 0 1 133864
box 0 0 1 1
use contact_8  contact_8_440
timestamp 1624857261
transform 1 0 1698 0 1 134200
box 0 0 1 1
use contact_8  contact_8_439
timestamp 1624857261
transform 1 0 1698 0 1 134536
box 0 0 1 1
use contact_8  contact_8_438
timestamp 1624857261
transform 1 0 1698 0 1 134872
box 0 0 1 1
use contact_8  contact_8_437
timestamp 1624857261
transform 1 0 1698 0 1 135208
box 0 0 1 1
use contact_8  contact_8_436
timestamp 1624857261
transform 1 0 1698 0 1 135544
box 0 0 1 1
use contact_8  contact_8_435
timestamp 1624857261
transform 1 0 1698 0 1 135880
box 0 0 1 1
use contact_8  contact_8_434
timestamp 1624857261
transform 1 0 1698 0 1 136216
box 0 0 1 1
use contact_8  contact_8_433
timestamp 1624857261
transform 1 0 1698 0 1 136552
box 0 0 1 1
use contact_8  contact_8_432
timestamp 1624857261
transform 1 0 1698 0 1 136888
box 0 0 1 1
use contact_8  contact_8_431
timestamp 1624857261
transform 1 0 1698 0 1 137224
box 0 0 1 1
use contact_8  contact_8_430
timestamp 1624857261
transform 1 0 1698 0 1 137560
box 0 0 1 1
use contact_8  contact_8_429
timestamp 1624857261
transform 1 0 1698 0 1 137896
box 0 0 1 1
use contact_8  contact_8_428
timestamp 1624857261
transform 1 0 1698 0 1 138232
box 0 0 1 1
use contact_8  contact_8_427
timestamp 1624857261
transform 1 0 1698 0 1 138568
box 0 0 1 1
use contact_8  contact_8_426
timestamp 1624857261
transform 1 0 1698 0 1 138904
box 0 0 1 1
use contact_8  contact_8_425
timestamp 1624857261
transform 1 0 1698 0 1 139240
box 0 0 1 1
use contact_8  contact_8_424
timestamp 1624857261
transform 1 0 1698 0 1 139576
box 0 0 1 1
use contact_8  contact_8_423
timestamp 1624857261
transform 1 0 1698 0 1 139912
box 0 0 1 1
use contact_8  contact_8_422
timestamp 1624857261
transform 1 0 1698 0 1 140248
box 0 0 1 1
use contact_8  contact_8_421
timestamp 1624857261
transform 1 0 1698 0 1 140584
box 0 0 1 1
use contact_8  contact_8_420
timestamp 1624857261
transform 1 0 1698 0 1 140920
box 0 0 1 1
use contact_8  contact_8_419
timestamp 1624857261
transform 1 0 1698 0 1 141256
box 0 0 1 1
use contact_8  contact_8_418
timestamp 1624857261
transform 1 0 1698 0 1 141592
box 0 0 1 1
use contact_8  contact_8_417
timestamp 1624857261
transform 1 0 1698 0 1 141928
box 0 0 1 1
use contact_8  contact_8_416
timestamp 1624857261
transform 1 0 216904 0 1 2152
box 0 0 1 1
use contact_8  contact_8_415
timestamp 1624857261
transform 1 0 216904 0 1 2488
box 0 0 1 1
use contact_8  contact_8_414
timestamp 1624857261
transform 1 0 216904 0 1 2824
box 0 0 1 1
use contact_8  contact_8_413
timestamp 1624857261
transform 1 0 216904 0 1 3160
box 0 0 1 1
use contact_8  contact_8_412
timestamp 1624857261
transform 1 0 216904 0 1 3496
box 0 0 1 1
use contact_8  contact_8_411
timestamp 1624857261
transform 1 0 216904 0 1 3832
box 0 0 1 1
use contact_8  contact_8_410
timestamp 1624857261
transform 1 0 216904 0 1 4168
box 0 0 1 1
use contact_8  contact_8_409
timestamp 1624857261
transform 1 0 216904 0 1 4504
box 0 0 1 1
use contact_8  contact_8_408
timestamp 1624857261
transform 1 0 216904 0 1 4840
box 0 0 1 1
use contact_8  contact_8_407
timestamp 1624857261
transform 1 0 216904 0 1 5176
box 0 0 1 1
use contact_8  contact_8_406
timestamp 1624857261
transform 1 0 216904 0 1 5512
box 0 0 1 1
use contact_8  contact_8_405
timestamp 1624857261
transform 1 0 216904 0 1 5848
box 0 0 1 1
use contact_8  contact_8_404
timestamp 1624857261
transform 1 0 216904 0 1 6184
box 0 0 1 1
use contact_8  contact_8_403
timestamp 1624857261
transform 1 0 216904 0 1 6520
box 0 0 1 1
use contact_8  contact_8_402
timestamp 1624857261
transform 1 0 216904 0 1 6856
box 0 0 1 1
use contact_8  contact_8_401
timestamp 1624857261
transform 1 0 216904 0 1 7192
box 0 0 1 1
use contact_8  contact_8_400
timestamp 1624857261
transform 1 0 216904 0 1 7528
box 0 0 1 1
use contact_8  contact_8_399
timestamp 1624857261
transform 1 0 216904 0 1 7864
box 0 0 1 1
use contact_8  contact_8_398
timestamp 1624857261
transform 1 0 216904 0 1 8200
box 0 0 1 1
use contact_8  contact_8_397
timestamp 1624857261
transform 1 0 216904 0 1 8536
box 0 0 1 1
use contact_8  contact_8_396
timestamp 1624857261
transform 1 0 216904 0 1 8872
box 0 0 1 1
use contact_8  contact_8_395
timestamp 1624857261
transform 1 0 216904 0 1 9208
box 0 0 1 1
use contact_8  contact_8_394
timestamp 1624857261
transform 1 0 216904 0 1 9544
box 0 0 1 1
use contact_8  contact_8_393
timestamp 1624857261
transform 1 0 216904 0 1 9880
box 0 0 1 1
use contact_8  contact_8_392
timestamp 1624857261
transform 1 0 216904 0 1 10216
box 0 0 1 1
use contact_8  contact_8_391
timestamp 1624857261
transform 1 0 216904 0 1 10552
box 0 0 1 1
use contact_8  contact_8_390
timestamp 1624857261
transform 1 0 216904 0 1 10888
box 0 0 1 1
use contact_8  contact_8_389
timestamp 1624857261
transform 1 0 216904 0 1 11224
box 0 0 1 1
use contact_8  contact_8_388
timestamp 1624857261
transform 1 0 216904 0 1 11560
box 0 0 1 1
use contact_8  contact_8_387
timestamp 1624857261
transform 1 0 216904 0 1 11896
box 0 0 1 1
use contact_8  contact_8_386
timestamp 1624857261
transform 1 0 216904 0 1 12232
box 0 0 1 1
use contact_8  contact_8_385
timestamp 1624857261
transform 1 0 216904 0 1 12568
box 0 0 1 1
use contact_8  contact_8_384
timestamp 1624857261
transform 1 0 216904 0 1 12904
box 0 0 1 1
use contact_8  contact_8_383
timestamp 1624857261
transform 1 0 216904 0 1 13240
box 0 0 1 1
use contact_8  contact_8_382
timestamp 1624857261
transform 1 0 216904 0 1 13576
box 0 0 1 1
use contact_8  contact_8_381
timestamp 1624857261
transform 1 0 216904 0 1 13912
box 0 0 1 1
use contact_8  contact_8_380
timestamp 1624857261
transform 1 0 216904 0 1 14248
box 0 0 1 1
use contact_8  contact_8_379
timestamp 1624857261
transform 1 0 216904 0 1 14584
box 0 0 1 1
use contact_8  contact_8_378
timestamp 1624857261
transform 1 0 216904 0 1 14920
box 0 0 1 1
use contact_8  contact_8_377
timestamp 1624857261
transform 1 0 216904 0 1 15256
box 0 0 1 1
use contact_8  contact_8_376
timestamp 1624857261
transform 1 0 216904 0 1 15592
box 0 0 1 1
use contact_8  contact_8_375
timestamp 1624857261
transform 1 0 216904 0 1 15928
box 0 0 1 1
use contact_8  contact_8_374
timestamp 1624857261
transform 1 0 216904 0 1 16264
box 0 0 1 1
use contact_8  contact_8_373
timestamp 1624857261
transform 1 0 216904 0 1 16600
box 0 0 1 1
use contact_8  contact_8_372
timestamp 1624857261
transform 1 0 216904 0 1 16936
box 0 0 1 1
use contact_8  contact_8_371
timestamp 1624857261
transform 1 0 216904 0 1 17272
box 0 0 1 1
use contact_8  contact_8_370
timestamp 1624857261
transform 1 0 216904 0 1 17608
box 0 0 1 1
use contact_8  contact_8_369
timestamp 1624857261
transform 1 0 216904 0 1 17944
box 0 0 1 1
use contact_8  contact_8_368
timestamp 1624857261
transform 1 0 216904 0 1 18280
box 0 0 1 1
use contact_8  contact_8_367
timestamp 1624857261
transform 1 0 216904 0 1 18616
box 0 0 1 1
use contact_8  contact_8_366
timestamp 1624857261
transform 1 0 216904 0 1 18952
box 0 0 1 1
use contact_8  contact_8_365
timestamp 1624857261
transform 1 0 216904 0 1 19288
box 0 0 1 1
use contact_8  contact_8_364
timestamp 1624857261
transform 1 0 216904 0 1 19624
box 0 0 1 1
use contact_8  contact_8_363
timestamp 1624857261
transform 1 0 216904 0 1 19960
box 0 0 1 1
use contact_8  contact_8_362
timestamp 1624857261
transform 1 0 216904 0 1 20296
box 0 0 1 1
use contact_8  contact_8_361
timestamp 1624857261
transform 1 0 216904 0 1 20632
box 0 0 1 1
use contact_8  contact_8_360
timestamp 1624857261
transform 1 0 216904 0 1 20968
box 0 0 1 1
use contact_8  contact_8_359
timestamp 1624857261
transform 1 0 216904 0 1 21304
box 0 0 1 1
use contact_8  contact_8_358
timestamp 1624857261
transform 1 0 216904 0 1 21640
box 0 0 1 1
use contact_8  contact_8_357
timestamp 1624857261
transform 1 0 216904 0 1 21976
box 0 0 1 1
use contact_8  contact_8_356
timestamp 1624857261
transform 1 0 216904 0 1 22312
box 0 0 1 1
use contact_8  contact_8_355
timestamp 1624857261
transform 1 0 216904 0 1 22648
box 0 0 1 1
use contact_8  contact_8_354
timestamp 1624857261
transform 1 0 216904 0 1 22984
box 0 0 1 1
use contact_8  contact_8_353
timestamp 1624857261
transform 1 0 216904 0 1 23320
box 0 0 1 1
use contact_8  contact_8_352
timestamp 1624857261
transform 1 0 216904 0 1 23656
box 0 0 1 1
use contact_8  contact_8_351
timestamp 1624857261
transform 1 0 216904 0 1 23992
box 0 0 1 1
use contact_8  contact_8_350
timestamp 1624857261
transform 1 0 216904 0 1 24328
box 0 0 1 1
use contact_8  contact_8_349
timestamp 1624857261
transform 1 0 216904 0 1 24664
box 0 0 1 1
use contact_8  contact_8_348
timestamp 1624857261
transform 1 0 216904 0 1 25000
box 0 0 1 1
use contact_8  contact_8_347
timestamp 1624857261
transform 1 0 216904 0 1 25336
box 0 0 1 1
use contact_8  contact_8_346
timestamp 1624857261
transform 1 0 216904 0 1 25672
box 0 0 1 1
use contact_8  contact_8_345
timestamp 1624857261
transform 1 0 216904 0 1 26008
box 0 0 1 1
use contact_8  contact_8_344
timestamp 1624857261
transform 1 0 216904 0 1 26344
box 0 0 1 1
use contact_8  contact_8_343
timestamp 1624857261
transform 1 0 216904 0 1 26680
box 0 0 1 1
use contact_8  contact_8_342
timestamp 1624857261
transform 1 0 216904 0 1 27016
box 0 0 1 1
use contact_8  contact_8_341
timestamp 1624857261
transform 1 0 216904 0 1 27352
box 0 0 1 1
use contact_8  contact_8_340
timestamp 1624857261
transform 1 0 216904 0 1 27688
box 0 0 1 1
use contact_8  contact_8_339
timestamp 1624857261
transform 1 0 216904 0 1 28024
box 0 0 1 1
use contact_8  contact_8_338
timestamp 1624857261
transform 1 0 216904 0 1 28360
box 0 0 1 1
use contact_8  contact_8_337
timestamp 1624857261
transform 1 0 216904 0 1 28696
box 0 0 1 1
use contact_8  contact_8_336
timestamp 1624857261
transform 1 0 216904 0 1 29032
box 0 0 1 1
use contact_8  contact_8_335
timestamp 1624857261
transform 1 0 216904 0 1 29368
box 0 0 1 1
use contact_8  contact_8_334
timestamp 1624857261
transform 1 0 216904 0 1 29704
box 0 0 1 1
use contact_8  contact_8_333
timestamp 1624857261
transform 1 0 216904 0 1 30040
box 0 0 1 1
use contact_8  contact_8_332
timestamp 1624857261
transform 1 0 216904 0 1 30376
box 0 0 1 1
use contact_8  contact_8_331
timestamp 1624857261
transform 1 0 216904 0 1 30712
box 0 0 1 1
use contact_8  contact_8_330
timestamp 1624857261
transform 1 0 216904 0 1 31048
box 0 0 1 1
use contact_8  contact_8_329
timestamp 1624857261
transform 1 0 216904 0 1 31384
box 0 0 1 1
use contact_8  contact_8_328
timestamp 1624857261
transform 1 0 216904 0 1 31720
box 0 0 1 1
use contact_8  contact_8_327
timestamp 1624857261
transform 1 0 216904 0 1 32056
box 0 0 1 1
use contact_8  contact_8_326
timestamp 1624857261
transform 1 0 216904 0 1 32392
box 0 0 1 1
use contact_8  contact_8_325
timestamp 1624857261
transform 1 0 216904 0 1 32728
box 0 0 1 1
use contact_8  contact_8_324
timestamp 1624857261
transform 1 0 216904 0 1 33064
box 0 0 1 1
use contact_8  contact_8_323
timestamp 1624857261
transform 1 0 216904 0 1 33400
box 0 0 1 1
use contact_8  contact_8_322
timestamp 1624857261
transform 1 0 216904 0 1 33736
box 0 0 1 1
use contact_8  contact_8_321
timestamp 1624857261
transform 1 0 216904 0 1 34072
box 0 0 1 1
use contact_8  contact_8_320
timestamp 1624857261
transform 1 0 216904 0 1 34408
box 0 0 1 1
use contact_8  contact_8_319
timestamp 1624857261
transform 1 0 216904 0 1 34744
box 0 0 1 1
use contact_8  contact_8_318
timestamp 1624857261
transform 1 0 216904 0 1 35080
box 0 0 1 1
use contact_8  contact_8_317
timestamp 1624857261
transform 1 0 216904 0 1 35416
box 0 0 1 1
use contact_8  contact_8_316
timestamp 1624857261
transform 1 0 216904 0 1 35752
box 0 0 1 1
use contact_8  contact_8_315
timestamp 1624857261
transform 1 0 216904 0 1 36088
box 0 0 1 1
use contact_8  contact_8_314
timestamp 1624857261
transform 1 0 216904 0 1 36424
box 0 0 1 1
use contact_8  contact_8_313
timestamp 1624857261
transform 1 0 216904 0 1 36760
box 0 0 1 1
use contact_8  contact_8_312
timestamp 1624857261
transform 1 0 216904 0 1 37096
box 0 0 1 1
use contact_8  contact_8_311
timestamp 1624857261
transform 1 0 216904 0 1 37432
box 0 0 1 1
use contact_8  contact_8_310
timestamp 1624857261
transform 1 0 216904 0 1 37768
box 0 0 1 1
use contact_8  contact_8_309
timestamp 1624857261
transform 1 0 216904 0 1 38104
box 0 0 1 1
use contact_8  contact_8_308
timestamp 1624857261
transform 1 0 216904 0 1 38440
box 0 0 1 1
use contact_8  contact_8_307
timestamp 1624857261
transform 1 0 216904 0 1 38776
box 0 0 1 1
use contact_8  contact_8_306
timestamp 1624857261
transform 1 0 216904 0 1 39112
box 0 0 1 1
use contact_8  contact_8_305
timestamp 1624857261
transform 1 0 216904 0 1 39448
box 0 0 1 1
use contact_8  contact_8_304
timestamp 1624857261
transform 1 0 216904 0 1 39784
box 0 0 1 1
use contact_8  contact_8_303
timestamp 1624857261
transform 1 0 216904 0 1 40120
box 0 0 1 1
use contact_8  contact_8_302
timestamp 1624857261
transform 1 0 216904 0 1 40456
box 0 0 1 1
use contact_8  contact_8_301
timestamp 1624857261
transform 1 0 216904 0 1 40792
box 0 0 1 1
use contact_8  contact_8_300
timestamp 1624857261
transform 1 0 216904 0 1 41128
box 0 0 1 1
use contact_8  contact_8_299
timestamp 1624857261
transform 1 0 216904 0 1 41464
box 0 0 1 1
use contact_8  contact_8_298
timestamp 1624857261
transform 1 0 216904 0 1 41800
box 0 0 1 1
use contact_8  contact_8_297
timestamp 1624857261
transform 1 0 216904 0 1 42136
box 0 0 1 1
use contact_8  contact_8_296
timestamp 1624857261
transform 1 0 216904 0 1 42472
box 0 0 1 1
use contact_8  contact_8_295
timestamp 1624857261
transform 1 0 216904 0 1 42808
box 0 0 1 1
use contact_8  contact_8_294
timestamp 1624857261
transform 1 0 216904 0 1 43144
box 0 0 1 1
use contact_8  contact_8_293
timestamp 1624857261
transform 1 0 216904 0 1 43480
box 0 0 1 1
use contact_8  contact_8_292
timestamp 1624857261
transform 1 0 216904 0 1 43816
box 0 0 1 1
use contact_8  contact_8_291
timestamp 1624857261
transform 1 0 216904 0 1 44152
box 0 0 1 1
use contact_8  contact_8_290
timestamp 1624857261
transform 1 0 216904 0 1 44488
box 0 0 1 1
use contact_8  contact_8_289
timestamp 1624857261
transform 1 0 216904 0 1 44824
box 0 0 1 1
use contact_8  contact_8_288
timestamp 1624857261
transform 1 0 216904 0 1 45160
box 0 0 1 1
use contact_8  contact_8_287
timestamp 1624857261
transform 1 0 216904 0 1 45496
box 0 0 1 1
use contact_8  contact_8_286
timestamp 1624857261
transform 1 0 216904 0 1 45832
box 0 0 1 1
use contact_8  contact_8_285
timestamp 1624857261
transform 1 0 216904 0 1 46168
box 0 0 1 1
use contact_8  contact_8_284
timestamp 1624857261
transform 1 0 216904 0 1 46504
box 0 0 1 1
use contact_8  contact_8_283
timestamp 1624857261
transform 1 0 216904 0 1 46840
box 0 0 1 1
use contact_8  contact_8_282
timestamp 1624857261
transform 1 0 216904 0 1 47176
box 0 0 1 1
use contact_8  contact_8_281
timestamp 1624857261
transform 1 0 216904 0 1 47512
box 0 0 1 1
use contact_8  contact_8_280
timestamp 1624857261
transform 1 0 216904 0 1 47848
box 0 0 1 1
use contact_8  contact_8_279
timestamp 1624857261
transform 1 0 216904 0 1 48184
box 0 0 1 1
use contact_8  contact_8_278
timestamp 1624857261
transform 1 0 216904 0 1 48520
box 0 0 1 1
use contact_8  contact_8_277
timestamp 1624857261
transform 1 0 216904 0 1 48856
box 0 0 1 1
use contact_8  contact_8_276
timestamp 1624857261
transform 1 0 216904 0 1 49192
box 0 0 1 1
use contact_8  contact_8_275
timestamp 1624857261
transform 1 0 216904 0 1 49528
box 0 0 1 1
use contact_8  contact_8_274
timestamp 1624857261
transform 1 0 216904 0 1 49864
box 0 0 1 1
use contact_8  contact_8_273
timestamp 1624857261
transform 1 0 216904 0 1 50200
box 0 0 1 1
use contact_8  contact_8_272
timestamp 1624857261
transform 1 0 216904 0 1 50536
box 0 0 1 1
use contact_8  contact_8_271
timestamp 1624857261
transform 1 0 216904 0 1 50872
box 0 0 1 1
use contact_8  contact_8_270
timestamp 1624857261
transform 1 0 216904 0 1 51208
box 0 0 1 1
use contact_8  contact_8_269
timestamp 1624857261
transform 1 0 216904 0 1 51544
box 0 0 1 1
use contact_8  contact_8_268
timestamp 1624857261
transform 1 0 216904 0 1 51880
box 0 0 1 1
use contact_8  contact_8_267
timestamp 1624857261
transform 1 0 216904 0 1 52216
box 0 0 1 1
use contact_8  contact_8_266
timestamp 1624857261
transform 1 0 216904 0 1 52552
box 0 0 1 1
use contact_8  contact_8_265
timestamp 1624857261
transform 1 0 216904 0 1 52888
box 0 0 1 1
use contact_8  contact_8_264
timestamp 1624857261
transform 1 0 216904 0 1 53224
box 0 0 1 1
use contact_8  contact_8_263
timestamp 1624857261
transform 1 0 216904 0 1 53560
box 0 0 1 1
use contact_8  contact_8_262
timestamp 1624857261
transform 1 0 216904 0 1 53896
box 0 0 1 1
use contact_8  contact_8_261
timestamp 1624857261
transform 1 0 216904 0 1 54232
box 0 0 1 1
use contact_8  contact_8_260
timestamp 1624857261
transform 1 0 216904 0 1 54568
box 0 0 1 1
use contact_8  contact_8_259
timestamp 1624857261
transform 1 0 216904 0 1 54904
box 0 0 1 1
use contact_8  contact_8_258
timestamp 1624857261
transform 1 0 216904 0 1 55240
box 0 0 1 1
use contact_8  contact_8_257
timestamp 1624857261
transform 1 0 216904 0 1 55576
box 0 0 1 1
use contact_8  contact_8_256
timestamp 1624857261
transform 1 0 216904 0 1 55912
box 0 0 1 1
use contact_8  contact_8_255
timestamp 1624857261
transform 1 0 216904 0 1 56248
box 0 0 1 1
use contact_8  contact_8_254
timestamp 1624857261
transform 1 0 216904 0 1 56584
box 0 0 1 1
use contact_8  contact_8_253
timestamp 1624857261
transform 1 0 216904 0 1 56920
box 0 0 1 1
use contact_8  contact_8_252
timestamp 1624857261
transform 1 0 216904 0 1 57256
box 0 0 1 1
use contact_8  contact_8_251
timestamp 1624857261
transform 1 0 216904 0 1 57592
box 0 0 1 1
use contact_8  contact_8_250
timestamp 1624857261
transform 1 0 216904 0 1 57928
box 0 0 1 1
use contact_8  contact_8_249
timestamp 1624857261
transform 1 0 216904 0 1 58264
box 0 0 1 1
use contact_8  contact_8_248
timestamp 1624857261
transform 1 0 216904 0 1 58600
box 0 0 1 1
use contact_8  contact_8_247
timestamp 1624857261
transform 1 0 216904 0 1 58936
box 0 0 1 1
use contact_8  contact_8_246
timestamp 1624857261
transform 1 0 216904 0 1 59272
box 0 0 1 1
use contact_8  contact_8_245
timestamp 1624857261
transform 1 0 216904 0 1 59608
box 0 0 1 1
use contact_8  contact_8_244
timestamp 1624857261
transform 1 0 216904 0 1 59944
box 0 0 1 1
use contact_8  contact_8_243
timestamp 1624857261
transform 1 0 216904 0 1 60280
box 0 0 1 1
use contact_8  contact_8_242
timestamp 1624857261
transform 1 0 216904 0 1 60616
box 0 0 1 1
use contact_8  contact_8_241
timestamp 1624857261
transform 1 0 216904 0 1 60952
box 0 0 1 1
use contact_8  contact_8_240
timestamp 1624857261
transform 1 0 216904 0 1 61288
box 0 0 1 1
use contact_8  contact_8_239
timestamp 1624857261
transform 1 0 216904 0 1 61624
box 0 0 1 1
use contact_8  contact_8_238
timestamp 1624857261
transform 1 0 216904 0 1 61960
box 0 0 1 1
use contact_8  contact_8_237
timestamp 1624857261
transform 1 0 216904 0 1 62296
box 0 0 1 1
use contact_8  contact_8_236
timestamp 1624857261
transform 1 0 216904 0 1 62632
box 0 0 1 1
use contact_8  contact_8_235
timestamp 1624857261
transform 1 0 216904 0 1 62968
box 0 0 1 1
use contact_8  contact_8_234
timestamp 1624857261
transform 1 0 216904 0 1 63304
box 0 0 1 1
use contact_8  contact_8_233
timestamp 1624857261
transform 1 0 216904 0 1 63640
box 0 0 1 1
use contact_8  contact_8_232
timestamp 1624857261
transform 1 0 216904 0 1 63976
box 0 0 1 1
use contact_8  contact_8_231
timestamp 1624857261
transform 1 0 216904 0 1 64312
box 0 0 1 1
use contact_8  contact_8_230
timestamp 1624857261
transform 1 0 216904 0 1 64648
box 0 0 1 1
use contact_8  contact_8_229
timestamp 1624857261
transform 1 0 216904 0 1 64984
box 0 0 1 1
use contact_8  contact_8_228
timestamp 1624857261
transform 1 0 216904 0 1 65320
box 0 0 1 1
use contact_8  contact_8_227
timestamp 1624857261
transform 1 0 216904 0 1 65656
box 0 0 1 1
use contact_8  contact_8_226
timestamp 1624857261
transform 1 0 216904 0 1 65992
box 0 0 1 1
use contact_8  contact_8_225
timestamp 1624857261
transform 1 0 216904 0 1 66328
box 0 0 1 1
use contact_8  contact_8_224
timestamp 1624857261
transform 1 0 216904 0 1 66664
box 0 0 1 1
use contact_8  contact_8_223
timestamp 1624857261
transform 1 0 216904 0 1 67000
box 0 0 1 1
use contact_8  contact_8_222
timestamp 1624857261
transform 1 0 216904 0 1 67336
box 0 0 1 1
use contact_8  contact_8_221
timestamp 1624857261
transform 1 0 216904 0 1 67672
box 0 0 1 1
use contact_8  contact_8_220
timestamp 1624857261
transform 1 0 216904 0 1 68008
box 0 0 1 1
use contact_8  contact_8_219
timestamp 1624857261
transform 1 0 216904 0 1 68344
box 0 0 1 1
use contact_8  contact_8_218
timestamp 1624857261
transform 1 0 216904 0 1 68680
box 0 0 1 1
use contact_8  contact_8_217
timestamp 1624857261
transform 1 0 216904 0 1 69016
box 0 0 1 1
use contact_8  contact_8_216
timestamp 1624857261
transform 1 0 216904 0 1 69352
box 0 0 1 1
use contact_8  contact_8_215
timestamp 1624857261
transform 1 0 216904 0 1 69688
box 0 0 1 1
use contact_8  contact_8_214
timestamp 1624857261
transform 1 0 216904 0 1 70024
box 0 0 1 1
use contact_8  contact_8_213
timestamp 1624857261
transform 1 0 216904 0 1 70360
box 0 0 1 1
use contact_8  contact_8_212
timestamp 1624857261
transform 1 0 216904 0 1 70696
box 0 0 1 1
use contact_8  contact_8_211
timestamp 1624857261
transform 1 0 216904 0 1 71032
box 0 0 1 1
use contact_8  contact_8_210
timestamp 1624857261
transform 1 0 216904 0 1 71368
box 0 0 1 1
use contact_8  contact_8_209
timestamp 1624857261
transform 1 0 216904 0 1 71704
box 0 0 1 1
use contact_8  contact_8_208
timestamp 1624857261
transform 1 0 216904 0 1 72040
box 0 0 1 1
use contact_8  contact_8_207
timestamp 1624857261
transform 1 0 216904 0 1 72376
box 0 0 1 1
use contact_8  contact_8_206
timestamp 1624857261
transform 1 0 216904 0 1 72712
box 0 0 1 1
use contact_8  contact_8_205
timestamp 1624857261
transform 1 0 216904 0 1 73048
box 0 0 1 1
use contact_8  contact_8_204
timestamp 1624857261
transform 1 0 216904 0 1 73384
box 0 0 1 1
use contact_8  contact_8_203
timestamp 1624857261
transform 1 0 216904 0 1 73720
box 0 0 1 1
use contact_8  contact_8_202
timestamp 1624857261
transform 1 0 216904 0 1 74056
box 0 0 1 1
use contact_8  contact_8_201
timestamp 1624857261
transform 1 0 216904 0 1 74392
box 0 0 1 1
use contact_8  contact_8_200
timestamp 1624857261
transform 1 0 216904 0 1 74728
box 0 0 1 1
use contact_8  contact_8_199
timestamp 1624857261
transform 1 0 216904 0 1 75064
box 0 0 1 1
use contact_8  contact_8_198
timestamp 1624857261
transform 1 0 216904 0 1 75400
box 0 0 1 1
use contact_8  contact_8_197
timestamp 1624857261
transform 1 0 216904 0 1 75736
box 0 0 1 1
use contact_8  contact_8_196
timestamp 1624857261
transform 1 0 216904 0 1 76072
box 0 0 1 1
use contact_8  contact_8_195
timestamp 1624857261
transform 1 0 216904 0 1 76408
box 0 0 1 1
use contact_8  contact_8_194
timestamp 1624857261
transform 1 0 216904 0 1 76744
box 0 0 1 1
use contact_8  contact_8_193
timestamp 1624857261
transform 1 0 216904 0 1 77080
box 0 0 1 1
use contact_8  contact_8_192
timestamp 1624857261
transform 1 0 216904 0 1 77416
box 0 0 1 1
use contact_8  contact_8_191
timestamp 1624857261
transform 1 0 216904 0 1 77752
box 0 0 1 1
use contact_8  contact_8_190
timestamp 1624857261
transform 1 0 216904 0 1 78088
box 0 0 1 1
use contact_8  contact_8_189
timestamp 1624857261
transform 1 0 216904 0 1 78424
box 0 0 1 1
use contact_8  contact_8_188
timestamp 1624857261
transform 1 0 216904 0 1 78760
box 0 0 1 1
use contact_8  contact_8_187
timestamp 1624857261
transform 1 0 216904 0 1 79096
box 0 0 1 1
use contact_8  contact_8_186
timestamp 1624857261
transform 1 0 216904 0 1 79432
box 0 0 1 1
use contact_8  contact_8_185
timestamp 1624857261
transform 1 0 216904 0 1 79768
box 0 0 1 1
use contact_8  contact_8_184
timestamp 1624857261
transform 1 0 216904 0 1 80104
box 0 0 1 1
use contact_8  contact_8_183
timestamp 1624857261
transform 1 0 216904 0 1 80440
box 0 0 1 1
use contact_8  contact_8_182
timestamp 1624857261
transform 1 0 216904 0 1 80776
box 0 0 1 1
use contact_8  contact_8_181
timestamp 1624857261
transform 1 0 216904 0 1 81112
box 0 0 1 1
use contact_8  contact_8_180
timestamp 1624857261
transform 1 0 216904 0 1 81448
box 0 0 1 1
use contact_8  contact_8_179
timestamp 1624857261
transform 1 0 216904 0 1 81784
box 0 0 1 1
use contact_8  contact_8_178
timestamp 1624857261
transform 1 0 216904 0 1 82120
box 0 0 1 1
use contact_8  contact_8_177
timestamp 1624857261
transform 1 0 216904 0 1 82456
box 0 0 1 1
use contact_8  contact_8_176
timestamp 1624857261
transform 1 0 216904 0 1 82792
box 0 0 1 1
use contact_8  contact_8_175
timestamp 1624857261
transform 1 0 216904 0 1 83128
box 0 0 1 1
use contact_8  contact_8_174
timestamp 1624857261
transform 1 0 216904 0 1 83464
box 0 0 1 1
use contact_8  contact_8_173
timestamp 1624857261
transform 1 0 216904 0 1 83800
box 0 0 1 1
use contact_8  contact_8_172
timestamp 1624857261
transform 1 0 216904 0 1 84136
box 0 0 1 1
use contact_8  contact_8_171
timestamp 1624857261
transform 1 0 216904 0 1 84472
box 0 0 1 1
use contact_8  contact_8_170
timestamp 1624857261
transform 1 0 216904 0 1 84808
box 0 0 1 1
use contact_8  contact_8_169
timestamp 1624857261
transform 1 0 216904 0 1 85144
box 0 0 1 1
use contact_8  contact_8_168
timestamp 1624857261
transform 1 0 216904 0 1 85480
box 0 0 1 1
use contact_8  contact_8_167
timestamp 1624857261
transform 1 0 216904 0 1 85816
box 0 0 1 1
use contact_8  contact_8_166
timestamp 1624857261
transform 1 0 216904 0 1 86152
box 0 0 1 1
use contact_8  contact_8_165
timestamp 1624857261
transform 1 0 216904 0 1 86488
box 0 0 1 1
use contact_8  contact_8_164
timestamp 1624857261
transform 1 0 216904 0 1 86824
box 0 0 1 1
use contact_8  contact_8_163
timestamp 1624857261
transform 1 0 216904 0 1 87160
box 0 0 1 1
use contact_8  contact_8_162
timestamp 1624857261
transform 1 0 216904 0 1 87496
box 0 0 1 1
use contact_8  contact_8_161
timestamp 1624857261
transform 1 0 216904 0 1 87832
box 0 0 1 1
use contact_8  contact_8_160
timestamp 1624857261
transform 1 0 216904 0 1 88168
box 0 0 1 1
use contact_8  contact_8_159
timestamp 1624857261
transform 1 0 216904 0 1 88504
box 0 0 1 1
use contact_8  contact_8_158
timestamp 1624857261
transform 1 0 216904 0 1 88840
box 0 0 1 1
use contact_8  contact_8_157
timestamp 1624857261
transform 1 0 216904 0 1 89176
box 0 0 1 1
use contact_8  contact_8_156
timestamp 1624857261
transform 1 0 216904 0 1 89512
box 0 0 1 1
use contact_8  contact_8_155
timestamp 1624857261
transform 1 0 216904 0 1 89848
box 0 0 1 1
use contact_8  contact_8_154
timestamp 1624857261
transform 1 0 216904 0 1 90184
box 0 0 1 1
use contact_8  contact_8_153
timestamp 1624857261
transform 1 0 216904 0 1 90520
box 0 0 1 1
use contact_8  contact_8_152
timestamp 1624857261
transform 1 0 216904 0 1 90856
box 0 0 1 1
use contact_8  contact_8_151
timestamp 1624857261
transform 1 0 216904 0 1 91192
box 0 0 1 1
use contact_8  contact_8_150
timestamp 1624857261
transform 1 0 216904 0 1 91528
box 0 0 1 1
use contact_8  contact_8_149
timestamp 1624857261
transform 1 0 216904 0 1 91864
box 0 0 1 1
use contact_8  contact_8_148
timestamp 1624857261
transform 1 0 216904 0 1 92200
box 0 0 1 1
use contact_8  contact_8_147
timestamp 1624857261
transform 1 0 216904 0 1 92536
box 0 0 1 1
use contact_8  contact_8_146
timestamp 1624857261
transform 1 0 216904 0 1 92872
box 0 0 1 1
use contact_8  contact_8_145
timestamp 1624857261
transform 1 0 216904 0 1 93208
box 0 0 1 1
use contact_8  contact_8_144
timestamp 1624857261
transform 1 0 216904 0 1 93544
box 0 0 1 1
use contact_8  contact_8_143
timestamp 1624857261
transform 1 0 216904 0 1 93880
box 0 0 1 1
use contact_8  contact_8_142
timestamp 1624857261
transform 1 0 216904 0 1 94216
box 0 0 1 1
use contact_8  contact_8_141
timestamp 1624857261
transform 1 0 216904 0 1 94552
box 0 0 1 1
use contact_8  contact_8_140
timestamp 1624857261
transform 1 0 216904 0 1 94888
box 0 0 1 1
use contact_8  contact_8_139
timestamp 1624857261
transform 1 0 216904 0 1 95224
box 0 0 1 1
use contact_8  contact_8_138
timestamp 1624857261
transform 1 0 216904 0 1 95560
box 0 0 1 1
use contact_8  contact_8_137
timestamp 1624857261
transform 1 0 216904 0 1 95896
box 0 0 1 1
use contact_8  contact_8_136
timestamp 1624857261
transform 1 0 216904 0 1 96232
box 0 0 1 1
use contact_8  contact_8_135
timestamp 1624857261
transform 1 0 216904 0 1 96568
box 0 0 1 1
use contact_8  contact_8_134
timestamp 1624857261
transform 1 0 216904 0 1 96904
box 0 0 1 1
use contact_8  contact_8_133
timestamp 1624857261
transform 1 0 216904 0 1 97240
box 0 0 1 1
use contact_8  contact_8_132
timestamp 1624857261
transform 1 0 216904 0 1 97576
box 0 0 1 1
use contact_8  contact_8_131
timestamp 1624857261
transform 1 0 216904 0 1 97912
box 0 0 1 1
use contact_8  contact_8_130
timestamp 1624857261
transform 1 0 216904 0 1 98248
box 0 0 1 1
use contact_8  contact_8_129
timestamp 1624857261
transform 1 0 216904 0 1 98584
box 0 0 1 1
use contact_8  contact_8_128
timestamp 1624857261
transform 1 0 216904 0 1 98920
box 0 0 1 1
use contact_8  contact_8_127
timestamp 1624857261
transform 1 0 216904 0 1 99256
box 0 0 1 1
use contact_8  contact_8_126
timestamp 1624857261
transform 1 0 216904 0 1 99592
box 0 0 1 1
use contact_8  contact_8_125
timestamp 1624857261
transform 1 0 216904 0 1 99928
box 0 0 1 1
use contact_8  contact_8_124
timestamp 1624857261
transform 1 0 216904 0 1 100264
box 0 0 1 1
use contact_8  contact_8_123
timestamp 1624857261
transform 1 0 216904 0 1 100600
box 0 0 1 1
use contact_8  contact_8_122
timestamp 1624857261
transform 1 0 216904 0 1 100936
box 0 0 1 1
use contact_8  contact_8_121
timestamp 1624857261
transform 1 0 216904 0 1 101272
box 0 0 1 1
use contact_8  contact_8_120
timestamp 1624857261
transform 1 0 216904 0 1 101608
box 0 0 1 1
use contact_8  contact_8_119
timestamp 1624857261
transform 1 0 216904 0 1 101944
box 0 0 1 1
use contact_8  contact_8_118
timestamp 1624857261
transform 1 0 216904 0 1 102280
box 0 0 1 1
use contact_8  contact_8_117
timestamp 1624857261
transform 1 0 216904 0 1 102616
box 0 0 1 1
use contact_8  contact_8_116
timestamp 1624857261
transform 1 0 216904 0 1 102952
box 0 0 1 1
use contact_8  contact_8_115
timestamp 1624857261
transform 1 0 216904 0 1 103288
box 0 0 1 1
use contact_8  contact_8_114
timestamp 1624857261
transform 1 0 216904 0 1 103624
box 0 0 1 1
use contact_8  contact_8_113
timestamp 1624857261
transform 1 0 216904 0 1 103960
box 0 0 1 1
use contact_8  contact_8_112
timestamp 1624857261
transform 1 0 216904 0 1 104296
box 0 0 1 1
use contact_8  contact_8_111
timestamp 1624857261
transform 1 0 216904 0 1 104632
box 0 0 1 1
use contact_8  contact_8_110
timestamp 1624857261
transform 1 0 216904 0 1 104968
box 0 0 1 1
use contact_8  contact_8_109
timestamp 1624857261
transform 1 0 216904 0 1 105304
box 0 0 1 1
use contact_8  contact_8_108
timestamp 1624857261
transform 1 0 216904 0 1 105640
box 0 0 1 1
use contact_8  contact_8_107
timestamp 1624857261
transform 1 0 216904 0 1 105976
box 0 0 1 1
use contact_8  contact_8_106
timestamp 1624857261
transform 1 0 216904 0 1 106312
box 0 0 1 1
use contact_8  contact_8_105
timestamp 1624857261
transform 1 0 216904 0 1 106648
box 0 0 1 1
use contact_8  contact_8_104
timestamp 1624857261
transform 1 0 216904 0 1 106984
box 0 0 1 1
use contact_8  contact_8_103
timestamp 1624857261
transform 1 0 216904 0 1 107320
box 0 0 1 1
use contact_8  contact_8_102
timestamp 1624857261
transform 1 0 216904 0 1 107656
box 0 0 1 1
use contact_8  contact_8_101
timestamp 1624857261
transform 1 0 216904 0 1 107992
box 0 0 1 1
use contact_8  contact_8_100
timestamp 1624857261
transform 1 0 216904 0 1 108328
box 0 0 1 1
use contact_8  contact_8_99
timestamp 1624857261
transform 1 0 216904 0 1 108664
box 0 0 1 1
use contact_8  contact_8_98
timestamp 1624857261
transform 1 0 216904 0 1 109000
box 0 0 1 1
use contact_8  contact_8_97
timestamp 1624857261
transform 1 0 216904 0 1 109336
box 0 0 1 1
use contact_8  contact_8_96
timestamp 1624857261
transform 1 0 216904 0 1 109672
box 0 0 1 1
use contact_8  contact_8_95
timestamp 1624857261
transform 1 0 216904 0 1 110008
box 0 0 1 1
use contact_8  contact_8_94
timestamp 1624857261
transform 1 0 216904 0 1 110344
box 0 0 1 1
use contact_8  contact_8_93
timestamp 1624857261
transform 1 0 216904 0 1 110680
box 0 0 1 1
use contact_8  contact_8_92
timestamp 1624857261
transform 1 0 216904 0 1 111016
box 0 0 1 1
use contact_8  contact_8_91
timestamp 1624857261
transform 1 0 216904 0 1 111352
box 0 0 1 1
use contact_8  contact_8_90
timestamp 1624857261
transform 1 0 216904 0 1 111688
box 0 0 1 1
use contact_8  contact_8_89
timestamp 1624857261
transform 1 0 216904 0 1 112024
box 0 0 1 1
use contact_8  contact_8_88
timestamp 1624857261
transform 1 0 216904 0 1 112360
box 0 0 1 1
use contact_8  contact_8_87
timestamp 1624857261
transform 1 0 216904 0 1 112696
box 0 0 1 1
use contact_8  contact_8_86
timestamp 1624857261
transform 1 0 216904 0 1 113032
box 0 0 1 1
use contact_8  contact_8_85
timestamp 1624857261
transform 1 0 216904 0 1 113368
box 0 0 1 1
use contact_8  contact_8_84
timestamp 1624857261
transform 1 0 216904 0 1 113704
box 0 0 1 1
use contact_8  contact_8_83
timestamp 1624857261
transform 1 0 216904 0 1 114040
box 0 0 1 1
use contact_8  contact_8_82
timestamp 1624857261
transform 1 0 216904 0 1 114376
box 0 0 1 1
use contact_8  contact_8_81
timestamp 1624857261
transform 1 0 216904 0 1 114712
box 0 0 1 1
use contact_8  contact_8_80
timestamp 1624857261
transform 1 0 216904 0 1 115048
box 0 0 1 1
use contact_8  contact_8_79
timestamp 1624857261
transform 1 0 216904 0 1 115384
box 0 0 1 1
use contact_8  contact_8_78
timestamp 1624857261
transform 1 0 216904 0 1 115720
box 0 0 1 1
use contact_8  contact_8_77
timestamp 1624857261
transform 1 0 216904 0 1 116056
box 0 0 1 1
use contact_8  contact_8_76
timestamp 1624857261
transform 1 0 216904 0 1 116392
box 0 0 1 1
use contact_8  contact_8_75
timestamp 1624857261
transform 1 0 216904 0 1 116728
box 0 0 1 1
use contact_8  contact_8_74
timestamp 1624857261
transform 1 0 216904 0 1 117064
box 0 0 1 1
use contact_8  contact_8_73
timestamp 1624857261
transform 1 0 216904 0 1 117400
box 0 0 1 1
use contact_8  contact_8_72
timestamp 1624857261
transform 1 0 216904 0 1 117736
box 0 0 1 1
use contact_8  contact_8_71
timestamp 1624857261
transform 1 0 216904 0 1 118072
box 0 0 1 1
use contact_8  contact_8_70
timestamp 1624857261
transform 1 0 216904 0 1 118408
box 0 0 1 1
use contact_8  contact_8_69
timestamp 1624857261
transform 1 0 216904 0 1 118744
box 0 0 1 1
use contact_8  contact_8_68
timestamp 1624857261
transform 1 0 216904 0 1 119080
box 0 0 1 1
use contact_8  contact_8_67
timestamp 1624857261
transform 1 0 216904 0 1 119416
box 0 0 1 1
use contact_8  contact_8_66
timestamp 1624857261
transform 1 0 216904 0 1 119752
box 0 0 1 1
use contact_8  contact_8_65
timestamp 1624857261
transform 1 0 216904 0 1 120088
box 0 0 1 1
use contact_8  contact_8_64
timestamp 1624857261
transform 1 0 216904 0 1 120424
box 0 0 1 1
use contact_8  contact_8_63
timestamp 1624857261
transform 1 0 216904 0 1 120760
box 0 0 1 1
use contact_8  contact_8_62
timestamp 1624857261
transform 1 0 216904 0 1 121096
box 0 0 1 1
use contact_8  contact_8_61
timestamp 1624857261
transform 1 0 216904 0 1 121432
box 0 0 1 1
use contact_8  contact_8_60
timestamp 1624857261
transform 1 0 216904 0 1 121768
box 0 0 1 1
use contact_8  contact_8_59
timestamp 1624857261
transform 1 0 216904 0 1 122104
box 0 0 1 1
use contact_8  contact_8_58
timestamp 1624857261
transform 1 0 216904 0 1 122440
box 0 0 1 1
use contact_8  contact_8_57
timestamp 1624857261
transform 1 0 216904 0 1 122776
box 0 0 1 1
use contact_8  contact_8_56
timestamp 1624857261
transform 1 0 216904 0 1 123112
box 0 0 1 1
use contact_8  contact_8_55
timestamp 1624857261
transform 1 0 216904 0 1 123448
box 0 0 1 1
use contact_8  contact_8_54
timestamp 1624857261
transform 1 0 216904 0 1 123784
box 0 0 1 1
use contact_8  contact_8_53
timestamp 1624857261
transform 1 0 216904 0 1 124120
box 0 0 1 1
use contact_8  contact_8_52
timestamp 1624857261
transform 1 0 216904 0 1 124456
box 0 0 1 1
use contact_8  contact_8_51
timestamp 1624857261
transform 1 0 216904 0 1 124792
box 0 0 1 1
use contact_8  contact_8_50
timestamp 1624857261
transform 1 0 216904 0 1 125128
box 0 0 1 1
use contact_8  contact_8_49
timestamp 1624857261
transform 1 0 216904 0 1 125464
box 0 0 1 1
use contact_8  contact_8_48
timestamp 1624857261
transform 1 0 216904 0 1 125800
box 0 0 1 1
use contact_8  contact_8_47
timestamp 1624857261
transform 1 0 216904 0 1 126136
box 0 0 1 1
use contact_8  contact_8_46
timestamp 1624857261
transform 1 0 216904 0 1 126472
box 0 0 1 1
use contact_8  contact_8_45
timestamp 1624857261
transform 1 0 216904 0 1 126808
box 0 0 1 1
use contact_8  contact_8_44
timestamp 1624857261
transform 1 0 216904 0 1 127144
box 0 0 1 1
use contact_8  contact_8_43
timestamp 1624857261
transform 1 0 216904 0 1 127480
box 0 0 1 1
use contact_8  contact_8_42
timestamp 1624857261
transform 1 0 216904 0 1 127816
box 0 0 1 1
use contact_8  contact_8_41
timestamp 1624857261
transform 1 0 216904 0 1 128152
box 0 0 1 1
use contact_8  contact_8_40
timestamp 1624857261
transform 1 0 216904 0 1 128488
box 0 0 1 1
use contact_8  contact_8_39
timestamp 1624857261
transform 1 0 216904 0 1 128824
box 0 0 1 1
use contact_8  contact_8_38
timestamp 1624857261
transform 1 0 216904 0 1 129160
box 0 0 1 1
use contact_8  contact_8_37
timestamp 1624857261
transform 1 0 216904 0 1 129496
box 0 0 1 1
use contact_8  contact_8_36
timestamp 1624857261
transform 1 0 216904 0 1 129832
box 0 0 1 1
use contact_8  contact_8_35
timestamp 1624857261
transform 1 0 216904 0 1 130168
box 0 0 1 1
use contact_8  contact_8_34
timestamp 1624857261
transform 1 0 216904 0 1 130504
box 0 0 1 1
use contact_8  contact_8_33
timestamp 1624857261
transform 1 0 216904 0 1 130840
box 0 0 1 1
use contact_8  contact_8_32
timestamp 1624857261
transform 1 0 216904 0 1 131176
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1624857261
transform 1 0 216904 0 1 131512
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1624857261
transform 1 0 216904 0 1 131848
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1624857261
transform 1 0 216904 0 1 132184
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1624857261
transform 1 0 216904 0 1 132520
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1624857261
transform 1 0 216904 0 1 132856
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1624857261
transform 1 0 216904 0 1 133192
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1624857261
transform 1 0 216904 0 1 133528
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1624857261
transform 1 0 216904 0 1 133864
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1624857261
transform 1 0 216904 0 1 134200
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1624857261
transform 1 0 216904 0 1 134536
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1624857261
transform 1 0 216904 0 1 134872
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1624857261
transform 1 0 216904 0 1 135208
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1624857261
transform 1 0 216904 0 1 135544
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1624857261
transform 1 0 216904 0 1 135880
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1624857261
transform 1 0 216904 0 1 136216
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1624857261
transform 1 0 216904 0 1 136552
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1624857261
transform 1 0 216904 0 1 136888
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1624857261
transform 1 0 216904 0 1 137224
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1624857261
transform 1 0 216904 0 1 137560
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1624857261
transform 1 0 216904 0 1 137896
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1624857261
transform 1 0 216904 0 1 138232
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1624857261
transform 1 0 216904 0 1 138568
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1624857261
transform 1 0 216904 0 1 138904
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1624857261
transform 1 0 216904 0 1 139240
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1624857261
transform 1 0 216904 0 1 139576
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1624857261
transform 1 0 216904 0 1 139912
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1624857261
transform 1 0 216904 0 1 140248
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1624857261
transform 1 0 216904 0 1 140584
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1624857261
transform 1 0 216904 0 1 140920
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1624857261
transform 1 0 216904 0 1 141256
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1624857261
transform 1 0 216904 0 1 141592
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1624857261
transform 1 0 216904 0 1 141928
box 0 0 1 1
use contact_7  contact_7_2111
timestamp 1624857261
transform 1 0 2037 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2110
timestamp 1624857261
transform 1 0 2373 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2109
timestamp 1624857261
transform 1 0 2709 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2108
timestamp 1624857261
transform 1 0 3045 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2107
timestamp 1624857261
transform 1 0 3381 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2106
timestamp 1624857261
transform 1 0 3717 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2105
timestamp 1624857261
transform 1 0 4053 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2104
timestamp 1624857261
transform 1 0 4389 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2103
timestamp 1624857261
transform 1 0 4725 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2102
timestamp 1624857261
transform 1 0 5061 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2101
timestamp 1624857261
transform 1 0 5397 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2100
timestamp 1624857261
transform 1 0 5733 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2099
timestamp 1624857261
transform 1 0 6069 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2098
timestamp 1624857261
transform 1 0 6405 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2097
timestamp 1624857261
transform 1 0 6741 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2096
timestamp 1624857261
transform 1 0 7077 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2095
timestamp 1624857261
transform 1 0 7413 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2094
timestamp 1624857261
transform 1 0 7749 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2093
timestamp 1624857261
transform 1 0 8085 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2092
timestamp 1624857261
transform 1 0 8421 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2091
timestamp 1624857261
transform 1 0 8757 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2090
timestamp 1624857261
transform 1 0 9093 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2089
timestamp 1624857261
transform 1 0 9429 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2088
timestamp 1624857261
transform 1 0 9765 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2087
timestamp 1624857261
transform 1 0 10101 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2086
timestamp 1624857261
transform 1 0 10437 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2085
timestamp 1624857261
transform 1 0 10773 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2084
timestamp 1624857261
transform 1 0 11109 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2083
timestamp 1624857261
transform 1 0 11445 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2082
timestamp 1624857261
transform 1 0 11781 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2081
timestamp 1624857261
transform 1 0 12117 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2080
timestamp 1624857261
transform 1 0 12453 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2079
timestamp 1624857261
transform 1 0 12789 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2078
timestamp 1624857261
transform 1 0 13125 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2077
timestamp 1624857261
transform 1 0 13461 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2076
timestamp 1624857261
transform 1 0 13797 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2075
timestamp 1624857261
transform 1 0 14133 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2074
timestamp 1624857261
transform 1 0 14469 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2073
timestamp 1624857261
transform 1 0 14805 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2072
timestamp 1624857261
transform 1 0 15141 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2071
timestamp 1624857261
transform 1 0 15477 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2070
timestamp 1624857261
transform 1 0 15813 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2069
timestamp 1624857261
transform 1 0 16149 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2068
timestamp 1624857261
transform 1 0 16485 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2067
timestamp 1624857261
transform 1 0 16821 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2066
timestamp 1624857261
transform 1 0 17157 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2065
timestamp 1624857261
transform 1 0 17493 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2064
timestamp 1624857261
transform 1 0 17829 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2063
timestamp 1624857261
transform 1 0 18165 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2062
timestamp 1624857261
transform 1 0 18501 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2061
timestamp 1624857261
transform 1 0 18837 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2060
timestamp 1624857261
transform 1 0 19173 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2059
timestamp 1624857261
transform 1 0 19509 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2058
timestamp 1624857261
transform 1 0 19845 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2057
timestamp 1624857261
transform 1 0 20181 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2056
timestamp 1624857261
transform 1 0 20517 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2055
timestamp 1624857261
transform 1 0 20853 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2054
timestamp 1624857261
transform 1 0 21189 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2053
timestamp 1624857261
transform 1 0 21525 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2052
timestamp 1624857261
transform 1 0 21861 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2051
timestamp 1624857261
transform 1 0 22197 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2050
timestamp 1624857261
transform 1 0 22533 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2049
timestamp 1624857261
transform 1 0 22869 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2048
timestamp 1624857261
transform 1 0 23205 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2047
timestamp 1624857261
transform 1 0 23541 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2046
timestamp 1624857261
transform 1 0 23877 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2045
timestamp 1624857261
transform 1 0 24213 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2044
timestamp 1624857261
transform 1 0 24549 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2043
timestamp 1624857261
transform 1 0 24885 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2042
timestamp 1624857261
transform 1 0 25221 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2041
timestamp 1624857261
transform 1 0 25557 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2040
timestamp 1624857261
transform 1 0 25893 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2039
timestamp 1624857261
transform 1 0 26229 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2038
timestamp 1624857261
transform 1 0 26565 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2037
timestamp 1624857261
transform 1 0 26901 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2036
timestamp 1624857261
transform 1 0 27237 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2035
timestamp 1624857261
transform 1 0 27573 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2034
timestamp 1624857261
transform 1 0 27909 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2033
timestamp 1624857261
transform 1 0 28245 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2032
timestamp 1624857261
transform 1 0 28581 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2031
timestamp 1624857261
transform 1 0 28917 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2030
timestamp 1624857261
transform 1 0 29253 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2029
timestamp 1624857261
transform 1 0 29589 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2028
timestamp 1624857261
transform 1 0 29925 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2027
timestamp 1624857261
transform 1 0 30261 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2026
timestamp 1624857261
transform 1 0 30597 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2025
timestamp 1624857261
transform 1 0 30933 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2024
timestamp 1624857261
transform 1 0 31269 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2023
timestamp 1624857261
transform 1 0 31605 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2022
timestamp 1624857261
transform 1 0 31941 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2021
timestamp 1624857261
transform 1 0 32277 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2020
timestamp 1624857261
transform 1 0 32613 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2019
timestamp 1624857261
transform 1 0 32949 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2018
timestamp 1624857261
transform 1 0 33285 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2017
timestamp 1624857261
transform 1 0 33621 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2016
timestamp 1624857261
transform 1 0 33957 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2015
timestamp 1624857261
transform 1 0 34293 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2014
timestamp 1624857261
transform 1 0 34629 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2013
timestamp 1624857261
transform 1 0 34965 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2012
timestamp 1624857261
transform 1 0 35301 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2011
timestamp 1624857261
transform 1 0 35637 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2010
timestamp 1624857261
transform 1 0 35973 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2009
timestamp 1624857261
transform 1 0 36309 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2008
timestamp 1624857261
transform 1 0 36645 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2007
timestamp 1624857261
transform 1 0 36981 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2006
timestamp 1624857261
transform 1 0 37317 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2005
timestamp 1624857261
transform 1 0 37653 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2004
timestamp 1624857261
transform 1 0 37989 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2003
timestamp 1624857261
transform 1 0 38325 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2002
timestamp 1624857261
transform 1 0 38661 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2001
timestamp 1624857261
transform 1 0 38997 0 1 1815
box 0 0 1 1
use contact_7  contact_7_2000
timestamp 1624857261
transform 1 0 39333 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1999
timestamp 1624857261
transform 1 0 39669 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1998
timestamp 1624857261
transform 1 0 40005 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1997
timestamp 1624857261
transform 1 0 40341 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1996
timestamp 1624857261
transform 1 0 40677 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1995
timestamp 1624857261
transform 1 0 41013 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1994
timestamp 1624857261
transform 1 0 41349 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1993
timestamp 1624857261
transform 1 0 41685 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1992
timestamp 1624857261
transform 1 0 42021 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1991
timestamp 1624857261
transform 1 0 42357 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1990
timestamp 1624857261
transform 1 0 42693 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1989
timestamp 1624857261
transform 1 0 43029 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1988
timestamp 1624857261
transform 1 0 43365 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1987
timestamp 1624857261
transform 1 0 43701 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1986
timestamp 1624857261
transform 1 0 44037 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1985
timestamp 1624857261
transform 1 0 44373 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1984
timestamp 1624857261
transform 1 0 44709 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1983
timestamp 1624857261
transform 1 0 45045 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1982
timestamp 1624857261
transform 1 0 45381 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1981
timestamp 1624857261
transform 1 0 45717 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1980
timestamp 1624857261
transform 1 0 46053 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1979
timestamp 1624857261
transform 1 0 46389 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1978
timestamp 1624857261
transform 1 0 46725 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1977
timestamp 1624857261
transform 1 0 47061 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1976
timestamp 1624857261
transform 1 0 47397 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1975
timestamp 1624857261
transform 1 0 47733 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1974
timestamp 1624857261
transform 1 0 48069 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1973
timestamp 1624857261
transform 1 0 48405 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1972
timestamp 1624857261
transform 1 0 48741 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1971
timestamp 1624857261
transform 1 0 49077 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1970
timestamp 1624857261
transform 1 0 49413 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1969
timestamp 1624857261
transform 1 0 49749 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1968
timestamp 1624857261
transform 1 0 50085 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1967
timestamp 1624857261
transform 1 0 50421 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1966
timestamp 1624857261
transform 1 0 50757 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1965
timestamp 1624857261
transform 1 0 51093 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1964
timestamp 1624857261
transform 1 0 51429 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1963
timestamp 1624857261
transform 1 0 51765 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1962
timestamp 1624857261
transform 1 0 52101 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1961
timestamp 1624857261
transform 1 0 52437 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1960
timestamp 1624857261
transform 1 0 52773 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1959
timestamp 1624857261
transform 1 0 53109 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1958
timestamp 1624857261
transform 1 0 53445 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1957
timestamp 1624857261
transform 1 0 53781 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1956
timestamp 1624857261
transform 1 0 54117 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1955
timestamp 1624857261
transform 1 0 54453 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1954
timestamp 1624857261
transform 1 0 54789 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1953
timestamp 1624857261
transform 1 0 55125 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1952
timestamp 1624857261
transform 1 0 55461 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1951
timestamp 1624857261
transform 1 0 55797 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1950
timestamp 1624857261
transform 1 0 56133 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1949
timestamp 1624857261
transform 1 0 56469 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1948
timestamp 1624857261
transform 1 0 56805 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1947
timestamp 1624857261
transform 1 0 57141 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1946
timestamp 1624857261
transform 1 0 57477 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1945
timestamp 1624857261
transform 1 0 57813 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1944
timestamp 1624857261
transform 1 0 58149 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1943
timestamp 1624857261
transform 1 0 58485 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1942
timestamp 1624857261
transform 1 0 58821 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1941
timestamp 1624857261
transform 1 0 59157 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1940
timestamp 1624857261
transform 1 0 59493 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1939
timestamp 1624857261
transform 1 0 59829 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1938
timestamp 1624857261
transform 1 0 60165 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1937
timestamp 1624857261
transform 1 0 60501 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1936
timestamp 1624857261
transform 1 0 60837 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1935
timestamp 1624857261
transform 1 0 61173 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1934
timestamp 1624857261
transform 1 0 61509 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1933
timestamp 1624857261
transform 1 0 61845 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1932
timestamp 1624857261
transform 1 0 62181 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1931
timestamp 1624857261
transform 1 0 62517 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1930
timestamp 1624857261
transform 1 0 62853 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1929
timestamp 1624857261
transform 1 0 63189 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1928
timestamp 1624857261
transform 1 0 63525 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1927
timestamp 1624857261
transform 1 0 63861 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1926
timestamp 1624857261
transform 1 0 64197 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1925
timestamp 1624857261
transform 1 0 64533 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1924
timestamp 1624857261
transform 1 0 64869 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1923
timestamp 1624857261
transform 1 0 65205 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1922
timestamp 1624857261
transform 1 0 65541 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1921
timestamp 1624857261
transform 1 0 65877 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1920
timestamp 1624857261
transform 1 0 66213 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1919
timestamp 1624857261
transform 1 0 66549 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1918
timestamp 1624857261
transform 1 0 66885 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1917
timestamp 1624857261
transform 1 0 67221 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1916
timestamp 1624857261
transform 1 0 67557 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1915
timestamp 1624857261
transform 1 0 67893 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1914
timestamp 1624857261
transform 1 0 68229 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1913
timestamp 1624857261
transform 1 0 68565 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1912
timestamp 1624857261
transform 1 0 68901 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1911
timestamp 1624857261
transform 1 0 69237 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1910
timestamp 1624857261
transform 1 0 69573 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1909
timestamp 1624857261
transform 1 0 69909 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1908
timestamp 1624857261
transform 1 0 70245 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1907
timestamp 1624857261
transform 1 0 70581 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1906
timestamp 1624857261
transform 1 0 70917 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1905
timestamp 1624857261
transform 1 0 71253 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1904
timestamp 1624857261
transform 1 0 71589 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1903
timestamp 1624857261
transform 1 0 71925 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1902
timestamp 1624857261
transform 1 0 72261 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1901
timestamp 1624857261
transform 1 0 72597 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1900
timestamp 1624857261
transform 1 0 72933 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1899
timestamp 1624857261
transform 1 0 73269 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1898
timestamp 1624857261
transform 1 0 73605 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1897
timestamp 1624857261
transform 1 0 73941 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1896
timestamp 1624857261
transform 1 0 74277 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1895
timestamp 1624857261
transform 1 0 74613 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1894
timestamp 1624857261
transform 1 0 74949 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1893
timestamp 1624857261
transform 1 0 75285 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1892
timestamp 1624857261
transform 1 0 75621 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1891
timestamp 1624857261
transform 1 0 75957 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1890
timestamp 1624857261
transform 1 0 76293 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1889
timestamp 1624857261
transform 1 0 76629 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1888
timestamp 1624857261
transform 1 0 76965 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1887
timestamp 1624857261
transform 1 0 77301 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1886
timestamp 1624857261
transform 1 0 77637 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1885
timestamp 1624857261
transform 1 0 77973 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1884
timestamp 1624857261
transform 1 0 78309 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1883
timestamp 1624857261
transform 1 0 78645 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1882
timestamp 1624857261
transform 1 0 78981 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1881
timestamp 1624857261
transform 1 0 79317 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1880
timestamp 1624857261
transform 1 0 79653 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1879
timestamp 1624857261
transform 1 0 79989 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1878
timestamp 1624857261
transform 1 0 80325 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1877
timestamp 1624857261
transform 1 0 80661 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1876
timestamp 1624857261
transform 1 0 80997 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1875
timestamp 1624857261
transform 1 0 81333 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1874
timestamp 1624857261
transform 1 0 81669 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1873
timestamp 1624857261
transform 1 0 82005 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1872
timestamp 1624857261
transform 1 0 82341 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1871
timestamp 1624857261
transform 1 0 82677 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1870
timestamp 1624857261
transform 1 0 83013 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1869
timestamp 1624857261
transform 1 0 83349 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1868
timestamp 1624857261
transform 1 0 83685 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1867
timestamp 1624857261
transform 1 0 84021 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1866
timestamp 1624857261
transform 1 0 84357 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1865
timestamp 1624857261
transform 1 0 84693 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1864
timestamp 1624857261
transform 1 0 85029 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1863
timestamp 1624857261
transform 1 0 85365 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1862
timestamp 1624857261
transform 1 0 85701 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1861
timestamp 1624857261
transform 1 0 86037 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1860
timestamp 1624857261
transform 1 0 86373 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1859
timestamp 1624857261
transform 1 0 86709 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1858
timestamp 1624857261
transform 1 0 87045 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1857
timestamp 1624857261
transform 1 0 87381 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1856
timestamp 1624857261
transform 1 0 87717 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1855
timestamp 1624857261
transform 1 0 88053 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1854
timestamp 1624857261
transform 1 0 88389 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1853
timestamp 1624857261
transform 1 0 88725 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1852
timestamp 1624857261
transform 1 0 89061 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1851
timestamp 1624857261
transform 1 0 89397 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1850
timestamp 1624857261
transform 1 0 89733 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1849
timestamp 1624857261
transform 1 0 90069 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1848
timestamp 1624857261
transform 1 0 90405 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1847
timestamp 1624857261
transform 1 0 90741 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1846
timestamp 1624857261
transform 1 0 91077 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1845
timestamp 1624857261
transform 1 0 91413 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1844
timestamp 1624857261
transform 1 0 91749 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1843
timestamp 1624857261
transform 1 0 92085 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1842
timestamp 1624857261
transform 1 0 92421 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1841
timestamp 1624857261
transform 1 0 92757 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1840
timestamp 1624857261
transform 1 0 93093 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1839
timestamp 1624857261
transform 1 0 93429 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1838
timestamp 1624857261
transform 1 0 93765 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1837
timestamp 1624857261
transform 1 0 94101 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1836
timestamp 1624857261
transform 1 0 94437 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1835
timestamp 1624857261
transform 1 0 94773 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1834
timestamp 1624857261
transform 1 0 95109 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1833
timestamp 1624857261
transform 1 0 95445 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1832
timestamp 1624857261
transform 1 0 95781 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1831
timestamp 1624857261
transform 1 0 96117 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1830
timestamp 1624857261
transform 1 0 96453 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1829
timestamp 1624857261
transform 1 0 96789 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1828
timestamp 1624857261
transform 1 0 97125 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1827
timestamp 1624857261
transform 1 0 97461 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1826
timestamp 1624857261
transform 1 0 97797 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1825
timestamp 1624857261
transform 1 0 98133 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1824
timestamp 1624857261
transform 1 0 98469 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1823
timestamp 1624857261
transform 1 0 98805 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1822
timestamp 1624857261
transform 1 0 99141 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1821
timestamp 1624857261
transform 1 0 99477 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1820
timestamp 1624857261
transform 1 0 99813 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1819
timestamp 1624857261
transform 1 0 100149 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1818
timestamp 1624857261
transform 1 0 100485 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1817
timestamp 1624857261
transform 1 0 100821 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1816
timestamp 1624857261
transform 1 0 101157 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1815
timestamp 1624857261
transform 1 0 101493 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1814
timestamp 1624857261
transform 1 0 101829 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1813
timestamp 1624857261
transform 1 0 102165 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1812
timestamp 1624857261
transform 1 0 102501 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1811
timestamp 1624857261
transform 1 0 102837 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1810
timestamp 1624857261
transform 1 0 103173 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1809
timestamp 1624857261
transform 1 0 103509 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1808
timestamp 1624857261
transform 1 0 103845 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1807
timestamp 1624857261
transform 1 0 104181 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1806
timestamp 1624857261
transform 1 0 104517 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1805
timestamp 1624857261
transform 1 0 104853 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1804
timestamp 1624857261
transform 1 0 105189 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1803
timestamp 1624857261
transform 1 0 105525 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1802
timestamp 1624857261
transform 1 0 105861 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1801
timestamp 1624857261
transform 1 0 106197 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1800
timestamp 1624857261
transform 1 0 106533 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1799
timestamp 1624857261
transform 1 0 106869 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1798
timestamp 1624857261
transform 1 0 107205 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1797
timestamp 1624857261
transform 1 0 107541 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1796
timestamp 1624857261
transform 1 0 107877 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1795
timestamp 1624857261
transform 1 0 108213 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1794
timestamp 1624857261
transform 1 0 108549 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1793
timestamp 1624857261
transform 1 0 108885 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1792
timestamp 1624857261
transform 1 0 109221 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1791
timestamp 1624857261
transform 1 0 109557 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1790
timestamp 1624857261
transform 1 0 109893 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1789
timestamp 1624857261
transform 1 0 110229 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1788
timestamp 1624857261
transform 1 0 110565 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1787
timestamp 1624857261
transform 1 0 110901 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1786
timestamp 1624857261
transform 1 0 111237 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1785
timestamp 1624857261
transform 1 0 111573 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1784
timestamp 1624857261
transform 1 0 111909 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1783
timestamp 1624857261
transform 1 0 112245 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1782
timestamp 1624857261
transform 1 0 112581 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1781
timestamp 1624857261
transform 1 0 112917 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1780
timestamp 1624857261
transform 1 0 113253 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1779
timestamp 1624857261
transform 1 0 113589 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1778
timestamp 1624857261
transform 1 0 113925 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1777
timestamp 1624857261
transform 1 0 114261 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1776
timestamp 1624857261
transform 1 0 114597 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1775
timestamp 1624857261
transform 1 0 114933 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1774
timestamp 1624857261
transform 1 0 115269 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1773
timestamp 1624857261
transform 1 0 115605 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1772
timestamp 1624857261
transform 1 0 115941 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1771
timestamp 1624857261
transform 1 0 116277 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1770
timestamp 1624857261
transform 1 0 116613 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1769
timestamp 1624857261
transform 1 0 116949 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1768
timestamp 1624857261
transform 1 0 117285 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1767
timestamp 1624857261
transform 1 0 117621 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1766
timestamp 1624857261
transform 1 0 117957 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1765
timestamp 1624857261
transform 1 0 118293 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1764
timestamp 1624857261
transform 1 0 118629 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1763
timestamp 1624857261
transform 1 0 118965 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1762
timestamp 1624857261
transform 1 0 119301 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1761
timestamp 1624857261
transform 1 0 119637 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1760
timestamp 1624857261
transform 1 0 119973 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1759
timestamp 1624857261
transform 1 0 120309 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1758
timestamp 1624857261
transform 1 0 120645 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1757
timestamp 1624857261
transform 1 0 120981 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1756
timestamp 1624857261
transform 1 0 121317 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1755
timestamp 1624857261
transform 1 0 121653 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1754
timestamp 1624857261
transform 1 0 121989 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1753
timestamp 1624857261
transform 1 0 122325 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1752
timestamp 1624857261
transform 1 0 122661 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1751
timestamp 1624857261
transform 1 0 122997 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1750
timestamp 1624857261
transform 1 0 123333 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1749
timestamp 1624857261
transform 1 0 123669 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1748
timestamp 1624857261
transform 1 0 124005 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1747
timestamp 1624857261
transform 1 0 124341 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1746
timestamp 1624857261
transform 1 0 124677 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1745
timestamp 1624857261
transform 1 0 125013 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1744
timestamp 1624857261
transform 1 0 125349 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1743
timestamp 1624857261
transform 1 0 125685 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1742
timestamp 1624857261
transform 1 0 126021 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1741
timestamp 1624857261
transform 1 0 126357 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1740
timestamp 1624857261
transform 1 0 126693 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1739
timestamp 1624857261
transform 1 0 127029 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1738
timestamp 1624857261
transform 1 0 127365 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1737
timestamp 1624857261
transform 1 0 127701 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1736
timestamp 1624857261
transform 1 0 128037 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1735
timestamp 1624857261
transform 1 0 128373 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1734
timestamp 1624857261
transform 1 0 128709 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1733
timestamp 1624857261
transform 1 0 129045 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1732
timestamp 1624857261
transform 1 0 129381 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1731
timestamp 1624857261
transform 1 0 129717 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1730
timestamp 1624857261
transform 1 0 130053 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1729
timestamp 1624857261
transform 1 0 130389 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1728
timestamp 1624857261
transform 1 0 130725 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1727
timestamp 1624857261
transform 1 0 131061 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1726
timestamp 1624857261
transform 1 0 131397 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1725
timestamp 1624857261
transform 1 0 131733 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1724
timestamp 1624857261
transform 1 0 132069 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1723
timestamp 1624857261
transform 1 0 132405 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1722
timestamp 1624857261
transform 1 0 132741 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1721
timestamp 1624857261
transform 1 0 133077 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1720
timestamp 1624857261
transform 1 0 133413 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1719
timestamp 1624857261
transform 1 0 133749 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1718
timestamp 1624857261
transform 1 0 134085 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1717
timestamp 1624857261
transform 1 0 134421 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1716
timestamp 1624857261
transform 1 0 134757 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1715
timestamp 1624857261
transform 1 0 135093 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1714
timestamp 1624857261
transform 1 0 135429 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1713
timestamp 1624857261
transform 1 0 135765 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1712
timestamp 1624857261
transform 1 0 136101 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1711
timestamp 1624857261
transform 1 0 136437 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1710
timestamp 1624857261
transform 1 0 136773 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1709
timestamp 1624857261
transform 1 0 137109 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1708
timestamp 1624857261
transform 1 0 137445 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1707
timestamp 1624857261
transform 1 0 137781 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1706
timestamp 1624857261
transform 1 0 138117 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1705
timestamp 1624857261
transform 1 0 138453 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1704
timestamp 1624857261
transform 1 0 138789 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1703
timestamp 1624857261
transform 1 0 139125 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1702
timestamp 1624857261
transform 1 0 139461 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1701
timestamp 1624857261
transform 1 0 139797 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1700
timestamp 1624857261
transform 1 0 140133 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1699
timestamp 1624857261
transform 1 0 140469 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1698
timestamp 1624857261
transform 1 0 140805 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1697
timestamp 1624857261
transform 1 0 141141 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1696
timestamp 1624857261
transform 1 0 141477 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1695
timestamp 1624857261
transform 1 0 141813 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1694
timestamp 1624857261
transform 1 0 142149 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1693
timestamp 1624857261
transform 1 0 142485 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1692
timestamp 1624857261
transform 1 0 142821 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1691
timestamp 1624857261
transform 1 0 143157 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1690
timestamp 1624857261
transform 1 0 143493 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1689
timestamp 1624857261
transform 1 0 143829 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1688
timestamp 1624857261
transform 1 0 144165 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1687
timestamp 1624857261
transform 1 0 144501 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1686
timestamp 1624857261
transform 1 0 144837 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1685
timestamp 1624857261
transform 1 0 145173 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1684
timestamp 1624857261
transform 1 0 145509 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1683
timestamp 1624857261
transform 1 0 145845 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1682
timestamp 1624857261
transform 1 0 146181 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1681
timestamp 1624857261
transform 1 0 146517 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1680
timestamp 1624857261
transform 1 0 146853 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1679
timestamp 1624857261
transform 1 0 147189 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1678
timestamp 1624857261
transform 1 0 147525 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1677
timestamp 1624857261
transform 1 0 147861 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1676
timestamp 1624857261
transform 1 0 148197 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1675
timestamp 1624857261
transform 1 0 148533 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1674
timestamp 1624857261
transform 1 0 148869 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1673
timestamp 1624857261
transform 1 0 149205 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1672
timestamp 1624857261
transform 1 0 149541 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1671
timestamp 1624857261
transform 1 0 149877 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1670
timestamp 1624857261
transform 1 0 150213 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1669
timestamp 1624857261
transform 1 0 150549 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1668
timestamp 1624857261
transform 1 0 150885 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1667
timestamp 1624857261
transform 1 0 151221 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1666
timestamp 1624857261
transform 1 0 151557 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1665
timestamp 1624857261
transform 1 0 151893 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1664
timestamp 1624857261
transform 1 0 152229 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1663
timestamp 1624857261
transform 1 0 152565 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1662
timestamp 1624857261
transform 1 0 152901 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1661
timestamp 1624857261
transform 1 0 153237 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1660
timestamp 1624857261
transform 1 0 153573 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1659
timestamp 1624857261
transform 1 0 153909 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1658
timestamp 1624857261
transform 1 0 154245 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1657
timestamp 1624857261
transform 1 0 154581 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1656
timestamp 1624857261
transform 1 0 154917 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1655
timestamp 1624857261
transform 1 0 155253 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1654
timestamp 1624857261
transform 1 0 155589 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1653
timestamp 1624857261
transform 1 0 155925 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1652
timestamp 1624857261
transform 1 0 156261 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1651
timestamp 1624857261
transform 1 0 156597 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1650
timestamp 1624857261
transform 1 0 156933 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1649
timestamp 1624857261
transform 1 0 157269 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1648
timestamp 1624857261
transform 1 0 157605 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1647
timestamp 1624857261
transform 1 0 157941 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1646
timestamp 1624857261
transform 1 0 158277 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1645
timestamp 1624857261
transform 1 0 158613 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1644
timestamp 1624857261
transform 1 0 158949 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1643
timestamp 1624857261
transform 1 0 159285 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1642
timestamp 1624857261
transform 1 0 159621 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1641
timestamp 1624857261
transform 1 0 159957 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1640
timestamp 1624857261
transform 1 0 160293 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1639
timestamp 1624857261
transform 1 0 160629 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1638
timestamp 1624857261
transform 1 0 160965 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1637
timestamp 1624857261
transform 1 0 161301 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1636
timestamp 1624857261
transform 1 0 161637 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1635
timestamp 1624857261
transform 1 0 161973 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1634
timestamp 1624857261
transform 1 0 162309 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1633
timestamp 1624857261
transform 1 0 162645 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1632
timestamp 1624857261
transform 1 0 162981 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1631
timestamp 1624857261
transform 1 0 163317 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1630
timestamp 1624857261
transform 1 0 163653 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1629
timestamp 1624857261
transform 1 0 163989 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1628
timestamp 1624857261
transform 1 0 164325 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1627
timestamp 1624857261
transform 1 0 164661 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1626
timestamp 1624857261
transform 1 0 164997 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1625
timestamp 1624857261
transform 1 0 165333 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1624
timestamp 1624857261
transform 1 0 165669 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1623
timestamp 1624857261
transform 1 0 166005 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1622
timestamp 1624857261
transform 1 0 166341 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1621
timestamp 1624857261
transform 1 0 166677 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1620
timestamp 1624857261
transform 1 0 167013 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1619
timestamp 1624857261
transform 1 0 167349 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1618
timestamp 1624857261
transform 1 0 167685 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1617
timestamp 1624857261
transform 1 0 168021 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1616
timestamp 1624857261
transform 1 0 168357 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1615
timestamp 1624857261
transform 1 0 168693 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1614
timestamp 1624857261
transform 1 0 169029 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1613
timestamp 1624857261
transform 1 0 169365 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1612
timestamp 1624857261
transform 1 0 169701 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1611
timestamp 1624857261
transform 1 0 170037 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1610
timestamp 1624857261
transform 1 0 170373 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1609
timestamp 1624857261
transform 1 0 170709 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1608
timestamp 1624857261
transform 1 0 171045 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1607
timestamp 1624857261
transform 1 0 171381 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1606
timestamp 1624857261
transform 1 0 171717 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1605
timestamp 1624857261
transform 1 0 172053 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1604
timestamp 1624857261
transform 1 0 172389 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1603
timestamp 1624857261
transform 1 0 172725 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1602
timestamp 1624857261
transform 1 0 173061 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1601
timestamp 1624857261
transform 1 0 173397 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1600
timestamp 1624857261
transform 1 0 173733 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1599
timestamp 1624857261
transform 1 0 174069 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1598
timestamp 1624857261
transform 1 0 174405 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1597
timestamp 1624857261
transform 1 0 174741 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1596
timestamp 1624857261
transform 1 0 175077 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1595
timestamp 1624857261
transform 1 0 175413 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1594
timestamp 1624857261
transform 1 0 175749 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1593
timestamp 1624857261
transform 1 0 176085 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1592
timestamp 1624857261
transform 1 0 176421 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1591
timestamp 1624857261
transform 1 0 176757 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1590
timestamp 1624857261
transform 1 0 177093 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1589
timestamp 1624857261
transform 1 0 177429 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1588
timestamp 1624857261
transform 1 0 177765 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1587
timestamp 1624857261
transform 1 0 178101 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1586
timestamp 1624857261
transform 1 0 178437 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1585
timestamp 1624857261
transform 1 0 178773 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1584
timestamp 1624857261
transform 1 0 179109 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1583
timestamp 1624857261
transform 1 0 179445 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1582
timestamp 1624857261
transform 1 0 179781 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1581
timestamp 1624857261
transform 1 0 180117 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1580
timestamp 1624857261
transform 1 0 180453 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1579
timestamp 1624857261
transform 1 0 180789 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1578
timestamp 1624857261
transform 1 0 181125 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1577
timestamp 1624857261
transform 1 0 181461 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1576
timestamp 1624857261
transform 1 0 181797 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1575
timestamp 1624857261
transform 1 0 182133 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1574
timestamp 1624857261
transform 1 0 182469 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1573
timestamp 1624857261
transform 1 0 182805 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1572
timestamp 1624857261
transform 1 0 183141 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1571
timestamp 1624857261
transform 1 0 183477 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1570
timestamp 1624857261
transform 1 0 183813 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1569
timestamp 1624857261
transform 1 0 184149 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1568
timestamp 1624857261
transform 1 0 184485 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1567
timestamp 1624857261
transform 1 0 184821 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1566
timestamp 1624857261
transform 1 0 185157 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1565
timestamp 1624857261
transform 1 0 185493 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1564
timestamp 1624857261
transform 1 0 185829 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1563
timestamp 1624857261
transform 1 0 186165 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1562
timestamp 1624857261
transform 1 0 186501 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1561
timestamp 1624857261
transform 1 0 186837 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1560
timestamp 1624857261
transform 1 0 187173 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1559
timestamp 1624857261
transform 1 0 187509 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1558
timestamp 1624857261
transform 1 0 187845 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1557
timestamp 1624857261
transform 1 0 188181 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1556
timestamp 1624857261
transform 1 0 188517 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1555
timestamp 1624857261
transform 1 0 188853 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1554
timestamp 1624857261
transform 1 0 189189 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1553
timestamp 1624857261
transform 1 0 189525 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1552
timestamp 1624857261
transform 1 0 189861 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1551
timestamp 1624857261
transform 1 0 190197 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1550
timestamp 1624857261
transform 1 0 190533 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1549
timestamp 1624857261
transform 1 0 190869 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1548
timestamp 1624857261
transform 1 0 191205 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1547
timestamp 1624857261
transform 1 0 191541 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1546
timestamp 1624857261
transform 1 0 191877 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1545
timestamp 1624857261
transform 1 0 192213 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1544
timestamp 1624857261
transform 1 0 192549 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1543
timestamp 1624857261
transform 1 0 192885 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1542
timestamp 1624857261
transform 1 0 193221 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1541
timestamp 1624857261
transform 1 0 193557 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1540
timestamp 1624857261
transform 1 0 193893 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1539
timestamp 1624857261
transform 1 0 194229 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1538
timestamp 1624857261
transform 1 0 194565 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1537
timestamp 1624857261
transform 1 0 194901 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1536
timestamp 1624857261
transform 1 0 195237 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1535
timestamp 1624857261
transform 1 0 195573 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1534
timestamp 1624857261
transform 1 0 195909 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1533
timestamp 1624857261
transform 1 0 196245 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1532
timestamp 1624857261
transform 1 0 196581 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1531
timestamp 1624857261
transform 1 0 196917 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1530
timestamp 1624857261
transform 1 0 197253 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1529
timestamp 1624857261
transform 1 0 197589 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1528
timestamp 1624857261
transform 1 0 197925 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1527
timestamp 1624857261
transform 1 0 198261 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1526
timestamp 1624857261
transform 1 0 198597 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1525
timestamp 1624857261
transform 1 0 198933 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1524
timestamp 1624857261
transform 1 0 199269 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1523
timestamp 1624857261
transform 1 0 199605 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1522
timestamp 1624857261
transform 1 0 199941 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1521
timestamp 1624857261
transform 1 0 200277 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1520
timestamp 1624857261
transform 1 0 200613 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1519
timestamp 1624857261
transform 1 0 200949 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1518
timestamp 1624857261
transform 1 0 201285 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1517
timestamp 1624857261
transform 1 0 201621 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1516
timestamp 1624857261
transform 1 0 201957 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1515
timestamp 1624857261
transform 1 0 202293 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1514
timestamp 1624857261
transform 1 0 202629 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1513
timestamp 1624857261
transform 1 0 202965 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1512
timestamp 1624857261
transform 1 0 203301 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1511
timestamp 1624857261
transform 1 0 203637 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1510
timestamp 1624857261
transform 1 0 203973 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1509
timestamp 1624857261
transform 1 0 204309 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1508
timestamp 1624857261
transform 1 0 204645 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1507
timestamp 1624857261
transform 1 0 204981 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1506
timestamp 1624857261
transform 1 0 205317 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1505
timestamp 1624857261
transform 1 0 205653 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1504
timestamp 1624857261
transform 1 0 205989 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1503
timestamp 1624857261
transform 1 0 206325 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1502
timestamp 1624857261
transform 1 0 206661 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1501
timestamp 1624857261
transform 1 0 206997 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1500
timestamp 1624857261
transform 1 0 207333 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1499
timestamp 1624857261
transform 1 0 207669 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1498
timestamp 1624857261
transform 1 0 208005 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1497
timestamp 1624857261
transform 1 0 208341 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1496
timestamp 1624857261
transform 1 0 208677 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1495
timestamp 1624857261
transform 1 0 209013 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1494
timestamp 1624857261
transform 1 0 209349 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1493
timestamp 1624857261
transform 1 0 209685 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1492
timestamp 1624857261
transform 1 0 210021 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1491
timestamp 1624857261
transform 1 0 210357 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1490
timestamp 1624857261
transform 1 0 210693 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1489
timestamp 1624857261
transform 1 0 211029 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1488
timestamp 1624857261
transform 1 0 211365 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1487
timestamp 1624857261
transform 1 0 211701 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1486
timestamp 1624857261
transform 1 0 212037 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1485
timestamp 1624857261
transform 1 0 212373 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1484
timestamp 1624857261
transform 1 0 212709 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1483
timestamp 1624857261
transform 1 0 213045 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1482
timestamp 1624857261
transform 1 0 213381 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1481
timestamp 1624857261
transform 1 0 213717 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1480
timestamp 1624857261
transform 1 0 214053 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1479
timestamp 1624857261
transform 1 0 214389 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1478
timestamp 1624857261
transform 1 0 214725 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1477
timestamp 1624857261
transform 1 0 215061 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1476
timestamp 1624857261
transform 1 0 215397 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1475
timestamp 1624857261
transform 1 0 215733 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1474
timestamp 1624857261
transform 1 0 216069 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1473
timestamp 1624857261
transform 1 0 216405 0 1 1815
box 0 0 1 1
use contact_7  contact_7_1472
timestamp 1624857261
transform 1 0 2037 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1471
timestamp 1624857261
transform 1 0 2373 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1470
timestamp 1624857261
transform 1 0 2709 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1469
timestamp 1624857261
transform 1 0 3045 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1468
timestamp 1624857261
transform 1 0 3381 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1467
timestamp 1624857261
transform 1 0 3717 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1466
timestamp 1624857261
transform 1 0 4053 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1465
timestamp 1624857261
transform 1 0 4389 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1464
timestamp 1624857261
transform 1 0 4725 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1463
timestamp 1624857261
transform 1 0 5061 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1462
timestamp 1624857261
transform 1 0 5397 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1461
timestamp 1624857261
transform 1 0 5733 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1460
timestamp 1624857261
transform 1 0 6069 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1459
timestamp 1624857261
transform 1 0 6405 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1458
timestamp 1624857261
transform 1 0 6741 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1457
timestamp 1624857261
transform 1 0 7077 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1456
timestamp 1624857261
transform 1 0 7413 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1455
timestamp 1624857261
transform 1 0 7749 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1454
timestamp 1624857261
transform 1 0 8085 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1453
timestamp 1624857261
transform 1 0 8421 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1452
timestamp 1624857261
transform 1 0 8757 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1451
timestamp 1624857261
transform 1 0 9093 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1450
timestamp 1624857261
transform 1 0 9429 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1449
timestamp 1624857261
transform 1 0 9765 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1448
timestamp 1624857261
transform 1 0 10101 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1447
timestamp 1624857261
transform 1 0 10437 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1446
timestamp 1624857261
transform 1 0 10773 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1445
timestamp 1624857261
transform 1 0 11109 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1444
timestamp 1624857261
transform 1 0 11445 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1443
timestamp 1624857261
transform 1 0 11781 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1442
timestamp 1624857261
transform 1 0 12117 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1441
timestamp 1624857261
transform 1 0 12453 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1440
timestamp 1624857261
transform 1 0 12789 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1439
timestamp 1624857261
transform 1 0 13125 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1438
timestamp 1624857261
transform 1 0 13461 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1437
timestamp 1624857261
transform 1 0 13797 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1436
timestamp 1624857261
transform 1 0 14133 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1435
timestamp 1624857261
transform 1 0 14469 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1434
timestamp 1624857261
transform 1 0 14805 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1433
timestamp 1624857261
transform 1 0 15141 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1432
timestamp 1624857261
transform 1 0 15477 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1431
timestamp 1624857261
transform 1 0 15813 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1430
timestamp 1624857261
transform 1 0 16149 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1429
timestamp 1624857261
transform 1 0 16485 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1428
timestamp 1624857261
transform 1 0 16821 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1427
timestamp 1624857261
transform 1 0 17157 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1426
timestamp 1624857261
transform 1 0 17493 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1425
timestamp 1624857261
transform 1 0 17829 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1424
timestamp 1624857261
transform 1 0 18165 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1423
timestamp 1624857261
transform 1 0 18501 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1422
timestamp 1624857261
transform 1 0 18837 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1421
timestamp 1624857261
transform 1 0 19173 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1420
timestamp 1624857261
transform 1 0 19509 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1419
timestamp 1624857261
transform 1 0 19845 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1418
timestamp 1624857261
transform 1 0 20181 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1417
timestamp 1624857261
transform 1 0 20517 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1416
timestamp 1624857261
transform 1 0 20853 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1415
timestamp 1624857261
transform 1 0 21189 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1414
timestamp 1624857261
transform 1 0 21525 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1413
timestamp 1624857261
transform 1 0 21861 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1412
timestamp 1624857261
transform 1 0 22197 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1411
timestamp 1624857261
transform 1 0 22533 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1410
timestamp 1624857261
transform 1 0 22869 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1409
timestamp 1624857261
transform 1 0 23205 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1408
timestamp 1624857261
transform 1 0 23541 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1407
timestamp 1624857261
transform 1 0 23877 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1406
timestamp 1624857261
transform 1 0 24213 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1405
timestamp 1624857261
transform 1 0 24549 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1404
timestamp 1624857261
transform 1 0 24885 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1403
timestamp 1624857261
transform 1 0 25221 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1402
timestamp 1624857261
transform 1 0 25557 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1401
timestamp 1624857261
transform 1 0 25893 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1400
timestamp 1624857261
transform 1 0 26229 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1399
timestamp 1624857261
transform 1 0 26565 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1398
timestamp 1624857261
transform 1 0 26901 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1397
timestamp 1624857261
transform 1 0 27237 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1396
timestamp 1624857261
transform 1 0 27573 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1395
timestamp 1624857261
transform 1 0 27909 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1394
timestamp 1624857261
transform 1 0 28245 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1393
timestamp 1624857261
transform 1 0 28581 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1392
timestamp 1624857261
transform 1 0 28917 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1391
timestamp 1624857261
transform 1 0 29253 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1390
timestamp 1624857261
transform 1 0 29589 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1389
timestamp 1624857261
transform 1 0 29925 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1388
timestamp 1624857261
transform 1 0 30261 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1387
timestamp 1624857261
transform 1 0 30597 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1386
timestamp 1624857261
transform 1 0 30933 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1385
timestamp 1624857261
transform 1 0 31269 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1384
timestamp 1624857261
transform 1 0 31605 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1383
timestamp 1624857261
transform 1 0 31941 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1382
timestamp 1624857261
transform 1 0 32277 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1381
timestamp 1624857261
transform 1 0 32613 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1380
timestamp 1624857261
transform 1 0 32949 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1379
timestamp 1624857261
transform 1 0 33285 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1378
timestamp 1624857261
transform 1 0 33621 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1377
timestamp 1624857261
transform 1 0 33957 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1376
timestamp 1624857261
transform 1 0 34293 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1375
timestamp 1624857261
transform 1 0 34629 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1374
timestamp 1624857261
transform 1 0 34965 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1373
timestamp 1624857261
transform 1 0 35301 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1372
timestamp 1624857261
transform 1 0 35637 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1371
timestamp 1624857261
transform 1 0 35973 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1370
timestamp 1624857261
transform 1 0 36309 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1369
timestamp 1624857261
transform 1 0 36645 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1368
timestamp 1624857261
transform 1 0 36981 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1367
timestamp 1624857261
transform 1 0 37317 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1366
timestamp 1624857261
transform 1 0 37653 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1365
timestamp 1624857261
transform 1 0 37989 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1364
timestamp 1624857261
transform 1 0 38325 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1363
timestamp 1624857261
transform 1 0 38661 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1362
timestamp 1624857261
transform 1 0 38997 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1361
timestamp 1624857261
transform 1 0 39333 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1360
timestamp 1624857261
transform 1 0 39669 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1359
timestamp 1624857261
transform 1 0 40005 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1358
timestamp 1624857261
transform 1 0 40341 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1357
timestamp 1624857261
transform 1 0 40677 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1356
timestamp 1624857261
transform 1 0 41013 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1355
timestamp 1624857261
transform 1 0 41349 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1354
timestamp 1624857261
transform 1 0 41685 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1353
timestamp 1624857261
transform 1 0 42021 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1352
timestamp 1624857261
transform 1 0 42357 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1351
timestamp 1624857261
transform 1 0 42693 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1350
timestamp 1624857261
transform 1 0 43029 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1349
timestamp 1624857261
transform 1 0 43365 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1348
timestamp 1624857261
transform 1 0 43701 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1347
timestamp 1624857261
transform 1 0 44037 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1346
timestamp 1624857261
transform 1 0 44373 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1345
timestamp 1624857261
transform 1 0 44709 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1344
timestamp 1624857261
transform 1 0 45045 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1343
timestamp 1624857261
transform 1 0 45381 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1342
timestamp 1624857261
transform 1 0 45717 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1341
timestamp 1624857261
transform 1 0 46053 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1340
timestamp 1624857261
transform 1 0 46389 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1339
timestamp 1624857261
transform 1 0 46725 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1338
timestamp 1624857261
transform 1 0 47061 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1337
timestamp 1624857261
transform 1 0 47397 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1336
timestamp 1624857261
transform 1 0 47733 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1335
timestamp 1624857261
transform 1 0 48069 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1334
timestamp 1624857261
transform 1 0 48405 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1333
timestamp 1624857261
transform 1 0 48741 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1332
timestamp 1624857261
transform 1 0 49077 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1331
timestamp 1624857261
transform 1 0 49413 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1330
timestamp 1624857261
transform 1 0 49749 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1329
timestamp 1624857261
transform 1 0 50085 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1328
timestamp 1624857261
transform 1 0 50421 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1327
timestamp 1624857261
transform 1 0 50757 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1326
timestamp 1624857261
transform 1 0 51093 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1325
timestamp 1624857261
transform 1 0 51429 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1324
timestamp 1624857261
transform 1 0 51765 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1323
timestamp 1624857261
transform 1 0 52101 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1322
timestamp 1624857261
transform 1 0 52437 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1321
timestamp 1624857261
transform 1 0 52773 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1320
timestamp 1624857261
transform 1 0 53109 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1319
timestamp 1624857261
transform 1 0 53445 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1318
timestamp 1624857261
transform 1 0 53781 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1317
timestamp 1624857261
transform 1 0 54117 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1316
timestamp 1624857261
transform 1 0 54453 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1315
timestamp 1624857261
transform 1 0 54789 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1314
timestamp 1624857261
transform 1 0 55125 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1313
timestamp 1624857261
transform 1 0 55461 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1312
timestamp 1624857261
transform 1 0 55797 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1311
timestamp 1624857261
transform 1 0 56133 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1310
timestamp 1624857261
transform 1 0 56469 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1309
timestamp 1624857261
transform 1 0 56805 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1308
timestamp 1624857261
transform 1 0 57141 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1307
timestamp 1624857261
transform 1 0 57477 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1306
timestamp 1624857261
transform 1 0 57813 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1305
timestamp 1624857261
transform 1 0 58149 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1304
timestamp 1624857261
transform 1 0 58485 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1303
timestamp 1624857261
transform 1 0 58821 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1302
timestamp 1624857261
transform 1 0 59157 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1301
timestamp 1624857261
transform 1 0 59493 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1300
timestamp 1624857261
transform 1 0 59829 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1299
timestamp 1624857261
transform 1 0 60165 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1298
timestamp 1624857261
transform 1 0 60501 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1297
timestamp 1624857261
transform 1 0 60837 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1296
timestamp 1624857261
transform 1 0 61173 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1295
timestamp 1624857261
transform 1 0 61509 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1294
timestamp 1624857261
transform 1 0 61845 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1293
timestamp 1624857261
transform 1 0 62181 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1292
timestamp 1624857261
transform 1 0 62517 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1291
timestamp 1624857261
transform 1 0 62853 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1290
timestamp 1624857261
transform 1 0 63189 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1289
timestamp 1624857261
transform 1 0 63525 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1288
timestamp 1624857261
transform 1 0 63861 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1287
timestamp 1624857261
transform 1 0 64197 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1286
timestamp 1624857261
transform 1 0 64533 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1285
timestamp 1624857261
transform 1 0 64869 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1284
timestamp 1624857261
transform 1 0 65205 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1283
timestamp 1624857261
transform 1 0 65541 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1282
timestamp 1624857261
transform 1 0 65877 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1281
timestamp 1624857261
transform 1 0 66213 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1280
timestamp 1624857261
transform 1 0 66549 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1279
timestamp 1624857261
transform 1 0 66885 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1278
timestamp 1624857261
transform 1 0 67221 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1277
timestamp 1624857261
transform 1 0 67557 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1276
timestamp 1624857261
transform 1 0 67893 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1275
timestamp 1624857261
transform 1 0 68229 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1274
timestamp 1624857261
transform 1 0 68565 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1273
timestamp 1624857261
transform 1 0 68901 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1272
timestamp 1624857261
transform 1 0 69237 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1271
timestamp 1624857261
transform 1 0 69573 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1270
timestamp 1624857261
transform 1 0 69909 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1269
timestamp 1624857261
transform 1 0 70245 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1268
timestamp 1624857261
transform 1 0 70581 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1267
timestamp 1624857261
transform 1 0 70917 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1266
timestamp 1624857261
transform 1 0 71253 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1265
timestamp 1624857261
transform 1 0 71589 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1264
timestamp 1624857261
transform 1 0 71925 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1263
timestamp 1624857261
transform 1 0 72261 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1262
timestamp 1624857261
transform 1 0 72597 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1261
timestamp 1624857261
transform 1 0 72933 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1260
timestamp 1624857261
transform 1 0 73269 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1259
timestamp 1624857261
transform 1 0 73605 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1258
timestamp 1624857261
transform 1 0 73941 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1257
timestamp 1624857261
transform 1 0 74277 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1256
timestamp 1624857261
transform 1 0 74613 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1255
timestamp 1624857261
transform 1 0 74949 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1254
timestamp 1624857261
transform 1 0 75285 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1253
timestamp 1624857261
transform 1 0 75621 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1252
timestamp 1624857261
transform 1 0 75957 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1251
timestamp 1624857261
transform 1 0 76293 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1250
timestamp 1624857261
transform 1 0 76629 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1249
timestamp 1624857261
transform 1 0 76965 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1248
timestamp 1624857261
transform 1 0 77301 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1247
timestamp 1624857261
transform 1 0 77637 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1246
timestamp 1624857261
transform 1 0 77973 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1245
timestamp 1624857261
transform 1 0 78309 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1244
timestamp 1624857261
transform 1 0 78645 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1243
timestamp 1624857261
transform 1 0 78981 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1242
timestamp 1624857261
transform 1 0 79317 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1241
timestamp 1624857261
transform 1 0 79653 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1240
timestamp 1624857261
transform 1 0 79989 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1239
timestamp 1624857261
transform 1 0 80325 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1238
timestamp 1624857261
transform 1 0 80661 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1237
timestamp 1624857261
transform 1 0 80997 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1236
timestamp 1624857261
transform 1 0 81333 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1235
timestamp 1624857261
transform 1 0 81669 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1234
timestamp 1624857261
transform 1 0 82005 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1233
timestamp 1624857261
transform 1 0 82341 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1232
timestamp 1624857261
transform 1 0 82677 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1231
timestamp 1624857261
transform 1 0 83013 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1230
timestamp 1624857261
transform 1 0 83349 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1229
timestamp 1624857261
transform 1 0 83685 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1228
timestamp 1624857261
transform 1 0 84021 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1227
timestamp 1624857261
transform 1 0 84357 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1226
timestamp 1624857261
transform 1 0 84693 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1225
timestamp 1624857261
transform 1 0 85029 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1224
timestamp 1624857261
transform 1 0 85365 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1223
timestamp 1624857261
transform 1 0 85701 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1222
timestamp 1624857261
transform 1 0 86037 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1221
timestamp 1624857261
transform 1 0 86373 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1220
timestamp 1624857261
transform 1 0 86709 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1219
timestamp 1624857261
transform 1 0 87045 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1218
timestamp 1624857261
transform 1 0 87381 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1217
timestamp 1624857261
transform 1 0 87717 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1216
timestamp 1624857261
transform 1 0 88053 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1215
timestamp 1624857261
transform 1 0 88389 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1214
timestamp 1624857261
transform 1 0 88725 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1213
timestamp 1624857261
transform 1 0 89061 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1212
timestamp 1624857261
transform 1 0 89397 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1211
timestamp 1624857261
transform 1 0 89733 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1210
timestamp 1624857261
transform 1 0 90069 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1209
timestamp 1624857261
transform 1 0 90405 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1208
timestamp 1624857261
transform 1 0 90741 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1207
timestamp 1624857261
transform 1 0 91077 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1206
timestamp 1624857261
transform 1 0 91413 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1205
timestamp 1624857261
transform 1 0 91749 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1204
timestamp 1624857261
transform 1 0 92085 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1203
timestamp 1624857261
transform 1 0 92421 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1202
timestamp 1624857261
transform 1 0 92757 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1201
timestamp 1624857261
transform 1 0 93093 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1200
timestamp 1624857261
transform 1 0 93429 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1199
timestamp 1624857261
transform 1 0 93765 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1198
timestamp 1624857261
transform 1 0 94101 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1197
timestamp 1624857261
transform 1 0 94437 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1196
timestamp 1624857261
transform 1 0 94773 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1195
timestamp 1624857261
transform 1 0 95109 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1194
timestamp 1624857261
transform 1 0 95445 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1193
timestamp 1624857261
transform 1 0 95781 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1192
timestamp 1624857261
transform 1 0 96117 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1191
timestamp 1624857261
transform 1 0 96453 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1190
timestamp 1624857261
transform 1 0 96789 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1189
timestamp 1624857261
transform 1 0 97125 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1188
timestamp 1624857261
transform 1 0 97461 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1187
timestamp 1624857261
transform 1 0 97797 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1186
timestamp 1624857261
transform 1 0 98133 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1185
timestamp 1624857261
transform 1 0 98469 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1184
timestamp 1624857261
transform 1 0 98805 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1183
timestamp 1624857261
transform 1 0 99141 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1182
timestamp 1624857261
transform 1 0 99477 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1181
timestamp 1624857261
transform 1 0 99813 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1180
timestamp 1624857261
transform 1 0 100149 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1179
timestamp 1624857261
transform 1 0 100485 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1178
timestamp 1624857261
transform 1 0 100821 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1177
timestamp 1624857261
transform 1 0 101157 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1176
timestamp 1624857261
transform 1 0 101493 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1175
timestamp 1624857261
transform 1 0 101829 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1174
timestamp 1624857261
transform 1 0 102165 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1173
timestamp 1624857261
transform 1 0 102501 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1172
timestamp 1624857261
transform 1 0 102837 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1171
timestamp 1624857261
transform 1 0 103173 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1170
timestamp 1624857261
transform 1 0 103509 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1169
timestamp 1624857261
transform 1 0 103845 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1168
timestamp 1624857261
transform 1 0 104181 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1167
timestamp 1624857261
transform 1 0 104517 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1166
timestamp 1624857261
transform 1 0 104853 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1165
timestamp 1624857261
transform 1 0 105189 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1164
timestamp 1624857261
transform 1 0 105525 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1163
timestamp 1624857261
transform 1 0 105861 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1162
timestamp 1624857261
transform 1 0 106197 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1161
timestamp 1624857261
transform 1 0 106533 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1160
timestamp 1624857261
transform 1 0 106869 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1159
timestamp 1624857261
transform 1 0 107205 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1158
timestamp 1624857261
transform 1 0 107541 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1157
timestamp 1624857261
transform 1 0 107877 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1156
timestamp 1624857261
transform 1 0 108213 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1155
timestamp 1624857261
transform 1 0 108549 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1154
timestamp 1624857261
transform 1 0 108885 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1153
timestamp 1624857261
transform 1 0 109221 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1152
timestamp 1624857261
transform 1 0 109557 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1151
timestamp 1624857261
transform 1 0 109893 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1150
timestamp 1624857261
transform 1 0 110229 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1149
timestamp 1624857261
transform 1 0 110565 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1148
timestamp 1624857261
transform 1 0 110901 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1147
timestamp 1624857261
transform 1 0 111237 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1146
timestamp 1624857261
transform 1 0 111573 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1145
timestamp 1624857261
transform 1 0 111909 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1144
timestamp 1624857261
transform 1 0 112245 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1143
timestamp 1624857261
transform 1 0 112581 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1142
timestamp 1624857261
transform 1 0 112917 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1141
timestamp 1624857261
transform 1 0 113253 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1140
timestamp 1624857261
transform 1 0 113589 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1139
timestamp 1624857261
transform 1 0 113925 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1138
timestamp 1624857261
transform 1 0 114261 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1137
timestamp 1624857261
transform 1 0 114597 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1136
timestamp 1624857261
transform 1 0 114933 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1135
timestamp 1624857261
transform 1 0 115269 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1134
timestamp 1624857261
transform 1 0 115605 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1133
timestamp 1624857261
transform 1 0 115941 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1132
timestamp 1624857261
transform 1 0 116277 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1131
timestamp 1624857261
transform 1 0 116613 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1130
timestamp 1624857261
transform 1 0 116949 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1129
timestamp 1624857261
transform 1 0 117285 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1128
timestamp 1624857261
transform 1 0 117621 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1127
timestamp 1624857261
transform 1 0 117957 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1126
timestamp 1624857261
transform 1 0 118293 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1125
timestamp 1624857261
transform 1 0 118629 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1124
timestamp 1624857261
transform 1 0 118965 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1123
timestamp 1624857261
transform 1 0 119301 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1122
timestamp 1624857261
transform 1 0 119637 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1121
timestamp 1624857261
transform 1 0 119973 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1120
timestamp 1624857261
transform 1 0 120309 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1119
timestamp 1624857261
transform 1 0 120645 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1118
timestamp 1624857261
transform 1 0 120981 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1117
timestamp 1624857261
transform 1 0 121317 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1116
timestamp 1624857261
transform 1 0 121653 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1115
timestamp 1624857261
transform 1 0 121989 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1114
timestamp 1624857261
transform 1 0 122325 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1113
timestamp 1624857261
transform 1 0 122661 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1112
timestamp 1624857261
transform 1 0 122997 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1111
timestamp 1624857261
transform 1 0 123333 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1110
timestamp 1624857261
transform 1 0 123669 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1109
timestamp 1624857261
transform 1 0 124005 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1108
timestamp 1624857261
transform 1 0 124341 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1107
timestamp 1624857261
transform 1 0 124677 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1106
timestamp 1624857261
transform 1 0 125013 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1105
timestamp 1624857261
transform 1 0 125349 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1104
timestamp 1624857261
transform 1 0 125685 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1103
timestamp 1624857261
transform 1 0 126021 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1102
timestamp 1624857261
transform 1 0 126357 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1101
timestamp 1624857261
transform 1 0 126693 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1100
timestamp 1624857261
transform 1 0 127029 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1099
timestamp 1624857261
transform 1 0 127365 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1098
timestamp 1624857261
transform 1 0 127701 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1097
timestamp 1624857261
transform 1 0 128037 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1096
timestamp 1624857261
transform 1 0 128373 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1095
timestamp 1624857261
transform 1 0 128709 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1094
timestamp 1624857261
transform 1 0 129045 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1093
timestamp 1624857261
transform 1 0 129381 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1092
timestamp 1624857261
transform 1 0 129717 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1091
timestamp 1624857261
transform 1 0 130053 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1090
timestamp 1624857261
transform 1 0 130389 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1089
timestamp 1624857261
transform 1 0 130725 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1088
timestamp 1624857261
transform 1 0 131061 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1087
timestamp 1624857261
transform 1 0 131397 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1086
timestamp 1624857261
transform 1 0 131733 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1085
timestamp 1624857261
transform 1 0 132069 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1084
timestamp 1624857261
transform 1 0 132405 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1083
timestamp 1624857261
transform 1 0 132741 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1082
timestamp 1624857261
transform 1 0 133077 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1081
timestamp 1624857261
transform 1 0 133413 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1080
timestamp 1624857261
transform 1 0 133749 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1079
timestamp 1624857261
transform 1 0 134085 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1078
timestamp 1624857261
transform 1 0 134421 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1077
timestamp 1624857261
transform 1 0 134757 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1076
timestamp 1624857261
transform 1 0 135093 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1075
timestamp 1624857261
transform 1 0 135429 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1074
timestamp 1624857261
transform 1 0 135765 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1073
timestamp 1624857261
transform 1 0 136101 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1072
timestamp 1624857261
transform 1 0 136437 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1071
timestamp 1624857261
transform 1 0 136773 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1070
timestamp 1624857261
transform 1 0 137109 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1069
timestamp 1624857261
transform 1 0 137445 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1068
timestamp 1624857261
transform 1 0 137781 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1067
timestamp 1624857261
transform 1 0 138117 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1066
timestamp 1624857261
transform 1 0 138453 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1065
timestamp 1624857261
transform 1 0 138789 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1064
timestamp 1624857261
transform 1 0 139125 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1063
timestamp 1624857261
transform 1 0 139461 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1062
timestamp 1624857261
transform 1 0 139797 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1061
timestamp 1624857261
transform 1 0 140133 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1060
timestamp 1624857261
transform 1 0 140469 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1059
timestamp 1624857261
transform 1 0 140805 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1058
timestamp 1624857261
transform 1 0 141141 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1057
timestamp 1624857261
transform 1 0 141477 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1056
timestamp 1624857261
transform 1 0 141813 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1055
timestamp 1624857261
transform 1 0 142149 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1054
timestamp 1624857261
transform 1 0 142485 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1053
timestamp 1624857261
transform 1 0 142821 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1052
timestamp 1624857261
transform 1 0 143157 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1051
timestamp 1624857261
transform 1 0 143493 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1050
timestamp 1624857261
transform 1 0 143829 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1049
timestamp 1624857261
transform 1 0 144165 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1048
timestamp 1624857261
transform 1 0 144501 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1047
timestamp 1624857261
transform 1 0 144837 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1046
timestamp 1624857261
transform 1 0 145173 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1045
timestamp 1624857261
transform 1 0 145509 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1044
timestamp 1624857261
transform 1 0 145845 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1043
timestamp 1624857261
transform 1 0 146181 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1042
timestamp 1624857261
transform 1 0 146517 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1041
timestamp 1624857261
transform 1 0 146853 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1040
timestamp 1624857261
transform 1 0 147189 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1039
timestamp 1624857261
transform 1 0 147525 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1038
timestamp 1624857261
transform 1 0 147861 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1037
timestamp 1624857261
transform 1 0 148197 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1036
timestamp 1624857261
transform 1 0 148533 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1035
timestamp 1624857261
transform 1 0 148869 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1034
timestamp 1624857261
transform 1 0 149205 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1033
timestamp 1624857261
transform 1 0 149541 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1032
timestamp 1624857261
transform 1 0 149877 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1031
timestamp 1624857261
transform 1 0 150213 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1030
timestamp 1624857261
transform 1 0 150549 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1029
timestamp 1624857261
transform 1 0 150885 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1028
timestamp 1624857261
transform 1 0 151221 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1027
timestamp 1624857261
transform 1 0 151557 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1026
timestamp 1624857261
transform 1 0 151893 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1025
timestamp 1624857261
transform 1 0 152229 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1024
timestamp 1624857261
transform 1 0 152565 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1023
timestamp 1624857261
transform 1 0 152901 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1022
timestamp 1624857261
transform 1 0 153237 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1021
timestamp 1624857261
transform 1 0 153573 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1020
timestamp 1624857261
transform 1 0 153909 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1019
timestamp 1624857261
transform 1 0 154245 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1018
timestamp 1624857261
transform 1 0 154581 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1017
timestamp 1624857261
transform 1 0 154917 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1016
timestamp 1624857261
transform 1 0 155253 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1015
timestamp 1624857261
transform 1 0 155589 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1014
timestamp 1624857261
transform 1 0 155925 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1013
timestamp 1624857261
transform 1 0 156261 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1012
timestamp 1624857261
transform 1 0 156597 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1011
timestamp 1624857261
transform 1 0 156933 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1010
timestamp 1624857261
transform 1 0 157269 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1009
timestamp 1624857261
transform 1 0 157605 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1008
timestamp 1624857261
transform 1 0 157941 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1007
timestamp 1624857261
transform 1 0 158277 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1006
timestamp 1624857261
transform 1 0 158613 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1005
timestamp 1624857261
transform 1 0 158949 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1004
timestamp 1624857261
transform 1 0 159285 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1003
timestamp 1624857261
transform 1 0 159621 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1002
timestamp 1624857261
transform 1 0 159957 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1001
timestamp 1624857261
transform 1 0 160293 0 1 142311
box 0 0 1 1
use contact_7  contact_7_1000
timestamp 1624857261
transform 1 0 160629 0 1 142311
box 0 0 1 1
use contact_7  contact_7_999
timestamp 1624857261
transform 1 0 160965 0 1 142311
box 0 0 1 1
use contact_7  contact_7_998
timestamp 1624857261
transform 1 0 161301 0 1 142311
box 0 0 1 1
use contact_7  contact_7_997
timestamp 1624857261
transform 1 0 161637 0 1 142311
box 0 0 1 1
use contact_7  contact_7_996
timestamp 1624857261
transform 1 0 161973 0 1 142311
box 0 0 1 1
use contact_7  contact_7_995
timestamp 1624857261
transform 1 0 162309 0 1 142311
box 0 0 1 1
use contact_7  contact_7_994
timestamp 1624857261
transform 1 0 162645 0 1 142311
box 0 0 1 1
use contact_7  contact_7_993
timestamp 1624857261
transform 1 0 162981 0 1 142311
box 0 0 1 1
use contact_7  contact_7_992
timestamp 1624857261
transform 1 0 163317 0 1 142311
box 0 0 1 1
use contact_7  contact_7_991
timestamp 1624857261
transform 1 0 163653 0 1 142311
box 0 0 1 1
use contact_7  contact_7_990
timestamp 1624857261
transform 1 0 163989 0 1 142311
box 0 0 1 1
use contact_7  contact_7_989
timestamp 1624857261
transform 1 0 164325 0 1 142311
box 0 0 1 1
use contact_7  contact_7_988
timestamp 1624857261
transform 1 0 164661 0 1 142311
box 0 0 1 1
use contact_7  contact_7_987
timestamp 1624857261
transform 1 0 164997 0 1 142311
box 0 0 1 1
use contact_7  contact_7_986
timestamp 1624857261
transform 1 0 165333 0 1 142311
box 0 0 1 1
use contact_7  contact_7_985
timestamp 1624857261
transform 1 0 165669 0 1 142311
box 0 0 1 1
use contact_7  contact_7_984
timestamp 1624857261
transform 1 0 166005 0 1 142311
box 0 0 1 1
use contact_7  contact_7_983
timestamp 1624857261
transform 1 0 166341 0 1 142311
box 0 0 1 1
use contact_7  contact_7_982
timestamp 1624857261
transform 1 0 166677 0 1 142311
box 0 0 1 1
use contact_7  contact_7_981
timestamp 1624857261
transform 1 0 167013 0 1 142311
box 0 0 1 1
use contact_7  contact_7_980
timestamp 1624857261
transform 1 0 167349 0 1 142311
box 0 0 1 1
use contact_7  contact_7_979
timestamp 1624857261
transform 1 0 167685 0 1 142311
box 0 0 1 1
use contact_7  contact_7_978
timestamp 1624857261
transform 1 0 168021 0 1 142311
box 0 0 1 1
use contact_7  contact_7_977
timestamp 1624857261
transform 1 0 168357 0 1 142311
box 0 0 1 1
use contact_7  contact_7_976
timestamp 1624857261
transform 1 0 168693 0 1 142311
box 0 0 1 1
use contact_7  contact_7_975
timestamp 1624857261
transform 1 0 169029 0 1 142311
box 0 0 1 1
use contact_7  contact_7_974
timestamp 1624857261
transform 1 0 169365 0 1 142311
box 0 0 1 1
use contact_7  contact_7_973
timestamp 1624857261
transform 1 0 169701 0 1 142311
box 0 0 1 1
use contact_7  contact_7_972
timestamp 1624857261
transform 1 0 170037 0 1 142311
box 0 0 1 1
use contact_7  contact_7_971
timestamp 1624857261
transform 1 0 170373 0 1 142311
box 0 0 1 1
use contact_7  contact_7_970
timestamp 1624857261
transform 1 0 170709 0 1 142311
box 0 0 1 1
use contact_7  contact_7_969
timestamp 1624857261
transform 1 0 171045 0 1 142311
box 0 0 1 1
use contact_7  contact_7_968
timestamp 1624857261
transform 1 0 171381 0 1 142311
box 0 0 1 1
use contact_7  contact_7_967
timestamp 1624857261
transform 1 0 171717 0 1 142311
box 0 0 1 1
use contact_7  contact_7_966
timestamp 1624857261
transform 1 0 172053 0 1 142311
box 0 0 1 1
use contact_7  contact_7_965
timestamp 1624857261
transform 1 0 172389 0 1 142311
box 0 0 1 1
use contact_7  contact_7_964
timestamp 1624857261
transform 1 0 172725 0 1 142311
box 0 0 1 1
use contact_7  contact_7_963
timestamp 1624857261
transform 1 0 173061 0 1 142311
box 0 0 1 1
use contact_7  contact_7_962
timestamp 1624857261
transform 1 0 173397 0 1 142311
box 0 0 1 1
use contact_7  contact_7_961
timestamp 1624857261
transform 1 0 173733 0 1 142311
box 0 0 1 1
use contact_7  contact_7_960
timestamp 1624857261
transform 1 0 174069 0 1 142311
box 0 0 1 1
use contact_7  contact_7_959
timestamp 1624857261
transform 1 0 174405 0 1 142311
box 0 0 1 1
use contact_7  contact_7_958
timestamp 1624857261
transform 1 0 174741 0 1 142311
box 0 0 1 1
use contact_7  contact_7_957
timestamp 1624857261
transform 1 0 175077 0 1 142311
box 0 0 1 1
use contact_7  contact_7_956
timestamp 1624857261
transform 1 0 175413 0 1 142311
box 0 0 1 1
use contact_7  contact_7_955
timestamp 1624857261
transform 1 0 175749 0 1 142311
box 0 0 1 1
use contact_7  contact_7_954
timestamp 1624857261
transform 1 0 176085 0 1 142311
box 0 0 1 1
use contact_7  contact_7_953
timestamp 1624857261
transform 1 0 176421 0 1 142311
box 0 0 1 1
use contact_7  contact_7_952
timestamp 1624857261
transform 1 0 176757 0 1 142311
box 0 0 1 1
use contact_7  contact_7_951
timestamp 1624857261
transform 1 0 177093 0 1 142311
box 0 0 1 1
use contact_7  contact_7_950
timestamp 1624857261
transform 1 0 177429 0 1 142311
box 0 0 1 1
use contact_7  contact_7_949
timestamp 1624857261
transform 1 0 177765 0 1 142311
box 0 0 1 1
use contact_7  contact_7_948
timestamp 1624857261
transform 1 0 178101 0 1 142311
box 0 0 1 1
use contact_7  contact_7_947
timestamp 1624857261
transform 1 0 178437 0 1 142311
box 0 0 1 1
use contact_7  contact_7_946
timestamp 1624857261
transform 1 0 178773 0 1 142311
box 0 0 1 1
use contact_7  contact_7_945
timestamp 1624857261
transform 1 0 179109 0 1 142311
box 0 0 1 1
use contact_7  contact_7_944
timestamp 1624857261
transform 1 0 179445 0 1 142311
box 0 0 1 1
use contact_7  contact_7_943
timestamp 1624857261
transform 1 0 179781 0 1 142311
box 0 0 1 1
use contact_7  contact_7_942
timestamp 1624857261
transform 1 0 180117 0 1 142311
box 0 0 1 1
use contact_7  contact_7_941
timestamp 1624857261
transform 1 0 180453 0 1 142311
box 0 0 1 1
use contact_7  contact_7_940
timestamp 1624857261
transform 1 0 180789 0 1 142311
box 0 0 1 1
use contact_7  contact_7_939
timestamp 1624857261
transform 1 0 181125 0 1 142311
box 0 0 1 1
use contact_7  contact_7_938
timestamp 1624857261
transform 1 0 181461 0 1 142311
box 0 0 1 1
use contact_7  contact_7_937
timestamp 1624857261
transform 1 0 181797 0 1 142311
box 0 0 1 1
use contact_7  contact_7_936
timestamp 1624857261
transform 1 0 182133 0 1 142311
box 0 0 1 1
use contact_7  contact_7_935
timestamp 1624857261
transform 1 0 182469 0 1 142311
box 0 0 1 1
use contact_7  contact_7_934
timestamp 1624857261
transform 1 0 182805 0 1 142311
box 0 0 1 1
use contact_7  contact_7_933
timestamp 1624857261
transform 1 0 183141 0 1 142311
box 0 0 1 1
use contact_7  contact_7_932
timestamp 1624857261
transform 1 0 183477 0 1 142311
box 0 0 1 1
use contact_7  contact_7_931
timestamp 1624857261
transform 1 0 183813 0 1 142311
box 0 0 1 1
use contact_7  contact_7_930
timestamp 1624857261
transform 1 0 184149 0 1 142311
box 0 0 1 1
use contact_7  contact_7_929
timestamp 1624857261
transform 1 0 184485 0 1 142311
box 0 0 1 1
use contact_7  contact_7_928
timestamp 1624857261
transform 1 0 184821 0 1 142311
box 0 0 1 1
use contact_7  contact_7_927
timestamp 1624857261
transform 1 0 185157 0 1 142311
box 0 0 1 1
use contact_7  contact_7_926
timestamp 1624857261
transform 1 0 185493 0 1 142311
box 0 0 1 1
use contact_7  contact_7_925
timestamp 1624857261
transform 1 0 185829 0 1 142311
box 0 0 1 1
use contact_7  contact_7_924
timestamp 1624857261
transform 1 0 186165 0 1 142311
box 0 0 1 1
use contact_7  contact_7_923
timestamp 1624857261
transform 1 0 186501 0 1 142311
box 0 0 1 1
use contact_7  contact_7_922
timestamp 1624857261
transform 1 0 186837 0 1 142311
box 0 0 1 1
use contact_7  contact_7_921
timestamp 1624857261
transform 1 0 187173 0 1 142311
box 0 0 1 1
use contact_7  contact_7_920
timestamp 1624857261
transform 1 0 187509 0 1 142311
box 0 0 1 1
use contact_7  contact_7_919
timestamp 1624857261
transform 1 0 187845 0 1 142311
box 0 0 1 1
use contact_7  contact_7_918
timestamp 1624857261
transform 1 0 188181 0 1 142311
box 0 0 1 1
use contact_7  contact_7_917
timestamp 1624857261
transform 1 0 188517 0 1 142311
box 0 0 1 1
use contact_7  contact_7_916
timestamp 1624857261
transform 1 0 188853 0 1 142311
box 0 0 1 1
use contact_7  contact_7_915
timestamp 1624857261
transform 1 0 189189 0 1 142311
box 0 0 1 1
use contact_7  contact_7_914
timestamp 1624857261
transform 1 0 189525 0 1 142311
box 0 0 1 1
use contact_7  contact_7_913
timestamp 1624857261
transform 1 0 189861 0 1 142311
box 0 0 1 1
use contact_7  contact_7_912
timestamp 1624857261
transform 1 0 190197 0 1 142311
box 0 0 1 1
use contact_7  contact_7_911
timestamp 1624857261
transform 1 0 190533 0 1 142311
box 0 0 1 1
use contact_7  contact_7_910
timestamp 1624857261
transform 1 0 190869 0 1 142311
box 0 0 1 1
use contact_7  contact_7_909
timestamp 1624857261
transform 1 0 191205 0 1 142311
box 0 0 1 1
use contact_7  contact_7_908
timestamp 1624857261
transform 1 0 191541 0 1 142311
box 0 0 1 1
use contact_7  contact_7_907
timestamp 1624857261
transform 1 0 191877 0 1 142311
box 0 0 1 1
use contact_7  contact_7_906
timestamp 1624857261
transform 1 0 192213 0 1 142311
box 0 0 1 1
use contact_7  contact_7_905
timestamp 1624857261
transform 1 0 192549 0 1 142311
box 0 0 1 1
use contact_7  contact_7_904
timestamp 1624857261
transform 1 0 192885 0 1 142311
box 0 0 1 1
use contact_7  contact_7_903
timestamp 1624857261
transform 1 0 193221 0 1 142311
box 0 0 1 1
use contact_7  contact_7_902
timestamp 1624857261
transform 1 0 193557 0 1 142311
box 0 0 1 1
use contact_7  contact_7_901
timestamp 1624857261
transform 1 0 193893 0 1 142311
box 0 0 1 1
use contact_7  contact_7_900
timestamp 1624857261
transform 1 0 194229 0 1 142311
box 0 0 1 1
use contact_7  contact_7_899
timestamp 1624857261
transform 1 0 194565 0 1 142311
box 0 0 1 1
use contact_7  contact_7_898
timestamp 1624857261
transform 1 0 194901 0 1 142311
box 0 0 1 1
use contact_7  contact_7_897
timestamp 1624857261
transform 1 0 195237 0 1 142311
box 0 0 1 1
use contact_7  contact_7_896
timestamp 1624857261
transform 1 0 195573 0 1 142311
box 0 0 1 1
use contact_7  contact_7_895
timestamp 1624857261
transform 1 0 195909 0 1 142311
box 0 0 1 1
use contact_7  contact_7_894
timestamp 1624857261
transform 1 0 196245 0 1 142311
box 0 0 1 1
use contact_7  contact_7_893
timestamp 1624857261
transform 1 0 196581 0 1 142311
box 0 0 1 1
use contact_7  contact_7_892
timestamp 1624857261
transform 1 0 196917 0 1 142311
box 0 0 1 1
use contact_7  contact_7_891
timestamp 1624857261
transform 1 0 197253 0 1 142311
box 0 0 1 1
use contact_7  contact_7_890
timestamp 1624857261
transform 1 0 197589 0 1 142311
box 0 0 1 1
use contact_7  contact_7_889
timestamp 1624857261
transform 1 0 197925 0 1 142311
box 0 0 1 1
use contact_7  contact_7_888
timestamp 1624857261
transform 1 0 198261 0 1 142311
box 0 0 1 1
use contact_7  contact_7_887
timestamp 1624857261
transform 1 0 198597 0 1 142311
box 0 0 1 1
use contact_7  contact_7_886
timestamp 1624857261
transform 1 0 198933 0 1 142311
box 0 0 1 1
use contact_7  contact_7_885
timestamp 1624857261
transform 1 0 199269 0 1 142311
box 0 0 1 1
use contact_7  contact_7_884
timestamp 1624857261
transform 1 0 199605 0 1 142311
box 0 0 1 1
use contact_7  contact_7_883
timestamp 1624857261
transform 1 0 199941 0 1 142311
box 0 0 1 1
use contact_7  contact_7_882
timestamp 1624857261
transform 1 0 200277 0 1 142311
box 0 0 1 1
use contact_7  contact_7_881
timestamp 1624857261
transform 1 0 200613 0 1 142311
box 0 0 1 1
use contact_7  contact_7_880
timestamp 1624857261
transform 1 0 200949 0 1 142311
box 0 0 1 1
use contact_7  contact_7_879
timestamp 1624857261
transform 1 0 201285 0 1 142311
box 0 0 1 1
use contact_7  contact_7_878
timestamp 1624857261
transform 1 0 201621 0 1 142311
box 0 0 1 1
use contact_7  contact_7_877
timestamp 1624857261
transform 1 0 201957 0 1 142311
box 0 0 1 1
use contact_7  contact_7_876
timestamp 1624857261
transform 1 0 202293 0 1 142311
box 0 0 1 1
use contact_7  contact_7_875
timestamp 1624857261
transform 1 0 202629 0 1 142311
box 0 0 1 1
use contact_7  contact_7_874
timestamp 1624857261
transform 1 0 202965 0 1 142311
box 0 0 1 1
use contact_7  contact_7_873
timestamp 1624857261
transform 1 0 203301 0 1 142311
box 0 0 1 1
use contact_7  contact_7_872
timestamp 1624857261
transform 1 0 203637 0 1 142311
box 0 0 1 1
use contact_7  contact_7_871
timestamp 1624857261
transform 1 0 203973 0 1 142311
box 0 0 1 1
use contact_7  contact_7_870
timestamp 1624857261
transform 1 0 204309 0 1 142311
box 0 0 1 1
use contact_7  contact_7_869
timestamp 1624857261
transform 1 0 204645 0 1 142311
box 0 0 1 1
use contact_7  contact_7_868
timestamp 1624857261
transform 1 0 204981 0 1 142311
box 0 0 1 1
use contact_7  contact_7_867
timestamp 1624857261
transform 1 0 205317 0 1 142311
box 0 0 1 1
use contact_7  contact_7_866
timestamp 1624857261
transform 1 0 205653 0 1 142311
box 0 0 1 1
use contact_7  contact_7_865
timestamp 1624857261
transform 1 0 205989 0 1 142311
box 0 0 1 1
use contact_7  contact_7_864
timestamp 1624857261
transform 1 0 206325 0 1 142311
box 0 0 1 1
use contact_7  contact_7_863
timestamp 1624857261
transform 1 0 206661 0 1 142311
box 0 0 1 1
use contact_7  contact_7_862
timestamp 1624857261
transform 1 0 206997 0 1 142311
box 0 0 1 1
use contact_7  contact_7_861
timestamp 1624857261
transform 1 0 207333 0 1 142311
box 0 0 1 1
use contact_7  contact_7_860
timestamp 1624857261
transform 1 0 207669 0 1 142311
box 0 0 1 1
use contact_7  contact_7_859
timestamp 1624857261
transform 1 0 208005 0 1 142311
box 0 0 1 1
use contact_7  contact_7_858
timestamp 1624857261
transform 1 0 208341 0 1 142311
box 0 0 1 1
use contact_7  contact_7_857
timestamp 1624857261
transform 1 0 208677 0 1 142311
box 0 0 1 1
use contact_7  contact_7_856
timestamp 1624857261
transform 1 0 209013 0 1 142311
box 0 0 1 1
use contact_7  contact_7_855
timestamp 1624857261
transform 1 0 209349 0 1 142311
box 0 0 1 1
use contact_7  contact_7_854
timestamp 1624857261
transform 1 0 209685 0 1 142311
box 0 0 1 1
use contact_7  contact_7_853
timestamp 1624857261
transform 1 0 210021 0 1 142311
box 0 0 1 1
use contact_7  contact_7_852
timestamp 1624857261
transform 1 0 210357 0 1 142311
box 0 0 1 1
use contact_7  contact_7_851
timestamp 1624857261
transform 1 0 210693 0 1 142311
box 0 0 1 1
use contact_7  contact_7_850
timestamp 1624857261
transform 1 0 211029 0 1 142311
box 0 0 1 1
use contact_7  contact_7_849
timestamp 1624857261
transform 1 0 211365 0 1 142311
box 0 0 1 1
use contact_7  contact_7_848
timestamp 1624857261
transform 1 0 211701 0 1 142311
box 0 0 1 1
use contact_7  contact_7_847
timestamp 1624857261
transform 1 0 212037 0 1 142311
box 0 0 1 1
use contact_7  contact_7_846
timestamp 1624857261
transform 1 0 212373 0 1 142311
box 0 0 1 1
use contact_7  contact_7_845
timestamp 1624857261
transform 1 0 212709 0 1 142311
box 0 0 1 1
use contact_7  contact_7_844
timestamp 1624857261
transform 1 0 213045 0 1 142311
box 0 0 1 1
use contact_7  contact_7_843
timestamp 1624857261
transform 1 0 213381 0 1 142311
box 0 0 1 1
use contact_7  contact_7_842
timestamp 1624857261
transform 1 0 213717 0 1 142311
box 0 0 1 1
use contact_7  contact_7_841
timestamp 1624857261
transform 1 0 214053 0 1 142311
box 0 0 1 1
use contact_7  contact_7_840
timestamp 1624857261
transform 1 0 214389 0 1 142311
box 0 0 1 1
use contact_7  contact_7_839
timestamp 1624857261
transform 1 0 214725 0 1 142311
box 0 0 1 1
use contact_7  contact_7_838
timestamp 1624857261
transform 1 0 215061 0 1 142311
box 0 0 1 1
use contact_7  contact_7_837
timestamp 1624857261
transform 1 0 215397 0 1 142311
box 0 0 1 1
use contact_7  contact_7_836
timestamp 1624857261
transform 1 0 215733 0 1 142311
box 0 0 1 1
use contact_7  contact_7_835
timestamp 1624857261
transform 1 0 216069 0 1 142311
box 0 0 1 1
use contact_7  contact_7_834
timestamp 1624857261
transform 1 0 216405 0 1 142311
box 0 0 1 1
use contact_7  contact_7_833
timestamp 1624857261
transform 1 0 1701 0 1 2151
box 0 0 1 1
use contact_7  contact_7_832
timestamp 1624857261
transform 1 0 1701 0 1 2487
box 0 0 1 1
use contact_7  contact_7_831
timestamp 1624857261
transform 1 0 1701 0 1 2823
box 0 0 1 1
use contact_7  contact_7_830
timestamp 1624857261
transform 1 0 1701 0 1 3159
box 0 0 1 1
use contact_7  contact_7_829
timestamp 1624857261
transform 1 0 1701 0 1 3495
box 0 0 1 1
use contact_7  contact_7_828
timestamp 1624857261
transform 1 0 1701 0 1 3831
box 0 0 1 1
use contact_7  contact_7_827
timestamp 1624857261
transform 1 0 1701 0 1 4167
box 0 0 1 1
use contact_7  contact_7_826
timestamp 1624857261
transform 1 0 1701 0 1 4503
box 0 0 1 1
use contact_7  contact_7_825
timestamp 1624857261
transform 1 0 1701 0 1 4839
box 0 0 1 1
use contact_7  contact_7_824
timestamp 1624857261
transform 1 0 1701 0 1 5175
box 0 0 1 1
use contact_7  contact_7_823
timestamp 1624857261
transform 1 0 1701 0 1 5511
box 0 0 1 1
use contact_7  contact_7_822
timestamp 1624857261
transform 1 0 1701 0 1 5847
box 0 0 1 1
use contact_7  contact_7_821
timestamp 1624857261
transform 1 0 1701 0 1 6183
box 0 0 1 1
use contact_7  contact_7_820
timestamp 1624857261
transform 1 0 1701 0 1 6519
box 0 0 1 1
use contact_7  contact_7_819
timestamp 1624857261
transform 1 0 1701 0 1 6855
box 0 0 1 1
use contact_7  contact_7_818
timestamp 1624857261
transform 1 0 1701 0 1 7191
box 0 0 1 1
use contact_7  contact_7_817
timestamp 1624857261
transform 1 0 1701 0 1 7527
box 0 0 1 1
use contact_7  contact_7_816
timestamp 1624857261
transform 1 0 1701 0 1 7863
box 0 0 1 1
use contact_7  contact_7_815
timestamp 1624857261
transform 1 0 1701 0 1 8199
box 0 0 1 1
use contact_7  contact_7_814
timestamp 1624857261
transform 1 0 1701 0 1 8535
box 0 0 1 1
use contact_7  contact_7_813
timestamp 1624857261
transform 1 0 1701 0 1 8871
box 0 0 1 1
use contact_7  contact_7_812
timestamp 1624857261
transform 1 0 1701 0 1 9207
box 0 0 1 1
use contact_7  contact_7_811
timestamp 1624857261
transform 1 0 1701 0 1 9543
box 0 0 1 1
use contact_7  contact_7_810
timestamp 1624857261
transform 1 0 1701 0 1 9879
box 0 0 1 1
use contact_7  contact_7_809
timestamp 1624857261
transform 1 0 1701 0 1 10215
box 0 0 1 1
use contact_7  contact_7_808
timestamp 1624857261
transform 1 0 1701 0 1 10551
box 0 0 1 1
use contact_7  contact_7_807
timestamp 1624857261
transform 1 0 1701 0 1 10887
box 0 0 1 1
use contact_7  contact_7_806
timestamp 1624857261
transform 1 0 1701 0 1 11223
box 0 0 1 1
use contact_7  contact_7_805
timestamp 1624857261
transform 1 0 1701 0 1 11559
box 0 0 1 1
use contact_7  contact_7_804
timestamp 1624857261
transform 1 0 1701 0 1 11895
box 0 0 1 1
use contact_7  contact_7_803
timestamp 1624857261
transform 1 0 1701 0 1 12231
box 0 0 1 1
use contact_7  contact_7_802
timestamp 1624857261
transform 1 0 1701 0 1 12567
box 0 0 1 1
use contact_7  contact_7_801
timestamp 1624857261
transform 1 0 1701 0 1 12903
box 0 0 1 1
use contact_7  contact_7_800
timestamp 1624857261
transform 1 0 1701 0 1 13239
box 0 0 1 1
use contact_7  contact_7_799
timestamp 1624857261
transform 1 0 1701 0 1 13575
box 0 0 1 1
use contact_7  contact_7_798
timestamp 1624857261
transform 1 0 1701 0 1 13911
box 0 0 1 1
use contact_7  contact_7_797
timestamp 1624857261
transform 1 0 1701 0 1 14247
box 0 0 1 1
use contact_7  contact_7_796
timestamp 1624857261
transform 1 0 1701 0 1 14583
box 0 0 1 1
use contact_7  contact_7_795
timestamp 1624857261
transform 1 0 1701 0 1 14919
box 0 0 1 1
use contact_7  contact_7_794
timestamp 1624857261
transform 1 0 1701 0 1 15255
box 0 0 1 1
use contact_7  contact_7_793
timestamp 1624857261
transform 1 0 1701 0 1 15591
box 0 0 1 1
use contact_7  contact_7_792
timestamp 1624857261
transform 1 0 1701 0 1 15927
box 0 0 1 1
use contact_7  contact_7_791
timestamp 1624857261
transform 1 0 1701 0 1 16263
box 0 0 1 1
use contact_7  contact_7_790
timestamp 1624857261
transform 1 0 1701 0 1 16599
box 0 0 1 1
use contact_7  contact_7_789
timestamp 1624857261
transform 1 0 1701 0 1 16935
box 0 0 1 1
use contact_7  contact_7_788
timestamp 1624857261
transform 1 0 1701 0 1 17271
box 0 0 1 1
use contact_7  contact_7_787
timestamp 1624857261
transform 1 0 1701 0 1 17607
box 0 0 1 1
use contact_7  contact_7_786
timestamp 1624857261
transform 1 0 1701 0 1 17943
box 0 0 1 1
use contact_7  contact_7_785
timestamp 1624857261
transform 1 0 1701 0 1 18279
box 0 0 1 1
use contact_7  contact_7_784
timestamp 1624857261
transform 1 0 1701 0 1 18615
box 0 0 1 1
use contact_7  contact_7_783
timestamp 1624857261
transform 1 0 1701 0 1 18951
box 0 0 1 1
use contact_7  contact_7_782
timestamp 1624857261
transform 1 0 1701 0 1 19287
box 0 0 1 1
use contact_7  contact_7_781
timestamp 1624857261
transform 1 0 1701 0 1 19623
box 0 0 1 1
use contact_7  contact_7_780
timestamp 1624857261
transform 1 0 1701 0 1 19959
box 0 0 1 1
use contact_7  contact_7_779
timestamp 1624857261
transform 1 0 1701 0 1 20295
box 0 0 1 1
use contact_7  contact_7_778
timestamp 1624857261
transform 1 0 1701 0 1 20631
box 0 0 1 1
use contact_7  contact_7_777
timestamp 1624857261
transform 1 0 1701 0 1 20967
box 0 0 1 1
use contact_7  contact_7_776
timestamp 1624857261
transform 1 0 1701 0 1 21303
box 0 0 1 1
use contact_7  contact_7_775
timestamp 1624857261
transform 1 0 1701 0 1 21639
box 0 0 1 1
use contact_7  contact_7_774
timestamp 1624857261
transform 1 0 1701 0 1 21975
box 0 0 1 1
use contact_7  contact_7_773
timestamp 1624857261
transform 1 0 1701 0 1 22311
box 0 0 1 1
use contact_7  contact_7_772
timestamp 1624857261
transform 1 0 1701 0 1 22647
box 0 0 1 1
use contact_7  contact_7_771
timestamp 1624857261
transform 1 0 1701 0 1 22983
box 0 0 1 1
use contact_7  contact_7_770
timestamp 1624857261
transform 1 0 1701 0 1 23319
box 0 0 1 1
use contact_7  contact_7_769
timestamp 1624857261
transform 1 0 1701 0 1 23655
box 0 0 1 1
use contact_7  contact_7_768
timestamp 1624857261
transform 1 0 1701 0 1 23991
box 0 0 1 1
use contact_7  contact_7_767
timestamp 1624857261
transform 1 0 1701 0 1 24327
box 0 0 1 1
use contact_7  contact_7_766
timestamp 1624857261
transform 1 0 1701 0 1 24663
box 0 0 1 1
use contact_7  contact_7_765
timestamp 1624857261
transform 1 0 1701 0 1 24999
box 0 0 1 1
use contact_7  contact_7_764
timestamp 1624857261
transform 1 0 1701 0 1 25335
box 0 0 1 1
use contact_7  contact_7_763
timestamp 1624857261
transform 1 0 1701 0 1 25671
box 0 0 1 1
use contact_7  contact_7_762
timestamp 1624857261
transform 1 0 1701 0 1 26007
box 0 0 1 1
use contact_7  contact_7_761
timestamp 1624857261
transform 1 0 1701 0 1 26343
box 0 0 1 1
use contact_7  contact_7_760
timestamp 1624857261
transform 1 0 1701 0 1 26679
box 0 0 1 1
use contact_7  contact_7_759
timestamp 1624857261
transform 1 0 1701 0 1 27015
box 0 0 1 1
use contact_7  contact_7_758
timestamp 1624857261
transform 1 0 1701 0 1 27351
box 0 0 1 1
use contact_7  contact_7_757
timestamp 1624857261
transform 1 0 1701 0 1 27687
box 0 0 1 1
use contact_7  contact_7_756
timestamp 1624857261
transform 1 0 1701 0 1 28023
box 0 0 1 1
use contact_7  contact_7_755
timestamp 1624857261
transform 1 0 1701 0 1 28359
box 0 0 1 1
use contact_7  contact_7_754
timestamp 1624857261
transform 1 0 1701 0 1 28695
box 0 0 1 1
use contact_7  contact_7_753
timestamp 1624857261
transform 1 0 1701 0 1 29031
box 0 0 1 1
use contact_7  contact_7_752
timestamp 1624857261
transform 1 0 1701 0 1 29367
box 0 0 1 1
use contact_7  contact_7_751
timestamp 1624857261
transform 1 0 1701 0 1 29703
box 0 0 1 1
use contact_7  contact_7_750
timestamp 1624857261
transform 1 0 1701 0 1 30039
box 0 0 1 1
use contact_7  contact_7_749
timestamp 1624857261
transform 1 0 1701 0 1 30375
box 0 0 1 1
use contact_7  contact_7_748
timestamp 1624857261
transform 1 0 1701 0 1 30711
box 0 0 1 1
use contact_7  contact_7_747
timestamp 1624857261
transform 1 0 1701 0 1 31047
box 0 0 1 1
use contact_7  contact_7_746
timestamp 1624857261
transform 1 0 1701 0 1 31383
box 0 0 1 1
use contact_7  contact_7_745
timestamp 1624857261
transform 1 0 1701 0 1 31719
box 0 0 1 1
use contact_7  contact_7_744
timestamp 1624857261
transform 1 0 1701 0 1 32055
box 0 0 1 1
use contact_7  contact_7_743
timestamp 1624857261
transform 1 0 1701 0 1 32391
box 0 0 1 1
use contact_7  contact_7_742
timestamp 1624857261
transform 1 0 1701 0 1 32727
box 0 0 1 1
use contact_7  contact_7_741
timestamp 1624857261
transform 1 0 1701 0 1 33063
box 0 0 1 1
use contact_7  contact_7_740
timestamp 1624857261
transform 1 0 1701 0 1 33399
box 0 0 1 1
use contact_7  contact_7_739
timestamp 1624857261
transform 1 0 1701 0 1 33735
box 0 0 1 1
use contact_7  contact_7_738
timestamp 1624857261
transform 1 0 1701 0 1 34071
box 0 0 1 1
use contact_7  contact_7_737
timestamp 1624857261
transform 1 0 1701 0 1 34407
box 0 0 1 1
use contact_7  contact_7_736
timestamp 1624857261
transform 1 0 1701 0 1 34743
box 0 0 1 1
use contact_7  contact_7_735
timestamp 1624857261
transform 1 0 1701 0 1 35079
box 0 0 1 1
use contact_7  contact_7_734
timestamp 1624857261
transform 1 0 1701 0 1 35415
box 0 0 1 1
use contact_7  contact_7_733
timestamp 1624857261
transform 1 0 1701 0 1 35751
box 0 0 1 1
use contact_7  contact_7_732
timestamp 1624857261
transform 1 0 1701 0 1 36087
box 0 0 1 1
use contact_7  contact_7_731
timestamp 1624857261
transform 1 0 1701 0 1 36423
box 0 0 1 1
use contact_7  contact_7_730
timestamp 1624857261
transform 1 0 1701 0 1 36759
box 0 0 1 1
use contact_7  contact_7_729
timestamp 1624857261
transform 1 0 1701 0 1 37095
box 0 0 1 1
use contact_7  contact_7_728
timestamp 1624857261
transform 1 0 1701 0 1 37431
box 0 0 1 1
use contact_7  contact_7_727
timestamp 1624857261
transform 1 0 1701 0 1 37767
box 0 0 1 1
use contact_7  contact_7_726
timestamp 1624857261
transform 1 0 1701 0 1 38103
box 0 0 1 1
use contact_7  contact_7_725
timestamp 1624857261
transform 1 0 1701 0 1 38439
box 0 0 1 1
use contact_7  contact_7_724
timestamp 1624857261
transform 1 0 1701 0 1 38775
box 0 0 1 1
use contact_7  contact_7_723
timestamp 1624857261
transform 1 0 1701 0 1 39111
box 0 0 1 1
use contact_7  contact_7_722
timestamp 1624857261
transform 1 0 1701 0 1 39447
box 0 0 1 1
use contact_7  contact_7_721
timestamp 1624857261
transform 1 0 1701 0 1 39783
box 0 0 1 1
use contact_7  contact_7_720
timestamp 1624857261
transform 1 0 1701 0 1 40119
box 0 0 1 1
use contact_7  contact_7_719
timestamp 1624857261
transform 1 0 1701 0 1 40455
box 0 0 1 1
use contact_7  contact_7_718
timestamp 1624857261
transform 1 0 1701 0 1 40791
box 0 0 1 1
use contact_7  contact_7_717
timestamp 1624857261
transform 1 0 1701 0 1 41127
box 0 0 1 1
use contact_7  contact_7_716
timestamp 1624857261
transform 1 0 1701 0 1 41463
box 0 0 1 1
use contact_7  contact_7_715
timestamp 1624857261
transform 1 0 1701 0 1 41799
box 0 0 1 1
use contact_7  contact_7_714
timestamp 1624857261
transform 1 0 1701 0 1 42135
box 0 0 1 1
use contact_7  contact_7_713
timestamp 1624857261
transform 1 0 1701 0 1 42471
box 0 0 1 1
use contact_7  contact_7_712
timestamp 1624857261
transform 1 0 1701 0 1 42807
box 0 0 1 1
use contact_7  contact_7_711
timestamp 1624857261
transform 1 0 1701 0 1 43143
box 0 0 1 1
use contact_7  contact_7_710
timestamp 1624857261
transform 1 0 1701 0 1 43479
box 0 0 1 1
use contact_7  contact_7_709
timestamp 1624857261
transform 1 0 1701 0 1 43815
box 0 0 1 1
use contact_7  contact_7_708
timestamp 1624857261
transform 1 0 1701 0 1 44151
box 0 0 1 1
use contact_7  contact_7_707
timestamp 1624857261
transform 1 0 1701 0 1 44487
box 0 0 1 1
use contact_7  contact_7_706
timestamp 1624857261
transform 1 0 1701 0 1 44823
box 0 0 1 1
use contact_7  contact_7_705
timestamp 1624857261
transform 1 0 1701 0 1 45159
box 0 0 1 1
use contact_7  contact_7_704
timestamp 1624857261
transform 1 0 1701 0 1 45495
box 0 0 1 1
use contact_7  contact_7_703
timestamp 1624857261
transform 1 0 1701 0 1 45831
box 0 0 1 1
use contact_7  contact_7_702
timestamp 1624857261
transform 1 0 1701 0 1 46167
box 0 0 1 1
use contact_7  contact_7_701
timestamp 1624857261
transform 1 0 1701 0 1 46503
box 0 0 1 1
use contact_7  contact_7_700
timestamp 1624857261
transform 1 0 1701 0 1 46839
box 0 0 1 1
use contact_7  contact_7_699
timestamp 1624857261
transform 1 0 1701 0 1 47175
box 0 0 1 1
use contact_7  contact_7_698
timestamp 1624857261
transform 1 0 1701 0 1 47511
box 0 0 1 1
use contact_7  contact_7_697
timestamp 1624857261
transform 1 0 1701 0 1 47847
box 0 0 1 1
use contact_7  contact_7_696
timestamp 1624857261
transform 1 0 1701 0 1 48183
box 0 0 1 1
use contact_7  contact_7_695
timestamp 1624857261
transform 1 0 1701 0 1 48519
box 0 0 1 1
use contact_7  contact_7_694
timestamp 1624857261
transform 1 0 1701 0 1 48855
box 0 0 1 1
use contact_7  contact_7_693
timestamp 1624857261
transform 1 0 1701 0 1 49191
box 0 0 1 1
use contact_7  contact_7_692
timestamp 1624857261
transform 1 0 1701 0 1 49527
box 0 0 1 1
use contact_7  contact_7_691
timestamp 1624857261
transform 1 0 1701 0 1 49863
box 0 0 1 1
use contact_7  contact_7_690
timestamp 1624857261
transform 1 0 1701 0 1 50199
box 0 0 1 1
use contact_7  contact_7_689
timestamp 1624857261
transform 1 0 1701 0 1 50535
box 0 0 1 1
use contact_7  contact_7_688
timestamp 1624857261
transform 1 0 1701 0 1 50871
box 0 0 1 1
use contact_7  contact_7_687
timestamp 1624857261
transform 1 0 1701 0 1 51207
box 0 0 1 1
use contact_7  contact_7_686
timestamp 1624857261
transform 1 0 1701 0 1 51543
box 0 0 1 1
use contact_7  contact_7_685
timestamp 1624857261
transform 1 0 1701 0 1 51879
box 0 0 1 1
use contact_7  contact_7_684
timestamp 1624857261
transform 1 0 1701 0 1 52215
box 0 0 1 1
use contact_7  contact_7_683
timestamp 1624857261
transform 1 0 1701 0 1 52551
box 0 0 1 1
use contact_7  contact_7_682
timestamp 1624857261
transform 1 0 1701 0 1 52887
box 0 0 1 1
use contact_7  contact_7_681
timestamp 1624857261
transform 1 0 1701 0 1 53223
box 0 0 1 1
use contact_7  contact_7_680
timestamp 1624857261
transform 1 0 1701 0 1 53559
box 0 0 1 1
use contact_7  contact_7_679
timestamp 1624857261
transform 1 0 1701 0 1 53895
box 0 0 1 1
use contact_7  contact_7_678
timestamp 1624857261
transform 1 0 1701 0 1 54231
box 0 0 1 1
use contact_7  contact_7_677
timestamp 1624857261
transform 1 0 1701 0 1 54567
box 0 0 1 1
use contact_7  contact_7_676
timestamp 1624857261
transform 1 0 1701 0 1 54903
box 0 0 1 1
use contact_7  contact_7_675
timestamp 1624857261
transform 1 0 1701 0 1 55239
box 0 0 1 1
use contact_7  contact_7_674
timestamp 1624857261
transform 1 0 1701 0 1 55575
box 0 0 1 1
use contact_7  contact_7_673
timestamp 1624857261
transform 1 0 1701 0 1 55911
box 0 0 1 1
use contact_7  contact_7_672
timestamp 1624857261
transform 1 0 1701 0 1 56247
box 0 0 1 1
use contact_7  contact_7_671
timestamp 1624857261
transform 1 0 1701 0 1 56583
box 0 0 1 1
use contact_7  contact_7_670
timestamp 1624857261
transform 1 0 1701 0 1 56919
box 0 0 1 1
use contact_7  contact_7_669
timestamp 1624857261
transform 1 0 1701 0 1 57255
box 0 0 1 1
use contact_7  contact_7_668
timestamp 1624857261
transform 1 0 1701 0 1 57591
box 0 0 1 1
use contact_7  contact_7_667
timestamp 1624857261
transform 1 0 1701 0 1 57927
box 0 0 1 1
use contact_7  contact_7_666
timestamp 1624857261
transform 1 0 1701 0 1 58263
box 0 0 1 1
use contact_7  contact_7_665
timestamp 1624857261
transform 1 0 1701 0 1 58599
box 0 0 1 1
use contact_7  contact_7_664
timestamp 1624857261
transform 1 0 1701 0 1 58935
box 0 0 1 1
use contact_7  contact_7_663
timestamp 1624857261
transform 1 0 1701 0 1 59271
box 0 0 1 1
use contact_7  contact_7_662
timestamp 1624857261
transform 1 0 1701 0 1 59607
box 0 0 1 1
use contact_7  contact_7_661
timestamp 1624857261
transform 1 0 1701 0 1 59943
box 0 0 1 1
use contact_7  contact_7_660
timestamp 1624857261
transform 1 0 1701 0 1 60279
box 0 0 1 1
use contact_7  contact_7_659
timestamp 1624857261
transform 1 0 1701 0 1 60615
box 0 0 1 1
use contact_7  contact_7_658
timestamp 1624857261
transform 1 0 1701 0 1 60951
box 0 0 1 1
use contact_7  contact_7_657
timestamp 1624857261
transform 1 0 1701 0 1 61287
box 0 0 1 1
use contact_7  contact_7_656
timestamp 1624857261
transform 1 0 1701 0 1 61623
box 0 0 1 1
use contact_7  contact_7_655
timestamp 1624857261
transform 1 0 1701 0 1 61959
box 0 0 1 1
use contact_7  contact_7_654
timestamp 1624857261
transform 1 0 1701 0 1 62295
box 0 0 1 1
use contact_7  contact_7_653
timestamp 1624857261
transform 1 0 1701 0 1 62631
box 0 0 1 1
use contact_7  contact_7_652
timestamp 1624857261
transform 1 0 1701 0 1 62967
box 0 0 1 1
use contact_7  contact_7_651
timestamp 1624857261
transform 1 0 1701 0 1 63303
box 0 0 1 1
use contact_7  contact_7_650
timestamp 1624857261
transform 1 0 1701 0 1 63639
box 0 0 1 1
use contact_7  contact_7_649
timestamp 1624857261
transform 1 0 1701 0 1 63975
box 0 0 1 1
use contact_7  contact_7_648
timestamp 1624857261
transform 1 0 1701 0 1 64311
box 0 0 1 1
use contact_7  contact_7_647
timestamp 1624857261
transform 1 0 1701 0 1 64647
box 0 0 1 1
use contact_7  contact_7_646
timestamp 1624857261
transform 1 0 1701 0 1 64983
box 0 0 1 1
use contact_7  contact_7_645
timestamp 1624857261
transform 1 0 1701 0 1 65319
box 0 0 1 1
use contact_7  contact_7_644
timestamp 1624857261
transform 1 0 1701 0 1 65655
box 0 0 1 1
use contact_7  contact_7_643
timestamp 1624857261
transform 1 0 1701 0 1 65991
box 0 0 1 1
use contact_7  contact_7_642
timestamp 1624857261
transform 1 0 1701 0 1 66327
box 0 0 1 1
use contact_7  contact_7_641
timestamp 1624857261
transform 1 0 1701 0 1 66663
box 0 0 1 1
use contact_7  contact_7_640
timestamp 1624857261
transform 1 0 1701 0 1 66999
box 0 0 1 1
use contact_7  contact_7_639
timestamp 1624857261
transform 1 0 1701 0 1 67335
box 0 0 1 1
use contact_7  contact_7_638
timestamp 1624857261
transform 1 0 1701 0 1 67671
box 0 0 1 1
use contact_7  contact_7_637
timestamp 1624857261
transform 1 0 1701 0 1 68007
box 0 0 1 1
use contact_7  contact_7_636
timestamp 1624857261
transform 1 0 1701 0 1 68343
box 0 0 1 1
use contact_7  contact_7_635
timestamp 1624857261
transform 1 0 1701 0 1 68679
box 0 0 1 1
use contact_7  contact_7_634
timestamp 1624857261
transform 1 0 1701 0 1 69015
box 0 0 1 1
use contact_7  contact_7_633
timestamp 1624857261
transform 1 0 1701 0 1 69351
box 0 0 1 1
use contact_7  contact_7_632
timestamp 1624857261
transform 1 0 1701 0 1 69687
box 0 0 1 1
use contact_7  contact_7_631
timestamp 1624857261
transform 1 0 1701 0 1 70023
box 0 0 1 1
use contact_7  contact_7_630
timestamp 1624857261
transform 1 0 1701 0 1 70359
box 0 0 1 1
use contact_7  contact_7_629
timestamp 1624857261
transform 1 0 1701 0 1 70695
box 0 0 1 1
use contact_7  contact_7_628
timestamp 1624857261
transform 1 0 1701 0 1 71031
box 0 0 1 1
use contact_7  contact_7_627
timestamp 1624857261
transform 1 0 1701 0 1 71367
box 0 0 1 1
use contact_7  contact_7_626
timestamp 1624857261
transform 1 0 1701 0 1 71703
box 0 0 1 1
use contact_7  contact_7_625
timestamp 1624857261
transform 1 0 1701 0 1 72039
box 0 0 1 1
use contact_7  contact_7_624
timestamp 1624857261
transform 1 0 1701 0 1 72375
box 0 0 1 1
use contact_7  contact_7_623
timestamp 1624857261
transform 1 0 1701 0 1 72711
box 0 0 1 1
use contact_7  contact_7_622
timestamp 1624857261
transform 1 0 1701 0 1 73047
box 0 0 1 1
use contact_7  contact_7_621
timestamp 1624857261
transform 1 0 1701 0 1 73383
box 0 0 1 1
use contact_7  contact_7_620
timestamp 1624857261
transform 1 0 1701 0 1 73719
box 0 0 1 1
use contact_7  contact_7_619
timestamp 1624857261
transform 1 0 1701 0 1 74055
box 0 0 1 1
use contact_7  contact_7_618
timestamp 1624857261
transform 1 0 1701 0 1 74391
box 0 0 1 1
use contact_7  contact_7_617
timestamp 1624857261
transform 1 0 1701 0 1 74727
box 0 0 1 1
use contact_7  contact_7_616
timestamp 1624857261
transform 1 0 1701 0 1 75063
box 0 0 1 1
use contact_7  contact_7_615
timestamp 1624857261
transform 1 0 1701 0 1 75399
box 0 0 1 1
use contact_7  contact_7_614
timestamp 1624857261
transform 1 0 1701 0 1 75735
box 0 0 1 1
use contact_7  contact_7_613
timestamp 1624857261
transform 1 0 1701 0 1 76071
box 0 0 1 1
use contact_7  contact_7_612
timestamp 1624857261
transform 1 0 1701 0 1 76407
box 0 0 1 1
use contact_7  contact_7_611
timestamp 1624857261
transform 1 0 1701 0 1 76743
box 0 0 1 1
use contact_7  contact_7_610
timestamp 1624857261
transform 1 0 1701 0 1 77079
box 0 0 1 1
use contact_7  contact_7_609
timestamp 1624857261
transform 1 0 1701 0 1 77415
box 0 0 1 1
use contact_7  contact_7_608
timestamp 1624857261
transform 1 0 1701 0 1 77751
box 0 0 1 1
use contact_7  contact_7_607
timestamp 1624857261
transform 1 0 1701 0 1 78087
box 0 0 1 1
use contact_7  contact_7_606
timestamp 1624857261
transform 1 0 1701 0 1 78423
box 0 0 1 1
use contact_7  contact_7_605
timestamp 1624857261
transform 1 0 1701 0 1 78759
box 0 0 1 1
use contact_7  contact_7_604
timestamp 1624857261
transform 1 0 1701 0 1 79095
box 0 0 1 1
use contact_7  contact_7_603
timestamp 1624857261
transform 1 0 1701 0 1 79431
box 0 0 1 1
use contact_7  contact_7_602
timestamp 1624857261
transform 1 0 1701 0 1 79767
box 0 0 1 1
use contact_7  contact_7_601
timestamp 1624857261
transform 1 0 1701 0 1 80103
box 0 0 1 1
use contact_7  contact_7_600
timestamp 1624857261
transform 1 0 1701 0 1 80439
box 0 0 1 1
use contact_7  contact_7_599
timestamp 1624857261
transform 1 0 1701 0 1 80775
box 0 0 1 1
use contact_7  contact_7_598
timestamp 1624857261
transform 1 0 1701 0 1 81111
box 0 0 1 1
use contact_7  contact_7_597
timestamp 1624857261
transform 1 0 1701 0 1 81447
box 0 0 1 1
use contact_7  contact_7_596
timestamp 1624857261
transform 1 0 1701 0 1 81783
box 0 0 1 1
use contact_7  contact_7_595
timestamp 1624857261
transform 1 0 1701 0 1 82119
box 0 0 1 1
use contact_7  contact_7_594
timestamp 1624857261
transform 1 0 1701 0 1 82455
box 0 0 1 1
use contact_7  contact_7_593
timestamp 1624857261
transform 1 0 1701 0 1 82791
box 0 0 1 1
use contact_7  contact_7_592
timestamp 1624857261
transform 1 0 1701 0 1 83127
box 0 0 1 1
use contact_7  contact_7_591
timestamp 1624857261
transform 1 0 1701 0 1 83463
box 0 0 1 1
use contact_7  contact_7_590
timestamp 1624857261
transform 1 0 1701 0 1 83799
box 0 0 1 1
use contact_7  contact_7_589
timestamp 1624857261
transform 1 0 1701 0 1 84135
box 0 0 1 1
use contact_7  contact_7_588
timestamp 1624857261
transform 1 0 1701 0 1 84471
box 0 0 1 1
use contact_7  contact_7_587
timestamp 1624857261
transform 1 0 1701 0 1 84807
box 0 0 1 1
use contact_7  contact_7_586
timestamp 1624857261
transform 1 0 1701 0 1 85143
box 0 0 1 1
use contact_7  contact_7_585
timestamp 1624857261
transform 1 0 1701 0 1 85479
box 0 0 1 1
use contact_7  contact_7_584
timestamp 1624857261
transform 1 0 1701 0 1 85815
box 0 0 1 1
use contact_7  contact_7_583
timestamp 1624857261
transform 1 0 1701 0 1 86151
box 0 0 1 1
use contact_7  contact_7_582
timestamp 1624857261
transform 1 0 1701 0 1 86487
box 0 0 1 1
use contact_7  contact_7_581
timestamp 1624857261
transform 1 0 1701 0 1 86823
box 0 0 1 1
use contact_7  contact_7_580
timestamp 1624857261
transform 1 0 1701 0 1 87159
box 0 0 1 1
use contact_7  contact_7_579
timestamp 1624857261
transform 1 0 1701 0 1 87495
box 0 0 1 1
use contact_7  contact_7_578
timestamp 1624857261
transform 1 0 1701 0 1 87831
box 0 0 1 1
use contact_7  contact_7_577
timestamp 1624857261
transform 1 0 1701 0 1 88167
box 0 0 1 1
use contact_7  contact_7_576
timestamp 1624857261
transform 1 0 1701 0 1 88503
box 0 0 1 1
use contact_7  contact_7_575
timestamp 1624857261
transform 1 0 1701 0 1 88839
box 0 0 1 1
use contact_7  contact_7_574
timestamp 1624857261
transform 1 0 1701 0 1 89175
box 0 0 1 1
use contact_7  contact_7_573
timestamp 1624857261
transform 1 0 1701 0 1 89511
box 0 0 1 1
use contact_7  contact_7_572
timestamp 1624857261
transform 1 0 1701 0 1 89847
box 0 0 1 1
use contact_7  contact_7_571
timestamp 1624857261
transform 1 0 1701 0 1 90183
box 0 0 1 1
use contact_7  contact_7_570
timestamp 1624857261
transform 1 0 1701 0 1 90519
box 0 0 1 1
use contact_7  contact_7_569
timestamp 1624857261
transform 1 0 1701 0 1 90855
box 0 0 1 1
use contact_7  contact_7_568
timestamp 1624857261
transform 1 0 1701 0 1 91191
box 0 0 1 1
use contact_7  contact_7_567
timestamp 1624857261
transform 1 0 1701 0 1 91527
box 0 0 1 1
use contact_7  contact_7_566
timestamp 1624857261
transform 1 0 1701 0 1 91863
box 0 0 1 1
use contact_7  contact_7_565
timestamp 1624857261
transform 1 0 1701 0 1 92199
box 0 0 1 1
use contact_7  contact_7_564
timestamp 1624857261
transform 1 0 1701 0 1 92535
box 0 0 1 1
use contact_7  contact_7_563
timestamp 1624857261
transform 1 0 1701 0 1 92871
box 0 0 1 1
use contact_7  contact_7_562
timestamp 1624857261
transform 1 0 1701 0 1 93207
box 0 0 1 1
use contact_7  contact_7_561
timestamp 1624857261
transform 1 0 1701 0 1 93543
box 0 0 1 1
use contact_7  contact_7_560
timestamp 1624857261
transform 1 0 1701 0 1 93879
box 0 0 1 1
use contact_7  contact_7_559
timestamp 1624857261
transform 1 0 1701 0 1 94215
box 0 0 1 1
use contact_7  contact_7_558
timestamp 1624857261
transform 1 0 1701 0 1 94551
box 0 0 1 1
use contact_7  contact_7_557
timestamp 1624857261
transform 1 0 1701 0 1 94887
box 0 0 1 1
use contact_7  contact_7_556
timestamp 1624857261
transform 1 0 1701 0 1 95223
box 0 0 1 1
use contact_7  contact_7_555
timestamp 1624857261
transform 1 0 1701 0 1 95559
box 0 0 1 1
use contact_7  contact_7_554
timestamp 1624857261
transform 1 0 1701 0 1 95895
box 0 0 1 1
use contact_7  contact_7_553
timestamp 1624857261
transform 1 0 1701 0 1 96231
box 0 0 1 1
use contact_7  contact_7_552
timestamp 1624857261
transform 1 0 1701 0 1 96567
box 0 0 1 1
use contact_7  contact_7_551
timestamp 1624857261
transform 1 0 1701 0 1 96903
box 0 0 1 1
use contact_7  contact_7_550
timestamp 1624857261
transform 1 0 1701 0 1 97239
box 0 0 1 1
use contact_7  contact_7_549
timestamp 1624857261
transform 1 0 1701 0 1 97575
box 0 0 1 1
use contact_7  contact_7_548
timestamp 1624857261
transform 1 0 1701 0 1 97911
box 0 0 1 1
use contact_7  contact_7_547
timestamp 1624857261
transform 1 0 1701 0 1 98247
box 0 0 1 1
use contact_7  contact_7_546
timestamp 1624857261
transform 1 0 1701 0 1 98583
box 0 0 1 1
use contact_7  contact_7_545
timestamp 1624857261
transform 1 0 1701 0 1 98919
box 0 0 1 1
use contact_7  contact_7_544
timestamp 1624857261
transform 1 0 1701 0 1 99255
box 0 0 1 1
use contact_7  contact_7_543
timestamp 1624857261
transform 1 0 1701 0 1 99591
box 0 0 1 1
use contact_7  contact_7_542
timestamp 1624857261
transform 1 0 1701 0 1 99927
box 0 0 1 1
use contact_7  contact_7_541
timestamp 1624857261
transform 1 0 1701 0 1 100263
box 0 0 1 1
use contact_7  contact_7_540
timestamp 1624857261
transform 1 0 1701 0 1 100599
box 0 0 1 1
use contact_7  contact_7_539
timestamp 1624857261
transform 1 0 1701 0 1 100935
box 0 0 1 1
use contact_7  contact_7_538
timestamp 1624857261
transform 1 0 1701 0 1 101271
box 0 0 1 1
use contact_7  contact_7_537
timestamp 1624857261
transform 1 0 1701 0 1 101607
box 0 0 1 1
use contact_7  contact_7_536
timestamp 1624857261
transform 1 0 1701 0 1 101943
box 0 0 1 1
use contact_7  contact_7_535
timestamp 1624857261
transform 1 0 1701 0 1 102279
box 0 0 1 1
use contact_7  contact_7_534
timestamp 1624857261
transform 1 0 1701 0 1 102615
box 0 0 1 1
use contact_7  contact_7_533
timestamp 1624857261
transform 1 0 1701 0 1 102951
box 0 0 1 1
use contact_7  contact_7_532
timestamp 1624857261
transform 1 0 1701 0 1 103287
box 0 0 1 1
use contact_7  contact_7_531
timestamp 1624857261
transform 1 0 1701 0 1 103623
box 0 0 1 1
use contact_7  contact_7_530
timestamp 1624857261
transform 1 0 1701 0 1 103959
box 0 0 1 1
use contact_7  contact_7_529
timestamp 1624857261
transform 1 0 1701 0 1 104295
box 0 0 1 1
use contact_7  contact_7_528
timestamp 1624857261
transform 1 0 1701 0 1 104631
box 0 0 1 1
use contact_7  contact_7_527
timestamp 1624857261
transform 1 0 1701 0 1 104967
box 0 0 1 1
use contact_7  contact_7_526
timestamp 1624857261
transform 1 0 1701 0 1 105303
box 0 0 1 1
use contact_7  contact_7_525
timestamp 1624857261
transform 1 0 1701 0 1 105639
box 0 0 1 1
use contact_7  contact_7_524
timestamp 1624857261
transform 1 0 1701 0 1 105975
box 0 0 1 1
use contact_7  contact_7_523
timestamp 1624857261
transform 1 0 1701 0 1 106311
box 0 0 1 1
use contact_7  contact_7_522
timestamp 1624857261
transform 1 0 1701 0 1 106647
box 0 0 1 1
use contact_7  contact_7_521
timestamp 1624857261
transform 1 0 1701 0 1 106983
box 0 0 1 1
use contact_7  contact_7_520
timestamp 1624857261
transform 1 0 1701 0 1 107319
box 0 0 1 1
use contact_7  contact_7_519
timestamp 1624857261
transform 1 0 1701 0 1 107655
box 0 0 1 1
use contact_7  contact_7_518
timestamp 1624857261
transform 1 0 1701 0 1 107991
box 0 0 1 1
use contact_7  contact_7_517
timestamp 1624857261
transform 1 0 1701 0 1 108327
box 0 0 1 1
use contact_7  contact_7_516
timestamp 1624857261
transform 1 0 1701 0 1 108663
box 0 0 1 1
use contact_7  contact_7_515
timestamp 1624857261
transform 1 0 1701 0 1 108999
box 0 0 1 1
use contact_7  contact_7_514
timestamp 1624857261
transform 1 0 1701 0 1 109335
box 0 0 1 1
use contact_7  contact_7_513
timestamp 1624857261
transform 1 0 1701 0 1 109671
box 0 0 1 1
use contact_7  contact_7_512
timestamp 1624857261
transform 1 0 1701 0 1 110007
box 0 0 1 1
use contact_7  contact_7_511
timestamp 1624857261
transform 1 0 1701 0 1 110343
box 0 0 1 1
use contact_7  contact_7_510
timestamp 1624857261
transform 1 0 1701 0 1 110679
box 0 0 1 1
use contact_7  contact_7_509
timestamp 1624857261
transform 1 0 1701 0 1 111015
box 0 0 1 1
use contact_7  contact_7_508
timestamp 1624857261
transform 1 0 1701 0 1 111351
box 0 0 1 1
use contact_7  contact_7_507
timestamp 1624857261
transform 1 0 1701 0 1 111687
box 0 0 1 1
use contact_7  contact_7_506
timestamp 1624857261
transform 1 0 1701 0 1 112023
box 0 0 1 1
use contact_7  contact_7_505
timestamp 1624857261
transform 1 0 1701 0 1 112359
box 0 0 1 1
use contact_7  contact_7_504
timestamp 1624857261
transform 1 0 1701 0 1 112695
box 0 0 1 1
use contact_7  contact_7_503
timestamp 1624857261
transform 1 0 1701 0 1 113031
box 0 0 1 1
use contact_7  contact_7_502
timestamp 1624857261
transform 1 0 1701 0 1 113367
box 0 0 1 1
use contact_7  contact_7_501
timestamp 1624857261
transform 1 0 1701 0 1 113703
box 0 0 1 1
use contact_7  contact_7_500
timestamp 1624857261
transform 1 0 1701 0 1 114039
box 0 0 1 1
use contact_7  contact_7_499
timestamp 1624857261
transform 1 0 1701 0 1 114375
box 0 0 1 1
use contact_7  contact_7_498
timestamp 1624857261
transform 1 0 1701 0 1 114711
box 0 0 1 1
use contact_7  contact_7_497
timestamp 1624857261
transform 1 0 1701 0 1 115047
box 0 0 1 1
use contact_7  contact_7_496
timestamp 1624857261
transform 1 0 1701 0 1 115383
box 0 0 1 1
use contact_7  contact_7_495
timestamp 1624857261
transform 1 0 1701 0 1 115719
box 0 0 1 1
use contact_7  contact_7_494
timestamp 1624857261
transform 1 0 1701 0 1 116055
box 0 0 1 1
use contact_7  contact_7_493
timestamp 1624857261
transform 1 0 1701 0 1 116391
box 0 0 1 1
use contact_7  contact_7_492
timestamp 1624857261
transform 1 0 1701 0 1 116727
box 0 0 1 1
use contact_7  contact_7_491
timestamp 1624857261
transform 1 0 1701 0 1 117063
box 0 0 1 1
use contact_7  contact_7_490
timestamp 1624857261
transform 1 0 1701 0 1 117399
box 0 0 1 1
use contact_7  contact_7_489
timestamp 1624857261
transform 1 0 1701 0 1 117735
box 0 0 1 1
use contact_7  contact_7_488
timestamp 1624857261
transform 1 0 1701 0 1 118071
box 0 0 1 1
use contact_7  contact_7_487
timestamp 1624857261
transform 1 0 1701 0 1 118407
box 0 0 1 1
use contact_7  contact_7_486
timestamp 1624857261
transform 1 0 1701 0 1 118743
box 0 0 1 1
use contact_7  contact_7_485
timestamp 1624857261
transform 1 0 1701 0 1 119079
box 0 0 1 1
use contact_7  contact_7_484
timestamp 1624857261
transform 1 0 1701 0 1 119415
box 0 0 1 1
use contact_7  contact_7_483
timestamp 1624857261
transform 1 0 1701 0 1 119751
box 0 0 1 1
use contact_7  contact_7_482
timestamp 1624857261
transform 1 0 1701 0 1 120087
box 0 0 1 1
use contact_7  contact_7_481
timestamp 1624857261
transform 1 0 1701 0 1 120423
box 0 0 1 1
use contact_7  contact_7_480
timestamp 1624857261
transform 1 0 1701 0 1 120759
box 0 0 1 1
use contact_7  contact_7_479
timestamp 1624857261
transform 1 0 1701 0 1 121095
box 0 0 1 1
use contact_7  contact_7_478
timestamp 1624857261
transform 1 0 1701 0 1 121431
box 0 0 1 1
use contact_7  contact_7_477
timestamp 1624857261
transform 1 0 1701 0 1 121767
box 0 0 1 1
use contact_7  contact_7_476
timestamp 1624857261
transform 1 0 1701 0 1 122103
box 0 0 1 1
use contact_7  contact_7_475
timestamp 1624857261
transform 1 0 1701 0 1 122439
box 0 0 1 1
use contact_7  contact_7_474
timestamp 1624857261
transform 1 0 1701 0 1 122775
box 0 0 1 1
use contact_7  contact_7_473
timestamp 1624857261
transform 1 0 1701 0 1 123111
box 0 0 1 1
use contact_7  contact_7_472
timestamp 1624857261
transform 1 0 1701 0 1 123447
box 0 0 1 1
use contact_7  contact_7_471
timestamp 1624857261
transform 1 0 1701 0 1 123783
box 0 0 1 1
use contact_7  contact_7_470
timestamp 1624857261
transform 1 0 1701 0 1 124119
box 0 0 1 1
use contact_7  contact_7_469
timestamp 1624857261
transform 1 0 1701 0 1 124455
box 0 0 1 1
use contact_7  contact_7_468
timestamp 1624857261
transform 1 0 1701 0 1 124791
box 0 0 1 1
use contact_7  contact_7_467
timestamp 1624857261
transform 1 0 1701 0 1 125127
box 0 0 1 1
use contact_7  contact_7_466
timestamp 1624857261
transform 1 0 1701 0 1 125463
box 0 0 1 1
use contact_7  contact_7_465
timestamp 1624857261
transform 1 0 1701 0 1 125799
box 0 0 1 1
use contact_7  contact_7_464
timestamp 1624857261
transform 1 0 1701 0 1 126135
box 0 0 1 1
use contact_7  contact_7_463
timestamp 1624857261
transform 1 0 1701 0 1 126471
box 0 0 1 1
use contact_7  contact_7_462
timestamp 1624857261
transform 1 0 1701 0 1 126807
box 0 0 1 1
use contact_7  contact_7_461
timestamp 1624857261
transform 1 0 1701 0 1 127143
box 0 0 1 1
use contact_7  contact_7_460
timestamp 1624857261
transform 1 0 1701 0 1 127479
box 0 0 1 1
use contact_7  contact_7_459
timestamp 1624857261
transform 1 0 1701 0 1 127815
box 0 0 1 1
use contact_7  contact_7_458
timestamp 1624857261
transform 1 0 1701 0 1 128151
box 0 0 1 1
use contact_7  contact_7_457
timestamp 1624857261
transform 1 0 1701 0 1 128487
box 0 0 1 1
use contact_7  contact_7_456
timestamp 1624857261
transform 1 0 1701 0 1 128823
box 0 0 1 1
use contact_7  contact_7_455
timestamp 1624857261
transform 1 0 1701 0 1 129159
box 0 0 1 1
use contact_7  contact_7_454
timestamp 1624857261
transform 1 0 1701 0 1 129495
box 0 0 1 1
use contact_7  contact_7_453
timestamp 1624857261
transform 1 0 1701 0 1 129831
box 0 0 1 1
use contact_7  contact_7_452
timestamp 1624857261
transform 1 0 1701 0 1 130167
box 0 0 1 1
use contact_7  contact_7_451
timestamp 1624857261
transform 1 0 1701 0 1 130503
box 0 0 1 1
use contact_7  contact_7_450
timestamp 1624857261
transform 1 0 1701 0 1 130839
box 0 0 1 1
use contact_7  contact_7_449
timestamp 1624857261
transform 1 0 1701 0 1 131175
box 0 0 1 1
use contact_7  contact_7_448
timestamp 1624857261
transform 1 0 1701 0 1 131511
box 0 0 1 1
use contact_7  contact_7_447
timestamp 1624857261
transform 1 0 1701 0 1 131847
box 0 0 1 1
use contact_7  contact_7_446
timestamp 1624857261
transform 1 0 1701 0 1 132183
box 0 0 1 1
use contact_7  contact_7_445
timestamp 1624857261
transform 1 0 1701 0 1 132519
box 0 0 1 1
use contact_7  contact_7_444
timestamp 1624857261
transform 1 0 1701 0 1 132855
box 0 0 1 1
use contact_7  contact_7_443
timestamp 1624857261
transform 1 0 1701 0 1 133191
box 0 0 1 1
use contact_7  contact_7_442
timestamp 1624857261
transform 1 0 1701 0 1 133527
box 0 0 1 1
use contact_7  contact_7_441
timestamp 1624857261
transform 1 0 1701 0 1 133863
box 0 0 1 1
use contact_7  contact_7_440
timestamp 1624857261
transform 1 0 1701 0 1 134199
box 0 0 1 1
use contact_7  contact_7_439
timestamp 1624857261
transform 1 0 1701 0 1 134535
box 0 0 1 1
use contact_7  contact_7_438
timestamp 1624857261
transform 1 0 1701 0 1 134871
box 0 0 1 1
use contact_7  contact_7_437
timestamp 1624857261
transform 1 0 1701 0 1 135207
box 0 0 1 1
use contact_7  contact_7_436
timestamp 1624857261
transform 1 0 1701 0 1 135543
box 0 0 1 1
use contact_7  contact_7_435
timestamp 1624857261
transform 1 0 1701 0 1 135879
box 0 0 1 1
use contact_7  contact_7_434
timestamp 1624857261
transform 1 0 1701 0 1 136215
box 0 0 1 1
use contact_7  contact_7_433
timestamp 1624857261
transform 1 0 1701 0 1 136551
box 0 0 1 1
use contact_7  contact_7_432
timestamp 1624857261
transform 1 0 1701 0 1 136887
box 0 0 1 1
use contact_7  contact_7_431
timestamp 1624857261
transform 1 0 1701 0 1 137223
box 0 0 1 1
use contact_7  contact_7_430
timestamp 1624857261
transform 1 0 1701 0 1 137559
box 0 0 1 1
use contact_7  contact_7_429
timestamp 1624857261
transform 1 0 1701 0 1 137895
box 0 0 1 1
use contact_7  contact_7_428
timestamp 1624857261
transform 1 0 1701 0 1 138231
box 0 0 1 1
use contact_7  contact_7_427
timestamp 1624857261
transform 1 0 1701 0 1 138567
box 0 0 1 1
use contact_7  contact_7_426
timestamp 1624857261
transform 1 0 1701 0 1 138903
box 0 0 1 1
use contact_7  contact_7_425
timestamp 1624857261
transform 1 0 1701 0 1 139239
box 0 0 1 1
use contact_7  contact_7_424
timestamp 1624857261
transform 1 0 1701 0 1 139575
box 0 0 1 1
use contact_7  contact_7_423
timestamp 1624857261
transform 1 0 1701 0 1 139911
box 0 0 1 1
use contact_7  contact_7_422
timestamp 1624857261
transform 1 0 1701 0 1 140247
box 0 0 1 1
use contact_7  contact_7_421
timestamp 1624857261
transform 1 0 1701 0 1 140583
box 0 0 1 1
use contact_7  contact_7_420
timestamp 1624857261
transform 1 0 1701 0 1 140919
box 0 0 1 1
use contact_7  contact_7_419
timestamp 1624857261
transform 1 0 1701 0 1 141255
box 0 0 1 1
use contact_7  contact_7_418
timestamp 1624857261
transform 1 0 1701 0 1 141591
box 0 0 1 1
use contact_7  contact_7_417
timestamp 1624857261
transform 1 0 1701 0 1 141927
box 0 0 1 1
use contact_7  contact_7_416
timestamp 1624857261
transform 1 0 216907 0 1 2151
box 0 0 1 1
use contact_7  contact_7_415
timestamp 1624857261
transform 1 0 216907 0 1 2487
box 0 0 1 1
use contact_7  contact_7_414
timestamp 1624857261
transform 1 0 216907 0 1 2823
box 0 0 1 1
use contact_7  contact_7_413
timestamp 1624857261
transform 1 0 216907 0 1 3159
box 0 0 1 1
use contact_7  contact_7_412
timestamp 1624857261
transform 1 0 216907 0 1 3495
box 0 0 1 1
use contact_7  contact_7_411
timestamp 1624857261
transform 1 0 216907 0 1 3831
box 0 0 1 1
use contact_7  contact_7_410
timestamp 1624857261
transform 1 0 216907 0 1 4167
box 0 0 1 1
use contact_7  contact_7_409
timestamp 1624857261
transform 1 0 216907 0 1 4503
box 0 0 1 1
use contact_7  contact_7_408
timestamp 1624857261
transform 1 0 216907 0 1 4839
box 0 0 1 1
use contact_7  contact_7_407
timestamp 1624857261
transform 1 0 216907 0 1 5175
box 0 0 1 1
use contact_7  contact_7_406
timestamp 1624857261
transform 1 0 216907 0 1 5511
box 0 0 1 1
use contact_7  contact_7_405
timestamp 1624857261
transform 1 0 216907 0 1 5847
box 0 0 1 1
use contact_7  contact_7_404
timestamp 1624857261
transform 1 0 216907 0 1 6183
box 0 0 1 1
use contact_7  contact_7_403
timestamp 1624857261
transform 1 0 216907 0 1 6519
box 0 0 1 1
use contact_7  contact_7_402
timestamp 1624857261
transform 1 0 216907 0 1 6855
box 0 0 1 1
use contact_7  contact_7_401
timestamp 1624857261
transform 1 0 216907 0 1 7191
box 0 0 1 1
use contact_7  contact_7_400
timestamp 1624857261
transform 1 0 216907 0 1 7527
box 0 0 1 1
use contact_7  contact_7_399
timestamp 1624857261
transform 1 0 216907 0 1 7863
box 0 0 1 1
use contact_7  contact_7_398
timestamp 1624857261
transform 1 0 216907 0 1 8199
box 0 0 1 1
use contact_7  contact_7_397
timestamp 1624857261
transform 1 0 216907 0 1 8535
box 0 0 1 1
use contact_7  contact_7_396
timestamp 1624857261
transform 1 0 216907 0 1 8871
box 0 0 1 1
use contact_7  contact_7_395
timestamp 1624857261
transform 1 0 216907 0 1 9207
box 0 0 1 1
use contact_7  contact_7_394
timestamp 1624857261
transform 1 0 216907 0 1 9543
box 0 0 1 1
use contact_7  contact_7_393
timestamp 1624857261
transform 1 0 216907 0 1 9879
box 0 0 1 1
use contact_7  contact_7_392
timestamp 1624857261
transform 1 0 216907 0 1 10215
box 0 0 1 1
use contact_7  contact_7_391
timestamp 1624857261
transform 1 0 216907 0 1 10551
box 0 0 1 1
use contact_7  contact_7_390
timestamp 1624857261
transform 1 0 216907 0 1 10887
box 0 0 1 1
use contact_7  contact_7_389
timestamp 1624857261
transform 1 0 216907 0 1 11223
box 0 0 1 1
use contact_7  contact_7_388
timestamp 1624857261
transform 1 0 216907 0 1 11559
box 0 0 1 1
use contact_7  contact_7_387
timestamp 1624857261
transform 1 0 216907 0 1 11895
box 0 0 1 1
use contact_7  contact_7_386
timestamp 1624857261
transform 1 0 216907 0 1 12231
box 0 0 1 1
use contact_7  contact_7_385
timestamp 1624857261
transform 1 0 216907 0 1 12567
box 0 0 1 1
use contact_7  contact_7_384
timestamp 1624857261
transform 1 0 216907 0 1 12903
box 0 0 1 1
use contact_7  contact_7_383
timestamp 1624857261
transform 1 0 216907 0 1 13239
box 0 0 1 1
use contact_7  contact_7_382
timestamp 1624857261
transform 1 0 216907 0 1 13575
box 0 0 1 1
use contact_7  contact_7_381
timestamp 1624857261
transform 1 0 216907 0 1 13911
box 0 0 1 1
use contact_7  contact_7_380
timestamp 1624857261
transform 1 0 216907 0 1 14247
box 0 0 1 1
use contact_7  contact_7_379
timestamp 1624857261
transform 1 0 216907 0 1 14583
box 0 0 1 1
use contact_7  contact_7_378
timestamp 1624857261
transform 1 0 216907 0 1 14919
box 0 0 1 1
use contact_7  contact_7_377
timestamp 1624857261
transform 1 0 216907 0 1 15255
box 0 0 1 1
use contact_7  contact_7_376
timestamp 1624857261
transform 1 0 216907 0 1 15591
box 0 0 1 1
use contact_7  contact_7_375
timestamp 1624857261
transform 1 0 216907 0 1 15927
box 0 0 1 1
use contact_7  contact_7_374
timestamp 1624857261
transform 1 0 216907 0 1 16263
box 0 0 1 1
use contact_7  contact_7_373
timestamp 1624857261
transform 1 0 216907 0 1 16599
box 0 0 1 1
use contact_7  contact_7_372
timestamp 1624857261
transform 1 0 216907 0 1 16935
box 0 0 1 1
use contact_7  contact_7_371
timestamp 1624857261
transform 1 0 216907 0 1 17271
box 0 0 1 1
use contact_7  contact_7_370
timestamp 1624857261
transform 1 0 216907 0 1 17607
box 0 0 1 1
use contact_7  contact_7_369
timestamp 1624857261
transform 1 0 216907 0 1 17943
box 0 0 1 1
use contact_7  contact_7_368
timestamp 1624857261
transform 1 0 216907 0 1 18279
box 0 0 1 1
use contact_7  contact_7_367
timestamp 1624857261
transform 1 0 216907 0 1 18615
box 0 0 1 1
use contact_7  contact_7_366
timestamp 1624857261
transform 1 0 216907 0 1 18951
box 0 0 1 1
use contact_7  contact_7_365
timestamp 1624857261
transform 1 0 216907 0 1 19287
box 0 0 1 1
use contact_7  contact_7_364
timestamp 1624857261
transform 1 0 216907 0 1 19623
box 0 0 1 1
use contact_7  contact_7_363
timestamp 1624857261
transform 1 0 216907 0 1 19959
box 0 0 1 1
use contact_7  contact_7_362
timestamp 1624857261
transform 1 0 216907 0 1 20295
box 0 0 1 1
use contact_7  contact_7_361
timestamp 1624857261
transform 1 0 216907 0 1 20631
box 0 0 1 1
use contact_7  contact_7_360
timestamp 1624857261
transform 1 0 216907 0 1 20967
box 0 0 1 1
use contact_7  contact_7_359
timestamp 1624857261
transform 1 0 216907 0 1 21303
box 0 0 1 1
use contact_7  contact_7_358
timestamp 1624857261
transform 1 0 216907 0 1 21639
box 0 0 1 1
use contact_7  contact_7_357
timestamp 1624857261
transform 1 0 216907 0 1 21975
box 0 0 1 1
use contact_7  contact_7_356
timestamp 1624857261
transform 1 0 216907 0 1 22311
box 0 0 1 1
use contact_7  contact_7_355
timestamp 1624857261
transform 1 0 216907 0 1 22647
box 0 0 1 1
use contact_7  contact_7_354
timestamp 1624857261
transform 1 0 216907 0 1 22983
box 0 0 1 1
use contact_7  contact_7_353
timestamp 1624857261
transform 1 0 216907 0 1 23319
box 0 0 1 1
use contact_7  contact_7_352
timestamp 1624857261
transform 1 0 216907 0 1 23655
box 0 0 1 1
use contact_7  contact_7_351
timestamp 1624857261
transform 1 0 216907 0 1 23991
box 0 0 1 1
use contact_7  contact_7_350
timestamp 1624857261
transform 1 0 216907 0 1 24327
box 0 0 1 1
use contact_7  contact_7_349
timestamp 1624857261
transform 1 0 216907 0 1 24663
box 0 0 1 1
use contact_7  contact_7_348
timestamp 1624857261
transform 1 0 216907 0 1 24999
box 0 0 1 1
use contact_7  contact_7_347
timestamp 1624857261
transform 1 0 216907 0 1 25335
box 0 0 1 1
use contact_7  contact_7_346
timestamp 1624857261
transform 1 0 216907 0 1 25671
box 0 0 1 1
use contact_7  contact_7_345
timestamp 1624857261
transform 1 0 216907 0 1 26007
box 0 0 1 1
use contact_7  contact_7_344
timestamp 1624857261
transform 1 0 216907 0 1 26343
box 0 0 1 1
use contact_7  contact_7_343
timestamp 1624857261
transform 1 0 216907 0 1 26679
box 0 0 1 1
use contact_7  contact_7_342
timestamp 1624857261
transform 1 0 216907 0 1 27015
box 0 0 1 1
use contact_7  contact_7_341
timestamp 1624857261
transform 1 0 216907 0 1 27351
box 0 0 1 1
use contact_7  contact_7_340
timestamp 1624857261
transform 1 0 216907 0 1 27687
box 0 0 1 1
use contact_7  contact_7_339
timestamp 1624857261
transform 1 0 216907 0 1 28023
box 0 0 1 1
use contact_7  contact_7_338
timestamp 1624857261
transform 1 0 216907 0 1 28359
box 0 0 1 1
use contact_7  contact_7_337
timestamp 1624857261
transform 1 0 216907 0 1 28695
box 0 0 1 1
use contact_7  contact_7_336
timestamp 1624857261
transform 1 0 216907 0 1 29031
box 0 0 1 1
use contact_7  contact_7_335
timestamp 1624857261
transform 1 0 216907 0 1 29367
box 0 0 1 1
use contact_7  contact_7_334
timestamp 1624857261
transform 1 0 216907 0 1 29703
box 0 0 1 1
use contact_7  contact_7_333
timestamp 1624857261
transform 1 0 216907 0 1 30039
box 0 0 1 1
use contact_7  contact_7_332
timestamp 1624857261
transform 1 0 216907 0 1 30375
box 0 0 1 1
use contact_7  contact_7_331
timestamp 1624857261
transform 1 0 216907 0 1 30711
box 0 0 1 1
use contact_7  contact_7_330
timestamp 1624857261
transform 1 0 216907 0 1 31047
box 0 0 1 1
use contact_7  contact_7_329
timestamp 1624857261
transform 1 0 216907 0 1 31383
box 0 0 1 1
use contact_7  contact_7_328
timestamp 1624857261
transform 1 0 216907 0 1 31719
box 0 0 1 1
use contact_7  contact_7_327
timestamp 1624857261
transform 1 0 216907 0 1 32055
box 0 0 1 1
use contact_7  contact_7_326
timestamp 1624857261
transform 1 0 216907 0 1 32391
box 0 0 1 1
use contact_7  contact_7_325
timestamp 1624857261
transform 1 0 216907 0 1 32727
box 0 0 1 1
use contact_7  contact_7_324
timestamp 1624857261
transform 1 0 216907 0 1 33063
box 0 0 1 1
use contact_7  contact_7_323
timestamp 1624857261
transform 1 0 216907 0 1 33399
box 0 0 1 1
use contact_7  contact_7_322
timestamp 1624857261
transform 1 0 216907 0 1 33735
box 0 0 1 1
use contact_7  contact_7_321
timestamp 1624857261
transform 1 0 216907 0 1 34071
box 0 0 1 1
use contact_7  contact_7_320
timestamp 1624857261
transform 1 0 216907 0 1 34407
box 0 0 1 1
use contact_7  contact_7_319
timestamp 1624857261
transform 1 0 216907 0 1 34743
box 0 0 1 1
use contact_7  contact_7_318
timestamp 1624857261
transform 1 0 216907 0 1 35079
box 0 0 1 1
use contact_7  contact_7_317
timestamp 1624857261
transform 1 0 216907 0 1 35415
box 0 0 1 1
use contact_7  contact_7_316
timestamp 1624857261
transform 1 0 216907 0 1 35751
box 0 0 1 1
use contact_7  contact_7_315
timestamp 1624857261
transform 1 0 216907 0 1 36087
box 0 0 1 1
use contact_7  contact_7_314
timestamp 1624857261
transform 1 0 216907 0 1 36423
box 0 0 1 1
use contact_7  contact_7_313
timestamp 1624857261
transform 1 0 216907 0 1 36759
box 0 0 1 1
use contact_7  contact_7_312
timestamp 1624857261
transform 1 0 216907 0 1 37095
box 0 0 1 1
use contact_7  contact_7_311
timestamp 1624857261
transform 1 0 216907 0 1 37431
box 0 0 1 1
use contact_7  contact_7_310
timestamp 1624857261
transform 1 0 216907 0 1 37767
box 0 0 1 1
use contact_7  contact_7_309
timestamp 1624857261
transform 1 0 216907 0 1 38103
box 0 0 1 1
use contact_7  contact_7_308
timestamp 1624857261
transform 1 0 216907 0 1 38439
box 0 0 1 1
use contact_7  contact_7_307
timestamp 1624857261
transform 1 0 216907 0 1 38775
box 0 0 1 1
use contact_7  contact_7_306
timestamp 1624857261
transform 1 0 216907 0 1 39111
box 0 0 1 1
use contact_7  contact_7_305
timestamp 1624857261
transform 1 0 216907 0 1 39447
box 0 0 1 1
use contact_7  contact_7_304
timestamp 1624857261
transform 1 0 216907 0 1 39783
box 0 0 1 1
use contact_7  contact_7_303
timestamp 1624857261
transform 1 0 216907 0 1 40119
box 0 0 1 1
use contact_7  contact_7_302
timestamp 1624857261
transform 1 0 216907 0 1 40455
box 0 0 1 1
use contact_7  contact_7_301
timestamp 1624857261
transform 1 0 216907 0 1 40791
box 0 0 1 1
use contact_7  contact_7_300
timestamp 1624857261
transform 1 0 216907 0 1 41127
box 0 0 1 1
use contact_7  contact_7_299
timestamp 1624857261
transform 1 0 216907 0 1 41463
box 0 0 1 1
use contact_7  contact_7_298
timestamp 1624857261
transform 1 0 216907 0 1 41799
box 0 0 1 1
use contact_7  contact_7_297
timestamp 1624857261
transform 1 0 216907 0 1 42135
box 0 0 1 1
use contact_7  contact_7_296
timestamp 1624857261
transform 1 0 216907 0 1 42471
box 0 0 1 1
use contact_7  contact_7_295
timestamp 1624857261
transform 1 0 216907 0 1 42807
box 0 0 1 1
use contact_7  contact_7_294
timestamp 1624857261
transform 1 0 216907 0 1 43143
box 0 0 1 1
use contact_7  contact_7_293
timestamp 1624857261
transform 1 0 216907 0 1 43479
box 0 0 1 1
use contact_7  contact_7_292
timestamp 1624857261
transform 1 0 216907 0 1 43815
box 0 0 1 1
use contact_7  contact_7_291
timestamp 1624857261
transform 1 0 216907 0 1 44151
box 0 0 1 1
use contact_7  contact_7_290
timestamp 1624857261
transform 1 0 216907 0 1 44487
box 0 0 1 1
use contact_7  contact_7_289
timestamp 1624857261
transform 1 0 216907 0 1 44823
box 0 0 1 1
use contact_7  contact_7_288
timestamp 1624857261
transform 1 0 216907 0 1 45159
box 0 0 1 1
use contact_7  contact_7_287
timestamp 1624857261
transform 1 0 216907 0 1 45495
box 0 0 1 1
use contact_7  contact_7_286
timestamp 1624857261
transform 1 0 216907 0 1 45831
box 0 0 1 1
use contact_7  contact_7_285
timestamp 1624857261
transform 1 0 216907 0 1 46167
box 0 0 1 1
use contact_7  contact_7_284
timestamp 1624857261
transform 1 0 216907 0 1 46503
box 0 0 1 1
use contact_7  contact_7_283
timestamp 1624857261
transform 1 0 216907 0 1 46839
box 0 0 1 1
use contact_7  contact_7_282
timestamp 1624857261
transform 1 0 216907 0 1 47175
box 0 0 1 1
use contact_7  contact_7_281
timestamp 1624857261
transform 1 0 216907 0 1 47511
box 0 0 1 1
use contact_7  contact_7_280
timestamp 1624857261
transform 1 0 216907 0 1 47847
box 0 0 1 1
use contact_7  contact_7_279
timestamp 1624857261
transform 1 0 216907 0 1 48183
box 0 0 1 1
use contact_7  contact_7_278
timestamp 1624857261
transform 1 0 216907 0 1 48519
box 0 0 1 1
use contact_7  contact_7_277
timestamp 1624857261
transform 1 0 216907 0 1 48855
box 0 0 1 1
use contact_7  contact_7_276
timestamp 1624857261
transform 1 0 216907 0 1 49191
box 0 0 1 1
use contact_7  contact_7_275
timestamp 1624857261
transform 1 0 216907 0 1 49527
box 0 0 1 1
use contact_7  contact_7_274
timestamp 1624857261
transform 1 0 216907 0 1 49863
box 0 0 1 1
use contact_7  contact_7_273
timestamp 1624857261
transform 1 0 216907 0 1 50199
box 0 0 1 1
use contact_7  contact_7_272
timestamp 1624857261
transform 1 0 216907 0 1 50535
box 0 0 1 1
use contact_7  contact_7_271
timestamp 1624857261
transform 1 0 216907 0 1 50871
box 0 0 1 1
use contact_7  contact_7_270
timestamp 1624857261
transform 1 0 216907 0 1 51207
box 0 0 1 1
use contact_7  contact_7_269
timestamp 1624857261
transform 1 0 216907 0 1 51543
box 0 0 1 1
use contact_7  contact_7_268
timestamp 1624857261
transform 1 0 216907 0 1 51879
box 0 0 1 1
use contact_7  contact_7_267
timestamp 1624857261
transform 1 0 216907 0 1 52215
box 0 0 1 1
use contact_7  contact_7_266
timestamp 1624857261
transform 1 0 216907 0 1 52551
box 0 0 1 1
use contact_7  contact_7_265
timestamp 1624857261
transform 1 0 216907 0 1 52887
box 0 0 1 1
use contact_7  contact_7_264
timestamp 1624857261
transform 1 0 216907 0 1 53223
box 0 0 1 1
use contact_7  contact_7_263
timestamp 1624857261
transform 1 0 216907 0 1 53559
box 0 0 1 1
use contact_7  contact_7_262
timestamp 1624857261
transform 1 0 216907 0 1 53895
box 0 0 1 1
use contact_7  contact_7_261
timestamp 1624857261
transform 1 0 216907 0 1 54231
box 0 0 1 1
use contact_7  contact_7_260
timestamp 1624857261
transform 1 0 216907 0 1 54567
box 0 0 1 1
use contact_7  contact_7_259
timestamp 1624857261
transform 1 0 216907 0 1 54903
box 0 0 1 1
use contact_7  contact_7_258
timestamp 1624857261
transform 1 0 216907 0 1 55239
box 0 0 1 1
use contact_7  contact_7_257
timestamp 1624857261
transform 1 0 216907 0 1 55575
box 0 0 1 1
use contact_7  contact_7_256
timestamp 1624857261
transform 1 0 216907 0 1 55911
box 0 0 1 1
use contact_7  contact_7_255
timestamp 1624857261
transform 1 0 216907 0 1 56247
box 0 0 1 1
use contact_7  contact_7_254
timestamp 1624857261
transform 1 0 216907 0 1 56583
box 0 0 1 1
use contact_7  contact_7_253
timestamp 1624857261
transform 1 0 216907 0 1 56919
box 0 0 1 1
use contact_7  contact_7_252
timestamp 1624857261
transform 1 0 216907 0 1 57255
box 0 0 1 1
use contact_7  contact_7_251
timestamp 1624857261
transform 1 0 216907 0 1 57591
box 0 0 1 1
use contact_7  contact_7_250
timestamp 1624857261
transform 1 0 216907 0 1 57927
box 0 0 1 1
use contact_7  contact_7_249
timestamp 1624857261
transform 1 0 216907 0 1 58263
box 0 0 1 1
use contact_7  contact_7_248
timestamp 1624857261
transform 1 0 216907 0 1 58599
box 0 0 1 1
use contact_7  contact_7_247
timestamp 1624857261
transform 1 0 216907 0 1 58935
box 0 0 1 1
use contact_7  contact_7_246
timestamp 1624857261
transform 1 0 216907 0 1 59271
box 0 0 1 1
use contact_7  contact_7_245
timestamp 1624857261
transform 1 0 216907 0 1 59607
box 0 0 1 1
use contact_7  contact_7_244
timestamp 1624857261
transform 1 0 216907 0 1 59943
box 0 0 1 1
use contact_7  contact_7_243
timestamp 1624857261
transform 1 0 216907 0 1 60279
box 0 0 1 1
use contact_7  contact_7_242
timestamp 1624857261
transform 1 0 216907 0 1 60615
box 0 0 1 1
use contact_7  contact_7_241
timestamp 1624857261
transform 1 0 216907 0 1 60951
box 0 0 1 1
use contact_7  contact_7_240
timestamp 1624857261
transform 1 0 216907 0 1 61287
box 0 0 1 1
use contact_7  contact_7_239
timestamp 1624857261
transform 1 0 216907 0 1 61623
box 0 0 1 1
use contact_7  contact_7_238
timestamp 1624857261
transform 1 0 216907 0 1 61959
box 0 0 1 1
use contact_7  contact_7_237
timestamp 1624857261
transform 1 0 216907 0 1 62295
box 0 0 1 1
use contact_7  contact_7_236
timestamp 1624857261
transform 1 0 216907 0 1 62631
box 0 0 1 1
use contact_7  contact_7_235
timestamp 1624857261
transform 1 0 216907 0 1 62967
box 0 0 1 1
use contact_7  contact_7_234
timestamp 1624857261
transform 1 0 216907 0 1 63303
box 0 0 1 1
use contact_7  contact_7_233
timestamp 1624857261
transform 1 0 216907 0 1 63639
box 0 0 1 1
use contact_7  contact_7_232
timestamp 1624857261
transform 1 0 216907 0 1 63975
box 0 0 1 1
use contact_7  contact_7_231
timestamp 1624857261
transform 1 0 216907 0 1 64311
box 0 0 1 1
use contact_7  contact_7_230
timestamp 1624857261
transform 1 0 216907 0 1 64647
box 0 0 1 1
use contact_7  contact_7_229
timestamp 1624857261
transform 1 0 216907 0 1 64983
box 0 0 1 1
use contact_7  contact_7_228
timestamp 1624857261
transform 1 0 216907 0 1 65319
box 0 0 1 1
use contact_7  contact_7_227
timestamp 1624857261
transform 1 0 216907 0 1 65655
box 0 0 1 1
use contact_7  contact_7_226
timestamp 1624857261
transform 1 0 216907 0 1 65991
box 0 0 1 1
use contact_7  contact_7_225
timestamp 1624857261
transform 1 0 216907 0 1 66327
box 0 0 1 1
use contact_7  contact_7_224
timestamp 1624857261
transform 1 0 216907 0 1 66663
box 0 0 1 1
use contact_7  contact_7_223
timestamp 1624857261
transform 1 0 216907 0 1 66999
box 0 0 1 1
use contact_7  contact_7_222
timestamp 1624857261
transform 1 0 216907 0 1 67335
box 0 0 1 1
use contact_7  contact_7_221
timestamp 1624857261
transform 1 0 216907 0 1 67671
box 0 0 1 1
use contact_7  contact_7_220
timestamp 1624857261
transform 1 0 216907 0 1 68007
box 0 0 1 1
use contact_7  contact_7_219
timestamp 1624857261
transform 1 0 216907 0 1 68343
box 0 0 1 1
use contact_7  contact_7_218
timestamp 1624857261
transform 1 0 216907 0 1 68679
box 0 0 1 1
use contact_7  contact_7_217
timestamp 1624857261
transform 1 0 216907 0 1 69015
box 0 0 1 1
use contact_7  contact_7_216
timestamp 1624857261
transform 1 0 216907 0 1 69351
box 0 0 1 1
use contact_7  contact_7_215
timestamp 1624857261
transform 1 0 216907 0 1 69687
box 0 0 1 1
use contact_7  contact_7_214
timestamp 1624857261
transform 1 0 216907 0 1 70023
box 0 0 1 1
use contact_7  contact_7_213
timestamp 1624857261
transform 1 0 216907 0 1 70359
box 0 0 1 1
use contact_7  contact_7_212
timestamp 1624857261
transform 1 0 216907 0 1 70695
box 0 0 1 1
use contact_7  contact_7_211
timestamp 1624857261
transform 1 0 216907 0 1 71031
box 0 0 1 1
use contact_7  contact_7_210
timestamp 1624857261
transform 1 0 216907 0 1 71367
box 0 0 1 1
use contact_7  contact_7_209
timestamp 1624857261
transform 1 0 216907 0 1 71703
box 0 0 1 1
use contact_7  contact_7_208
timestamp 1624857261
transform 1 0 216907 0 1 72039
box 0 0 1 1
use contact_7  contact_7_207
timestamp 1624857261
transform 1 0 216907 0 1 72375
box 0 0 1 1
use contact_7  contact_7_206
timestamp 1624857261
transform 1 0 216907 0 1 72711
box 0 0 1 1
use contact_7  contact_7_205
timestamp 1624857261
transform 1 0 216907 0 1 73047
box 0 0 1 1
use contact_7  contact_7_204
timestamp 1624857261
transform 1 0 216907 0 1 73383
box 0 0 1 1
use contact_7  contact_7_203
timestamp 1624857261
transform 1 0 216907 0 1 73719
box 0 0 1 1
use contact_7  contact_7_202
timestamp 1624857261
transform 1 0 216907 0 1 74055
box 0 0 1 1
use contact_7  contact_7_201
timestamp 1624857261
transform 1 0 216907 0 1 74391
box 0 0 1 1
use contact_7  contact_7_200
timestamp 1624857261
transform 1 0 216907 0 1 74727
box 0 0 1 1
use contact_7  contact_7_199
timestamp 1624857261
transform 1 0 216907 0 1 75063
box 0 0 1 1
use contact_7  contact_7_198
timestamp 1624857261
transform 1 0 216907 0 1 75399
box 0 0 1 1
use contact_7  contact_7_197
timestamp 1624857261
transform 1 0 216907 0 1 75735
box 0 0 1 1
use contact_7  contact_7_196
timestamp 1624857261
transform 1 0 216907 0 1 76071
box 0 0 1 1
use contact_7  contact_7_195
timestamp 1624857261
transform 1 0 216907 0 1 76407
box 0 0 1 1
use contact_7  contact_7_194
timestamp 1624857261
transform 1 0 216907 0 1 76743
box 0 0 1 1
use contact_7  contact_7_193
timestamp 1624857261
transform 1 0 216907 0 1 77079
box 0 0 1 1
use contact_7  contact_7_192
timestamp 1624857261
transform 1 0 216907 0 1 77415
box 0 0 1 1
use contact_7  contact_7_191
timestamp 1624857261
transform 1 0 216907 0 1 77751
box 0 0 1 1
use contact_7  contact_7_190
timestamp 1624857261
transform 1 0 216907 0 1 78087
box 0 0 1 1
use contact_7  contact_7_189
timestamp 1624857261
transform 1 0 216907 0 1 78423
box 0 0 1 1
use contact_7  contact_7_188
timestamp 1624857261
transform 1 0 216907 0 1 78759
box 0 0 1 1
use contact_7  contact_7_187
timestamp 1624857261
transform 1 0 216907 0 1 79095
box 0 0 1 1
use contact_7  contact_7_186
timestamp 1624857261
transform 1 0 216907 0 1 79431
box 0 0 1 1
use contact_7  contact_7_185
timestamp 1624857261
transform 1 0 216907 0 1 79767
box 0 0 1 1
use contact_7  contact_7_184
timestamp 1624857261
transform 1 0 216907 0 1 80103
box 0 0 1 1
use contact_7  contact_7_183
timestamp 1624857261
transform 1 0 216907 0 1 80439
box 0 0 1 1
use contact_7  contact_7_182
timestamp 1624857261
transform 1 0 216907 0 1 80775
box 0 0 1 1
use contact_7  contact_7_181
timestamp 1624857261
transform 1 0 216907 0 1 81111
box 0 0 1 1
use contact_7  contact_7_180
timestamp 1624857261
transform 1 0 216907 0 1 81447
box 0 0 1 1
use contact_7  contact_7_179
timestamp 1624857261
transform 1 0 216907 0 1 81783
box 0 0 1 1
use contact_7  contact_7_178
timestamp 1624857261
transform 1 0 216907 0 1 82119
box 0 0 1 1
use contact_7  contact_7_177
timestamp 1624857261
transform 1 0 216907 0 1 82455
box 0 0 1 1
use contact_7  contact_7_176
timestamp 1624857261
transform 1 0 216907 0 1 82791
box 0 0 1 1
use contact_7  contact_7_175
timestamp 1624857261
transform 1 0 216907 0 1 83127
box 0 0 1 1
use contact_7  contact_7_174
timestamp 1624857261
transform 1 0 216907 0 1 83463
box 0 0 1 1
use contact_7  contact_7_173
timestamp 1624857261
transform 1 0 216907 0 1 83799
box 0 0 1 1
use contact_7  contact_7_172
timestamp 1624857261
transform 1 0 216907 0 1 84135
box 0 0 1 1
use contact_7  contact_7_171
timestamp 1624857261
transform 1 0 216907 0 1 84471
box 0 0 1 1
use contact_7  contact_7_170
timestamp 1624857261
transform 1 0 216907 0 1 84807
box 0 0 1 1
use contact_7  contact_7_169
timestamp 1624857261
transform 1 0 216907 0 1 85143
box 0 0 1 1
use contact_7  contact_7_168
timestamp 1624857261
transform 1 0 216907 0 1 85479
box 0 0 1 1
use contact_7  contact_7_167
timestamp 1624857261
transform 1 0 216907 0 1 85815
box 0 0 1 1
use contact_7  contact_7_166
timestamp 1624857261
transform 1 0 216907 0 1 86151
box 0 0 1 1
use contact_7  contact_7_165
timestamp 1624857261
transform 1 0 216907 0 1 86487
box 0 0 1 1
use contact_7  contact_7_164
timestamp 1624857261
transform 1 0 216907 0 1 86823
box 0 0 1 1
use contact_7  contact_7_163
timestamp 1624857261
transform 1 0 216907 0 1 87159
box 0 0 1 1
use contact_7  contact_7_162
timestamp 1624857261
transform 1 0 216907 0 1 87495
box 0 0 1 1
use contact_7  contact_7_161
timestamp 1624857261
transform 1 0 216907 0 1 87831
box 0 0 1 1
use contact_7  contact_7_160
timestamp 1624857261
transform 1 0 216907 0 1 88167
box 0 0 1 1
use contact_7  contact_7_159
timestamp 1624857261
transform 1 0 216907 0 1 88503
box 0 0 1 1
use contact_7  contact_7_158
timestamp 1624857261
transform 1 0 216907 0 1 88839
box 0 0 1 1
use contact_7  contact_7_157
timestamp 1624857261
transform 1 0 216907 0 1 89175
box 0 0 1 1
use contact_7  contact_7_156
timestamp 1624857261
transform 1 0 216907 0 1 89511
box 0 0 1 1
use contact_7  contact_7_155
timestamp 1624857261
transform 1 0 216907 0 1 89847
box 0 0 1 1
use contact_7  contact_7_154
timestamp 1624857261
transform 1 0 216907 0 1 90183
box 0 0 1 1
use contact_7  contact_7_153
timestamp 1624857261
transform 1 0 216907 0 1 90519
box 0 0 1 1
use contact_7  contact_7_152
timestamp 1624857261
transform 1 0 216907 0 1 90855
box 0 0 1 1
use contact_7  contact_7_151
timestamp 1624857261
transform 1 0 216907 0 1 91191
box 0 0 1 1
use contact_7  contact_7_150
timestamp 1624857261
transform 1 0 216907 0 1 91527
box 0 0 1 1
use contact_7  contact_7_149
timestamp 1624857261
transform 1 0 216907 0 1 91863
box 0 0 1 1
use contact_7  contact_7_148
timestamp 1624857261
transform 1 0 216907 0 1 92199
box 0 0 1 1
use contact_7  contact_7_147
timestamp 1624857261
transform 1 0 216907 0 1 92535
box 0 0 1 1
use contact_7  contact_7_146
timestamp 1624857261
transform 1 0 216907 0 1 92871
box 0 0 1 1
use contact_7  contact_7_145
timestamp 1624857261
transform 1 0 216907 0 1 93207
box 0 0 1 1
use contact_7  contact_7_144
timestamp 1624857261
transform 1 0 216907 0 1 93543
box 0 0 1 1
use contact_7  contact_7_143
timestamp 1624857261
transform 1 0 216907 0 1 93879
box 0 0 1 1
use contact_7  contact_7_142
timestamp 1624857261
transform 1 0 216907 0 1 94215
box 0 0 1 1
use contact_7  contact_7_141
timestamp 1624857261
transform 1 0 216907 0 1 94551
box 0 0 1 1
use contact_7  contact_7_140
timestamp 1624857261
transform 1 0 216907 0 1 94887
box 0 0 1 1
use contact_7  contact_7_139
timestamp 1624857261
transform 1 0 216907 0 1 95223
box 0 0 1 1
use contact_7  contact_7_138
timestamp 1624857261
transform 1 0 216907 0 1 95559
box 0 0 1 1
use contact_7  contact_7_137
timestamp 1624857261
transform 1 0 216907 0 1 95895
box 0 0 1 1
use contact_7  contact_7_136
timestamp 1624857261
transform 1 0 216907 0 1 96231
box 0 0 1 1
use contact_7  contact_7_135
timestamp 1624857261
transform 1 0 216907 0 1 96567
box 0 0 1 1
use contact_7  contact_7_134
timestamp 1624857261
transform 1 0 216907 0 1 96903
box 0 0 1 1
use contact_7  contact_7_133
timestamp 1624857261
transform 1 0 216907 0 1 97239
box 0 0 1 1
use contact_7  contact_7_132
timestamp 1624857261
transform 1 0 216907 0 1 97575
box 0 0 1 1
use contact_7  contact_7_131
timestamp 1624857261
transform 1 0 216907 0 1 97911
box 0 0 1 1
use contact_7  contact_7_130
timestamp 1624857261
transform 1 0 216907 0 1 98247
box 0 0 1 1
use contact_7  contact_7_129
timestamp 1624857261
transform 1 0 216907 0 1 98583
box 0 0 1 1
use contact_7  contact_7_128
timestamp 1624857261
transform 1 0 216907 0 1 98919
box 0 0 1 1
use contact_7  contact_7_127
timestamp 1624857261
transform 1 0 216907 0 1 99255
box 0 0 1 1
use contact_7  contact_7_126
timestamp 1624857261
transform 1 0 216907 0 1 99591
box 0 0 1 1
use contact_7  contact_7_125
timestamp 1624857261
transform 1 0 216907 0 1 99927
box 0 0 1 1
use contact_7  contact_7_124
timestamp 1624857261
transform 1 0 216907 0 1 100263
box 0 0 1 1
use contact_7  contact_7_123
timestamp 1624857261
transform 1 0 216907 0 1 100599
box 0 0 1 1
use contact_7  contact_7_122
timestamp 1624857261
transform 1 0 216907 0 1 100935
box 0 0 1 1
use contact_7  contact_7_121
timestamp 1624857261
transform 1 0 216907 0 1 101271
box 0 0 1 1
use contact_7  contact_7_120
timestamp 1624857261
transform 1 0 216907 0 1 101607
box 0 0 1 1
use contact_7  contact_7_119
timestamp 1624857261
transform 1 0 216907 0 1 101943
box 0 0 1 1
use contact_7  contact_7_118
timestamp 1624857261
transform 1 0 216907 0 1 102279
box 0 0 1 1
use contact_7  contact_7_117
timestamp 1624857261
transform 1 0 216907 0 1 102615
box 0 0 1 1
use contact_7  contact_7_116
timestamp 1624857261
transform 1 0 216907 0 1 102951
box 0 0 1 1
use contact_7  contact_7_115
timestamp 1624857261
transform 1 0 216907 0 1 103287
box 0 0 1 1
use contact_7  contact_7_114
timestamp 1624857261
transform 1 0 216907 0 1 103623
box 0 0 1 1
use contact_7  contact_7_113
timestamp 1624857261
transform 1 0 216907 0 1 103959
box 0 0 1 1
use contact_7  contact_7_112
timestamp 1624857261
transform 1 0 216907 0 1 104295
box 0 0 1 1
use contact_7  contact_7_111
timestamp 1624857261
transform 1 0 216907 0 1 104631
box 0 0 1 1
use contact_7  contact_7_110
timestamp 1624857261
transform 1 0 216907 0 1 104967
box 0 0 1 1
use contact_7  contact_7_109
timestamp 1624857261
transform 1 0 216907 0 1 105303
box 0 0 1 1
use contact_7  contact_7_108
timestamp 1624857261
transform 1 0 216907 0 1 105639
box 0 0 1 1
use contact_7  contact_7_107
timestamp 1624857261
transform 1 0 216907 0 1 105975
box 0 0 1 1
use contact_7  contact_7_106
timestamp 1624857261
transform 1 0 216907 0 1 106311
box 0 0 1 1
use contact_7  contact_7_105
timestamp 1624857261
transform 1 0 216907 0 1 106647
box 0 0 1 1
use contact_7  contact_7_104
timestamp 1624857261
transform 1 0 216907 0 1 106983
box 0 0 1 1
use contact_7  contact_7_103
timestamp 1624857261
transform 1 0 216907 0 1 107319
box 0 0 1 1
use contact_7  contact_7_102
timestamp 1624857261
transform 1 0 216907 0 1 107655
box 0 0 1 1
use contact_7  contact_7_101
timestamp 1624857261
transform 1 0 216907 0 1 107991
box 0 0 1 1
use contact_7  contact_7_100
timestamp 1624857261
transform 1 0 216907 0 1 108327
box 0 0 1 1
use contact_7  contact_7_99
timestamp 1624857261
transform 1 0 216907 0 1 108663
box 0 0 1 1
use contact_7  contact_7_98
timestamp 1624857261
transform 1 0 216907 0 1 108999
box 0 0 1 1
use contact_7  contact_7_97
timestamp 1624857261
transform 1 0 216907 0 1 109335
box 0 0 1 1
use contact_7  contact_7_96
timestamp 1624857261
transform 1 0 216907 0 1 109671
box 0 0 1 1
use contact_7  contact_7_95
timestamp 1624857261
transform 1 0 216907 0 1 110007
box 0 0 1 1
use contact_7  contact_7_94
timestamp 1624857261
transform 1 0 216907 0 1 110343
box 0 0 1 1
use contact_7  contact_7_93
timestamp 1624857261
transform 1 0 216907 0 1 110679
box 0 0 1 1
use contact_7  contact_7_92
timestamp 1624857261
transform 1 0 216907 0 1 111015
box 0 0 1 1
use contact_7  contact_7_91
timestamp 1624857261
transform 1 0 216907 0 1 111351
box 0 0 1 1
use contact_7  contact_7_90
timestamp 1624857261
transform 1 0 216907 0 1 111687
box 0 0 1 1
use contact_7  contact_7_89
timestamp 1624857261
transform 1 0 216907 0 1 112023
box 0 0 1 1
use contact_7  contact_7_88
timestamp 1624857261
transform 1 0 216907 0 1 112359
box 0 0 1 1
use contact_7  contact_7_87
timestamp 1624857261
transform 1 0 216907 0 1 112695
box 0 0 1 1
use contact_7  contact_7_86
timestamp 1624857261
transform 1 0 216907 0 1 113031
box 0 0 1 1
use contact_7  contact_7_85
timestamp 1624857261
transform 1 0 216907 0 1 113367
box 0 0 1 1
use contact_7  contact_7_84
timestamp 1624857261
transform 1 0 216907 0 1 113703
box 0 0 1 1
use contact_7  contact_7_83
timestamp 1624857261
transform 1 0 216907 0 1 114039
box 0 0 1 1
use contact_7  contact_7_82
timestamp 1624857261
transform 1 0 216907 0 1 114375
box 0 0 1 1
use contact_7  contact_7_81
timestamp 1624857261
transform 1 0 216907 0 1 114711
box 0 0 1 1
use contact_7  contact_7_80
timestamp 1624857261
transform 1 0 216907 0 1 115047
box 0 0 1 1
use contact_7  contact_7_79
timestamp 1624857261
transform 1 0 216907 0 1 115383
box 0 0 1 1
use contact_7  contact_7_78
timestamp 1624857261
transform 1 0 216907 0 1 115719
box 0 0 1 1
use contact_7  contact_7_77
timestamp 1624857261
transform 1 0 216907 0 1 116055
box 0 0 1 1
use contact_7  contact_7_76
timestamp 1624857261
transform 1 0 216907 0 1 116391
box 0 0 1 1
use contact_7  contact_7_75
timestamp 1624857261
transform 1 0 216907 0 1 116727
box 0 0 1 1
use contact_7  contact_7_74
timestamp 1624857261
transform 1 0 216907 0 1 117063
box 0 0 1 1
use contact_7  contact_7_73
timestamp 1624857261
transform 1 0 216907 0 1 117399
box 0 0 1 1
use contact_7  contact_7_72
timestamp 1624857261
transform 1 0 216907 0 1 117735
box 0 0 1 1
use contact_7  contact_7_71
timestamp 1624857261
transform 1 0 216907 0 1 118071
box 0 0 1 1
use contact_7  contact_7_70
timestamp 1624857261
transform 1 0 216907 0 1 118407
box 0 0 1 1
use contact_7  contact_7_69
timestamp 1624857261
transform 1 0 216907 0 1 118743
box 0 0 1 1
use contact_7  contact_7_68
timestamp 1624857261
transform 1 0 216907 0 1 119079
box 0 0 1 1
use contact_7  contact_7_67
timestamp 1624857261
transform 1 0 216907 0 1 119415
box 0 0 1 1
use contact_7  contact_7_66
timestamp 1624857261
transform 1 0 216907 0 1 119751
box 0 0 1 1
use contact_7  contact_7_65
timestamp 1624857261
transform 1 0 216907 0 1 120087
box 0 0 1 1
use contact_7  contact_7_64
timestamp 1624857261
transform 1 0 216907 0 1 120423
box 0 0 1 1
use contact_7  contact_7_63
timestamp 1624857261
transform 1 0 216907 0 1 120759
box 0 0 1 1
use contact_7  contact_7_62
timestamp 1624857261
transform 1 0 216907 0 1 121095
box 0 0 1 1
use contact_7  contact_7_61
timestamp 1624857261
transform 1 0 216907 0 1 121431
box 0 0 1 1
use contact_7  contact_7_60
timestamp 1624857261
transform 1 0 216907 0 1 121767
box 0 0 1 1
use contact_7  contact_7_59
timestamp 1624857261
transform 1 0 216907 0 1 122103
box 0 0 1 1
use contact_7  contact_7_58
timestamp 1624857261
transform 1 0 216907 0 1 122439
box 0 0 1 1
use contact_7  contact_7_57
timestamp 1624857261
transform 1 0 216907 0 1 122775
box 0 0 1 1
use contact_7  contact_7_56
timestamp 1624857261
transform 1 0 216907 0 1 123111
box 0 0 1 1
use contact_7  contact_7_55
timestamp 1624857261
transform 1 0 216907 0 1 123447
box 0 0 1 1
use contact_7  contact_7_54
timestamp 1624857261
transform 1 0 216907 0 1 123783
box 0 0 1 1
use contact_7  contact_7_53
timestamp 1624857261
transform 1 0 216907 0 1 124119
box 0 0 1 1
use contact_7  contact_7_52
timestamp 1624857261
transform 1 0 216907 0 1 124455
box 0 0 1 1
use contact_7  contact_7_51
timestamp 1624857261
transform 1 0 216907 0 1 124791
box 0 0 1 1
use contact_7  contact_7_50
timestamp 1624857261
transform 1 0 216907 0 1 125127
box 0 0 1 1
use contact_7  contact_7_49
timestamp 1624857261
transform 1 0 216907 0 1 125463
box 0 0 1 1
use contact_7  contact_7_48
timestamp 1624857261
transform 1 0 216907 0 1 125799
box 0 0 1 1
use contact_7  contact_7_47
timestamp 1624857261
transform 1 0 216907 0 1 126135
box 0 0 1 1
use contact_7  contact_7_46
timestamp 1624857261
transform 1 0 216907 0 1 126471
box 0 0 1 1
use contact_7  contact_7_45
timestamp 1624857261
transform 1 0 216907 0 1 126807
box 0 0 1 1
use contact_7  contact_7_44
timestamp 1624857261
transform 1 0 216907 0 1 127143
box 0 0 1 1
use contact_7  contact_7_43
timestamp 1624857261
transform 1 0 216907 0 1 127479
box 0 0 1 1
use contact_7  contact_7_42
timestamp 1624857261
transform 1 0 216907 0 1 127815
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1624857261
transform 1 0 216907 0 1 128151
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1624857261
transform 1 0 216907 0 1 128487
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1624857261
transform 1 0 216907 0 1 128823
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1624857261
transform 1 0 216907 0 1 129159
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1624857261
transform 1 0 216907 0 1 129495
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1624857261
transform 1 0 216907 0 1 129831
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1624857261
transform 1 0 216907 0 1 130167
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1624857261
transform 1 0 216907 0 1 130503
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1624857261
transform 1 0 216907 0 1 130839
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1624857261
transform 1 0 216907 0 1 131175
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1624857261
transform 1 0 216907 0 1 131511
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1624857261
transform 1 0 216907 0 1 131847
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1624857261
transform 1 0 216907 0 1 132183
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1624857261
transform 1 0 216907 0 1 132519
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1624857261
transform 1 0 216907 0 1 132855
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1624857261
transform 1 0 216907 0 1 133191
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1624857261
transform 1 0 216907 0 1 133527
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1624857261
transform 1 0 216907 0 1 133863
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1624857261
transform 1 0 216907 0 1 134199
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1624857261
transform 1 0 216907 0 1 134535
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1624857261
transform 1 0 216907 0 1 134871
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1624857261
transform 1 0 216907 0 1 135207
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1624857261
transform 1 0 216907 0 1 135543
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1624857261
transform 1 0 216907 0 1 135879
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1624857261
transform 1 0 216907 0 1 136215
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1624857261
transform 1 0 216907 0 1 136551
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1624857261
transform 1 0 216907 0 1 136887
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1624857261
transform 1 0 216907 0 1 137223
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1624857261
transform 1 0 216907 0 1 137559
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1624857261
transform 1 0 216907 0 1 137895
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1624857261
transform 1 0 216907 0 1 138231
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1624857261
transform 1 0 216907 0 1 138567
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1624857261
transform 1 0 216907 0 1 138903
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1624857261
transform 1 0 216907 0 1 139239
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1624857261
transform 1 0 216907 0 1 139575
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1624857261
transform 1 0 216907 0 1 139911
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1624857261
transform 1 0 216907 0 1 140247
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1624857261
transform 1 0 216907 0 1 140583
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1624857261
transform 1 0 216907 0 1 140919
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1624857261
transform 1 0 216907 0 1 141255
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1624857261
transform 1 0 216907 0 1 141591
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1624857261
transform 1 0 216907 0 1 141927
box 0 0 1 1
use contact_38  contact_38_71
timestamp 1624857261
transform 1 0 218416 0 1 143621
box 0 0 192 192
use contact_38  contact_38_70
timestamp 1624857261
transform 1 0 218144 0 1 277
box 0 0 192 192
use contact_38  contact_38_69
timestamp 1624857261
transform 1 0 218416 0 1 549
box 0 0 192 192
use contact_38  contact_38_68
timestamp 1624857261
transform 1 0 272 0 1 549
box 0 0 192 192
use contact_38  contact_38_67
timestamp 1624857261
transform 1 0 272 0 1 143621
box 0 0 192 192
use contact_38  contact_38_66
timestamp 1624857261
transform 1 0 544 0 1 413
box 0 0 192 192
use contact_38  contact_38_65
timestamp 1624857261
transform 1 0 544 0 1 549
box 0 0 192 192
use contact_38  contact_38_64
timestamp 1624857261
transform 1 0 218144 0 1 143485
box 0 0 192 192
use contact_38  contact_38_63
timestamp 1624857261
transform 1 0 218144 0 1 143621
box 0 0 192 192
use contact_38  contact_38_62
timestamp 1624857261
transform 1 0 218416 0 1 413
box 0 0 192 192
use contact_38  contact_38_61
timestamp 1624857261
transform 1 0 272 0 1 277
box 0 0 192 192
use contact_38  contact_38_60
timestamp 1624857261
transform 1 0 544 0 1 143757
box 0 0 192 192
use contact_38  contact_38_59
timestamp 1624857261
transform 1 0 218416 0 1 143485
box 0 0 192 192
use contact_38  contact_38_58
timestamp 1624857261
transform 1 0 218280 0 1 277
box 0 0 192 192
use contact_38  contact_38_57
timestamp 1624857261
transform 1 0 408 0 1 143621
box 0 0 192 192
use contact_38  contact_38_56
timestamp 1624857261
transform 1 0 408 0 1 143485
box 0 0 192 192
use contact_38  contact_38_55
timestamp 1624857261
transform 1 0 218280 0 1 143621
box 0 0 192 192
use contact_38  contact_38_54
timestamp 1624857261
transform 1 0 218280 0 1 549
box 0 0 192 192
use contact_38  contact_38_53
timestamp 1624857261
transform 1 0 544 0 1 277
box 0 0 192 192
use contact_38  contact_38_52
timestamp 1624857261
transform 1 0 408 0 1 277
box 0 0 192 192
use contact_38  contact_38_51
timestamp 1624857261
transform 1 0 218416 0 1 143757
box 0 0 192 192
use contact_38  contact_38_50
timestamp 1624857261
transform 1 0 218144 0 1 413
box 0 0 192 192
use contact_38  contact_38_49
timestamp 1624857261
transform 1 0 218416 0 1 277
box 0 0 192 192
use contact_38  contact_38_48
timestamp 1624857261
transform 1 0 544 0 1 143485
box 0 0 192 192
use contact_38  contact_38_47
timestamp 1624857261
transform 1 0 218144 0 1 549
box 0 0 192 192
use contact_38  contact_38_46
timestamp 1624857261
transform 1 0 544 0 1 143621
box 0 0 192 192
use contact_38  contact_38_45
timestamp 1624857261
transform 1 0 272 0 1 143757
box 0 0 192 192
use contact_38  contact_38_44
timestamp 1624857261
transform 1 0 272 0 1 143485
box 0 0 192 192
use contact_38  contact_38_43
timestamp 1624857261
transform 1 0 218280 0 1 413
box 0 0 192 192
use contact_38  contact_38_42
timestamp 1624857261
transform 1 0 218144 0 1 143757
box 0 0 192 192
use contact_38  contact_38_41
timestamp 1624857261
transform 1 0 408 0 1 143757
box 0 0 192 192
use contact_38  contact_38_40
timestamp 1624857261
transform 1 0 272 0 1 413
box 0 0 192 192
use contact_38  contact_38_39
timestamp 1624857261
transform 1 0 218280 0 1 143485
box 0 0 192 192
use contact_38  contact_38_38
timestamp 1624857261
transform 1 0 218280 0 1 143757
box 0 0 192 192
use contact_38  contact_38_37
timestamp 1624857261
transform 1 0 408 0 1 549
box 0 0 192 192
use contact_38  contact_38_36
timestamp 1624857261
transform 1 0 408 0 1 413
box 0 0 192 192
use contact_38  contact_38_35
timestamp 1624857261
transform 1 0 217464 0 1 142941
box 0 0 192 192
use contact_38  contact_38_34
timestamp 1624857261
transform 1 0 1224 0 1 957
box 0 0 192 192
use contact_38  contact_38_33
timestamp 1624857261
transform 1 0 952 0 1 1229
box 0 0 192 192
use contact_38  contact_38_32
timestamp 1624857261
transform 1 0 217736 0 1 957
box 0 0 192 192
use contact_38  contact_38_31
timestamp 1624857261
transform 1 0 952 0 1 957
box 0 0 192 192
use contact_38  contact_38_30
timestamp 1624857261
transform 1 0 217736 0 1 142805
box 0 0 192 192
use contact_38  contact_38_29
timestamp 1624857261
transform 1 0 1088 0 1 1093
box 0 0 192 192
use contact_38  contact_38_28
timestamp 1624857261
transform 1 0 1224 0 1 142805
box 0 0 192 192
use contact_38  contact_38_27
timestamp 1624857261
transform 1 0 1224 0 1 1093
box 0 0 192 192
use contact_38  contact_38_26
timestamp 1624857261
transform 1 0 1088 0 1 142941
box 0 0 192 192
use contact_38  contact_38_25
timestamp 1624857261
transform 1 0 217464 0 1 1229
box 0 0 192 192
use contact_38  contact_38_24
timestamp 1624857261
transform 1 0 952 0 1 142941
box 0 0 192 192
use contact_38  contact_38_23
timestamp 1624857261
transform 1 0 217600 0 1 142805
box 0 0 192 192
use contact_38  contact_38_22
timestamp 1624857261
transform 1 0 217600 0 1 1093
box 0 0 192 192
use contact_38  contact_38_21
timestamp 1624857261
transform 1 0 217736 0 1 1093
box 0 0 192 192
use contact_38  contact_38_20
timestamp 1624857261
transform 1 0 217464 0 1 957
box 0 0 192 192
use contact_38  contact_38_19
timestamp 1624857261
transform 1 0 217464 0 1 143077
box 0 0 192 192
use contact_38  contact_38_18
timestamp 1624857261
transform 1 0 217600 0 1 143077
box 0 0 192 192
use contact_38  contact_38_17
timestamp 1624857261
transform 1 0 217736 0 1 142941
box 0 0 192 192
use contact_38  contact_38_16
timestamp 1624857261
transform 1 0 1088 0 1 957
box 0 0 192 192
use contact_38  contact_38_15
timestamp 1624857261
transform 1 0 217464 0 1 142805
box 0 0 192 192
use contact_38  contact_38_14
timestamp 1624857261
transform 1 0 1224 0 1 142941
box 0 0 192 192
use contact_38  contact_38_13
timestamp 1624857261
transform 1 0 1224 0 1 1229
box 0 0 192 192
use contact_38  contact_38_12
timestamp 1624857261
transform 1 0 952 0 1 1093
box 0 0 192 192
use contact_38  contact_38_11
timestamp 1624857261
transform 1 0 1088 0 1 142805
box 0 0 192 192
use contact_38  contact_38_10
timestamp 1624857261
transform 1 0 952 0 1 143077
box 0 0 192 192
use contact_38  contact_38_9
timestamp 1624857261
transform 1 0 1088 0 1 1229
box 0 0 192 192
use contact_38  contact_38_8
timestamp 1624857261
transform 1 0 217736 0 1 143077
box 0 0 192 192
use contact_38  contact_38_7
timestamp 1624857261
transform 1 0 1224 0 1 143077
box 0 0 192 192
use contact_38  contact_38_6
timestamp 1624857261
transform 1 0 217736 0 1 1229
box 0 0 192 192
use contact_38  contact_38_5
timestamp 1624857261
transform 1 0 217464 0 1 1093
box 0 0 192 192
use contact_38  contact_38_4
timestamp 1624857261
transform 1 0 1088 0 1 143077
box 0 0 192 192
use contact_38  contact_38_3
timestamp 1624857261
transform 1 0 217600 0 1 957
box 0 0 192 192
use contact_38  contact_38_2
timestamp 1624857261
transform 1 0 952 0 1 142805
box 0 0 192 192
use contact_38  contact_38_1
timestamp 1624857261
transform 1 0 217600 0 1 142941
box 0 0 192 192
use contact_38  contact_38_0
timestamp 1624857261
transform 1 0 217600 0 1 1229
box 0 0 192 192
use contact_32  contact_32_6047
timestamp 1624857261
transform 1 0 2103 0 1 22884
box 0 0 1 1
use contact_32  contact_32_6046
timestamp 1624857261
transform 1 0 2103 0 1 30291
box 0 0 1 1
use contact_32  contact_32_6045
timestamp 1624857261
transform 1 0 216487 0 1 127844
box 0 0 1 1
use contact_32  contact_32_6044
timestamp 1624857261
transform 1 0 216487 0 1 117609
box 0 0 1 1
use contact_32  contact_32_6043
timestamp 1624857261
transform 1 0 24616 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6042
timestamp 1624857261
transform 1 0 25976 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6041
timestamp 1624857261
transform 1 0 27064 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6040
timestamp 1624857261
transform 1 0 28288 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6039
timestamp 1624857261
transform 1 0 29240 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6038
timestamp 1624857261
transform 1 0 30600 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6037
timestamp 1624857261
transform 1 0 31688 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6036
timestamp 1624857261
transform 1 0 32776 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6035
timestamp 1624857261
transform 1 0 34000 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6034
timestamp 1624857261
transform 1 0 35088 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6033
timestamp 1624857261
transform 1 0 36448 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6032
timestamp 1624857261
transform 1 0 37536 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6031
timestamp 1624857261
transform 1 0 38624 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6030
timestamp 1624857261
transform 1 0 39848 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6029
timestamp 1624857261
transform 1 0 40936 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6028
timestamp 1624857261
transform 1 0 42296 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6027
timestamp 1624857261
transform 1 0 43384 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6026
timestamp 1624857261
transform 1 0 44608 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6025
timestamp 1624857261
transform 1 0 45832 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6024
timestamp 1624857261
transform 1 0 46920 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6023
timestamp 1624857261
transform 1 0 48008 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6022
timestamp 1624857261
transform 1 0 49096 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6021
timestamp 1624857261
transform 1 0 50320 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6020
timestamp 1624857261
transform 1 0 51544 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6019
timestamp 1624857261
transform 1 0 52768 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6018
timestamp 1624857261
transform 1 0 53856 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6017
timestamp 1624857261
transform 1 0 54944 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6016
timestamp 1624857261
transform 1 0 56168 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6015
timestamp 1624857261
transform 1 0 57392 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6014
timestamp 1624857261
transform 1 0 58616 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6013
timestamp 1624857261
transform 1 0 59840 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6012
timestamp 1624857261
transform 1 0 60792 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6011
timestamp 1624857261
transform 1 0 16456 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6010
timestamp 1624857261
transform 1 0 17680 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6009
timestamp 1624857261
transform 1 0 18768 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6008
timestamp 1624857261
transform 1 0 19992 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6007
timestamp 1624857261
transform 1 0 21080 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6006
timestamp 1624857261
transform 1 0 22304 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6005
timestamp 1624857261
transform 1 0 23528 0 1 2589
box 0 0 1 1
use contact_32  contact_32_6004
timestamp 1624857261
transform 1 0 201008 0 1 141445
box 0 0 1 1
use contact_32  contact_32_6003
timestamp 1624857261
transform 1 0 199920 0 1 141445
box 0 0 1 1
use contact_32  contact_32_6002
timestamp 1624857261
transform 1 0 198560 0 1 141445
box 0 0 1 1
use contact_32  contact_32_6001
timestamp 1624857261
transform 1 0 29512 0 1 133149
box 0 0 1 1
use contact_32  contact_32_6000
timestamp 1624857261
transform 1 0 34408 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5999
timestamp 1624857261
transform 1 0 39440 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5998
timestamp 1624857261
transform 1 0 44472 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5997
timestamp 1624857261
transform 1 0 49504 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5996
timestamp 1624857261
transform 1 0 54536 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5995
timestamp 1624857261
transform 1 0 59432 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5994
timestamp 1624857261
transform 1 0 64464 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5993
timestamp 1624857261
transform 1 0 69496 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5992
timestamp 1624857261
transform 1 0 74528 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5991
timestamp 1624857261
transform 1 0 79560 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5990
timestamp 1624857261
transform 1 0 84320 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5989
timestamp 1624857261
transform 1 0 89352 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5988
timestamp 1624857261
transform 1 0 94520 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5987
timestamp 1624857261
transform 1 0 99416 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5986
timestamp 1624857261
transform 1 0 104312 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5985
timestamp 1624857261
transform 1 0 109344 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5984
timestamp 1624857261
transform 1 0 114376 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5983
timestamp 1624857261
transform 1 0 119272 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5982
timestamp 1624857261
transform 1 0 124304 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5981
timestamp 1624857261
transform 1 0 129336 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5980
timestamp 1624857261
transform 1 0 134368 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5979
timestamp 1624857261
transform 1 0 139400 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5978
timestamp 1624857261
transform 1 0 144296 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5977
timestamp 1624857261
transform 1 0 149328 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5976
timestamp 1624857261
transform 1 0 154360 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5975
timestamp 1624857261
transform 1 0 159392 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5974
timestamp 1624857261
transform 1 0 164424 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5973
timestamp 1624857261
transform 1 0 169184 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5972
timestamp 1624857261
transform 1 0 174216 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5971
timestamp 1624857261
transform 1 0 179384 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5970
timestamp 1624857261
transform 1 0 184280 0 1 133149
box 0 0 1 1
use contact_32  contact_32_5969
timestamp 1624857261
transform 1 0 28968 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5968
timestamp 1624857261
transform 1 0 34544 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5967
timestamp 1624857261
transform 1 0 39440 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5966
timestamp 1624857261
transform 1 0 44200 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5965
timestamp 1624857261
transform 1 0 49504 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5964
timestamp 1624857261
transform 1 0 54536 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5963
timestamp 1624857261
transform 1 0 59296 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5962
timestamp 1624857261
transform 1 0 64464 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5961
timestamp 1624857261
transform 1 0 69496 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5960
timestamp 1624857261
transform 1 0 74392 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5959
timestamp 1624857261
transform 1 0 79424 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5958
timestamp 1624857261
transform 1 0 84320 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5957
timestamp 1624857261
transform 1 0 89352 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5956
timestamp 1624857261
transform 1 0 94384 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5955
timestamp 1624857261
transform 1 0 99416 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5954
timestamp 1624857261
transform 1 0 104312 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5953
timestamp 1624857261
transform 1 0 109072 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5952
timestamp 1624857261
transform 1 0 114376 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5951
timestamp 1624857261
transform 1 0 119272 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5950
timestamp 1624857261
transform 1 0 124304 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5949
timestamp 1624857261
transform 1 0 129336 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5948
timestamp 1624857261
transform 1 0 134368 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5947
timestamp 1624857261
transform 1 0 139264 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5946
timestamp 1624857261
transform 1 0 144296 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5945
timestamp 1624857261
transform 1 0 149056 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5944
timestamp 1624857261
transform 1 0 154224 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5943
timestamp 1624857261
transform 1 0 159256 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5942
timestamp 1624857261
transform 1 0 164288 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5941
timestamp 1624857261
transform 1 0 169184 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5940
timestamp 1624857261
transform 1 0 174216 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5939
timestamp 1624857261
transform 1 0 179248 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5938
timestamp 1624857261
transform 1 0 184280 0 1 17549
box 0 0 1 1
use contact_32  contact_32_5937
timestamp 1624857261
transform 1 0 544 0 1 14149
box 0 0 1 1
use contact_32  contact_32_5936
timestamp 1624857261
transform 1 0 544 0 1 18365
box 0 0 1 1
use contact_32  contact_32_5935
timestamp 1624857261
transform 1 0 544 0 1 26661
box 0 0 1 1
use contact_32  contact_32_5934
timestamp 1624857261
transform 1 0 544 0 1 23805
box 0 0 1 1
use contact_32  contact_32_5933
timestamp 1624857261
transform 1 0 544 0 1 20949
box 0 0 1 1
use contact_32  contact_32_5932
timestamp 1624857261
transform 1 0 544 0 1 29653
box 0 0 1 1
use contact_32  contact_32_5931
timestamp 1624857261
transform 1 0 14552 0 1 41485
box 0 0 1 1
use contact_32  contact_32_5930
timestamp 1624857261
transform 1 0 14552 0 1 44069
box 0 0 1 1
use contact_32  contact_32_5929
timestamp 1624857261
transform 1 0 14552 0 1 41213
box 0 0 1 1
use contact_32  contact_32_5928
timestamp 1624857261
transform 1 0 14552 0 1 38629
box 0 0 1 1
use contact_32  contact_32_5927
timestamp 1624857261
transform 1 0 14552 0 1 35773
box 0 0 1 1
use contact_32  contact_32_5926
timestamp 1624857261
transform 1 0 14552 0 1 38493
box 0 0 1 1
use contact_32  contact_32_5925
timestamp 1624857261
transform 1 0 18496 0 1 35637
box 0 0 1 1
use contact_32  contact_32_5924
timestamp 1624857261
transform 1 0 18496 0 1 34005
box 0 0 1 1
use contact_32  contact_32_5923
timestamp 1624857261
transform 1 0 15096 0 1 19725
box 0 0 1 1
use contact_32  contact_32_5922
timestamp 1624857261
transform 1 0 15096 0 1 22445
box 0 0 1 1
use contact_32  contact_32_5921
timestamp 1624857261
transform 1 0 15096 0 1 19589
box 0 0 1 1
use contact_32  contact_32_5920
timestamp 1624857261
transform 1 0 15096 0 1 16869
box 0 0 1 1
use contact_32  contact_32_5919
timestamp 1624857261
transform 1 0 15096 0 1 14013
box 0 0 1 1
use contact_32  contact_32_5918
timestamp 1624857261
transform 1 0 15096 0 1 16733
box 0 0 1 1
use contact_32  contact_32_5917
timestamp 1624857261
transform 1 0 17544 0 1 22581
box 0 0 1 1
use contact_32  contact_32_5916
timestamp 1624857261
transform 1 0 17544 0 1 25165
box 0 0 1 1
use contact_32  contact_32_5915
timestamp 1624857261
transform 1 0 16864 0 1 3541
box 0 0 1 1
use contact_32  contact_32_5914
timestamp 1624857261
transform 1 0 16864 0 1 549
box 0 0 1 1
use contact_32  contact_32_5913
timestamp 1624857261
transform 1 0 18904 0 1 28565
box 0 0 1 1
use contact_32  contact_32_5912
timestamp 1624857261
transform 1 0 18904 0 1 29109
box 0 0 1 1
use contact_32  contact_32_5911
timestamp 1624857261
transform 1 0 18768 0 1 29925
box 0 0 1 1
use contact_32  contact_32_5910
timestamp 1624857261
transform 1 0 18904 0 1 29245
box 0 0 1 1
use contact_32  contact_32_5909
timestamp 1624857261
transform 1 0 18768 0 1 33053
box 0 0 1 1
use contact_32  contact_32_5908
timestamp 1624857261
transform 1 0 18904 0 1 32373
box 0 0 1 1
use contact_32  contact_32_5907
timestamp 1624857261
transform 1 0 19040 0 1 28293
box 0 0 1 1
use contact_32  contact_32_5906
timestamp 1624857261
transform 1 0 19040 0 1 27613
box 0 0 1 1
use contact_32  contact_32_5905
timestamp 1624857261
transform 1 0 18904 0 1 32237
box 0 0 1 1
use contact_32  contact_32_5904
timestamp 1624857261
transform 1 0 18904 0 1 31557
box 0 0 1 1
use contact_32  contact_32_5903
timestamp 1624857261
transform 1 0 18904 0 1 30061
box 0 0 1 1
use contact_32  contact_32_5902
timestamp 1624857261
transform 1 0 18904 0 1 31421
box 0 0 1 1
use contact_32  contact_32_5901
timestamp 1624857261
transform 1 0 18904 0 1 33189
box 0 0 1 1
use contact_32  contact_32_5900
timestamp 1624857261
transform 1 0 18904 0 1 33869
box 0 0 1 1
use contact_32  contact_32_5899
timestamp 1624857261
transform 1 0 19720 0 1 25437
box 0 0 1 1
use contact_32  contact_32_5898
timestamp 1624857261
transform 1 0 19720 0 1 25845
box 0 0 1 1
use contact_32  contact_32_5897
timestamp 1624857261
transform 1 0 19856 0 1 31557
box 0 0 1 1
use contact_32  contact_32_5896
timestamp 1624857261
transform 1 0 19856 0 1 32237
box 0 0 1 1
use contact_32  contact_32_5895
timestamp 1624857261
transform 1 0 19720 0 1 26117
box 0 0 1 1
use contact_32  contact_32_5894
timestamp 1624857261
transform 1 0 19720 0 1 27477
box 0 0 1 1
use contact_32  contact_32_5893
timestamp 1624857261
transform 1 0 19856 0 1 28293
box 0 0 1 1
use contact_32  contact_32_5892
timestamp 1624857261
transform 1 0 19856 0 1 27613
box 0 0 1 1
use contact_32  contact_32_5891
timestamp 1624857261
transform 1 0 19856 0 1 29925
box 0 0 1 1
use contact_32  contact_32_5890
timestamp 1624857261
transform 1 0 19856 0 1 29245
box 0 0 1 1
use contact_32  contact_32_5889
timestamp 1624857261
transform 1 0 22032 0 1 30197
box 0 0 1 1
use contact_32  contact_32_5888
timestamp 1624857261
transform 1 0 22032 0 1 30605
box 0 0 1 1
use contact_32  contact_32_5887
timestamp 1624857261
transform 1 0 20536 0 1 20813
box 0 0 1 1
use contact_32  contact_32_5886
timestamp 1624857261
transform 1 0 20536 0 1 18093
box 0 0 1 1
use contact_32  contact_32_5885
timestamp 1624857261
transform 1 0 20400 0 1 17957
box 0 0 1 1
use contact_32  contact_32_5884
timestamp 1624857261
transform 1 0 20400 0 1 15237
box 0 0 1 1
use contact_32  contact_32_5883
timestamp 1624857261
transform 1 0 21896 0 1 12381
box 0 0 1 1
use contact_32  contact_32_5882
timestamp 1624857261
transform 1 0 21896 0 1 15101
box 0 0 1 1
use contact_32  contact_32_5881
timestamp 1624857261
transform 1 0 23120 0 1 20949
box 0 0 1 1
use contact_32  contact_32_5880
timestamp 1624857261
transform 1 0 23120 0 1 24485
box 0 0 1 1
use contact_32  contact_32_5879
timestamp 1624857261
transform 1 0 22440 0 1 41757
box 0 0 1 1
use contact_32  contact_32_5878
timestamp 1624857261
transform 1 0 22440 0 1 41485
box 0 0 1 1
use contact_32  contact_32_5877
timestamp 1624857261
transform 1 0 22440 0 1 117645
box 0 0 1 1
use contact_32  contact_32_5876
timestamp 1624857261
transform 1 0 22440 0 1 117917
box 0 0 1 1
use contact_32  contact_32_5875
timestamp 1624857261
transform 1 0 22168 0 1 44205
box 0 0 1 1
use contact_32  contact_32_5874
timestamp 1624857261
transform 1 0 22168 0 1 44477
box 0 0 1 1
use contact_32  contact_32_5873
timestamp 1624857261
transform 1 0 22304 0 1 50053
box 0 0 1 1
use contact_32  contact_32_5872
timestamp 1624857261
transform 1 0 22304 0 1 49781
box 0 0 1 1
use contact_32  contact_32_5871
timestamp 1624857261
transform 1 0 22304 0 1 44885
box 0 0 1 1
use contact_32  contact_32_5870
timestamp 1624857261
transform 1 0 22304 0 1 44613
box 0 0 1 1
use contact_32  contact_32_5869
timestamp 1624857261
transform 1 0 22168 0 1 78205
box 0 0 1 1
use contact_32  contact_32_5868
timestamp 1624857261
transform 1 0 22168 0 1 78477
box 0 0 1 1
use contact_32  contact_32_5867
timestamp 1624857261
transform 1 0 22304 0 1 116557
box 0 0 1 1
use contact_32  contact_32_5866
timestamp 1624857261
transform 1 0 22304 0 1 116829
box 0 0 1 1
use contact_32  contact_32_5865
timestamp 1624857261
transform 1 0 22440 0 1 116557
box 0 0 1 1
use contact_32  contact_32_5864
timestamp 1624857261
transform 1 0 22440 0 1 116829
box 0 0 1 1
use contact_32  contact_32_5863
timestamp 1624857261
transform 1 0 22440 0 1 121997
box 0 0 1 1
use contact_32  contact_32_5862
timestamp 1624857261
transform 1 0 22440 0 1 121725
box 0 0 1 1
use contact_32  contact_32_5861
timestamp 1624857261
transform 1 0 22304 0 1 112069
box 0 0 1 1
use contact_32  contact_32_5860
timestamp 1624857261
transform 1 0 22304 0 1 111797
box 0 0 1 1
use contact_32  contact_32_5859
timestamp 1624857261
transform 1 0 22440 0 1 112069
box 0 0 1 1
use contact_32  contact_32_5858
timestamp 1624857261
transform 1 0 22440 0 1 111797
box 0 0 1 1
use contact_32  contact_32_5857
timestamp 1624857261
transform 1 0 22304 0 1 48149
box 0 0 1 1
use contact_32  contact_32_5856
timestamp 1624857261
transform 1 0 22304 0 1 48421
box 0 0 1 1
use contact_32  contact_32_5855
timestamp 1624857261
transform 1 0 22304 0 1 90309
box 0 0 1 1
use contact_32  contact_32_5854
timestamp 1624857261
transform 1 0 22304 0 1 90037
box 0 0 1 1
use contact_32  contact_32_5853
timestamp 1624857261
transform 1 0 22168 0 1 25709
box 0 0 1 1
use contact_32  contact_32_5852
timestamp 1624857261
transform 1 0 22168 0 1 25981
box 0 0 1 1
use contact_32  contact_32_5851
timestamp 1624857261
transform 1 0 22304 0 1 63109
box 0 0 1 1
use contact_32  contact_32_5850
timestamp 1624857261
transform 1 0 22304 0 1 62837
box 0 0 1 1
use contact_32  contact_32_5849
timestamp 1624857261
transform 1 0 22440 0 1 63109
box 0 0 1 1
use contact_32  contact_32_5848
timestamp 1624857261
transform 1 0 22440 0 1 62837
box 0 0 1 1
use contact_32  contact_32_5847
timestamp 1624857261
transform 1 0 22440 0 1 53181
box 0 0 1 1
use contact_32  contact_32_5846
timestamp 1624857261
transform 1 0 22440 0 1 52909
box 0 0 1 1
use contact_32  contact_32_5845
timestamp 1624857261
transform 1 0 22304 0 1 84053
box 0 0 1 1
use contact_32  contact_32_5844
timestamp 1624857261
transform 1 0 22304 0 1 84325
box 0 0 1 1
use contact_32  contact_32_5843
timestamp 1624857261
transform 1 0 22440 0 1 84053
box 0 0 1 1
use contact_32  contact_32_5842
timestamp 1624857261
transform 1 0 22440 0 1 84325
box 0 0 1 1
use contact_32  contact_32_5841
timestamp 1624857261
transform 1 0 22168 0 1 60797
box 0 0 1 1
use contact_32  contact_32_5840
timestamp 1624857261
transform 1 0 22168 0 1 61069
box 0 0 1 1
use contact_32  contact_32_5839
timestamp 1624857261
transform 1 0 22168 0 1 111661
box 0 0 1 1
use contact_32  contact_32_5838
timestamp 1624857261
transform 1 0 22168 0 1 111389
box 0 0 1 1
use contact_32  contact_32_5837
timestamp 1624857261
transform 1 0 22440 0 1 124309
box 0 0 1 1
use contact_32  contact_32_5836
timestamp 1624857261
transform 1 0 22440 0 1 124037
box 0 0 1 1
use contact_32  contact_32_5835
timestamp 1624857261
transform 1 0 22168 0 1 32237
box 0 0 1 1
use contact_32  contact_32_5834
timestamp 1624857261
transform 1 0 22168 0 1 31965
box 0 0 1 1
use contact_32  contact_32_5833
timestamp 1624857261
transform 1 0 22168 0 1 123629
box 0 0 1 1
use contact_32  contact_32_5832
timestamp 1624857261
transform 1 0 22168 0 1 123901
box 0 0 1 1
use contact_32  contact_32_5831
timestamp 1624857261
transform 1 0 22304 0 1 102685
box 0 0 1 1
use contact_32  contact_32_5830
timestamp 1624857261
transform 1 0 22304 0 1 102957
box 0 0 1 1
use contact_32  contact_32_5829
timestamp 1624857261
transform 1 0 22440 0 1 102549
box 0 0 1 1
use contact_32  contact_32_5828
timestamp 1624857261
transform 1 0 22440 0 1 102277
box 0 0 1 1
use contact_32  contact_32_5827
timestamp 1624857261
transform 1 0 22440 0 1 33053
box 0 0 1 1
use contact_32  contact_32_5826
timestamp 1624857261
transform 1 0 22440 0 1 32781
box 0 0 1 1
use contact_32  contact_32_5825
timestamp 1624857261
transform 1 0 22168 0 1 116013
box 0 0 1 1
use contact_32  contact_32_5824
timestamp 1624857261
transform 1 0 22168 0 1 115741
box 0 0 1 1
use contact_32  contact_32_5823
timestamp 1624857261
transform 1 0 22168 0 1 105405
box 0 0 1 1
use contact_32  contact_32_5822
timestamp 1624857261
transform 1 0 22168 0 1 105677
box 0 0 1 1
use contact_32  contact_32_5821
timestamp 1624857261
transform 1 0 22168 0 1 34413
box 0 0 1 1
use contact_32  contact_32_5820
timestamp 1624857261
transform 1 0 22168 0 1 34685
box 0 0 1 1
use contact_32  contact_32_5819
timestamp 1624857261
transform 1 0 22304 0 1 86365
box 0 0 1 1
use contact_32  contact_32_5818
timestamp 1624857261
transform 1 0 22304 0 1 86093
box 0 0 1 1
use contact_32  contact_32_5817
timestamp 1624857261
transform 1 0 22304 0 1 94661
box 0 0 1 1
use contact_32  contact_32_5816
timestamp 1624857261
transform 1 0 22304 0 1 94389
box 0 0 1 1
use contact_32  contact_32_5815
timestamp 1624857261
transform 1 0 22440 0 1 94661
box 0 0 1 1
use contact_32  contact_32_5814
timestamp 1624857261
transform 1 0 22440 0 1 94389
box 0 0 1 1
use contact_32  contact_32_5813
timestamp 1624857261
transform 1 0 22168 0 1 61613
box 0 0 1 1
use contact_32  contact_32_5812
timestamp 1624857261
transform 1 0 22168 0 1 61885
box 0 0 1 1
use contact_32  contact_32_5811
timestamp 1624857261
transform 1 0 22168 0 1 27885
box 0 0 1 1
use contact_32  contact_32_5810
timestamp 1624857261
transform 1 0 22168 0 1 27613
box 0 0 1 1
use contact_32  contact_32_5809
timestamp 1624857261
transform 1 0 22440 0 1 42981
box 0 0 1 1
use contact_32  contact_32_5808
timestamp 1624857261
transform 1 0 22440 0 1 43253
box 0 0 1 1
use contact_32  contact_32_5807
timestamp 1624857261
transform 1 0 22168 0 1 48557
box 0 0 1 1
use contact_32  contact_32_5806
timestamp 1624857261
transform 1 0 22168 0 1 48829
box 0 0 1 1
use contact_32  contact_32_5805
timestamp 1624857261
transform 1 0 22168 0 1 110845
box 0 0 1 1
use contact_32  contact_32_5804
timestamp 1624857261
transform 1 0 22168 0 1 110573
box 0 0 1 1
use contact_32  contact_32_5803
timestamp 1624857261
transform 1 0 22168 0 1 33597
box 0 0 1 1
use contact_32  contact_32_5802
timestamp 1624857261
transform 1 0 22168 0 1 33869
box 0 0 1 1
use contact_32  contact_32_5801
timestamp 1624857261
transform 1 0 22168 0 1 85549
box 0 0 1 1
use contact_32  contact_32_5800
timestamp 1624857261
transform 1 0 22168 0 1 85277
box 0 0 1 1
use contact_32  contact_32_5799
timestamp 1624857261
transform 1 0 22168 0 1 75757
box 0 0 1 1
use contact_32  contact_32_5798
timestamp 1624857261
transform 1 0 22168 0 1 75485
box 0 0 1 1
use contact_32  contact_32_5797
timestamp 1624857261
transform 1 0 22304 0 1 40533
box 0 0 1 1
use contact_32  contact_32_5796
timestamp 1624857261
transform 1 0 22304 0 1 40261
box 0 0 1 1
use contact_32  contact_32_5795
timestamp 1624857261
transform 1 0 22168 0 1 97517
box 0 0 1 1
use contact_32  contact_32_5794
timestamp 1624857261
transform 1 0 22168 0 1 97789
box 0 0 1 1
use contact_32  contact_32_5793
timestamp 1624857261
transform 1 0 22304 0 1 81605
box 0 0 1 1
use contact_32  contact_32_5792
timestamp 1624857261
transform 1 0 22304 0 1 81333
box 0 0 1 1
use contact_32  contact_32_5791
timestamp 1624857261
transform 1 0 22440 0 1 81605
box 0 0 1 1
use contact_32  contact_32_5790
timestamp 1624857261
transform 1 0 22440 0 1 81333
box 0 0 1 1
use contact_32  contact_32_5789
timestamp 1624857261
transform 1 0 22440 0 1 91533
box 0 0 1 1
use contact_32  contact_32_5788
timestamp 1624857261
transform 1 0 22440 0 1 91805
box 0 0 1 1
use contact_32  contact_32_5787
timestamp 1624857261
transform 1 0 22304 0 1 79701
box 0 0 1 1
use contact_32  contact_32_5786
timestamp 1624857261
transform 1 0 22304 0 1 79429
box 0 0 1 1
use contact_32  contact_32_5785
timestamp 1624857261
transform 1 0 22440 0 1 79701
box 0 0 1 1
use contact_32  contact_32_5784
timestamp 1624857261
transform 1 0 22440 0 1 79429
box 0 0 1 1
use contact_32  contact_32_5783
timestamp 1624857261
transform 1 0 22168 0 1 107309
box 0 0 1 1
use contact_32  contact_32_5782
timestamp 1624857261
transform 1 0 22168 0 1 107037
box 0 0 1 1
use contact_32  contact_32_5781
timestamp 1624857261
transform 1 0 22304 0 1 83645
box 0 0 1 1
use contact_32  contact_32_5780
timestamp 1624857261
transform 1 0 22304 0 1 83373
box 0 0 1 1
use contact_32  contact_32_5779
timestamp 1624857261
transform 1 0 22168 0 1 37541
box 0 0 1 1
use contact_32  contact_32_5778
timestamp 1624857261
transform 1 0 22168 0 1 37813
box 0 0 1 1
use contact_32  contact_32_5777
timestamp 1624857261
transform 1 0 22168 0 1 26661
box 0 0 1 1
use contact_32  contact_32_5776
timestamp 1624857261
transform 1 0 22168 0 1 26389
box 0 0 1 1
use contact_32  contact_32_5775
timestamp 1624857261
transform 1 0 22168 0 1 30333
box 0 0 1 1
use contact_32  contact_32_5774
timestamp 1624857261
transform 1 0 22168 0 1 30605
box 0 0 1 1
use contact_32  contact_32_5773
timestamp 1624857261
transform 1 0 22168 0 1 49645
box 0 0 1 1
use contact_32  contact_32_5772
timestamp 1624857261
transform 1 0 22168 0 1 49373
box 0 0 1 1
use contact_32  contact_32_5771
timestamp 1624857261
transform 1 0 22168 0 1 57261
box 0 0 1 1
use contact_32  contact_32_5770
timestamp 1624857261
transform 1 0 22168 0 1 57533
box 0 0 1 1
use contact_32  contact_32_5769
timestamp 1624857261
transform 1 0 22304 0 1 31557
box 0 0 1 1
use contact_32  contact_32_5768
timestamp 1624857261
transform 1 0 22304 0 1 31829
box 0 0 1 1
use contact_32  contact_32_5767
timestamp 1624857261
transform 1 0 22440 0 1 31557
box 0 0 1 1
use contact_32  contact_32_5766
timestamp 1624857261
transform 1 0 22440 0 1 31829
box 0 0 1 1
use contact_32  contact_32_5765
timestamp 1624857261
transform 1 0 22304 0 1 35093
box 0 0 1 1
use contact_32  contact_32_5764
timestamp 1624857261
transform 1 0 22304 0 1 35365
box 0 0 1 1
use contact_32  contact_32_5763
timestamp 1624857261
transform 1 0 22440 0 1 35093
box 0 0 1 1
use contact_32  contact_32_5762
timestamp 1624857261
transform 1 0 22440 0 1 35365
box 0 0 1 1
use contact_32  contact_32_5761
timestamp 1624857261
transform 1 0 22304 0 1 101461
box 0 0 1 1
use contact_32  contact_32_5760
timestamp 1624857261
transform 1 0 22304 0 1 101733
box 0 0 1 1
use contact_32  contact_32_5759
timestamp 1624857261
transform 1 0 22440 0 1 101461
box 0 0 1 1
use contact_32  contact_32_5758
timestamp 1624857261
transform 1 0 22440 0 1 101733
box 0 0 1 1
use contact_32  contact_32_5757
timestamp 1624857261
transform 1 0 22440 0 1 109757
box 0 0 1 1
use contact_32  contact_32_5756
timestamp 1624857261
transform 1 0 22440 0 1 110029
box 0 0 1 1
use contact_32  contact_32_5755
timestamp 1624857261
transform 1 0 22440 0 1 43797
box 0 0 1 1
use contact_32  contact_32_5754
timestamp 1624857261
transform 1 0 22440 0 1 44069
box 0 0 1 1
use contact_32  contact_32_5753
timestamp 1624857261
transform 1 0 22168 0 1 114925
box 0 0 1 1
use contact_32  contact_32_5752
timestamp 1624857261
transform 1 0 22168 0 1 115197
box 0 0 1 1
use contact_32  contact_32_5751
timestamp 1624857261
transform 1 0 22304 0 1 77253
box 0 0 1 1
use contact_32  contact_32_5750
timestamp 1624857261
transform 1 0 22304 0 1 76981
box 0 0 1 1
use contact_32  contact_32_5749
timestamp 1624857261
transform 1 0 22168 0 1 98605
box 0 0 1 1
use contact_32  contact_32_5748
timestamp 1624857261
transform 1 0 22168 0 1 98333
box 0 0 1 1
use contact_32  contact_32_5747
timestamp 1624857261
transform 1 0 22168 0 1 73853
box 0 0 1 1
use contact_32  contact_32_5746
timestamp 1624857261
transform 1 0 22168 0 1 74125
box 0 0 1 1
use contact_32  contact_32_5745
timestamp 1624857261
transform 1 0 22168 0 1 40125
box 0 0 1 1
use contact_32  contact_32_5744
timestamp 1624857261
transform 1 0 22168 0 1 39853
box 0 0 1 1
use contact_32  contact_32_5743
timestamp 1624857261
transform 1 0 22440 0 1 40125
box 0 0 1 1
use contact_32  contact_32_5742
timestamp 1624857261
transform 1 0 22440 0 1 39853
box 0 0 1 1
use contact_32  contact_32_5741
timestamp 1624857261
transform 1 0 22304 0 1 36997
box 0 0 1 1
use contact_32  contact_32_5740
timestamp 1624857261
transform 1 0 22304 0 1 36725
box 0 0 1 1
use contact_32  contact_32_5739
timestamp 1624857261
transform 1 0 22168 0 1 89901
box 0 0 1 1
use contact_32  contact_32_5738
timestamp 1624857261
transform 1 0 22168 0 1 89629
box 0 0 1 1
use contact_32  contact_32_5737
timestamp 1624857261
transform 1 0 22304 0 1 49237
box 0 0 1 1
use contact_32  contact_32_5736
timestamp 1624857261
transform 1 0 22304 0 1 48965
box 0 0 1 1
use contact_32  contact_32_5735
timestamp 1624857261
transform 1 0 22304 0 1 69773
box 0 0 1 1
use contact_32  contact_32_5734
timestamp 1624857261
transform 1 0 22304 0 1 69501
box 0 0 1 1
use contact_32  contact_32_5733
timestamp 1624857261
transform 1 0 22304 0 1 69909
box 0 0 1 1
use contact_32  contact_32_5732
timestamp 1624857261
transform 1 0 22304 0 1 70181
box 0 0 1 1
use contact_32  contact_32_5731
timestamp 1624857261
transform 1 0 22304 0 1 52501
box 0 0 1 1
use contact_32  contact_32_5730
timestamp 1624857261
transform 1 0 22304 0 1 52773
box 0 0 1 1
use contact_32  contact_32_5729
timestamp 1624857261
transform 1 0 22304 0 1 118869
box 0 0 1 1
use contact_32  contact_32_5728
timestamp 1624857261
transform 1 0 22304 0 1 119141
box 0 0 1 1
use contact_32  contact_32_5727
timestamp 1624857261
transform 1 0 22304 0 1 41349
box 0 0 1 1
use contact_32  contact_32_5726
timestamp 1624857261
transform 1 0 22304 0 1 41077
box 0 0 1 1
use contact_32  contact_32_5725
timestamp 1624857261
transform 1 0 22168 0 1 120365
box 0 0 1 1
use contact_32  contact_32_5724
timestamp 1624857261
transform 1 0 22168 0 1 120093
box 0 0 1 1
use contact_32  contact_32_5723
timestamp 1624857261
transform 1 0 22440 0 1 108941
box 0 0 1 1
use contact_32  contact_32_5722
timestamp 1624857261
transform 1 0 22440 0 1 108669
box 0 0 1 1
use contact_32  contact_32_5721
timestamp 1624857261
transform 1 0 22168 0 1 73309
box 0 0 1 1
use contact_32  contact_32_5720
timestamp 1624857261
transform 1 0 22168 0 1 73037
box 0 0 1 1
use contact_32  contact_32_5719
timestamp 1624857261
transform 1 0 22304 0 1 53725
box 0 0 1 1
use contact_32  contact_32_5718
timestamp 1624857261
transform 1 0 22304 0 1 53997
box 0 0 1 1
use contact_32  contact_32_5717
timestamp 1624857261
transform 1 0 22304 0 1 125261
box 0 0 1 1
use contact_32  contact_32_5716
timestamp 1624857261
transform 1 0 22304 0 1 125533
box 0 0 1 1
use contact_32  contact_32_5715
timestamp 1624857261
transform 1 0 22440 0 1 125261
box 0 0 1 1
use contact_32  contact_32_5714
timestamp 1624857261
transform 1 0 22440 0 1 125533
box 0 0 1 1
use contact_32  contact_32_5713
timestamp 1624857261
transform 1 0 22304 0 1 106901
box 0 0 1 1
use contact_32  contact_32_5712
timestamp 1624857261
transform 1 0 22304 0 1 106629
box 0 0 1 1
use contact_32  contact_32_5711
timestamp 1624857261
transform 1 0 22304 0 1 96021
box 0 0 1 1
use contact_32  contact_32_5710
timestamp 1624857261
transform 1 0 22304 0 1 96293
box 0 0 1 1
use contact_32  contact_32_5709
timestamp 1624857261
transform 1 0 22304 0 1 93845
box 0 0 1 1
use contact_32  contact_32_5708
timestamp 1624857261
transform 1 0 22304 0 1 93573
box 0 0 1 1
use contact_32  contact_32_5707
timestamp 1624857261
transform 1 0 22304 0 1 71813
box 0 0 1 1
use contact_32  contact_32_5706
timestamp 1624857261
transform 1 0 22304 0 1 71541
box 0 0 1 1
use contact_32  contact_32_5705
timestamp 1624857261
transform 1 0 22440 0 1 71813
box 0 0 1 1
use contact_32  contact_32_5704
timestamp 1624857261
transform 1 0 22440 0 1 71541
box 0 0 1 1
use contact_32  contact_32_5703
timestamp 1624857261
transform 1 0 22168 0 1 86909
box 0 0 1 1
use contact_32  contact_32_5702
timestamp 1624857261
transform 1 0 22168 0 1 87181
box 0 0 1 1
use contact_32  contact_32_5701
timestamp 1624857261
transform 1 0 22440 0 1 36181
box 0 0 1 1
use contact_32  contact_32_5700
timestamp 1624857261
transform 1 0 22440 0 1 35909
box 0 0 1 1
use contact_32  contact_32_5699
timestamp 1624857261
transform 1 0 22304 0 1 119957
box 0 0 1 1
use contact_32  contact_32_5698
timestamp 1624857261
transform 1 0 22304 0 1 119685
box 0 0 1 1
use contact_32  contact_32_5697
timestamp 1624857261
transform 1 0 22168 0 1 110437
box 0 0 1 1
use contact_32  contact_32_5696
timestamp 1624857261
transform 1 0 22168 0 1 110165
box 0 0 1 1
use contact_32  contact_32_5695
timestamp 1624857261
transform 1 0 22304 0 1 98197
box 0 0 1 1
use contact_32  contact_32_5694
timestamp 1624857261
transform 1 0 22304 0 1 97925
box 0 0 1 1
use contact_32  contact_32_5693
timestamp 1624857261
transform 1 0 22440 0 1 98197
box 0 0 1 1
use contact_32  contact_32_5692
timestamp 1624857261
transform 1 0 22440 0 1 97925
box 0 0 1 1
use contact_32  contact_32_5691
timestamp 1624857261
transform 1 0 22168 0 1 114109
box 0 0 1 1
use contact_32  contact_32_5690
timestamp 1624857261
transform 1 0 22168 0 1 114381
box 0 0 1 1
use contact_32  contact_32_5689
timestamp 1624857261
transform 1 0 22168 0 1 65965
box 0 0 1 1
use contact_32  contact_32_5688
timestamp 1624857261
transform 1 0 22168 0 1 66237
box 0 0 1 1
use contact_32  contact_32_5687
timestamp 1624857261
transform 1 0 22304 0 1 68549
box 0 0 1 1
use contact_32  contact_32_5686
timestamp 1624857261
transform 1 0 22304 0 1 68277
box 0 0 1 1
use contact_32  contact_32_5685
timestamp 1624857261
transform 1 0 22168 0 1 65149
box 0 0 1 1
use contact_32  contact_32_5684
timestamp 1624857261
transform 1 0 22168 0 1 65421
box 0 0 1 1
use contact_32  contact_32_5683
timestamp 1624857261
transform 1 0 22168 0 1 56445
box 0 0 1 1
use contact_32  contact_32_5682
timestamp 1624857261
transform 1 0 22168 0 1 56717
box 0 0 1 1
use contact_32  contact_32_5681
timestamp 1624857261
transform 1 0 22440 0 1 26389
box 0 0 1 1
use contact_32  contact_32_5680
timestamp 1624857261
transform 1 0 22440 0 1 26661
box 0 0 1 1
use contact_32  contact_32_5679
timestamp 1624857261
transform 1 0 22168 0 1 39037
box 0 0 1 1
use contact_32  contact_32_5678
timestamp 1624857261
transform 1 0 22168 0 1 39309
box 0 0 1 1
use contact_32  contact_32_5677
timestamp 1624857261
transform 1 0 22440 0 1 77661
box 0 0 1 1
use contact_32  contact_32_5676
timestamp 1624857261
transform 1 0 22440 0 1 77389
box 0 0 1 1
use contact_32  contact_32_5675
timestamp 1624857261
transform 1 0 22168 0 1 45429
box 0 0 1 1
use contact_32  contact_32_5674
timestamp 1624857261
transform 1 0 22168 0 1 45701
box 0 0 1 1
use contact_32  contact_32_5673
timestamp 1624857261
transform 1 0 22168 0 1 90853
box 0 0 1 1
use contact_32  contact_32_5672
timestamp 1624857261
transform 1 0 22168 0 1 91125
box 0 0 1 1
use contact_32  contact_32_5671
timestamp 1624857261
transform 1 0 22168 0 1 88133
box 0 0 1 1
use contact_32  contact_32_5670
timestamp 1624857261
transform 1 0 22168 0 1 88405
box 0 0 1 1
use contact_32  contact_32_5669
timestamp 1624857261
transform 1 0 22440 0 1 88133
box 0 0 1 1
use contact_32  contact_32_5668
timestamp 1624857261
transform 1 0 22440 0 1 88405
box 0 0 1 1
use contact_32  contact_32_5667
timestamp 1624857261
transform 1 0 22168 0 1 100917
box 0 0 1 1
use contact_32  contact_32_5666
timestamp 1624857261
transform 1 0 22168 0 1 100645
box 0 0 1 1
use contact_32  contact_32_5665
timestamp 1624857261
transform 1 0 22304 0 1 29517
box 0 0 1 1
use contact_32  contact_32_5664
timestamp 1624857261
transform 1 0 22304 0 1 29245
box 0 0 1 1
use contact_32  contact_32_5663
timestamp 1624857261
transform 1 0 22440 0 1 29653
box 0 0 1 1
use contact_32  contact_32_5662
timestamp 1624857261
transform 1 0 22440 0 1 29925
box 0 0 1 1
use contact_32  contact_32_5661
timestamp 1624857261
transform 1 0 22304 0 1 27477
box 0 0 1 1
use contact_32  contact_32_5660
timestamp 1624857261
transform 1 0 22304 0 1 27205
box 0 0 1 1
use contact_32  contact_32_5659
timestamp 1624857261
transform 1 0 22304 0 1 122405
box 0 0 1 1
use contact_32  contact_32_5658
timestamp 1624857261
transform 1 0 22304 0 1 122677
box 0 0 1 1
use contact_32  contact_32_5657
timestamp 1624857261
transform 1 0 22304 0 1 85141
box 0 0 1 1
use contact_32  contact_32_5656
timestamp 1624857261
transform 1 0 22304 0 1 84869
box 0 0 1 1
use contact_32  contact_32_5655
timestamp 1624857261
transform 1 0 22168 0 1 106221
box 0 0 1 1
use contact_32  contact_32_5654
timestamp 1624857261
transform 1 0 22168 0 1 106493
box 0 0 1 1
use contact_32  contact_32_5653
timestamp 1624857261
transform 1 0 22440 0 1 104725
box 0 0 1 1
use contact_32  contact_32_5652
timestamp 1624857261
transform 1 0 22440 0 1 104997
box 0 0 1 1
use contact_32  contact_32_5651
timestamp 1624857261
transform 1 0 22168 0 1 118053
box 0 0 1 1
use contact_32  contact_32_5650
timestamp 1624857261
transform 1 0 22168 0 1 118325
box 0 0 1 1
use contact_32  contact_32_5649
timestamp 1624857261
transform 1 0 22440 0 1 114517
box 0 0 1 1
use contact_32  contact_32_5648
timestamp 1624857261
transform 1 0 22440 0 1 114789
box 0 0 1 1
use contact_32  contact_32_5647
timestamp 1624857261
transform 1 0 22440 0 1 107717
box 0 0 1 1
use contact_32  contact_32_5646
timestamp 1624857261
transform 1 0 22440 0 1 107445
box 0 0 1 1
use contact_32  contact_32_5645
timestamp 1624857261
transform 1 0 22440 0 1 92349
box 0 0 1 1
use contact_32  contact_32_5644
timestamp 1624857261
transform 1 0 22440 0 1 92077
box 0 0 1 1
use contact_32  contact_32_5643
timestamp 1624857261
transform 1 0 22440 0 1 110165
box 0 0 1 1
use contact_32  contact_32_5642
timestamp 1624857261
transform 1 0 22440 0 1 110437
box 0 0 1 1
use contact_32  contact_32_5641
timestamp 1624857261
transform 1 0 22304 0 1 87317
box 0 0 1 1
use contact_32  contact_32_5640
timestamp 1624857261
transform 1 0 22304 0 1 87589
box 0 0 1 1
use contact_32  contact_32_5639
timestamp 1624857261
transform 1 0 22440 0 1 87317
box 0 0 1 1
use contact_32  contact_32_5638
timestamp 1624857261
transform 1 0 22440 0 1 87589
box 0 0 1 1
use contact_32  contact_32_5637
timestamp 1624857261
transform 1 0 22440 0 1 87181
box 0 0 1 1
use contact_32  contact_32_5636
timestamp 1624857261
transform 1 0 22440 0 1 86909
box 0 0 1 1
use contact_32  contact_32_5635
timestamp 1624857261
transform 1 0 22440 0 1 39309
box 0 0 1 1
use contact_32  contact_32_5634
timestamp 1624857261
transform 1 0 22440 0 1 39037
box 0 0 1 1
use contact_32  contact_32_5633
timestamp 1624857261
transform 1 0 22304 0 1 123085
box 0 0 1 1
use contact_32  contact_32_5632
timestamp 1624857261
transform 1 0 22304 0 1 122813
box 0 0 1 1
use contact_32  contact_32_5631
timestamp 1624857261
transform 1 0 22440 0 1 123221
box 0 0 1 1
use contact_32  contact_32_5630
timestamp 1624857261
transform 1 0 22440 0 1 123493
box 0 0 1 1
use contact_32  contact_32_5629
timestamp 1624857261
transform 1 0 22440 0 1 123085
box 0 0 1 1
use contact_32  contact_32_5628
timestamp 1624857261
transform 1 0 22440 0 1 122813
box 0 0 1 1
use contact_32  contact_32_5627
timestamp 1624857261
transform 1 0 22304 0 1 76437
box 0 0 1 1
use contact_32  contact_32_5626
timestamp 1624857261
transform 1 0 22304 0 1 76165
box 0 0 1 1
use contact_32  contact_32_5625
timestamp 1624857261
transform 1 0 22440 0 1 76437
box 0 0 1 1
use contact_32  contact_32_5624
timestamp 1624857261
transform 1 0 22440 0 1 76165
box 0 0 1 1
use contact_32  contact_32_5623
timestamp 1624857261
transform 1 0 22440 0 1 80109
box 0 0 1 1
use contact_32  contact_32_5622
timestamp 1624857261
transform 1 0 22440 0 1 80381
box 0 0 1 1
use contact_32  contact_32_5621
timestamp 1624857261
transform 1 0 22440 0 1 65421
box 0 0 1 1
use contact_32  contact_32_5620
timestamp 1624857261
transform 1 0 22440 0 1 65149
box 0 0 1 1
use contact_32  contact_32_5619
timestamp 1624857261
transform 1 0 22440 0 1 64605
box 0 0 1 1
use contact_32  contact_32_5618
timestamp 1624857261
transform 1 0 22440 0 1 64333
box 0 0 1 1
use contact_32  contact_32_5617
timestamp 1624857261
transform 1 0 22440 0 1 54405
box 0 0 1 1
use contact_32  contact_32_5616
timestamp 1624857261
transform 1 0 22440 0 1 54133
box 0 0 1 1
use contact_32  contact_32_5615
timestamp 1624857261
transform 1 0 22304 0 1 28429
box 0 0 1 1
use contact_32  contact_32_5614
timestamp 1624857261
transform 1 0 22304 0 1 28701
box 0 0 1 1
use contact_32  contact_32_5613
timestamp 1624857261
transform 1 0 22440 0 1 28293
box 0 0 1 1
use contact_32  contact_32_5612
timestamp 1624857261
transform 1 0 22440 0 1 28021
box 0 0 1 1
use contact_32  contact_32_5611
timestamp 1624857261
transform 1 0 22440 0 1 120773
box 0 0 1 1
use contact_32  contact_32_5610
timestamp 1624857261
transform 1 0 22440 0 1 120501
box 0 0 1 1
use contact_32  contact_32_5609
timestamp 1624857261
transform 1 0 22440 0 1 67597
box 0 0 1 1
use contact_32  contact_32_5608
timestamp 1624857261
transform 1 0 22440 0 1 67869
box 0 0 1 1
use contact_32  contact_32_5607
timestamp 1624857261
transform 1 0 22440 0 1 111253
box 0 0 1 1
use contact_32  contact_32_5606
timestamp 1624857261
transform 1 0 22440 0 1 110981
box 0 0 1 1
use contact_32  contact_32_5605
timestamp 1624857261
transform 1 0 22440 0 1 100237
box 0 0 1 1
use contact_32  contact_32_5604
timestamp 1624857261
transform 1 0 22440 0 1 99965
box 0 0 1 1
use contact_32  contact_32_5603
timestamp 1624857261
transform 1 0 22168 0 1 89085
box 0 0 1 1
use contact_32  contact_32_5602
timestamp 1624857261
transform 1 0 22168 0 1 88813
box 0 0 1 1
use contact_32  contact_32_5601
timestamp 1624857261
transform 1 0 22168 0 1 121589
box 0 0 1 1
use contact_32  contact_32_5600
timestamp 1624857261
transform 1 0 22168 0 1 121317
box 0 0 1 1
use contact_32  contact_32_5599
timestamp 1624857261
transform 1 0 22168 0 1 113565
box 0 0 1 1
use contact_32  contact_32_5598
timestamp 1624857261
transform 1 0 22168 0 1 113293
box 0 0 1 1
use contact_32  contact_32_5597
timestamp 1624857261
transform 1 0 22440 0 1 103365
box 0 0 1 1
use contact_32  contact_32_5596
timestamp 1624857261
transform 1 0 22440 0 1 103093
box 0 0 1 1
use contact_32  contact_32_5595
timestamp 1624857261
transform 1 0 22440 0 1 46925
box 0 0 1 1
use contact_32  contact_32_5594
timestamp 1624857261
transform 1 0 22440 0 1 47197
box 0 0 1 1
use contact_32  contact_32_5593
timestamp 1624857261
transform 1 0 22304 0 1 46789
box 0 0 1 1
use contact_32  contact_32_5592
timestamp 1624857261
transform 1 0 22440 0 1 46653
box 0 0 1 1
use contact_32  contact_32_5591
timestamp 1624857261
transform 1 0 22440 0 1 75485
box 0 0 1 1
use contact_32  contact_32_5590
timestamp 1624857261
transform 1 0 22440 0 1 75757
box 0 0 1 1
use contact_32  contact_32_5589
timestamp 1624857261
transform 1 0 22168 0 1 74669
box 0 0 1 1
use contact_32  contact_32_5588
timestamp 1624857261
transform 1 0 22168 0 1 74941
box 0 0 1 1
use contact_32  contact_32_5587
timestamp 1624857261
transform 1 0 22304 0 1 66645
box 0 0 1 1
use contact_32  contact_32_5586
timestamp 1624857261
transform 1 0 22304 0 1 66373
box 0 0 1 1
use contact_32  contact_32_5585
timestamp 1624857261
transform 1 0 22304 0 1 115605
box 0 0 1 1
use contact_32  contact_32_5584
timestamp 1624857261
transform 1 0 22304 0 1 115333
box 0 0 1 1
use contact_32  contact_32_5583
timestamp 1624857261
transform 1 0 22440 0 1 115605
box 0 0 1 1
use contact_32  contact_32_5582
timestamp 1624857261
transform 1 0 22440 0 1 115333
box 0 0 1 1
use contact_32  contact_32_5581
timestamp 1624857261
transform 1 0 22440 0 1 51685
box 0 0 1 1
use contact_32  contact_32_5580
timestamp 1624857261
transform 1 0 22440 0 1 51957
box 0 0 1 1
use contact_32  contact_32_5579
timestamp 1624857261
transform 1 0 22440 0 1 80925
box 0 0 1 1
use contact_32  contact_32_5578
timestamp 1624857261
transform 1 0 22440 0 1 80653
box 0 0 1 1
use contact_32  contact_32_5577
timestamp 1624857261
transform 1 0 22440 0 1 42573
box 0 0 1 1
use contact_32  contact_32_5576
timestamp 1624857261
transform 1 0 22440 0 1 42845
box 0 0 1 1
use contact_32  contact_32_5575
timestamp 1624857261
transform 1 0 22440 0 1 115197
box 0 0 1 1
use contact_32  contact_32_5574
timestamp 1624857261
transform 1 0 22440 0 1 114925
box 0 0 1 1
use contact_32  contact_32_5573
timestamp 1624857261
transform 1 0 22168 0 1 82149
box 0 0 1 1
use contact_32  contact_32_5572
timestamp 1624857261
transform 1 0 22168 0 1 82421
box 0 0 1 1
use contact_32  contact_32_5571
timestamp 1624857261
transform 1 0 22440 0 1 66237
box 0 0 1 1
use contact_32  contact_32_5570
timestamp 1624857261
transform 1 0 22440 0 1 65965
box 0 0 1 1
use contact_32  contact_32_5569
timestamp 1624857261
transform 1 0 22440 0 1 119549
box 0 0 1 1
use contact_32  contact_32_5568
timestamp 1624857261
transform 1 0 22440 0 1 119277
box 0 0 1 1
use contact_32  contact_32_5567
timestamp 1624857261
transform 1 0 22440 0 1 70317
box 0 0 1 1
use contact_32  contact_32_5566
timestamp 1624857261
transform 1 0 22440 0 1 70589
box 0 0 1 1
use contact_32  contact_32_5565
timestamp 1624857261
transform 1 0 22712 0 1 41485
box 0 0 1 1
use contact_32  contact_32_5564
timestamp 1624857261
transform 1 0 22712 0 1 41757
box 0 0 1 1
use contact_32  contact_32_5563
timestamp 1624857261
transform 1 0 22576 0 1 82149
box 0 0 1 1
use contact_32  contact_32_5562
timestamp 1624857261
transform 1 0 22576 0 1 82421
box 0 0 1 1
use contact_32  contact_32_5561
timestamp 1624857261
transform 1 0 22712 0 1 82013
box 0 0 1 1
use contact_32  contact_32_5560
timestamp 1624857261
transform 1 0 22712 0 1 81741
box 0 0 1 1
use contact_32  contact_32_5559
timestamp 1624857261
transform 1 0 22576 0 1 33461
box 0 0 1 1
use contact_32  contact_32_5558
timestamp 1624857261
transform 1 0 22576 0 1 33189
box 0 0 1 1
use contact_32  contact_32_5557
timestamp 1624857261
transform 1 0 22576 0 1 33597
box 0 0 1 1
use contact_32  contact_32_5556
timestamp 1624857261
transform 1 0 22576 0 1 33869
box 0 0 1 1
use contact_32  contact_32_5555
timestamp 1624857261
transform 1 0 22576 0 1 44205
box 0 0 1 1
use contact_32  contact_32_5554
timestamp 1624857261
transform 1 0 22576 0 1 44477
box 0 0 1 1
use contact_32  contact_32_5553
timestamp 1624857261
transform 1 0 22712 0 1 108125
box 0 0 1 1
use contact_32  contact_32_5552
timestamp 1624857261
transform 1 0 22712 0 1 107853
box 0 0 1 1
use contact_32  contact_32_5551
timestamp 1624857261
transform 1 0 22712 0 1 93981
box 0 0 1 1
use contact_32  contact_32_5550
timestamp 1624857261
transform 1 0 22712 0 1 94253
box 0 0 1 1
use contact_32  contact_32_5549
timestamp 1624857261
transform 1 0 22576 0 1 123629
box 0 0 1 1
use contact_32  contact_32_5548
timestamp 1624857261
transform 1 0 22576 0 1 123901
box 0 0 1 1
use contact_32  contact_32_5547
timestamp 1624857261
transform 1 0 22576 0 1 123493
box 0 0 1 1
use contact_32  contact_32_5546
timestamp 1624857261
transform 1 0 22576 0 1 123221
box 0 0 1 1
use contact_32  contact_32_5545
timestamp 1624857261
transform 1 0 22576 0 1 31149
box 0 0 1 1
use contact_32  contact_32_5544
timestamp 1624857261
transform 1 0 22576 0 1 31421
box 0 0 1 1
use contact_32  contact_32_5543
timestamp 1624857261
transform 1 0 22576 0 1 117237
box 0 0 1 1
use contact_32  contact_32_5542
timestamp 1624857261
transform 1 0 22576 0 1 117509
box 0 0 1 1
use contact_32  contact_32_5541
timestamp 1624857261
transform 1 0 22576 0 1 69501
box 0 0 1 1
use contact_32  contact_32_5540
timestamp 1624857261
transform 1 0 22576 0 1 69773
box 0 0 1 1
use contact_32  contact_32_5539
timestamp 1624857261
transform 1 0 22576 0 1 69365
box 0 0 1 1
use contact_32  contact_32_5538
timestamp 1624857261
transform 1 0 22576 0 1 69093
box 0 0 1 1
use contact_32  contact_32_5537
timestamp 1624857261
transform 1 0 22576 0 1 58349
box 0 0 1 1
use contact_32  contact_32_5536
timestamp 1624857261
transform 1 0 22576 0 1 58077
box 0 0 1 1
use contact_32  contact_32_5535
timestamp 1624857261
transform 1 0 22576 0 1 70181
box 0 0 1 1
use contact_32  contact_32_5534
timestamp 1624857261
transform 1 0 22576 0 1 69909
box 0 0 1 1
use contact_32  contact_32_5533
timestamp 1624857261
transform 1 0 22576 0 1 67053
box 0 0 1 1
use contact_32  contact_32_5532
timestamp 1624857261
transform 1 0 22576 0 1 66781
box 0 0 1 1
use contact_32  contact_32_5531
timestamp 1624857261
transform 1 0 22576 0 1 86501
box 0 0 1 1
use contact_32  contact_32_5530
timestamp 1624857261
transform 1 0 22576 0 1 86773
box 0 0 1 1
use contact_32  contact_32_5529
timestamp 1624857261
transform 1 0 22712 0 1 73037
box 0 0 1 1
use contact_32  contact_32_5528
timestamp 1624857261
transform 1 0 22712 0 1 73309
box 0 0 1 1
use contact_32  contact_32_5527
timestamp 1624857261
transform 1 0 22576 0 1 87589
box 0 0 1 1
use contact_32  contact_32_5526
timestamp 1624857261
transform 1 0 22576 0 1 87317
box 0 0 1 1
use contact_32  contact_32_5525
timestamp 1624857261
transform 1 0 22576 0 1 107309
box 0 0 1 1
use contact_32  contact_32_5524
timestamp 1624857261
transform 1 0 22576 0 1 107037
box 0 0 1 1
use contact_32  contact_32_5523
timestamp 1624857261
transform 1 0 22712 0 1 49373
box 0 0 1 1
use contact_32  contact_32_5522
timestamp 1624857261
transform 1 0 22712 0 1 49645
box 0 0 1 1
use contact_32  contact_32_5521
timestamp 1624857261
transform 1 0 22576 0 1 111661
box 0 0 1 1
use contact_32  contact_32_5520
timestamp 1624857261
transform 1 0 22576 0 1 111389
box 0 0 1 1
use contact_32  contact_32_5519
timestamp 1624857261
transform 1 0 22712 0 1 37133
box 0 0 1 1
use contact_32  contact_32_5518
timestamp 1624857261
transform 1 0 22712 0 1 37405
box 0 0 1 1
use contact_32  contact_32_5517
timestamp 1624857261
transform 1 0 22712 0 1 124445
box 0 0 1 1
use contact_32  contact_32_5516
timestamp 1624857261
transform 1 0 22712 0 1 124717
box 0 0 1 1
use contact_32  contact_32_5515
timestamp 1624857261
transform 1 0 22712 0 1 118733
box 0 0 1 1
use contact_32  contact_32_5514
timestamp 1624857261
transform 1 0 22712 0 1 118461
box 0 0 1 1
use contact_32  contact_32_5513
timestamp 1624857261
transform 1 0 22576 0 1 25709
box 0 0 1 1
use contact_32  contact_32_5512
timestamp 1624857261
transform 1 0 22576 0 1 25981
box 0 0 1 1
use contact_32  contact_32_5511
timestamp 1624857261
transform 1 0 22712 0 1 89629
box 0 0 1 1
use contact_32  contact_32_5510
timestamp 1624857261
transform 1 0 22712 0 1 89901
box 0 0 1 1
use contact_32  contact_32_5509
timestamp 1624857261
transform 1 0 22712 0 1 72493
box 0 0 1 1
use contact_32  contact_32_5508
timestamp 1624857261
transform 1 0 22712 0 1 72221
box 0 0 1 1
use contact_32  contact_32_5507
timestamp 1624857261
transform 1 0 22576 0 1 65013
box 0 0 1 1
use contact_32  contact_32_5506
timestamp 1624857261
transform 1 0 22576 0 1 64741
box 0 0 1 1
use contact_32  contact_32_5505
timestamp 1624857261
transform 1 0 22712 0 1 102685
box 0 0 1 1
use contact_32  contact_32_5504
timestamp 1624857261
transform 1 0 22712 0 1 102957
box 0 0 1 1
use contact_32  contact_32_5503
timestamp 1624857261
transform 1 0 22576 0 1 95205
box 0 0 1 1
use contact_32  contact_32_5502
timestamp 1624857261
transform 1 0 22576 0 1 95477
box 0 0 1 1
use contact_32  contact_32_5501
timestamp 1624857261
transform 1 0 22712 0 1 95069
box 0 0 1 1
use contact_32  contact_32_5500
timestamp 1624857261
transform 1 0 22712 0 1 94797
box 0 0 1 1
use contact_32  contact_32_5499
timestamp 1624857261
transform 1 0 22712 0 1 31965
box 0 0 1 1
use contact_32  contact_32_5498
timestamp 1624857261
transform 1 0 22712 0 1 32237
box 0 0 1 1
use contact_32  contact_32_5497
timestamp 1624857261
transform 1 0 22712 0 1 51005
box 0 0 1 1
use contact_32  contact_32_5496
timestamp 1624857261
transform 1 0 22712 0 1 51277
box 0 0 1 1
use contact_32  contact_32_5495
timestamp 1624857261
transform 1 0 22712 0 1 55629
box 0 0 1 1
use contact_32  contact_32_5494
timestamp 1624857261
transform 1 0 22712 0 1 55901
box 0 0 1 1
use contact_32  contact_32_5493
timestamp 1624857261
transform 1 0 22576 0 1 118325
box 0 0 1 1
use contact_32  contact_32_5492
timestamp 1624857261
transform 1 0 22576 0 1 118053
box 0 0 1 1
use contact_32  contact_32_5491
timestamp 1624857261
transform 1 0 22576 0 1 105405
box 0 0 1 1
use contact_32  contact_32_5490
timestamp 1624857261
transform 1 0 22576 0 1 105677
box 0 0 1 1
use contact_32  contact_32_5489
timestamp 1624857261
transform 1 0 22576 0 1 65829
box 0 0 1 1
use contact_32  contact_32_5488
timestamp 1624857261
transform 1 0 22576 0 1 65557
box 0 0 1 1
use contact_32  contact_32_5487
timestamp 1624857261
transform 1 0 22712 0 1 63517
box 0 0 1 1
use contact_32  contact_32_5486
timestamp 1624857261
transform 1 0 22712 0 1 63789
box 0 0 1 1
use contact_32  contact_32_5485
timestamp 1624857261
transform 1 0 22576 0 1 90853
box 0 0 1 1
use contact_32  contact_32_5484
timestamp 1624857261
transform 1 0 22576 0 1 91125
box 0 0 1 1
use contact_32  contact_32_5483
timestamp 1624857261
transform 1 0 22712 0 1 90717
box 0 0 1 1
use contact_32  contact_32_5482
timestamp 1624857261
transform 1 0 22712 0 1 90445
box 0 0 1 1
use contact_32  contact_32_5481
timestamp 1624857261
transform 1 0 22712 0 1 74125
box 0 0 1 1
use contact_32  contact_32_5480
timestamp 1624857261
transform 1 0 22712 0 1 73853
box 0 0 1 1
use contact_32  contact_32_5479
timestamp 1624857261
transform 1 0 22576 0 1 38357
box 0 0 1 1
use contact_32  contact_32_5478
timestamp 1624857261
transform 1 0 22576 0 1 38629
box 0 0 1 1
use contact_32  contact_32_5477
timestamp 1624857261
transform 1 0 22712 0 1 91533
box 0 0 1 1
use contact_32  contact_32_5476
timestamp 1624857261
transform 1 0 22712 0 1 91261
box 0 0 1 1
use contact_32  contact_32_5475
timestamp 1624857261
transform 1 0 22576 0 1 48421
box 0 0 1 1
use contact_32  contact_32_5474
timestamp 1624857261
transform 1 0 22576 0 1 48149
box 0 0 1 1
use contact_32  contact_32_5473
timestamp 1624857261
transform 1 0 22712 0 1 64333
box 0 0 1 1
use contact_32  contact_32_5472
timestamp 1624857261
transform 1 0 22712 0 1 64605
box 0 0 1 1
use contact_32  contact_32_5471
timestamp 1624857261
transform 1 0 22576 0 1 36589
box 0 0 1 1
use contact_32  contact_32_5470
timestamp 1624857261
transform 1 0 22576 0 1 36317
box 0 0 1 1
use contact_32  contact_32_5469
timestamp 1624857261
transform 1 0 22576 0 1 78885
box 0 0 1 1
use contact_32  contact_32_5468
timestamp 1624857261
transform 1 0 22576 0 1 78613
box 0 0 1 1
use contact_32  contact_32_5467
timestamp 1624857261
transform 1 0 22576 0 1 116013
box 0 0 1 1
use contact_32  contact_32_5466
timestamp 1624857261
transform 1 0 22576 0 1 115741
box 0 0 1 1
use contact_32  contact_32_5465
timestamp 1624857261
transform 1 0 22712 0 1 29517
box 0 0 1 1
use contact_32  contact_32_5464
timestamp 1624857261
transform 1 0 22712 0 1 29245
box 0 0 1 1
use contact_32  contact_32_5463
timestamp 1624857261
transform 1 0 22576 0 1 40941
box 0 0 1 1
use contact_32  contact_32_5462
timestamp 1624857261
transform 1 0 22576 0 1 40669
box 0 0 1 1
use contact_32  contact_32_5461
timestamp 1624857261
transform 1 0 22712 0 1 62021
box 0 0 1 1
use contact_32  contact_32_5460
timestamp 1624857261
transform 1 0 22712 0 1 62293
box 0 0 1 1
use contact_32  contact_32_5459
timestamp 1624857261
transform 1 0 22576 0 1 61885
box 0 0 1 1
use contact_32  contact_32_5458
timestamp 1624857261
transform 1 0 22576 0 1 61613
box 0 0 1 1
use contact_32  contact_32_5457
timestamp 1624857261
transform 1 0 22576 0 1 27885
box 0 0 1 1
use contact_32  contact_32_5456
timestamp 1624857261
transform 1 0 22576 0 1 27613
box 0 0 1 1
use contact_32  contact_32_5455
timestamp 1624857261
transform 1 0 22712 0 1 99149
box 0 0 1 1
use contact_32  contact_32_5454
timestamp 1624857261
transform 1 0 22712 0 1 99421
box 0 0 1 1
use contact_32  contact_32_5453
timestamp 1624857261
transform 1 0 22712 0 1 66373
box 0 0 1 1
use contact_32  contact_32_5452
timestamp 1624857261
transform 1 0 22712 0 1 66645
box 0 0 1 1
use contact_32  contact_32_5451
timestamp 1624857261
transform 1 0 22576 0 1 55221
box 0 0 1 1
use contact_32  contact_32_5450
timestamp 1624857261
transform 1 0 22576 0 1 54949
box 0 0 1 1
use contact_32  contact_32_5449
timestamp 1624857261
transform 1 0 22576 0 1 77797
box 0 0 1 1
use contact_32  contact_32_5448
timestamp 1624857261
transform 1 0 22576 0 1 78069
box 0 0 1 1
use contact_32  contact_32_5447
timestamp 1624857261
transform 1 0 22576 0 1 30605
box 0 0 1 1
use contact_32  contact_32_5446
timestamp 1624857261
transform 1 0 22576 0 1 30333
box 0 0 1 1
use contact_32  contact_32_5445
timestamp 1624857261
transform 1 0 22712 0 1 96973
box 0 0 1 1
use contact_32  contact_32_5444
timestamp 1624857261
transform 1 0 22712 0 1 96701
box 0 0 1 1
use contact_32  contact_32_5443
timestamp 1624857261
transform 1 0 22712 0 1 68685
box 0 0 1 1
use contact_32  contact_32_5442
timestamp 1624857261
transform 1 0 22712 0 1 68957
box 0 0 1 1
use contact_32  contact_32_5441
timestamp 1624857261
transform 1 0 22576 0 1 100645
box 0 0 1 1
use contact_32  contact_32_5440
timestamp 1624857261
transform 1 0 22576 0 1 100917
box 0 0 1 1
use contact_32  contact_32_5439
timestamp 1624857261
transform 1 0 22576 0 1 103909
box 0 0 1 1
use contact_32  contact_32_5438
timestamp 1624857261
transform 1 0 22576 0 1 104181
box 0 0 1 1
use contact_32  contact_32_5437
timestamp 1624857261
transform 1 0 22712 0 1 35909
box 0 0 1 1
use contact_32  contact_32_5436
timestamp 1624857261
transform 1 0 22712 0 1 36181
box 0 0 1 1
use contact_32  contact_32_5435
timestamp 1624857261
transform 1 0 22576 0 1 110845
box 0 0 1 1
use contact_32  contact_32_5434
timestamp 1624857261
transform 1 0 22576 0 1 110573
box 0 0 1 1
use contact_32  contact_32_5433
timestamp 1624857261
transform 1 0 22712 0 1 122269
box 0 0 1 1
use contact_32  contact_32_5432
timestamp 1624857261
transform 1 0 22712 0 1 121997
box 0 0 1 1
use contact_32  contact_32_5431
timestamp 1624857261
transform 1 0 22576 0 1 122405
box 0 0 1 1
use contact_32  contact_32_5430
timestamp 1624857261
transform 1 0 22576 0 1 122677
box 0 0 1 1
use contact_32  contact_32_5429
timestamp 1624857261
transform 1 0 22576 0 1 73445
box 0 0 1 1
use contact_32  contact_32_5428
timestamp 1624857261
transform 1 0 22576 0 1 73717
box 0 0 1 1
use contact_32  contact_32_5427
timestamp 1624857261
transform 1 0 22576 0 1 34685
box 0 0 1 1
use contact_32  contact_32_5426
timestamp 1624857261
transform 1 0 22576 0 1 34413
box 0 0 1 1
use contact_32  contact_32_5425
timestamp 1624857261
transform 1 0 22712 0 1 120093
box 0 0 1 1
use contact_32  contact_32_5424
timestamp 1624857261
transform 1 0 22712 0 1 120365
box 0 0 1 1
use contact_32  contact_32_5423
timestamp 1624857261
transform 1 0 22576 0 1 112885
box 0 0 1 1
use contact_32  contact_32_5422
timestamp 1624857261
transform 1 0 22576 0 1 112613
box 0 0 1 1
use contact_32  contact_32_5421
timestamp 1624857261
transform 1 0 22576 0 1 46245
box 0 0 1 1
use contact_32  contact_32_5420
timestamp 1624857261
transform 1 0 22576 0 1 46517
box 0 0 1 1
use contact_32  contact_32_5419
timestamp 1624857261
transform 1 0 22576 0 1 58893
box 0 0 1 1
use contact_32  contact_32_5418
timestamp 1624857261
transform 1 0 22576 0 1 59165
box 0 0 1 1
use contact_32  contact_32_5417
timestamp 1624857261
transform 1 0 22712 0 1 82829
box 0 0 1 1
use contact_32  contact_32_5416
timestamp 1624857261
transform 1 0 22712 0 1 82557
box 0 0 1 1
use contact_32  contact_32_5415
timestamp 1624857261
transform 1 0 22576 0 1 109621
box 0 0 1 1
use contact_32  contact_32_5414
timestamp 1624857261
transform 1 0 22576 0 1 109349
box 0 0 1 1
use contact_32  contact_32_5413
timestamp 1624857261
transform 1 0 22576 0 1 59845
box 0 0 1 1
use contact_32  contact_32_5412
timestamp 1624857261
transform 1 0 22576 0 1 59573
box 0 0 1 1
use contact_32  contact_32_5411
timestamp 1624857261
transform 1 0 22712 0 1 45021
box 0 0 1 1
use contact_32  contact_32_5410
timestamp 1624857261
transform 1 0 22712 0 1 45293
box 0 0 1 1
use contact_32  contact_32_5409
timestamp 1624857261
transform 1 0 22712 0 1 50461
box 0 0 1 1
use contact_32  contact_32_5408
timestamp 1624857261
transform 1 0 22712 0 1 50189
box 0 0 1 1
use contact_32  contact_32_5407
timestamp 1624857261
transform 1 0 22576 0 1 60389
box 0 0 1 1
use contact_32  contact_32_5406
timestamp 1624857261
transform 1 0 22576 0 1 60661
box 0 0 1 1
use contact_32  contact_32_5405
timestamp 1624857261
transform 1 0 22576 0 1 83645
box 0 0 1 1
use contact_32  contact_32_5404
timestamp 1624857261
transform 1 0 22576 0 1 83373
box 0 0 1 1
use contact_32  contact_32_5403
timestamp 1624857261
transform 1 0 22712 0 1 61069
box 0 0 1 1
use contact_32  contact_32_5402
timestamp 1624857261
transform 1 0 22712 0 1 60797
box 0 0 1 1
use contact_32  contact_32_5401
timestamp 1624857261
transform 1 0 22712 0 1 78477
box 0 0 1 1
use contact_32  contact_32_5400
timestamp 1624857261
transform 1 0 22712 0 1 78205
box 0 0 1 1
use contact_32  contact_32_5399
timestamp 1624857261
transform 1 0 22712 0 1 42573
box 0 0 1 1
use contact_32  contact_32_5398
timestamp 1624857261
transform 1 0 22712 0 1 42301
box 0 0 1 1
use contact_32  contact_32_5397
timestamp 1624857261
transform 1 0 22712 0 1 98333
box 0 0 1 1
use contact_32  contact_32_5396
timestamp 1624857261
transform 1 0 22712 0 1 98605
box 0 0 1 1
use contact_32  contact_32_5395
timestamp 1624857261
transform 1 0 22712 0 1 53725
box 0 0 1 1
use contact_32  contact_32_5394
timestamp 1624857261
transform 1 0 22712 0 1 53997
box 0 0 1 1
use contact_32  contact_32_5393
timestamp 1624857261
transform 1 0 22576 0 1 85549
box 0 0 1 1
use contact_32  contact_32_5392
timestamp 1624857261
transform 1 0 22576 0 1 85277
box 0 0 1 1
use contact_32  contact_32_5391
timestamp 1624857261
transform 1 0 22712 0 1 56717
box 0 0 1 1
use contact_32  contact_32_5390
timestamp 1624857261
transform 1 0 22712 0 1 56445
box 0 0 1 1
use contact_32  contact_32_5389
timestamp 1624857261
transform 1 0 22576 0 1 104997
box 0 0 1 1
use contact_32  contact_32_5388
timestamp 1624857261
transform 1 0 22576 0 1 104725
box 0 0 1 1
use contact_32  contact_32_5387
timestamp 1624857261
transform 1 0 22576 0 1 81197
box 0 0 1 1
use contact_32  contact_32_5386
timestamp 1624857261
transform 1 0 22576 0 1 80925
box 0 0 1 1
use contact_32  contact_32_5385
timestamp 1624857261
transform 1 0 22576 0 1 57261
box 0 0 1 1
use contact_32  contact_32_5384
timestamp 1624857261
transform 1 0 22576 0 1 57533
box 0 0 1 1
use contact_32  contact_32_5383
timestamp 1624857261
transform 1 0 22576 0 1 29109
box 0 0 1 1
use contact_32  contact_32_5382
timestamp 1624857261
transform 1 0 22576 0 1 28837
box 0 0 1 1
use contact_32  contact_32_5381
timestamp 1624857261
transform 1 0 22712 0 1 48013
box 0 0 1 1
use contact_32  contact_32_5380
timestamp 1624857261
transform 1 0 22712 0 1 47741
box 0 0 1 1
use contact_32  contact_32_5379
timestamp 1624857261
transform 1 0 22712 0 1 28429
box 0 0 1 1
use contact_32  contact_32_5378
timestamp 1624857261
transform 1 0 22712 0 1 28701
box 0 0 1 1
use contact_32  contact_32_5377
timestamp 1624857261
transform 1 0 22576 0 1 37813
box 0 0 1 1
use contact_32  contact_32_5376
timestamp 1624857261
transform 1 0 22576 0 1 37541
box 0 0 1 1
use contact_32  contact_32_5375
timestamp 1624857261
transform 1 0 23392 0 1 100237
box 0 0 1 1
use contact_32  contact_32_5374
timestamp 1624857261
transform 1 0 23392 0 1 99965
box 0 0 1 1
use contact_32  contact_32_5373
timestamp 1624857261
transform 1 0 23528 0 1 48557
box 0 0 1 1
use contact_32  contact_32_5372
timestamp 1624857261
transform 1 0 23528 0 1 48829
box 0 0 1 1
use contact_32  contact_32_5371
timestamp 1624857261
transform 1 0 23528 0 1 48421
box 0 0 1 1
use contact_32  contact_32_5370
timestamp 1624857261
transform 1 0 23528 0 1 48149
box 0 0 1 1
use contact_32  contact_32_5369
timestamp 1624857261
transform 1 0 23528 0 1 81197
box 0 0 1 1
use contact_32  contact_32_5368
timestamp 1624857261
transform 1 0 23528 0 1 80925
box 0 0 1 1
use contact_32  contact_32_5367
timestamp 1624857261
transform 1 0 23528 0 1 81333
box 0 0 1 1
use contact_32  contact_32_5366
timestamp 1624857261
transform 1 0 23528 0 1 81605
box 0 0 1 1
use contact_32  contact_32_5365
timestamp 1624857261
transform 1 0 23528 0 1 57533
box 0 0 1 1
use contact_32  contact_32_5364
timestamp 1624857261
transform 1 0 23528 0 1 57261
box 0 0 1 1
use contact_32  contact_32_5363
timestamp 1624857261
transform 1 0 23392 0 1 57669
box 0 0 1 1
use contact_32  contact_32_5362
timestamp 1624857261
transform 1 0 23392 0 1 57941
box 0 0 1 1
use contact_32  contact_32_5361
timestamp 1624857261
transform 1 0 23528 0 1 76981
box 0 0 1 1
use contact_32  contact_32_5360
timestamp 1624857261
transform 1 0 23528 0 1 77253
box 0 0 1 1
use contact_32  contact_32_5359
timestamp 1624857261
transform 1 0 23528 0 1 76845
box 0 0 1 1
use contact_32  contact_32_5358
timestamp 1624857261
transform 1 0 23528 0 1 76573
box 0 0 1 1
use contact_32  contact_32_5357
timestamp 1624857261
transform 1 0 23392 0 1 52365
box 0 0 1 1
use contact_32  contact_32_5356
timestamp 1624857261
transform 1 0 23392 0 1 52093
box 0 0 1 1
use contact_32  contact_32_5355
timestamp 1624857261
transform 1 0 23392 0 1 52501
box 0 0 1 1
use contact_32  contact_32_5354
timestamp 1624857261
transform 1 0 23392 0 1 52773
box 0 0 1 1
use contact_32  contact_32_5353
timestamp 1624857261
transform 1 0 23392 0 1 107037
box 0 0 1 1
use contact_32  contact_32_5352
timestamp 1624857261
transform 1 0 23392 0 1 107309
box 0 0 1 1
use contact_32  contact_32_5351
timestamp 1624857261
transform 1 0 23392 0 1 106901
box 0 0 1 1
use contact_32  contact_32_5350
timestamp 1624857261
transform 1 0 23392 0 1 106629
box 0 0 1 1
use contact_32  contact_32_5349
timestamp 1624857261
transform 1 0 23392 0 1 75077
box 0 0 1 1
use contact_32  contact_32_5348
timestamp 1624857261
transform 1 0 23392 0 1 75349
box 0 0 1 1
use contact_32  contact_32_5347
timestamp 1624857261
transform 1 0 23528 0 1 74941
box 0 0 1 1
use contact_32  contact_32_5346
timestamp 1624857261
transform 1 0 23528 0 1 74669
box 0 0 1 1
use contact_32  contact_32_5345
timestamp 1624857261
transform 1 0 23528 0 1 91941
box 0 0 1 1
use contact_32  contact_32_5344
timestamp 1624857261
transform 1 0 23528 0 1 91669
box 0 0 1 1
use contact_32  contact_32_5343
timestamp 1624857261
transform 1 0 23528 0 1 113973
box 0 0 1 1
use contact_32  contact_32_5342
timestamp 1624857261
transform 1 0 23528 0 1 113701
box 0 0 1 1
use contact_32  contact_32_5341
timestamp 1624857261
transform 1 0 23528 0 1 114109
box 0 0 1 1
use contact_32  contact_32_5340
timestamp 1624857261
transform 1 0 23528 0 1 114381
box 0 0 1 1
use contact_32  contact_32_5339
timestamp 1624857261
transform 1 0 23392 0 1 124445
box 0 0 1 1
use contact_32  contact_32_5338
timestamp 1624857261
transform 1 0 23392 0 1 124717
box 0 0 1 1
use contact_32  contact_32_5337
timestamp 1624857261
transform 1 0 23392 0 1 124309
box 0 0 1 1
use contact_32  contact_32_5336
timestamp 1624857261
transform 1 0 23392 0 1 124037
box 0 0 1 1
use contact_32  contact_32_5335
timestamp 1624857261
transform 1 0 23392 0 1 102685
box 0 0 1 1
use contact_32  contact_32_5334
timestamp 1624857261
transform 1 0 23392 0 1 102957
box 0 0 1 1
use contact_32  contact_32_5333
timestamp 1624857261
transform 1 0 23392 0 1 102549
box 0 0 1 1
use contact_32  contact_32_5332
timestamp 1624857261
transform 1 0 23392 0 1 102277
box 0 0 1 1
use contact_32  contact_32_5331
timestamp 1624857261
transform 1 0 23528 0 1 45293
box 0 0 1 1
use contact_32  contact_32_5330
timestamp 1624857261
transform 1 0 23528 0 1 45021
box 0 0 1 1
use contact_32  contact_32_5329
timestamp 1624857261
transform 1 0 23528 0 1 45429
box 0 0 1 1
use contact_32  contact_32_5328
timestamp 1624857261
transform 1 0 23528 0 1 45701
box 0 0 1 1
use contact_32  contact_32_5327
timestamp 1624857261
transform 1 0 23392 0 1 33053
box 0 0 1 1
use contact_32  contact_32_5326
timestamp 1624857261
transform 1 0 23392 0 1 32781
box 0 0 1 1
use contact_32  contact_32_5325
timestamp 1624857261
transform 1 0 23528 0 1 33189
box 0 0 1 1
use contact_32  contact_32_5324
timestamp 1624857261
transform 1 0 23528 0 1 33461
box 0 0 1 1
use contact_32  contact_32_5323
timestamp 1624857261
transform 1 0 23392 0 1 37405
box 0 0 1 1
use contact_32  contact_32_5322
timestamp 1624857261
transform 1 0 23392 0 1 37133
box 0 0 1 1
use contact_32  contact_32_5321
timestamp 1624857261
transform 1 0 23528 0 1 37541
box 0 0 1 1
use contact_32  contact_32_5320
timestamp 1624857261
transform 1 0 23528 0 1 37813
box 0 0 1 1
use contact_32  contact_32_5319
timestamp 1624857261
transform 1 0 23528 0 1 61477
box 0 0 1 1
use contact_32  contact_32_5318
timestamp 1624857261
transform 1 0 23528 0 1 61205
box 0 0 1 1
use contact_32  contact_32_5317
timestamp 1624857261
transform 1 0 23528 0 1 61613
box 0 0 1 1
use contact_32  contact_32_5316
timestamp 1624857261
transform 1 0 23528 0 1 61885
box 0 0 1 1
use contact_32  contact_32_5315
timestamp 1624857261
transform 1 0 23528 0 1 110437
box 0 0 1 1
use contact_32  contact_32_5314
timestamp 1624857261
transform 1 0 23528 0 1 110165
box 0 0 1 1
use contact_32  contact_32_5313
timestamp 1624857261
transform 1 0 23528 0 1 110573
box 0 0 1 1
use contact_32  contact_32_5312
timestamp 1624857261
transform 1 0 23528 0 1 110845
box 0 0 1 1
use contact_32  contact_32_5311
timestamp 1624857261
transform 1 0 23528 0 1 69093
box 0 0 1 1
use contact_32  contact_32_5310
timestamp 1624857261
transform 1 0 23528 0 1 69365
box 0 0 1 1
use contact_32  contact_32_5309
timestamp 1624857261
transform 1 0 23392 0 1 68957
box 0 0 1 1
use contact_32  contact_32_5308
timestamp 1624857261
transform 1 0 23392 0 1 68685
box 0 0 1 1
use contact_32  contact_32_5307
timestamp 1624857261
transform 1 0 23528 0 1 119141
box 0 0 1 1
use contact_32  contact_32_5306
timestamp 1624857261
transform 1 0 23528 0 1 118869
box 0 0 1 1
use contact_32  contact_32_5305
timestamp 1624857261
transform 1 0 23528 0 1 119277
box 0 0 1 1
use contact_32  contact_32_5304
timestamp 1624857261
transform 1 0 23528 0 1 119549
box 0 0 1 1
use contact_32  contact_32_5303
timestamp 1624857261
transform 1 0 23392 0 1 46109
box 0 0 1 1
use contact_32  contact_32_5302
timestamp 1624857261
transform 1 0 23392 0 1 45837
box 0 0 1 1
use contact_32  contact_32_5301
timestamp 1624857261
transform 1 0 23528 0 1 46245
box 0 0 1 1
use contact_32  contact_32_5300
timestamp 1624857261
transform 1 0 23528 0 1 46517
box 0 0 1 1
use contact_32  contact_32_5299
timestamp 1624857261
transform 1 0 23528 0 1 82421
box 0 0 1 1
use contact_32  contact_32_5298
timestamp 1624857261
transform 1 0 23528 0 1 82149
box 0 0 1 1
use contact_32  contact_32_5297
timestamp 1624857261
transform 1 0 23528 0 1 82557
box 0 0 1 1
use contact_32  contact_32_5296
timestamp 1624857261
transform 1 0 23528 0 1 82829
box 0 0 1 1
use contact_32  contact_32_5295
timestamp 1624857261
transform 1 0 23528 0 1 47333
box 0 0 1 1
use contact_32  contact_32_5294
timestamp 1624857261
transform 1 0 23528 0 1 47605
box 0 0 1 1
use contact_32  contact_32_5293
timestamp 1624857261
transform 1 0 23528 0 1 60797
box 0 0 1 1
use contact_32  contact_32_5292
timestamp 1624857261
transform 1 0 23528 0 1 61069
box 0 0 1 1
use contact_32  contact_32_5291
timestamp 1624857261
transform 1 0 23528 0 1 60661
box 0 0 1 1
use contact_32  contact_32_5290
timestamp 1624857261
transform 1 0 23528 0 1 60389
box 0 0 1 1
use contact_32  contact_32_5289
timestamp 1624857261
transform 1 0 23528 0 1 98741
box 0 0 1 1
use contact_32  contact_32_5288
timestamp 1624857261
transform 1 0 23528 0 1 99013
box 0 0 1 1
use contact_32  contact_32_5287
timestamp 1624857261
transform 1 0 23528 0 1 98605
box 0 0 1 1
use contact_32  contact_32_5286
timestamp 1624857261
transform 1 0 23528 0 1 98333
box 0 0 1 1
use contact_32  contact_32_5285
timestamp 1624857261
transform 1 0 23392 0 1 92757
box 0 0 1 1
use contact_32  contact_32_5284
timestamp 1624857261
transform 1 0 23392 0 1 93029
box 0 0 1 1
use contact_32  contact_32_5283
timestamp 1624857261
transform 1 0 23392 0 1 107717
box 0 0 1 1
use contact_32  contact_32_5282
timestamp 1624857261
transform 1 0 23392 0 1 107445
box 0 0 1 1
use contact_32  contact_32_5281
timestamp 1624857261
transform 1 0 23392 0 1 107853
box 0 0 1 1
use contact_32  contact_32_5280
timestamp 1624857261
transform 1 0 23392 0 1 108125
box 0 0 1 1
use contact_32  contact_32_5279
timestamp 1624857261
transform 1 0 23392 0 1 120773
box 0 0 1 1
use contact_32  contact_32_5278
timestamp 1624857261
transform 1 0 23392 0 1 120501
box 0 0 1 1
use contact_32  contact_32_5277
timestamp 1624857261
transform 1 0 23392 0 1 39309
box 0 0 1 1
use contact_32  contact_32_5276
timestamp 1624857261
transform 1 0 23392 0 1 39037
box 0 0 1 1
use contact_32  contact_32_5275
timestamp 1624857261
transform 1 0 23392 0 1 39445
box 0 0 1 1
use contact_32  contact_32_5274
timestamp 1624857261
transform 1 0 23392 0 1 39717
box 0 0 1 1
use contact_32  contact_32_5273
timestamp 1624857261
transform 1 0 23392 0 1 110029
box 0 0 1 1
use contact_32  contact_32_5272
timestamp 1624857261
transform 1 0 23392 0 1 109757
box 0 0 1 1
use contact_32  contact_32_5271
timestamp 1624857261
transform 1 0 23392 0 1 64197
box 0 0 1 1
use contact_32  contact_32_5270
timestamp 1624857261
transform 1 0 23392 0 1 63925
box 0 0 1 1
use contact_32  contact_32_5269
timestamp 1624857261
transform 1 0 23392 0 1 64333
box 0 0 1 1
use contact_32  contact_32_5268
timestamp 1624857261
transform 1 0 23392 0 1 64605
box 0 0 1 1
use contact_32  contact_32_5267
timestamp 1624857261
transform 1 0 23392 0 1 53317
box 0 0 1 1
use contact_32  contact_32_5266
timestamp 1624857261
transform 1 0 23392 0 1 53589
box 0 0 1 1
use contact_32  contact_32_5265
timestamp 1624857261
transform 1 0 23528 0 1 53181
box 0 0 1 1
use contact_32  contact_32_5264
timestamp 1624857261
transform 1 0 23528 0 1 52909
box 0 0 1 1
use contact_32  contact_32_5263
timestamp 1624857261
transform 1 0 23392 0 1 35093
box 0 0 1 1
use contact_32  contact_32_5262
timestamp 1624857261
transform 1 0 23392 0 1 35365
box 0 0 1 1
use contact_32  contact_32_5261
timestamp 1624857261
transform 1 0 23392 0 1 103365
box 0 0 1 1
use contact_32  contact_32_5260
timestamp 1624857261
transform 1 0 23392 0 1 103093
box 0 0 1 1
use contact_32  contact_32_5259
timestamp 1624857261
transform 1 0 23392 0 1 103501
box 0 0 1 1
use contact_32  contact_32_5258
timestamp 1624857261
transform 1 0 23392 0 1 103773
box 0 0 1 1
use contact_32  contact_32_5257
timestamp 1624857261
transform 1 0 23392 0 1 62293
box 0 0 1 1
use contact_32  contact_32_5256
timestamp 1624857261
transform 1 0 23392 0 1 62021
box 0 0 1 1
use contact_32  contact_32_5255
timestamp 1624857261
transform 1 0 23392 0 1 62429
box 0 0 1 1
use contact_32  contact_32_5254
timestamp 1624857261
transform 1 0 23392 0 1 62701
box 0 0 1 1
use contact_32  contact_32_5253
timestamp 1624857261
transform 1 0 23528 0 1 94253
box 0 0 1 1
use contact_32  contact_32_5252
timestamp 1624857261
transform 1 0 23528 0 1 93981
box 0 0 1 1
use contact_32  contact_32_5251
timestamp 1624857261
transform 1 0 23528 0 1 94389
box 0 0 1 1
use contact_32  contact_32_5250
timestamp 1624857261
transform 1 0 23528 0 1 94661
box 0 0 1 1
use contact_32  contact_32_5249
timestamp 1624857261
transform 1 0 23392 0 1 120093
box 0 0 1 1
use contact_32  contact_32_5248
timestamp 1624857261
transform 1 0 23392 0 1 120365
box 0 0 1 1
use contact_32  contact_32_5247
timestamp 1624857261
transform 1 0 23392 0 1 119957
box 0 0 1 1
use contact_32  contact_32_5246
timestamp 1624857261
transform 1 0 23392 0 1 119685
box 0 0 1 1
use contact_32  contact_32_5245
timestamp 1624857261
transform 1 0 23392 0 1 65557
box 0 0 1 1
use contact_32  contact_32_5244
timestamp 1624857261
transform 1 0 23392 0 1 65829
box 0 0 1 1
use contact_32  contact_32_5243
timestamp 1624857261
transform 1 0 23392 0 1 65421
box 0 0 1 1
use contact_32  contact_32_5242
timestamp 1624857261
transform 1 0 23392 0 1 65149
box 0 0 1 1
use contact_32  contact_32_5241
timestamp 1624857261
transform 1 0 23392 0 1 41349
box 0 0 1 1
use contact_32  contact_32_5240
timestamp 1624857261
transform 1 0 23392 0 1 41077
box 0 0 1 1
use contact_32  contact_32_5239
timestamp 1624857261
transform 1 0 23392 0 1 41485
box 0 0 1 1
use contact_32  contact_32_5238
timestamp 1624857261
transform 1 0 23392 0 1 41757
box 0 0 1 1
use contact_32  contact_32_5237
timestamp 1624857261
transform 1 0 23392 0 1 115605
box 0 0 1 1
use contact_32  contact_32_5236
timestamp 1624857261
transform 1 0 23392 0 1 115333
box 0 0 1 1
use contact_32  contact_32_5235
timestamp 1624857261
transform 1 0 23392 0 1 115741
box 0 0 1 1
use contact_32  contact_32_5234
timestamp 1624857261
transform 1 0 23392 0 1 116013
box 0 0 1 1
use contact_32  contact_32_5233
timestamp 1624857261
transform 1 0 23528 0 1 70589
box 0 0 1 1
use contact_32  contact_32_5232
timestamp 1624857261
transform 1 0 23528 0 1 70317
box 0 0 1 1
use contact_32  contact_32_5231
timestamp 1624857261
transform 1 0 23392 0 1 70725
box 0 0 1 1
use contact_32  contact_32_5230
timestamp 1624857261
transform 1 0 23392 0 1 70997
box 0 0 1 1
use contact_32  contact_32_5229
timestamp 1624857261
transform 1 0 23392 0 1 99421
box 0 0 1 1
use contact_32  contact_32_5228
timestamp 1624857261
transform 1 0 23392 0 1 99149
box 0 0 1 1
use contact_32  contact_32_5227
timestamp 1624857261
transform 1 0 23528 0 1 99557
box 0 0 1 1
use contact_32  contact_32_5226
timestamp 1624857261
transform 1 0 23528 0 1 99829
box 0 0 1 1
use contact_32  contact_32_5225
timestamp 1624857261
transform 1 0 23392 0 1 82013
box 0 0 1 1
use contact_32  contact_32_5224
timestamp 1624857261
transform 1 0 23392 0 1 81741
box 0 0 1 1
use contact_32  contact_32_5223
timestamp 1624857261
transform 1 0 23528 0 1 36589
box 0 0 1 1
use contact_32  contact_32_5222
timestamp 1624857261
transform 1 0 23528 0 1 36317
box 0 0 1 1
use contact_32  contact_32_5221
timestamp 1624857261
transform 1 0 23528 0 1 36725
box 0 0 1 1
use contact_32  contact_32_5220
timestamp 1624857261
transform 1 0 23528 0 1 36997
box 0 0 1 1
use contact_32  contact_32_5219
timestamp 1624857261
transform 1 0 23528 0 1 83373
box 0 0 1 1
use contact_32  contact_32_5218
timestamp 1624857261
transform 1 0 23528 0 1 83645
box 0 0 1 1
use contact_32  contact_32_5217
timestamp 1624857261
transform 1 0 23528 0 1 83237
box 0 0 1 1
use contact_32  contact_32_5216
timestamp 1624857261
transform 1 0 23528 0 1 82965
box 0 0 1 1
use contact_32  contact_32_5215
timestamp 1624857261
transform 1 0 23528 0 1 115197
box 0 0 1 1
use contact_32  contact_32_5214
timestamp 1624857261
transform 1 0 23528 0 1 114925
box 0 0 1 1
use contact_32  contact_32_5213
timestamp 1624857261
transform 1 0 23528 0 1 79293
box 0 0 1 1
use contact_32  contact_32_5212
timestamp 1624857261
transform 1 0 23528 0 1 79021
box 0 0 1 1
use contact_32  contact_32_5211
timestamp 1624857261
transform 1 0 23528 0 1 101053
box 0 0 1 1
use contact_32  contact_32_5210
timestamp 1624857261
transform 1 0 23528 0 1 101325
box 0 0 1 1
use contact_32  contact_32_5209
timestamp 1624857261
transform 1 0 23392 0 1 86093
box 0 0 1 1
use contact_32  contact_32_5208
timestamp 1624857261
transform 1 0 23392 0 1 86365
box 0 0 1 1
use contact_32  contact_32_5207
timestamp 1624857261
transform 1 0 23392 0 1 85957
box 0 0 1 1
use contact_32  contact_32_5206
timestamp 1624857261
transform 1 0 23392 0 1 85685
box 0 0 1 1
use contact_32  contact_32_5205
timestamp 1624857261
transform 1 0 23392 0 1 32645
box 0 0 1 1
use contact_32  contact_32_5204
timestamp 1624857261
transform 1 0 23392 0 1 32373
box 0 0 1 1
use contact_32  contact_32_5203
timestamp 1624857261
transform 1 0 23528 0 1 88813
box 0 0 1 1
use contact_32  contact_32_5202
timestamp 1624857261
transform 1 0 23528 0 1 89085
box 0 0 1 1
use contact_32  contact_32_5201
timestamp 1624857261
transform 1 0 23528 0 1 47741
box 0 0 1 1
use contact_32  contact_32_5200
timestamp 1624857261
transform 1 0 23528 0 1 48013
box 0 0 1 1
use contact_32  contact_32_5199
timestamp 1624857261
transform 1 0 23528 0 1 42165
box 0 0 1 1
use contact_32  contact_32_5198
timestamp 1624857261
transform 1 0 23528 0 1 41893
box 0 0 1 1
use contact_32  contact_32_5197
timestamp 1624857261
transform 1 0 23392 0 1 60253
box 0 0 1 1
use contact_32  contact_32_5196
timestamp 1624857261
transform 1 0 23392 0 1 59981
box 0 0 1 1
use contact_32  contact_32_5195
timestamp 1624857261
transform 1 0 23392 0 1 77389
box 0 0 1 1
use contact_32  contact_32_5194
timestamp 1624857261
transform 1 0 23392 0 1 77661
box 0 0 1 1
use contact_32  contact_32_5193
timestamp 1624857261
transform 1 0 23528 0 1 105405
box 0 0 1 1
use contact_32  contact_32_5192
timestamp 1624857261
transform 1 0 23528 0 1 105677
box 0 0 1 1
use contact_32  contact_32_5191
timestamp 1624857261
transform 1 0 23392 0 1 122269
box 0 0 1 1
use contact_32  contact_32_5190
timestamp 1624857261
transform 1 0 23392 0 1 121997
box 0 0 1 1
use contact_32  contact_32_5189
timestamp 1624857261
transform 1 0 23528 0 1 122405
box 0 0 1 1
use contact_32  contact_32_5188
timestamp 1624857261
transform 1 0 23528 0 1 122677
box 0 0 1 1
use contact_32  contact_32_5187
timestamp 1624857261
transform 1 0 23392 0 1 95885
box 0 0 1 1
use contact_32  contact_32_5186
timestamp 1624857261
transform 1 0 23392 0 1 95613
box 0 0 1 1
use contact_32  contact_32_5185
timestamp 1624857261
transform 1 0 23392 0 1 118733
box 0 0 1 1
use contact_32  contact_32_5184
timestamp 1624857261
transform 1 0 23392 0 1 118461
box 0 0 1 1
use contact_32  contact_32_5183
timestamp 1624857261
transform 1 0 23392 0 1 78613
box 0 0 1 1
use contact_32  contact_32_5182
timestamp 1624857261
transform 1 0 23392 0 1 78885
box 0 0 1 1
use contact_32  contact_32_5181
timestamp 1624857261
transform 1 0 23392 0 1 78477
box 0 0 1 1
use contact_32  contact_32_5180
timestamp 1624857261
transform 1 0 23392 0 1 78205
box 0 0 1 1
use contact_32  contact_32_5179
timestamp 1624857261
transform 1 0 23392 0 1 72221
box 0 0 1 1
use contact_32  contact_32_5178
timestamp 1624857261
transform 1 0 23392 0 1 72493
box 0 0 1 1
use contact_32  contact_32_5177
timestamp 1624857261
transform 1 0 23392 0 1 80789
box 0 0 1 1
use contact_32  contact_32_5176
timestamp 1624857261
transform 1 0 23392 0 1 80517
box 0 0 1 1
use contact_32  contact_32_5175
timestamp 1624857261
transform 1 0 23528 0 1 90853
box 0 0 1 1
use contact_32  contact_32_5174
timestamp 1624857261
transform 1 0 23528 0 1 91125
box 0 0 1 1
use contact_32  contact_32_5173
timestamp 1624857261
transform 1 0 23392 0 1 90717
box 0 0 1 1
use contact_32  contact_32_5172
timestamp 1624857261
transform 1 0 23392 0 1 90445
box 0 0 1 1
use contact_32  contact_32_5171
timestamp 1624857261
transform 1 0 23392 0 1 114517
box 0 0 1 1
use contact_32  contact_32_5170
timestamp 1624857261
transform 1 0 23392 0 1 114789
box 0 0 1 1
use contact_32  contact_32_5169
timestamp 1624857261
transform 1 0 23392 0 1 53725
box 0 0 1 1
use contact_32  contact_32_5168
timestamp 1624857261
transform 1 0 23392 0 1 53997
box 0 0 1 1
use contact_32  contact_32_5167
timestamp 1624857261
transform 1 0 23528 0 1 118325
box 0 0 1 1
use contact_32  contact_32_5166
timestamp 1624857261
transform 1 0 23528 0 1 118053
box 0 0 1 1
use contact_32  contact_32_5165
timestamp 1624857261
transform 1 0 23528 0 1 101869
box 0 0 1 1
use contact_32  contact_32_5164
timestamp 1624857261
transform 1 0 23528 0 1 102141
box 0 0 1 1
use contact_32  contact_32_5163
timestamp 1624857261
transform 1 0 23528 0 1 101733
box 0 0 1 1
use contact_32  contact_32_5162
timestamp 1624857261
transform 1 0 23528 0 1 101461
box 0 0 1 1
use contact_32  contact_32_5161
timestamp 1624857261
transform 1 0 23528 0 1 116149
box 0 0 1 1
use contact_32  contact_32_5160
timestamp 1624857261
transform 1 0 23528 0 1 116421
box 0 0 1 1
use contact_32  contact_32_5159
timestamp 1624857261
transform 1 0 23528 0 1 97517
box 0 0 1 1
use contact_32  contact_32_5158
timestamp 1624857261
transform 1 0 23528 0 1 97789
box 0 0 1 1
use contact_32  contact_32_5157
timestamp 1624857261
transform 1 0 23528 0 1 97381
box 0 0 1 1
use contact_32  contact_32_5156
timestamp 1624857261
transform 1 0 23528 0 1 97109
box 0 0 1 1
use contact_32  contact_32_5155
timestamp 1624857261
transform 1 0 23528 0 1 72629
box 0 0 1 1
use contact_32  contact_32_5154
timestamp 1624857261
transform 1 0 23528 0 1 72901
box 0 0 1 1
use contact_32  contact_32_5153
timestamp 1624857261
transform 1 0 23528 0 1 31013
box 0 0 1 1
use contact_32  contact_32_5152
timestamp 1624857261
transform 1 0 23528 0 1 30741
box 0 0 1 1
use contact_32  contact_32_5151
timestamp 1624857261
transform 1 0 23528 0 1 31149
box 0 0 1 1
use contact_32  contact_32_5150
timestamp 1624857261
transform 1 0 23528 0 1 31421
box 0 0 1 1
use contact_32  contact_32_5149
timestamp 1624857261
transform 1 0 23392 0 1 93845
box 0 0 1 1
use contact_32  contact_32_5148
timestamp 1624857261
transform 1 0 23392 0 1 93573
box 0 0 1 1
use contact_32  contact_32_5147
timestamp 1624857261
transform 1 0 23528 0 1 95205
box 0 0 1 1
use contact_32  contact_32_5146
timestamp 1624857261
transform 1 0 23528 0 1 95477
box 0 0 1 1
use contact_32  contact_32_5145
timestamp 1624857261
transform 1 0 23392 0 1 95069
box 0 0 1 1
use contact_32  contact_32_5144
timestamp 1624857261
transform 1 0 23392 0 1 94797
box 0 0 1 1
use contact_32  contact_32_5143
timestamp 1624857261
transform 1 0 23392 0 1 50461
box 0 0 1 1
use contact_32  contact_32_5142
timestamp 1624857261
transform 1 0 23392 0 1 50189
box 0 0 1 1
use contact_32  contact_32_5141
timestamp 1624857261
transform 1 0 23528 0 1 86501
box 0 0 1 1
use contact_32  contact_32_5140
timestamp 1624857261
transform 1 0 23528 0 1 86773
box 0 0 1 1
use contact_32  contact_32_5139
timestamp 1624857261
transform 1 0 23528 0 1 44205
box 0 0 1 1
use contact_32  contact_32_5138
timestamp 1624857261
transform 1 0 23528 0 1 44477
box 0 0 1 1
use contact_32  contact_32_5137
timestamp 1624857261
transform 1 0 23528 0 1 44069
box 0 0 1 1
use contact_32  contact_32_5136
timestamp 1624857261
transform 1 0 23528 0 1 43797
box 0 0 1 1
use contact_32  contact_32_5135
timestamp 1624857261
transform 1 0 23528 0 1 56309
box 0 0 1 1
use contact_32  contact_32_5134
timestamp 1624857261
transform 1 0 23528 0 1 56037
box 0 0 1 1
use contact_32  contact_32_5133
timestamp 1624857261
transform 1 0 23528 0 1 56445
box 0 0 1 1
use contact_32  contact_32_5132
timestamp 1624857261
transform 1 0 23528 0 1 56717
box 0 0 1 1
use contact_32  contact_32_5131
timestamp 1624857261
transform 1 0 23392 0 1 110981
box 0 0 1 1
use contact_32  contact_32_5130
timestamp 1624857261
transform 1 0 23392 0 1 111253
box 0 0 1 1
use contact_32  contact_32_5129
timestamp 1624857261
transform 1 0 23528 0 1 89901
box 0 0 1 1
use contact_32  contact_32_5128
timestamp 1624857261
transform 1 0 23528 0 1 89629
box 0 0 1 1
use contact_32  contact_32_5127
timestamp 1624857261
transform 1 0 23528 0 1 90037
box 0 0 1 1
use contact_32  contact_32_5126
timestamp 1624857261
transform 1 0 23528 0 1 90309
box 0 0 1 1
use contact_32  contact_32_5125
timestamp 1624857261
transform 1 0 23392 0 1 35909
box 0 0 1 1
use contact_32  contact_32_5124
timestamp 1624857261
transform 1 0 23392 0 1 36181
box 0 0 1 1
use contact_32  contact_32_5123
timestamp 1624857261
transform 1 0 23528 0 1 35773
box 0 0 1 1
use contact_32  contact_32_5122
timestamp 1624857261
transform 1 0 23528 0 1 35501
box 0 0 1 1
use contact_32  contact_32_5121
timestamp 1624857261
transform 1 0 23528 0 1 58485
box 0 0 1 1
use contact_32  contact_32_5120
timestamp 1624857261
transform 1 0 23528 0 1 58757
box 0 0 1 1
use contact_32  contact_32_5119
timestamp 1624857261
transform 1 0 23528 0 1 58349
box 0 0 1 1
use contact_32  contact_32_5118
timestamp 1624857261
transform 1 0 23528 0 1 58077
box 0 0 1 1
use contact_32  contact_32_5117
timestamp 1624857261
transform 1 0 23392 0 1 49237
box 0 0 1 1
use contact_32  contact_32_5116
timestamp 1624857261
transform 1 0 23392 0 1 48965
box 0 0 1 1
use contact_32  contact_32_5115
timestamp 1624857261
transform 1 0 23392 0 1 49373
box 0 0 1 1
use contact_32  contact_32_5114
timestamp 1624857261
transform 1 0 23392 0 1 49645
box 0 0 1 1
use contact_32  contact_32_5113
timestamp 1624857261
transform 1 0 23392 0 1 55901
box 0 0 1 1
use contact_32  contact_32_5112
timestamp 1624857261
transform 1 0 23392 0 1 55629
box 0 0 1 1
use contact_32  contact_32_5111
timestamp 1624857261
transform 1 0 23392 0 1 50053
box 0 0 1 1
use contact_32  contact_32_5110
timestamp 1624857261
transform 1 0 23392 0 1 49781
box 0 0 1 1
use contact_32  contact_32_5109
timestamp 1624857261
transform 1 0 23528 0 1 106493
box 0 0 1 1
use contact_32  contact_32_5108
timestamp 1624857261
transform 1 0 23528 0 1 106221
box 0 0 1 1
use contact_32  contact_32_5107
timestamp 1624857261
transform 1 0 23528 0 1 40125
box 0 0 1 1
use contact_32  contact_32_5106
timestamp 1624857261
transform 1 0 23528 0 1 39853
box 0 0 1 1
use contact_32  contact_32_5105
timestamp 1624857261
transform 1 0 23392 0 1 40261
box 0 0 1 1
use contact_32  contact_32_5104
timestamp 1624857261
transform 1 0 23392 0 1 40533
box 0 0 1 1
use contact_32  contact_32_5103
timestamp 1624857261
transform 1 0 23528 0 1 109349
box 0 0 1 1
use contact_32  contact_32_5102
timestamp 1624857261
transform 1 0 23528 0 1 109621
box 0 0 1 1
use contact_32  contact_32_5101
timestamp 1624857261
transform 1 0 23528 0 1 57125
box 0 0 1 1
use contact_32  contact_32_5100
timestamp 1624857261
transform 1 0 23528 0 1 56853
box 0 0 1 1
use contact_32  contact_32_5099
timestamp 1624857261
transform 1 0 23528 0 1 65965
box 0 0 1 1
use contact_32  contact_32_5098
timestamp 1624857261
transform 1 0 23528 0 1 66237
box 0 0 1 1
use contact_32  contact_32_5097
timestamp 1624857261
transform 1 0 23392 0 1 112069
box 0 0 1 1
use contact_32  contact_32_5096
timestamp 1624857261
transform 1 0 23392 0 1 111797
box 0 0 1 1
use contact_32  contact_32_5095
timestamp 1624857261
transform 1 0 23392 0 1 112205
box 0 0 1 1
use contact_32  contact_32_5094
timestamp 1624857261
transform 1 0 23392 0 1 112477
box 0 0 1 1
use contact_32  contact_32_5093
timestamp 1624857261
transform 1 0 23528 0 1 69501
box 0 0 1 1
use contact_32  contact_32_5092
timestamp 1624857261
transform 1 0 23528 0 1 69773
box 0 0 1 1
use contact_32  contact_32_5091
timestamp 1624857261
transform 1 0 23528 0 1 26797
box 0 0 1 1
use contact_32  contact_32_5090
timestamp 1624857261
transform 1 0 23528 0 1 27069
box 0 0 1 1
use contact_32  contact_32_5089
timestamp 1624857261
transform 1 0 23528 0 1 103909
box 0 0 1 1
use contact_32  contact_32_5088
timestamp 1624857261
transform 1 0 23528 0 1 104181
box 0 0 1 1
use contact_32  contact_32_5087
timestamp 1624857261
transform 1 0 23528 0 1 51685
box 0 0 1 1
use contact_32  contact_32_5086
timestamp 1624857261
transform 1 0 23528 0 1 51957
box 0 0 1 1
use contact_32  contact_32_5085
timestamp 1624857261
transform 1 0 23392 0 1 44613
box 0 0 1 1
use contact_32  contact_32_5084
timestamp 1624857261
transform 1 0 23392 0 1 44885
box 0 0 1 1
use contact_32  contact_32_5083
timestamp 1624857261
transform 1 0 23392 0 1 27613
box 0 0 1 1
use contact_32  contact_32_5082
timestamp 1624857261
transform 1 0 23392 0 1 27885
box 0 0 1 1
use contact_32  contact_32_5081
timestamp 1624857261
transform 1 0 23392 0 1 27477
box 0 0 1 1
use contact_32  contact_32_5080
timestamp 1624857261
transform 1 0 23392 0 1 27205
box 0 0 1 1
use contact_32  contact_32_5079
timestamp 1624857261
transform 1 0 23528 0 1 73717
box 0 0 1 1
use contact_32  contact_32_5078
timestamp 1624857261
transform 1 0 23528 0 1 73445
box 0 0 1 1
use contact_32  contact_32_5077
timestamp 1624857261
transform 1 0 23528 0 1 73853
box 0 0 1 1
use contact_32  contact_32_5076
timestamp 1624857261
transform 1 0 23528 0 1 74125
box 0 0 1 1
use contact_32  contact_32_5075
timestamp 1624857261
transform 1 0 23392 0 1 28293
box 0 0 1 1
use contact_32  contact_32_5074
timestamp 1624857261
transform 1 0 23392 0 1 28021
box 0 0 1 1
use contact_32  contact_32_5073
timestamp 1624857261
transform 1 0 23392 0 1 28429
box 0 0 1 1
use contact_32  contact_32_5072
timestamp 1624857261
transform 1 0 23392 0 1 28701
box 0 0 1 1
use contact_32  contact_32_5071
timestamp 1624857261
transform 1 0 23528 0 1 87589
box 0 0 1 1
use contact_32  contact_32_5070
timestamp 1624857261
transform 1 0 23528 0 1 87317
box 0 0 1 1
use contact_32  contact_32_5069
timestamp 1624857261
transform 1 0 23392 0 1 117917
box 0 0 1 1
use contact_32  contact_32_5068
timestamp 1624857261
transform 1 0 23392 0 1 117645
box 0 0 1 1
use contact_32  contact_32_5067
timestamp 1624857261
transform 1 0 23392 0 1 25301
box 0 0 1 1
use contact_32  contact_32_5066
timestamp 1624857261
transform 1 0 23392 0 1 25573
box 0 0 1 1
use contact_32  contact_32_5065
timestamp 1624857261
transform 1 0 23392 0 1 25165
box 0 0 1 1
use contact_32  contact_32_5064
timestamp 1624857261
transform 1 0 23392 0 1 24757
box 0 0 1 1
use contact_32  contact_32_5063
timestamp 1624857261
transform 1 0 23528 0 1 65013
box 0 0 1 1
use contact_32  contact_32_5062
timestamp 1624857261
transform 1 0 23528 0 1 64741
box 0 0 1 1
use contact_32  contact_32_5061
timestamp 1624857261
transform 1 0 23528 0 1 93165
box 0 0 1 1
use contact_32  contact_32_5060
timestamp 1624857261
transform 1 0 23528 0 1 93437
box 0 0 1 1
use contact_32  contact_32_5059
timestamp 1624857261
transform 1 0 23392 0 1 43661
box 0 0 1 1
use contact_32  contact_32_5058
timestamp 1624857261
transform 1 0 23392 0 1 43389
box 0 0 1 1
use contact_32  contact_32_5057
timestamp 1624857261
transform 1 0 23392 0 1 29517
box 0 0 1 1
use contact_32  contact_32_5056
timestamp 1624857261
transform 1 0 23392 0 1 29245
box 0 0 1 1
use contact_32  contact_32_5055
timestamp 1624857261
transform 1 0 23392 0 1 29653
box 0 0 1 1
use contact_32  contact_32_5054
timestamp 1624857261
transform 1 0 23392 0 1 29925
box 0 0 1 1
use contact_32  contact_32_5053
timestamp 1624857261
transform 1 0 23392 0 1 87181
box 0 0 1 1
use contact_32  contact_32_5052
timestamp 1624857261
transform 1 0 23392 0 1 86909
box 0 0 1 1
use contact_32  contact_32_5051
timestamp 1624857261
transform 1 0 23528 0 1 123901
box 0 0 1 1
use contact_32  contact_32_5050
timestamp 1624857261
transform 1 0 23528 0 1 123629
box 0 0 1 1
use contact_32  contact_32_5049
timestamp 1624857261
transform 1 0 23392 0 1 73309
box 0 0 1 1
use contact_32  contact_32_5048
timestamp 1624857261
transform 1 0 23392 0 1 73037
box 0 0 1 1
use contact_32  contact_32_5047
timestamp 1624857261
transform 1 0 23392 0 1 54405
box 0 0 1 1
use contact_32  contact_32_5046
timestamp 1624857261
transform 1 0 23392 0 1 54133
box 0 0 1 1
use contact_32  contact_32_5045
timestamp 1624857261
transform 1 0 23528 0 1 84733
box 0 0 1 1
use contact_32  contact_32_5044
timestamp 1624857261
transform 1 0 23528 0 1 84461
box 0 0 1 1
use contact_32  contact_32_5043
timestamp 1624857261
transform 1 0 23392 0 1 84869
box 0 0 1 1
use contact_32  contact_32_5042
timestamp 1624857261
transform 1 0 23392 0 1 85141
box 0 0 1 1
use contact_32  contact_32_5041
timestamp 1624857261
transform 1 0 23528 0 1 68277
box 0 0 1 1
use contact_32  contact_32_5040
timestamp 1624857261
transform 1 0 23528 0 1 68549
box 0 0 1 1
use contact_32  contact_32_5039
timestamp 1624857261
transform 1 0 23392 0 1 89221
box 0 0 1 1
use contact_32  contact_32_5038
timestamp 1624857261
transform 1 0 23392 0 1 89493
box 0 0 1 1
use contact_32  contact_32_5037
timestamp 1624857261
transform 1 0 23392 0 1 97925
box 0 0 1 1
use contact_32  contact_32_5036
timestamp 1624857261
transform 1 0 23392 0 1 98197
box 0 0 1 1
use contact_32  contact_32_5035
timestamp 1624857261
transform 1 0 23528 0 1 77797
box 0 0 1 1
use contact_32  contact_32_5034
timestamp 1624857261
transform 1 0 23528 0 1 78069
box 0 0 1 1
use contact_32  contact_32_5033
timestamp 1624857261
transform 1 0 23528 0 1 70181
box 0 0 1 1
use contact_32  contact_32_5032
timestamp 1624857261
transform 1 0 23528 0 1 69909
box 0 0 1 1
use contact_32  contact_32_5031
timestamp 1624857261
transform 1 0 23392 0 1 66781
box 0 0 1 1
use contact_32  contact_32_5030
timestamp 1624857261
transform 1 0 23392 0 1 67053
box 0 0 1 1
use contact_32  contact_32_5029
timestamp 1624857261
transform 1 0 23392 0 1 66645
box 0 0 1 1
use contact_32  contact_32_5028
timestamp 1624857261
transform 1 0 23392 0 1 66373
box 0 0 1 1
use contact_32  contact_32_5027
timestamp 1624857261
transform 1 0 23528 0 1 111661
box 0 0 1 1
use contact_32  contact_32_5026
timestamp 1624857261
transform 1 0 23528 0 1 111389
box 0 0 1 1
use contact_32  contact_32_5025
timestamp 1624857261
transform 1 0 23528 0 1 123493
box 0 0 1 1
use contact_32  contact_32_5024
timestamp 1624857261
transform 1 0 23528 0 1 123221
box 0 0 1 1
use contact_32  contact_32_5023
timestamp 1624857261
transform 1 0 23528 0 1 91261
box 0 0 1 1
use contact_32  contact_32_5022
timestamp 1624857261
transform 1 0 23528 0 1 91533
box 0 0 1 1
use contact_32  contact_32_5021
timestamp 1624857261
transform 1 0 23528 0 1 29109
box 0 0 1 1
use contact_32  contact_32_5020
timestamp 1624857261
transform 1 0 23528 0 1 28837
box 0 0 1 1
use contact_32  contact_32_5019
timestamp 1624857261
transform 1 0 23528 0 1 33597
box 0 0 1 1
use contact_32  contact_32_5018
timestamp 1624857261
transform 1 0 23528 0 1 33869
box 0 0 1 1
use contact_32  contact_32_5017
timestamp 1624857261
transform 1 0 23528 0 1 40941
box 0 0 1 1
use contact_32  contact_32_5016
timestamp 1624857261
transform 1 0 23528 0 1 40669
box 0 0 1 1
use contact_32  contact_32_5015
timestamp 1624857261
transform 1 0 23528 0 1 32237
box 0 0 1 1
use contact_32  contact_32_5014
timestamp 1624857261
transform 1 0 23528 0 1 31965
box 0 0 1 1
use contact_32  contact_32_5013
timestamp 1624857261
transform 1 0 23392 0 1 31829
box 0 0 1 1
use contact_32  contact_32_5012
timestamp 1624857261
transform 1 0 23392 0 1 31557
box 0 0 1 1
use contact_32  contact_32_5011
timestamp 1624857261
transform 1 0 23392 0 1 123085
box 0 0 1 1
use contact_32  contact_32_5010
timestamp 1624857261
transform 1 0 23392 0 1 122813
box 0 0 1 1
use contact_32  contact_32_5009
timestamp 1624857261
transform 1 0 23528 0 1 74533
box 0 0 1 1
use contact_32  contact_32_5008
timestamp 1624857261
transform 1 0 23528 0 1 74261
box 0 0 1 1
use contact_32  contact_32_5007
timestamp 1624857261
transform 1 0 23392 0 1 38221
box 0 0 1 1
use contact_32  contact_32_5006
timestamp 1624857261
transform 1 0 23392 0 1 37949
box 0 0 1 1
use contact_32  contact_32_5005
timestamp 1624857261
transform 1 0 23528 0 1 106085
box 0 0 1 1
use contact_32  contact_32_5004
timestamp 1624857261
transform 1 0 23528 0 1 105813
box 0 0 1 1
use contact_32  contact_32_5003
timestamp 1624857261
transform 1 0 23392 0 1 85277
box 0 0 1 1
use contact_32  contact_32_5002
timestamp 1624857261
transform 1 0 23392 0 1 85549
box 0 0 1 1
use contact_32  contact_32_5001
timestamp 1624857261
transform 1 0 29512 0 1 15101
box 0 0 1 1
use contact_32  contact_32_5000
timestamp 1624857261
transform 1 0 29512 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4999
timestamp 1624857261
transform 1 0 29376 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4998
timestamp 1624857261
transform 1 0 29376 0 1 24349
box 0 0 1 1
use contact_32  contact_32_4997
timestamp 1624857261
transform 1 0 29648 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4996
timestamp 1624857261
transform 1 0 29648 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4995
timestamp 1624857261
transform 1 0 29648 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4994
timestamp 1624857261
transform 1 0 29648 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4993
timestamp 1624857261
transform 1 0 29648 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4992
timestamp 1624857261
transform 1 0 29648 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4991
timestamp 1624857261
transform 1 0 29648 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4990
timestamp 1624857261
transform 1 0 29648 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4989
timestamp 1624857261
transform 1 0 29920 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4988
timestamp 1624857261
transform 1 0 29920 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4987
timestamp 1624857261
transform 1 0 29784 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4986
timestamp 1624857261
transform 1 0 29784 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4985
timestamp 1624857261
transform 1 0 29784 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4984
timestamp 1624857261
transform 1 0 29784 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4983
timestamp 1624857261
transform 1 0 30600 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4982
timestamp 1624857261
transform 1 0 30600 0 1 24349
box 0 0 1 1
use contact_32  contact_32_4981
timestamp 1624857261
transform 1 0 30872 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4980
timestamp 1624857261
transform 1 0 30872 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4979
timestamp 1624857261
transform 1 0 31688 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4978
timestamp 1624857261
transform 1 0 31688 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4977
timestamp 1624857261
transform 1 0 32232 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4976
timestamp 1624857261
transform 1 0 32232 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4975
timestamp 1624857261
transform 1 0 32912 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4974
timestamp 1624857261
transform 1 0 32912 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4973
timestamp 1624857261
transform 1 0 32912 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4972
timestamp 1624857261
transform 1 0 32912 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4971
timestamp 1624857261
transform 1 0 33456 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4970
timestamp 1624857261
transform 1 0 33456 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4969
timestamp 1624857261
transform 1 0 33456 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4968
timestamp 1624857261
transform 1 0 33456 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4967
timestamp 1624857261
transform 1 0 34136 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4966
timestamp 1624857261
transform 1 0 34136 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4965
timestamp 1624857261
transform 1 0 34136 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4964
timestamp 1624857261
transform 1 0 34136 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4963
timestamp 1624857261
transform 1 0 34680 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4962
timestamp 1624857261
transform 1 0 34680 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4961
timestamp 1624857261
transform 1 0 34680 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4960
timestamp 1624857261
transform 1 0 34680 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4959
timestamp 1624857261
transform 1 0 34816 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4958
timestamp 1624857261
transform 1 0 34816 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4957
timestamp 1624857261
transform 1 0 34816 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4956
timestamp 1624857261
transform 1 0 34816 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4955
timestamp 1624857261
transform 1 0 34680 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4954
timestamp 1624857261
transform 1 0 34680 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4953
timestamp 1624857261
transform 1 0 35768 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4952
timestamp 1624857261
transform 1 0 35768 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4951
timestamp 1624857261
transform 1 0 34680 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4950
timestamp 1624857261
transform 1 0 34680 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4949
timestamp 1624857261
transform 1 0 35496 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4948
timestamp 1624857261
transform 1 0 35496 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4947
timestamp 1624857261
transform 1 0 35904 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4946
timestamp 1624857261
transform 1 0 35904 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4945
timestamp 1624857261
transform 1 0 36584 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4944
timestamp 1624857261
transform 1 0 36584 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4943
timestamp 1624857261
transform 1 0 37128 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4942
timestamp 1624857261
transform 1 0 37128 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4941
timestamp 1624857261
transform 1 0 37128 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4940
timestamp 1624857261
transform 1 0 37128 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4939
timestamp 1624857261
transform 1 0 38080 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4938
timestamp 1624857261
transform 1 0 38080 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4937
timestamp 1624857261
transform 1 0 38488 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4936
timestamp 1624857261
transform 1 0 38488 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4935
timestamp 1624857261
transform 1 0 39304 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4934
timestamp 1624857261
transform 1 0 39304 0 1 24349
box 0 0 1 1
use contact_32  contact_32_4933
timestamp 1624857261
transform 1 0 39440 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4932
timestamp 1624857261
transform 1 0 39440 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4931
timestamp 1624857261
transform 1 0 39712 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4930
timestamp 1624857261
transform 1 0 39712 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4929
timestamp 1624857261
transform 1 0 39712 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4928
timestamp 1624857261
transform 1 0 39712 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4927
timestamp 1624857261
transform 1 0 39712 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4926
timestamp 1624857261
transform 1 0 39712 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4925
timestamp 1624857261
transform 1 0 39712 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4924
timestamp 1624857261
transform 1 0 39712 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4923
timestamp 1624857261
transform 1 0 39712 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4922
timestamp 1624857261
transform 1 0 39712 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4921
timestamp 1624857261
transform 1 0 39712 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4920
timestamp 1624857261
transform 1 0 39712 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4919
timestamp 1624857261
transform 1 0 40392 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4918
timestamp 1624857261
transform 1 0 40392 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4917
timestamp 1624857261
transform 1 0 40936 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4916
timestamp 1624857261
transform 1 0 40936 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4915
timestamp 1624857261
transform 1 0 41616 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4914
timestamp 1624857261
transform 1 0 41616 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4913
timestamp 1624857261
transform 1 0 41616 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4912
timestamp 1624857261
transform 1 0 41616 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4911
timestamp 1624857261
transform 1 0 42160 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4910
timestamp 1624857261
transform 1 0 42160 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4909
timestamp 1624857261
transform 1 0 42976 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4908
timestamp 1624857261
transform 1 0 42976 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4907
timestamp 1624857261
transform 1 0 43248 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4906
timestamp 1624857261
transform 1 0 43248 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4905
timestamp 1624857261
transform 1 0 42840 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4904
timestamp 1624857261
transform 1 0 42840 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4903
timestamp 1624857261
transform 1 0 44336 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4902
timestamp 1624857261
transform 1 0 44336 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4901
timestamp 1624857261
transform 1 0 44608 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4900
timestamp 1624857261
transform 1 0 44608 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4899
timestamp 1624857261
transform 1 0 44608 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4898
timestamp 1624857261
transform 1 0 44608 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4897
timestamp 1624857261
transform 1 0 44744 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4896
timestamp 1624857261
transform 1 0 44744 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4895
timestamp 1624857261
transform 1 0 44880 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4894
timestamp 1624857261
transform 1 0 44880 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4893
timestamp 1624857261
transform 1 0 44744 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4892
timestamp 1624857261
transform 1 0 44744 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4891
timestamp 1624857261
transform 1 0 44744 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4890
timestamp 1624857261
transform 1 0 44744 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4889
timestamp 1624857261
transform 1 0 45424 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4888
timestamp 1624857261
transform 1 0 45424 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4887
timestamp 1624857261
transform 1 0 45424 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4886
timestamp 1624857261
transform 1 0 45424 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4885
timestamp 1624857261
transform 1 0 45424 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4884
timestamp 1624857261
transform 1 0 45424 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4883
timestamp 1624857261
transform 1 0 45968 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4882
timestamp 1624857261
transform 1 0 45968 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4881
timestamp 1624857261
transform 1 0 46648 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4880
timestamp 1624857261
transform 1 0 46648 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4879
timestamp 1624857261
transform 1 0 46784 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4878
timestamp 1624857261
transform 1 0 46784 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4877
timestamp 1624857261
transform 1 0 47192 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4876
timestamp 1624857261
transform 1 0 47192 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4875
timestamp 1624857261
transform 1 0 48008 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4874
timestamp 1624857261
transform 1 0 48008 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4873
timestamp 1624857261
transform 1 0 48416 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4872
timestamp 1624857261
transform 1 0 48416 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4871
timestamp 1624857261
transform 1 0 49096 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4870
timestamp 1624857261
transform 1 0 49096 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4869
timestamp 1624857261
transform 1 0 49368 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4868
timestamp 1624857261
transform 1 0 49368 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4867
timestamp 1624857261
transform 1 0 49640 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4866
timestamp 1624857261
transform 1 0 49640 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4865
timestamp 1624857261
transform 1 0 49776 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4864
timestamp 1624857261
transform 1 0 49776 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4863
timestamp 1624857261
transform 1 0 49776 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4862
timestamp 1624857261
transform 1 0 49776 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4861
timestamp 1624857261
transform 1 0 49640 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4860
timestamp 1624857261
transform 1 0 49640 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4859
timestamp 1624857261
transform 1 0 50728 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4858
timestamp 1624857261
transform 1 0 50728 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4857
timestamp 1624857261
transform 1 0 49640 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4856
timestamp 1624857261
transform 1 0 49640 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4855
timestamp 1624857261
transform 1 0 50456 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4854
timestamp 1624857261
transform 1 0 50456 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4853
timestamp 1624857261
transform 1 0 50320 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4852
timestamp 1624857261
transform 1 0 50320 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4851
timestamp 1624857261
transform 1 0 50864 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4850
timestamp 1624857261
transform 1 0 50864 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4849
timestamp 1624857261
transform 1 0 50864 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4848
timestamp 1624857261
transform 1 0 50864 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4847
timestamp 1624857261
transform 1 0 51680 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4846
timestamp 1624857261
transform 1 0 51680 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4845
timestamp 1624857261
transform 1 0 52224 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4844
timestamp 1624857261
transform 1 0 52224 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4843
timestamp 1624857261
transform 1 0 52768 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4842
timestamp 1624857261
transform 1 0 52768 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4841
timestamp 1624857261
transform 1 0 52904 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4840
timestamp 1624857261
transform 1 0 52904 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4839
timestamp 1624857261
transform 1 0 53312 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4838
timestamp 1624857261
transform 1 0 53312 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4837
timestamp 1624857261
transform 1 0 54128 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4836
timestamp 1624857261
transform 1 0 54128 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4835
timestamp 1624857261
transform 1 0 54264 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4834
timestamp 1624857261
transform 1 0 54264 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4833
timestamp 1624857261
transform 1 0 54672 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4832
timestamp 1624857261
transform 1 0 54672 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4831
timestamp 1624857261
transform 1 0 54672 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4830
timestamp 1624857261
transform 1 0 54672 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4829
timestamp 1624857261
transform 1 0 54672 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4828
timestamp 1624857261
transform 1 0 54672 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4827
timestamp 1624857261
transform 1 0 54808 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4826
timestamp 1624857261
transform 1 0 54808 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4825
timestamp 1624857261
transform 1 0 54808 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4824
timestamp 1624857261
transform 1 0 54808 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4823
timestamp 1624857261
transform 1 0 54672 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4822
timestamp 1624857261
transform 1 0 54672 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4821
timestamp 1624857261
transform 1 0 54672 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4820
timestamp 1624857261
transform 1 0 54672 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4819
timestamp 1624857261
transform 1 0 55352 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4818
timestamp 1624857261
transform 1 0 55352 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4817
timestamp 1624857261
transform 1 0 55352 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4816
timestamp 1624857261
transform 1 0 55352 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4815
timestamp 1624857261
transform 1 0 55896 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4814
timestamp 1624857261
transform 1 0 55896 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4813
timestamp 1624857261
transform 1 0 56576 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4812
timestamp 1624857261
transform 1 0 56576 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4811
timestamp 1624857261
transform 1 0 57120 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4810
timestamp 1624857261
transform 1 0 57120 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4809
timestamp 1624857261
transform 1 0 57800 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4808
timestamp 1624857261
transform 1 0 57800 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4807
timestamp 1624857261
transform 1 0 58072 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4806
timestamp 1624857261
transform 1 0 58072 0 1 24349
box 0 0 1 1
use contact_32  contact_32_4805
timestamp 1624857261
transform 1 0 59704 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4804
timestamp 1624857261
transform 1 0 59704 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4803
timestamp 1624857261
transform 1 0 59568 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4802
timestamp 1624857261
transform 1 0 59568 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4801
timestamp 1624857261
transform 1 0 59704 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4800
timestamp 1624857261
transform 1 0 59704 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4799
timestamp 1624857261
transform 1 0 59840 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4798
timestamp 1624857261
transform 1 0 59840 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4797
timestamp 1624857261
transform 1 0 59704 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4796
timestamp 1624857261
transform 1 0 59704 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4795
timestamp 1624857261
transform 1 0 60792 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4794
timestamp 1624857261
transform 1 0 60792 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4793
timestamp 1624857261
transform 1 0 59704 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4792
timestamp 1624857261
transform 1 0 59704 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4791
timestamp 1624857261
transform 1 0 60792 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4790
timestamp 1624857261
transform 1 0 60792 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4789
timestamp 1624857261
transform 1 0 60384 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4788
timestamp 1624857261
transform 1 0 60384 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4787
timestamp 1624857261
transform 1 0 60928 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4786
timestamp 1624857261
transform 1 0 60928 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4785
timestamp 1624857261
transform 1 0 61472 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4784
timestamp 1624857261
transform 1 0 61472 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4783
timestamp 1624857261
transform 1 0 61608 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4782
timestamp 1624857261
transform 1 0 61608 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4781
timestamp 1624857261
transform 1 0 61608 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4780
timestamp 1624857261
transform 1 0 61608 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4779
timestamp 1624857261
transform 1 0 62152 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4778
timestamp 1624857261
transform 1 0 62152 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4777
timestamp 1624857261
transform 1 0 62152 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4776
timestamp 1624857261
transform 1 0 62152 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4775
timestamp 1624857261
transform 1 0 62832 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4774
timestamp 1624857261
transform 1 0 62832 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4773
timestamp 1624857261
transform 1 0 62832 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4772
timestamp 1624857261
transform 1 0 62832 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4771
timestamp 1624857261
transform 1 0 63376 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4770
timestamp 1624857261
transform 1 0 63376 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4769
timestamp 1624857261
transform 1 0 64056 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4768
timestamp 1624857261
transform 1 0 64056 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4767
timestamp 1624857261
transform 1 0 64056 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4766
timestamp 1624857261
transform 1 0 64056 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4765
timestamp 1624857261
transform 1 0 64600 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4764
timestamp 1624857261
transform 1 0 64600 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4763
timestamp 1624857261
transform 1 0 64600 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4762
timestamp 1624857261
transform 1 0 64600 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4761
timestamp 1624857261
transform 1 0 64736 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4760
timestamp 1624857261
transform 1 0 64736 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4759
timestamp 1624857261
transform 1 0 64736 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4758
timestamp 1624857261
transform 1 0 64736 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4757
timestamp 1624857261
transform 1 0 64872 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4756
timestamp 1624857261
transform 1 0 64872 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4755
timestamp 1624857261
transform 1 0 64872 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4754
timestamp 1624857261
transform 1 0 64872 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4753
timestamp 1624857261
transform 1 0 65688 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4752
timestamp 1624857261
transform 1 0 65688 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4751
timestamp 1624857261
transform 1 0 66640 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4750
timestamp 1624857261
transform 1 0 66640 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4749
timestamp 1624857261
transform 1 0 66640 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4748
timestamp 1624857261
transform 1 0 66640 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4747
timestamp 1624857261
transform 1 0 67184 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4746
timestamp 1624857261
transform 1 0 67184 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4745
timestamp 1624857261
transform 1 0 67320 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4744
timestamp 1624857261
transform 1 0 67320 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4743
timestamp 1624857261
transform 1 0 67864 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4742
timestamp 1624857261
transform 1 0 67864 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4741
timestamp 1624857261
transform 1 0 68408 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4740
timestamp 1624857261
transform 1 0 68408 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4739
timestamp 1624857261
transform 1 0 68408 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4738
timestamp 1624857261
transform 1 0 68408 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4737
timestamp 1624857261
transform 1 0 69088 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4736
timestamp 1624857261
transform 1 0 69088 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4735
timestamp 1624857261
transform 1 0 69088 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4734
timestamp 1624857261
transform 1 0 69088 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4733
timestamp 1624857261
transform 1 0 69224 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4732
timestamp 1624857261
transform 1 0 69224 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4731
timestamp 1624857261
transform 1 0 69632 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4730
timestamp 1624857261
transform 1 0 69632 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4729
timestamp 1624857261
transform 1 0 69632 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4728
timestamp 1624857261
transform 1 0 69632 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4727
timestamp 1624857261
transform 1 0 69768 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4726
timestamp 1624857261
transform 1 0 69768 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4725
timestamp 1624857261
transform 1 0 69768 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4724
timestamp 1624857261
transform 1 0 69768 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4723
timestamp 1624857261
transform 1 0 69768 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4722
timestamp 1624857261
transform 1 0 69768 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4721
timestamp 1624857261
transform 1 0 69768 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4720
timestamp 1624857261
transform 1 0 69768 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4719
timestamp 1624857261
transform 1 0 70312 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4718
timestamp 1624857261
transform 1 0 70312 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4717
timestamp 1624857261
transform 1 0 70312 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4716
timestamp 1624857261
transform 1 0 70312 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4715
timestamp 1624857261
transform 1 0 70312 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4714
timestamp 1624857261
transform 1 0 70312 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4713
timestamp 1624857261
transform 1 0 70856 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4712
timestamp 1624857261
transform 1 0 70856 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4711
timestamp 1624857261
transform 1 0 70856 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4710
timestamp 1624857261
transform 1 0 70856 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4709
timestamp 1624857261
transform 1 0 71672 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4708
timestamp 1624857261
transform 1 0 71672 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4707
timestamp 1624857261
transform 1 0 71944 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4706
timestamp 1624857261
transform 1 0 71944 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4705
timestamp 1624857261
transform 1 0 72896 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4704
timestamp 1624857261
transform 1 0 72896 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4703
timestamp 1624857261
transform 1 0 73440 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4702
timestamp 1624857261
transform 1 0 73440 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4701
timestamp 1624857261
transform 1 0 74120 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4700
timestamp 1624857261
transform 1 0 74120 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4699
timestamp 1624857261
transform 1 0 74664 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4698
timestamp 1624857261
transform 1 0 74664 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4697
timestamp 1624857261
transform 1 0 75208 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4696
timestamp 1624857261
transform 1 0 75208 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4695
timestamp 1624857261
transform 1 0 74664 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4694
timestamp 1624857261
transform 1 0 74664 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4693
timestamp 1624857261
transform 1 0 75208 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4692
timestamp 1624857261
transform 1 0 75208 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4691
timestamp 1624857261
transform 1 0 74528 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4690
timestamp 1624857261
transform 1 0 74528 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4689
timestamp 1624857261
transform 1 0 74800 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4688
timestamp 1624857261
transform 1 0 74800 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4687
timestamp 1624857261
transform 1 0 74664 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4686
timestamp 1624857261
transform 1 0 74664 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4685
timestamp 1624857261
transform 1 0 75344 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4684
timestamp 1624857261
transform 1 0 75344 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4683
timestamp 1624857261
transform 1 0 74664 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4682
timestamp 1624857261
transform 1 0 74664 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4681
timestamp 1624857261
transform 1 0 75344 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4680
timestamp 1624857261
transform 1 0 75344 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4679
timestamp 1624857261
transform 1 0 75888 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4678
timestamp 1624857261
transform 1 0 75888 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4677
timestamp 1624857261
transform 1 0 75888 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4676
timestamp 1624857261
transform 1 0 75888 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4675
timestamp 1624857261
transform 1 0 76568 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4674
timestamp 1624857261
transform 1 0 76568 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4673
timestamp 1624857261
transform 1 0 76568 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4672
timestamp 1624857261
transform 1 0 76568 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4671
timestamp 1624857261
transform 1 0 77112 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4670
timestamp 1624857261
transform 1 0 77112 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4669
timestamp 1624857261
transform 1 0 77792 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4668
timestamp 1624857261
transform 1 0 77792 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4667
timestamp 1624857261
transform 1 0 78336 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4666
timestamp 1624857261
transform 1 0 78336 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4665
timestamp 1624857261
transform 1 0 78336 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4664
timestamp 1624857261
transform 1 0 78336 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4663
timestamp 1624857261
transform 1 0 79288 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4662
timestamp 1624857261
transform 1 0 79288 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4661
timestamp 1624857261
transform 1 0 79560 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4660
timestamp 1624857261
transform 1 0 79560 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4659
timestamp 1624857261
transform 1 0 79560 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4658
timestamp 1624857261
transform 1 0 79560 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4657
timestamp 1624857261
transform 1 0 79696 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4656
timestamp 1624857261
transform 1 0 79696 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4655
timestamp 1624857261
transform 1 0 79832 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4654
timestamp 1624857261
transform 1 0 79832 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4653
timestamp 1624857261
transform 1 0 79696 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4652
timestamp 1624857261
transform 1 0 79696 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4651
timestamp 1624857261
transform 1 0 79696 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4650
timestamp 1624857261
transform 1 0 79696 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4649
timestamp 1624857261
transform 1 0 80512 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4648
timestamp 1624857261
transform 1 0 80512 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4647
timestamp 1624857261
transform 1 0 80920 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4646
timestamp 1624857261
transform 1 0 80920 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4645
timestamp 1624857261
transform 1 0 81464 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4644
timestamp 1624857261
transform 1 0 81464 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4643
timestamp 1624857261
transform 1 0 81600 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4642
timestamp 1624857261
transform 1 0 81600 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4641
timestamp 1624857261
transform 1 0 82008 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4640
timestamp 1624857261
transform 1 0 82008 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4639
timestamp 1624857261
transform 1 0 82008 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4638
timestamp 1624857261
transform 1 0 82008 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4637
timestamp 1624857261
transform 1 0 82824 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4636
timestamp 1624857261
transform 1 0 82824 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4635
timestamp 1624857261
transform 1 0 83368 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4634
timestamp 1624857261
transform 1 0 83368 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4633
timestamp 1624857261
transform 1 0 84048 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4632
timestamp 1624857261
transform 1 0 84048 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4631
timestamp 1624857261
transform 1 0 84184 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4630
timestamp 1624857261
transform 1 0 84184 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4629
timestamp 1624857261
transform 1 0 84184 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4628
timestamp 1624857261
transform 1 0 84184 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4627
timestamp 1624857261
transform 1 0 84592 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4626
timestamp 1624857261
transform 1 0 84592 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4625
timestamp 1624857261
transform 1 0 84592 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4624
timestamp 1624857261
transform 1 0 84592 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4623
timestamp 1624857261
transform 1 0 84592 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4622
timestamp 1624857261
transform 1 0 84592 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4621
timestamp 1624857261
transform 1 0 84728 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4620
timestamp 1624857261
transform 1 0 84728 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4619
timestamp 1624857261
transform 1 0 84728 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4618
timestamp 1624857261
transform 1 0 84728 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4617
timestamp 1624857261
transform 1 0 84728 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4616
timestamp 1624857261
transform 1 0 84728 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4615
timestamp 1624857261
transform 1 0 85680 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4614
timestamp 1624857261
transform 1 0 85680 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4613
timestamp 1624857261
transform 1 0 85272 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4612
timestamp 1624857261
transform 1 0 85272 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4611
timestamp 1624857261
transform 1 0 85816 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4610
timestamp 1624857261
transform 1 0 85816 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4609
timestamp 1624857261
transform 1 0 86496 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4608
timestamp 1624857261
transform 1 0 86496 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4607
timestamp 1624857261
transform 1 0 86496 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4606
timestamp 1624857261
transform 1 0 86496 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4605
timestamp 1624857261
transform 1 0 87040 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4604
timestamp 1624857261
transform 1 0 87040 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4603
timestamp 1624857261
transform 1 0 88400 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4602
timestamp 1624857261
transform 1 0 88400 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4601
timestamp 1624857261
transform 1 0 88400 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4600
timestamp 1624857261
transform 1 0 88400 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4599
timestamp 1624857261
transform 1 0 89080 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4598
timestamp 1624857261
transform 1 0 89080 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4597
timestamp 1624857261
transform 1 0 89216 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4596
timestamp 1624857261
transform 1 0 89216 0 1 126485
box 0 0 1 1
use contact_32  contact_32_4595
timestamp 1624857261
transform 1 0 89624 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4594
timestamp 1624857261
transform 1 0 89624 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4593
timestamp 1624857261
transform 1 0 89624 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4592
timestamp 1624857261
transform 1 0 89624 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4591
timestamp 1624857261
transform 1 0 89488 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4590
timestamp 1624857261
transform 1 0 89488 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4589
timestamp 1624857261
transform 1 0 89760 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4588
timestamp 1624857261
transform 1 0 89760 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4587
timestamp 1624857261
transform 1 0 89760 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4586
timestamp 1624857261
transform 1 0 89760 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4585
timestamp 1624857261
transform 1 0 89760 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4584
timestamp 1624857261
transform 1 0 89760 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4583
timestamp 1624857261
transform 1 0 89760 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4582
timestamp 1624857261
transform 1 0 89760 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4581
timestamp 1624857261
transform 1 0 90304 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4580
timestamp 1624857261
transform 1 0 90304 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4579
timestamp 1624857261
transform 1 0 90848 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4578
timestamp 1624857261
transform 1 0 90848 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4577
timestamp 1624857261
transform 1 0 91528 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4576
timestamp 1624857261
transform 1 0 91528 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4575
timestamp 1624857261
transform 1 0 92072 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4574
timestamp 1624857261
transform 1 0 92072 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4573
timestamp 1624857261
transform 1 0 92752 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4572
timestamp 1624857261
transform 1 0 92752 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4571
timestamp 1624857261
transform 1 0 93296 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4570
timestamp 1624857261
transform 1 0 93296 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4569
timestamp 1624857261
transform 1 0 94656 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4568
timestamp 1624857261
transform 1 0 94656 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4567
timestamp 1624857261
transform 1 0 94656 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4566
timestamp 1624857261
transform 1 0 94656 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4565
timestamp 1624857261
transform 1 0 94656 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4564
timestamp 1624857261
transform 1 0 94656 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4563
timestamp 1624857261
transform 1 0 94656 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4562
timestamp 1624857261
transform 1 0 94656 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4561
timestamp 1624857261
transform 1 0 94792 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4560
timestamp 1624857261
transform 1 0 94792 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4559
timestamp 1624857261
transform 1 0 94792 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4558
timestamp 1624857261
transform 1 0 94792 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4557
timestamp 1624857261
transform 1 0 95336 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4556
timestamp 1624857261
transform 1 0 95336 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4555
timestamp 1624857261
transform 1 0 94792 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4554
timestamp 1624857261
transform 1 0 94792 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4553
timestamp 1624857261
transform 1 0 95336 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4552
timestamp 1624857261
transform 1 0 95336 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4551
timestamp 1624857261
transform 1 0 95336 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4550
timestamp 1624857261
transform 1 0 95336 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4549
timestamp 1624857261
transform 1 0 95744 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4548
timestamp 1624857261
transform 1 0 95744 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4547
timestamp 1624857261
transform 1 0 95744 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4546
timestamp 1624857261
transform 1 0 95744 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4545
timestamp 1624857261
transform 1 0 96560 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4544
timestamp 1624857261
transform 1 0 96560 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4543
timestamp 1624857261
transform 1 0 97104 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4542
timestamp 1624857261
transform 1 0 97104 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4541
timestamp 1624857261
transform 1 0 97104 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4540
timestamp 1624857261
transform 1 0 97104 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4539
timestamp 1624857261
transform 1 0 97784 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4538
timestamp 1624857261
transform 1 0 97784 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4537
timestamp 1624857261
transform 1 0 97920 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4536
timestamp 1624857261
transform 1 0 97920 0 1 126485
box 0 0 1 1
use contact_32  contact_32_4535
timestamp 1624857261
transform 1 0 99552 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4534
timestamp 1624857261
transform 1 0 99552 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4533
timestamp 1624857261
transform 1 0 99552 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4532
timestamp 1624857261
transform 1 0 99552 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4531
timestamp 1624857261
transform 1 0 99552 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4530
timestamp 1624857261
transform 1 0 99552 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4529
timestamp 1624857261
transform 1 0 99552 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4528
timestamp 1624857261
transform 1 0 99552 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4527
timestamp 1624857261
transform 1 0 99552 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4526
timestamp 1624857261
transform 1 0 99552 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4525
timestamp 1624857261
transform 1 0 99688 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4524
timestamp 1624857261
transform 1 0 99688 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4523
timestamp 1624857261
transform 1 0 99688 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4522
timestamp 1624857261
transform 1 0 99688 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4521
timestamp 1624857261
transform 1 0 100232 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4520
timestamp 1624857261
transform 1 0 100232 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4519
timestamp 1624857261
transform 1 0 100504 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4518
timestamp 1624857261
transform 1 0 100504 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4517
timestamp 1624857261
transform 1 0 100776 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4516
timestamp 1624857261
transform 1 0 100776 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4515
timestamp 1624857261
transform 1 0 101592 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4514
timestamp 1624857261
transform 1 0 101592 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4513
timestamp 1624857261
transform 1 0 102000 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4512
timestamp 1624857261
transform 1 0 102000 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4511
timestamp 1624857261
transform 1 0 102136 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4510
timestamp 1624857261
transform 1 0 102136 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4509
timestamp 1624857261
transform 1 0 103360 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4508
timestamp 1624857261
transform 1 0 103360 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4507
timestamp 1624857261
transform 1 0 103360 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4506
timestamp 1624857261
transform 1 0 103360 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4505
timestamp 1624857261
transform 1 0 104040 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4504
timestamp 1624857261
transform 1 0 104040 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4503
timestamp 1624857261
transform 1 0 104040 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4502
timestamp 1624857261
transform 1 0 104040 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4501
timestamp 1624857261
transform 1 0 104312 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4500
timestamp 1624857261
transform 1 0 104312 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4499
timestamp 1624857261
transform 1 0 104584 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4498
timestamp 1624857261
transform 1 0 104584 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4497
timestamp 1624857261
transform 1 0 104584 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4496
timestamp 1624857261
transform 1 0 104584 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4495
timestamp 1624857261
transform 1 0 104584 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4494
timestamp 1624857261
transform 1 0 104584 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4493
timestamp 1624857261
transform 1 0 104720 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4492
timestamp 1624857261
transform 1 0 104720 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4491
timestamp 1624857261
transform 1 0 104584 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4490
timestamp 1624857261
transform 1 0 104584 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4489
timestamp 1624857261
transform 1 0 105264 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4488
timestamp 1624857261
transform 1 0 105264 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4487
timestamp 1624857261
transform 1 0 104584 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4486
timestamp 1624857261
transform 1 0 104584 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4485
timestamp 1624857261
transform 1 0 105264 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4484
timestamp 1624857261
transform 1 0 105264 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4483
timestamp 1624857261
transform 1 0 105264 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4482
timestamp 1624857261
transform 1 0 105264 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4481
timestamp 1624857261
transform 1 0 105808 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4480
timestamp 1624857261
transform 1 0 105808 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4479
timestamp 1624857261
transform 1 0 106488 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4478
timestamp 1624857261
transform 1 0 106488 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4477
timestamp 1624857261
transform 1 0 108120 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4476
timestamp 1624857261
transform 1 0 108120 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4475
timestamp 1624857261
transform 1 0 109208 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4474
timestamp 1624857261
transform 1 0 109208 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4473
timestamp 1624857261
transform 1 0 109616 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4472
timestamp 1624857261
transform 1 0 109616 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4471
timestamp 1624857261
transform 1 0 109616 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4470
timestamp 1624857261
transform 1 0 109616 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4469
timestamp 1624857261
transform 1 0 109616 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4468
timestamp 1624857261
transform 1 0 109616 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4467
timestamp 1624857261
transform 1 0 109752 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4466
timestamp 1624857261
transform 1 0 109752 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4465
timestamp 1624857261
transform 1 0 109752 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4464
timestamp 1624857261
transform 1 0 109752 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4463
timestamp 1624857261
transform 1 0 109752 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4462
timestamp 1624857261
transform 1 0 109752 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4461
timestamp 1624857261
transform 1 0 110296 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4460
timestamp 1624857261
transform 1 0 110296 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4459
timestamp 1624857261
transform 1 0 110296 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4458
timestamp 1624857261
transform 1 0 110296 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4457
timestamp 1624857261
transform 1 0 110296 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4456
timestamp 1624857261
transform 1 0 110296 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4455
timestamp 1624857261
transform 1 0 110840 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4454
timestamp 1624857261
transform 1 0 110840 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4453
timestamp 1624857261
transform 1 0 110840 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4452
timestamp 1624857261
transform 1 0 110840 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4451
timestamp 1624857261
transform 1 0 111520 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4450
timestamp 1624857261
transform 1 0 111520 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4449
timestamp 1624857261
transform 1 0 111520 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4448
timestamp 1624857261
transform 1 0 111520 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4447
timestamp 1624857261
transform 1 0 112064 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4446
timestamp 1624857261
transform 1 0 112064 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4445
timestamp 1624857261
transform 1 0 112744 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4444
timestamp 1624857261
transform 1 0 112744 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4443
timestamp 1624857261
transform 1 0 112744 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4442
timestamp 1624857261
transform 1 0 112744 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4441
timestamp 1624857261
transform 1 0 113288 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4440
timestamp 1624857261
transform 1 0 113288 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4439
timestamp 1624857261
transform 1 0 113288 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4438
timestamp 1624857261
transform 1 0 113288 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4437
timestamp 1624857261
transform 1 0 114240 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4436
timestamp 1624857261
transform 1 0 114240 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4435
timestamp 1624857261
transform 1 0 114240 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4434
timestamp 1624857261
transform 1 0 114240 0 1 24349
box 0 0 1 1
use contact_32  contact_32_4433
timestamp 1624857261
transform 1 0 114512 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4432
timestamp 1624857261
transform 1 0 114512 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4431
timestamp 1624857261
transform 1 0 114512 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4430
timestamp 1624857261
transform 1 0 114512 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4429
timestamp 1624857261
transform 1 0 114512 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4428
timestamp 1624857261
transform 1 0 114512 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4427
timestamp 1624857261
transform 1 0 114784 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4426
timestamp 1624857261
transform 1 0 114784 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4425
timestamp 1624857261
transform 1 0 114784 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4424
timestamp 1624857261
transform 1 0 114784 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4423
timestamp 1624857261
transform 1 0 114784 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4422
timestamp 1624857261
transform 1 0 114784 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4421
timestamp 1624857261
transform 1 0 115328 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4420
timestamp 1624857261
transform 1 0 115328 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4419
timestamp 1624857261
transform 1 0 115736 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4418
timestamp 1624857261
transform 1 0 115736 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4417
timestamp 1624857261
transform 1 0 116552 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4416
timestamp 1624857261
transform 1 0 116552 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4415
timestamp 1624857261
transform 1 0 117096 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4414
timestamp 1624857261
transform 1 0 117096 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4413
timestamp 1624857261
transform 1 0 117640 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4412
timestamp 1624857261
transform 1 0 117640 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4411
timestamp 1624857261
transform 1 0 117640 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4410
timestamp 1624857261
transform 1 0 117640 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4409
timestamp 1624857261
transform 1 0 117776 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4408
timestamp 1624857261
transform 1 0 117776 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4407
timestamp 1624857261
transform 1 0 118320 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4406
timestamp 1624857261
transform 1 0 118320 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4405
timestamp 1624857261
transform 1 0 119000 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4404
timestamp 1624857261
transform 1 0 119000 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4403
timestamp 1624857261
transform 1 0 119000 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4402
timestamp 1624857261
transform 1 0 119000 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4401
timestamp 1624857261
transform 1 0 119272 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4400
timestamp 1624857261
transform 1 0 119272 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4399
timestamp 1624857261
transform 1 0 119544 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4398
timestamp 1624857261
transform 1 0 119544 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4397
timestamp 1624857261
transform 1 0 119680 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4396
timestamp 1624857261
transform 1 0 119680 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4395
timestamp 1624857261
transform 1 0 119680 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4394
timestamp 1624857261
transform 1 0 119680 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4393
timestamp 1624857261
transform 1 0 119544 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4392
timestamp 1624857261
transform 1 0 119544 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4391
timestamp 1624857261
transform 1 0 120224 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4390
timestamp 1624857261
transform 1 0 120224 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4389
timestamp 1624857261
transform 1 0 119544 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4388
timestamp 1624857261
transform 1 0 119544 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4387
timestamp 1624857261
transform 1 0 120224 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4386
timestamp 1624857261
transform 1 0 120224 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4385
timestamp 1624857261
transform 1 0 120768 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4384
timestamp 1624857261
transform 1 0 120768 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4383
timestamp 1624857261
transform 1 0 121448 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4382
timestamp 1624857261
transform 1 0 121448 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4381
timestamp 1624857261
transform 1 0 121992 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4380
timestamp 1624857261
transform 1 0 121992 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4379
timestamp 1624857261
transform 1 0 121992 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4378
timestamp 1624857261
transform 1 0 121992 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4377
timestamp 1624857261
transform 1 0 122944 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4376
timestamp 1624857261
transform 1 0 122944 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4375
timestamp 1624857261
transform 1 0 122944 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4374
timestamp 1624857261
transform 1 0 122944 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4373
timestamp 1624857261
transform 1 0 123896 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4372
timestamp 1624857261
transform 1 0 123896 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4371
timestamp 1624857261
transform 1 0 123896 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4370
timestamp 1624857261
transform 1 0 123896 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4369
timestamp 1624857261
transform 1 0 124304 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4368
timestamp 1624857261
transform 1 0 124440 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4367
timestamp 1624857261
transform 1 0 124440 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4366
timestamp 1624857261
transform 1 0 124440 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4365
timestamp 1624857261
transform 1 0 124576 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4364
timestamp 1624857261
transform 1 0 124576 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4363
timestamp 1624857261
transform 1 0 124576 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4362
timestamp 1624857261
transform 1 0 124576 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4361
timestamp 1624857261
transform 1 0 124576 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4360
timestamp 1624857261
transform 1 0 124576 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4359
timestamp 1624857261
transform 1 0 124712 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4358
timestamp 1624857261
transform 1 0 124712 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4357
timestamp 1624857261
transform 1 0 124576 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4356
timestamp 1624857261
transform 1 0 124576 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4355
timestamp 1624857261
transform 1 0 124576 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4354
timestamp 1624857261
transform 1 0 124576 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4353
timestamp 1624857261
transform 1 0 125256 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4352
timestamp 1624857261
transform 1 0 125256 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4351
timestamp 1624857261
transform 1 0 125800 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4350
timestamp 1624857261
transform 1 0 125800 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4349
timestamp 1624857261
transform 1 0 125800 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4348
timestamp 1624857261
transform 1 0 125800 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4347
timestamp 1624857261
transform 1 0 126480 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4346
timestamp 1624857261
transform 1 0 126480 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4345
timestamp 1624857261
transform 1 0 127024 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4344
timestamp 1624857261
transform 1 0 127024 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4343
timestamp 1624857261
transform 1 0 127024 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4342
timestamp 1624857261
transform 1 0 127024 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4341
timestamp 1624857261
transform 1 0 128248 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4340
timestamp 1624857261
transform 1 0 128248 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4339
timestamp 1624857261
transform 1 0 128928 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4338
timestamp 1624857261
transform 1 0 128928 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4337
timestamp 1624857261
transform 1 0 128928 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4336
timestamp 1624857261
transform 1 0 128928 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4335
timestamp 1624857261
transform 1 0 129200 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4334
timestamp 1624857261
transform 1 0 129200 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4333
timestamp 1624857261
transform 1 0 129472 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4332
timestamp 1624857261
transform 1 0 129472 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4331
timestamp 1624857261
transform 1 0 129608 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4330
timestamp 1624857261
transform 1 0 129608 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4329
timestamp 1624857261
transform 1 0 129744 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4328
timestamp 1624857261
transform 1 0 129744 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4327
timestamp 1624857261
transform 1 0 129608 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4326
timestamp 1624857261
transform 1 0 129608 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4325
timestamp 1624857261
transform 1 0 130288 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4324
timestamp 1624857261
transform 1 0 130288 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4323
timestamp 1624857261
transform 1 0 129608 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4322
timestamp 1624857261
transform 1 0 129608 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4321
timestamp 1624857261
transform 1 0 130288 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4320
timestamp 1624857261
transform 1 0 130288 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4319
timestamp 1624857261
transform 1 0 130288 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4318
timestamp 1624857261
transform 1 0 130288 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4317
timestamp 1624857261
transform 1 0 130832 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4316
timestamp 1624857261
transform 1 0 130832 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4315
timestamp 1624857261
transform 1 0 131648 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4314
timestamp 1624857261
transform 1 0 131648 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4313
timestamp 1624857261
transform 1 0 132056 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4312
timestamp 1624857261
transform 1 0 132056 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4311
timestamp 1624857261
transform 1 0 133280 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4310
timestamp 1624857261
transform 1 0 133280 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4309
timestamp 1624857261
transform 1 0 133280 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4308
timestamp 1624857261
transform 1 0 133280 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4307
timestamp 1624857261
transform 1 0 133960 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4306
timestamp 1624857261
transform 1 0 133960 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4305
timestamp 1624857261
transform 1 0 134096 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4304
timestamp 1624857261
transform 1 0 134096 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4303
timestamp 1624857261
transform 1 0 134504 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4302
timestamp 1624857261
transform 1 0 134504 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4301
timestamp 1624857261
transform 1 0 134504 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4300
timestamp 1624857261
transform 1 0 134504 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4299
timestamp 1624857261
transform 1 0 134640 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4298
timestamp 1624857261
transform 1 0 134640 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4297
timestamp 1624857261
transform 1 0 134640 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4296
timestamp 1624857261
transform 1 0 134640 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4295
timestamp 1624857261
transform 1 0 134504 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4294
timestamp 1624857261
transform 1 0 134504 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4293
timestamp 1624857261
transform 1 0 134640 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4292
timestamp 1624857261
transform 1 0 134640 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4291
timestamp 1624857261
transform 1 0 135592 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4290
timestamp 1624857261
transform 1 0 135592 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4289
timestamp 1624857261
transform 1 0 135184 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4288
timestamp 1624857261
transform 1 0 135184 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4287
timestamp 1624857261
transform 1 0 135184 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4286
timestamp 1624857261
transform 1 0 135184 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4285
timestamp 1624857261
transform 1 0 135456 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4284
timestamp 1624857261
transform 1 0 135456 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4283
timestamp 1624857261
transform 1 0 135728 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4282
timestamp 1624857261
transform 1 0 135728 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4281
timestamp 1624857261
transform 1 0 136680 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4280
timestamp 1624857261
transform 1 0 136680 0 1 24349
box 0 0 1 1
use contact_32  contact_32_4279
timestamp 1624857261
transform 1 0 137088 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4278
timestamp 1624857261
transform 1 0 137088 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4277
timestamp 1624857261
transform 1 0 138176 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4276
timestamp 1624857261
transform 1 0 138176 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4275
timestamp 1624857261
transform 1 0 138176 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4274
timestamp 1624857261
transform 1 0 138176 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4273
timestamp 1624857261
transform 1 0 139128 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4272
timestamp 1624857261
transform 1 0 139128 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4271
timestamp 1624857261
transform 1 0 139536 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4270
timestamp 1624857261
transform 1 0 139536 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4269
timestamp 1624857261
transform 1 0 139536 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4268
timestamp 1624857261
transform 1 0 139536 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4267
timestamp 1624857261
transform 1 0 139536 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4266
timestamp 1624857261
transform 1 0 139536 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4265
timestamp 1624857261
transform 1 0 139536 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4264
timestamp 1624857261
transform 1 0 139536 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4263
timestamp 1624857261
transform 1 0 139672 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4262
timestamp 1624857261
transform 1 0 139672 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4261
timestamp 1624857261
transform 1 0 139536 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4260
timestamp 1624857261
transform 1 0 139536 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4259
timestamp 1624857261
transform 1 0 139536 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4258
timestamp 1624857261
transform 1 0 139536 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4257
timestamp 1624857261
transform 1 0 140216 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4256
timestamp 1624857261
transform 1 0 140216 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4255
timestamp 1624857261
transform 1 0 140352 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4254
timestamp 1624857261
transform 1 0 140352 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4253
timestamp 1624857261
transform 1 0 141440 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4252
timestamp 1624857261
transform 1 0 141440 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4251
timestamp 1624857261
transform 1 0 141848 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4250
timestamp 1624857261
transform 1 0 141848 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4249
timestamp 1624857261
transform 1 0 141984 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4248
timestamp 1624857261
transform 1 0 141984 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4247
timestamp 1624857261
transform 1 0 142664 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4246
timestamp 1624857261
transform 1 0 142664 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4245
timestamp 1624857261
transform 1 0 143208 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4244
timestamp 1624857261
transform 1 0 143208 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4243
timestamp 1624857261
transform 1 0 144024 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4242
timestamp 1624857261
transform 1 0 144024 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4241
timestamp 1624857261
transform 1 0 144432 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4240
timestamp 1624857261
transform 1 0 144432 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4239
timestamp 1624857261
transform 1 0 144568 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4238
timestamp 1624857261
transform 1 0 144568 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4237
timestamp 1624857261
transform 1 0 144704 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4236
timestamp 1624857261
transform 1 0 144704 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4235
timestamp 1624857261
transform 1 0 144568 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4234
timestamp 1624857261
transform 1 0 144568 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4233
timestamp 1624857261
transform 1 0 145656 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4232
timestamp 1624857261
transform 1 0 145656 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4231
timestamp 1624857261
transform 1 0 144568 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4230
timestamp 1624857261
transform 1 0 144568 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4229
timestamp 1624857261
transform 1 0 145248 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4228
timestamp 1624857261
transform 1 0 145248 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4227
timestamp 1624857261
transform 1 0 145248 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4226
timestamp 1624857261
transform 1 0 145248 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4225
timestamp 1624857261
transform 1 0 145384 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4224
timestamp 1624857261
transform 1 0 145384 0 1 24349
box 0 0 1 1
use contact_32  contact_32_4223
timestamp 1624857261
transform 1 0 146472 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4222
timestamp 1624857261
transform 1 0 146472 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4221
timestamp 1624857261
transform 1 0 146472 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4220
timestamp 1624857261
transform 1 0 146472 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4219
timestamp 1624857261
transform 1 0 147016 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4218
timestamp 1624857261
transform 1 0 147016 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4217
timestamp 1624857261
transform 1 0 147016 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4216
timestamp 1624857261
transform 1 0 147016 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4215
timestamp 1624857261
transform 1 0 147696 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4214
timestamp 1624857261
transform 1 0 147696 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4213
timestamp 1624857261
transform 1 0 147696 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4212
timestamp 1624857261
transform 1 0 147696 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4211
timestamp 1624857261
transform 1 0 148240 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4210
timestamp 1624857261
transform 1 0 148240 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4209
timestamp 1624857261
transform 1 0 149056 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4208
timestamp 1624857261
transform 1 0 149056 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4207
timestamp 1624857261
transform 1 0 149464 0 1 126893
box 0 0 1 1
use contact_32  contact_32_4206
timestamp 1624857261
transform 1 0 149464 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4205
timestamp 1624857261
transform 1 0 149464 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4204
timestamp 1624857261
transform 1 0 149464 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4203
timestamp 1624857261
transform 1 0 149464 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4202
timestamp 1624857261
transform 1 0 149464 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4201
timestamp 1624857261
transform 1 0 149600 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4200
timestamp 1624857261
transform 1 0 149600 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4199
timestamp 1624857261
transform 1 0 149736 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4198
timestamp 1624857261
transform 1 0 149736 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4197
timestamp 1624857261
transform 1 0 149600 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4196
timestamp 1624857261
transform 1 0 149600 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4195
timestamp 1624857261
transform 1 0 149600 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4194
timestamp 1624857261
transform 1 0 149600 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4193
timestamp 1624857261
transform 1 0 150144 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4192
timestamp 1624857261
transform 1 0 150144 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4191
timestamp 1624857261
transform 1 0 150416 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4190
timestamp 1624857261
transform 1 0 150416 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4189
timestamp 1624857261
transform 1 0 151504 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4188
timestamp 1624857261
transform 1 0 151504 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4187
timestamp 1624857261
transform 1 0 152048 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4186
timestamp 1624857261
transform 1 0 152048 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4185
timestamp 1624857261
transform 1 0 151912 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4184
timestamp 1624857261
transform 1 0 151912 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4183
timestamp 1624857261
transform 1 0 152728 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4182
timestamp 1624857261
transform 1 0 152728 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4181
timestamp 1624857261
transform 1 0 153272 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4180
timestamp 1624857261
transform 1 0 153272 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4179
timestamp 1624857261
transform 1 0 153272 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4178
timestamp 1624857261
transform 1 0 153272 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4177
timestamp 1624857261
transform 1 0 153952 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4176
timestamp 1624857261
transform 1 0 153952 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4175
timestamp 1624857261
transform 1 0 154088 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4174
timestamp 1624857261
transform 1 0 154088 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4173
timestamp 1624857261
transform 1 0 154496 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4172
timestamp 1624857261
transform 1 0 154496 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4171
timestamp 1624857261
transform 1 0 154496 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4170
timestamp 1624857261
transform 1 0 154496 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4169
timestamp 1624857261
transform 1 0 154496 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4168
timestamp 1624857261
transform 1 0 154496 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4167
timestamp 1624857261
transform 1 0 154632 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4166
timestamp 1624857261
transform 1 0 154632 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4165
timestamp 1624857261
transform 1 0 154632 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4164
timestamp 1624857261
transform 1 0 154632 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4163
timestamp 1624857261
transform 1 0 154632 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4162
timestamp 1624857261
transform 1 0 154632 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4161
timestamp 1624857261
transform 1 0 155176 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4160
timestamp 1624857261
transform 1 0 155176 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4159
timestamp 1624857261
transform 1 0 155176 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4158
timestamp 1624857261
transform 1 0 155176 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4157
timestamp 1624857261
transform 1 0 155176 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4156
timestamp 1624857261
transform 1 0 155176 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4155
timestamp 1624857261
transform 1 0 155720 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4154
timestamp 1624857261
transform 1 0 155720 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4153
timestamp 1624857261
transform 1 0 155720 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4152
timestamp 1624857261
transform 1 0 155720 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4151
timestamp 1624857261
transform 1 0 156672 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4150
timestamp 1624857261
transform 1 0 156672 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4149
timestamp 1624857261
transform 1 0 156944 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4148
timestamp 1624857261
transform 1 0 156944 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4147
timestamp 1624857261
transform 1 0 157896 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4146
timestamp 1624857261
transform 1 0 157896 0 1 126485
box 0 0 1 1
use contact_32  contact_32_4145
timestamp 1624857261
transform 1 0 158168 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4144
timestamp 1624857261
transform 1 0 158168 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4143
timestamp 1624857261
transform 1 0 158984 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4142
timestamp 1624857261
transform 1 0 158984 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4141
timestamp 1624857261
transform 1 0 159528 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4140
timestamp 1624857261
transform 1 0 159528 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4139
timestamp 1624857261
transform 1 0 159392 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4138
timestamp 1624857261
transform 1 0 159392 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4137
timestamp 1624857261
transform 1 0 159664 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4136
timestamp 1624857261
transform 1 0 159664 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4135
timestamp 1624857261
transform 1 0 159664 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4134
timestamp 1624857261
transform 1 0 159664 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4133
timestamp 1624857261
transform 1 0 160208 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4132
timestamp 1624857261
transform 1 0 160208 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4131
timestamp 1624857261
transform 1 0 159528 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4130
timestamp 1624857261
transform 1 0 159528 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4129
timestamp 1624857261
transform 1 0 160208 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4128
timestamp 1624857261
transform 1 0 160208 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4127
timestamp 1624857261
transform 1 0 160208 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4126
timestamp 1624857261
transform 1 0 160208 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4125
timestamp 1624857261
transform 1 0 160208 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4124
timestamp 1624857261
transform 1 0 160208 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4123
timestamp 1624857261
transform 1 0 160752 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4122
timestamp 1624857261
transform 1 0 160752 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4121
timestamp 1624857261
transform 1 0 160752 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4120
timestamp 1624857261
transform 1 0 160752 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4119
timestamp 1624857261
transform 1 0 161432 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4118
timestamp 1624857261
transform 1 0 161432 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4117
timestamp 1624857261
transform 1 0 161976 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4116
timestamp 1624857261
transform 1 0 161976 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4115
timestamp 1624857261
transform 1 0 163200 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4114
timestamp 1624857261
transform 1 0 163200 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4113
timestamp 1624857261
transform 1 0 163200 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4112
timestamp 1624857261
transform 1 0 163200 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4111
timestamp 1624857261
transform 1 0 163880 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4110
timestamp 1624857261
transform 1 0 163880 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4109
timestamp 1624857261
transform 1 0 164152 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4108
timestamp 1624857261
transform 1 0 164152 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4107
timestamp 1624857261
transform 1 0 164424 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4106
timestamp 1624857261
transform 1 0 164424 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4105
timestamp 1624857261
transform 1 0 164424 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4104
timestamp 1624857261
transform 1 0 164424 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4103
timestamp 1624857261
transform 1 0 164560 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4102
timestamp 1624857261
transform 1 0 164560 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4101
timestamp 1624857261
transform 1 0 164560 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4100
timestamp 1624857261
transform 1 0 164560 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4099
timestamp 1624857261
transform 1 0 164560 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4098
timestamp 1624857261
transform 1 0 164560 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4097
timestamp 1624857261
transform 1 0 164560 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4096
timestamp 1624857261
transform 1 0 164560 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4095
timestamp 1624857261
transform 1 0 165512 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4094
timestamp 1624857261
transform 1 0 165512 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4093
timestamp 1624857261
transform 1 0 165376 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4092
timestamp 1624857261
transform 1 0 165376 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4091
timestamp 1624857261
transform 1 0 165376 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4090
timestamp 1624857261
transform 1 0 165376 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4089
timestamp 1624857261
transform 1 0 166328 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4088
timestamp 1624857261
transform 1 0 166328 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4087
timestamp 1624857261
transform 1 0 166464 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4086
timestamp 1624857261
transform 1 0 166464 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4085
timestamp 1624857261
transform 1 0 166872 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4084
timestamp 1624857261
transform 1 0 166872 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4083
timestamp 1624857261
transform 1 0 168232 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4082
timestamp 1624857261
transform 1 0 168232 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4081
timestamp 1624857261
transform 1 0 168232 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4080
timestamp 1624857261
transform 1 0 168232 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4079
timestamp 1624857261
transform 1 0 168912 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4078
timestamp 1624857261
transform 1 0 168912 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4077
timestamp 1624857261
transform 1 0 169456 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4076
timestamp 1624857261
transform 1 0 169456 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4075
timestamp 1624857261
transform 1 0 169456 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4074
timestamp 1624857261
transform 1 0 169456 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4073
timestamp 1624857261
transform 1 0 169592 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4072
timestamp 1624857261
transform 1 0 169592 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4071
timestamp 1624857261
transform 1 0 169592 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4070
timestamp 1624857261
transform 1 0 169592 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4069
timestamp 1624857261
transform 1 0 169592 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4068
timestamp 1624857261
transform 1 0 169592 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4067
timestamp 1624857261
transform 1 0 170136 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4066
timestamp 1624857261
transform 1 0 170136 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4065
timestamp 1624857261
transform 1 0 169592 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4064
timestamp 1624857261
transform 1 0 169592 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4063
timestamp 1624857261
transform 1 0 170136 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4062
timestamp 1624857261
transform 1 0 170136 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4061
timestamp 1624857261
transform 1 0 170544 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4060
timestamp 1624857261
transform 1 0 170544 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4059
timestamp 1624857261
transform 1 0 170680 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4058
timestamp 1624857261
transform 1 0 170680 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4057
timestamp 1624857261
transform 1 0 171360 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4056
timestamp 1624857261
transform 1 0 171360 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4055
timestamp 1624857261
transform 1 0 171360 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4054
timestamp 1624857261
transform 1 0 171360 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4053
timestamp 1624857261
transform 1 0 171904 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4052
timestamp 1624857261
transform 1 0 171904 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4051
timestamp 1624857261
transform 1 0 171904 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4050
timestamp 1624857261
transform 1 0 171904 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4049
timestamp 1624857261
transform 1 0 173128 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4048
timestamp 1624857261
transform 1 0 173128 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4047
timestamp 1624857261
transform 1 0 173264 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4046
timestamp 1624857261
transform 1 0 173264 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4045
timestamp 1624857261
transform 1 0 174488 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4044
timestamp 1624857261
transform 1 0 174488 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4043
timestamp 1624857261
transform 1 0 174488 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4042
timestamp 1624857261
transform 1 0 174488 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4041
timestamp 1624857261
transform 1 0 174488 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4040
timestamp 1624857261
transform 1 0 174488 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4039
timestamp 1624857261
transform 1 0 174488 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4038
timestamp 1624857261
transform 1 0 174488 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4037
timestamp 1624857261
transform 1 0 174624 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4036
timestamp 1624857261
transform 1 0 174624 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4035
timestamp 1624857261
transform 1 0 174624 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4034
timestamp 1624857261
transform 1 0 174624 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4033
timestamp 1624857261
transform 1 0 174624 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4032
timestamp 1624857261
transform 1 0 174624 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4031
timestamp 1624857261
transform 1 0 175168 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4030
timestamp 1624857261
transform 1 0 175168 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4029
timestamp 1624857261
transform 1 0 175168 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4028
timestamp 1624857261
transform 1 0 175168 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4027
timestamp 1624857261
transform 1 0 175712 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4026
timestamp 1624857261
transform 1 0 175712 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4025
timestamp 1624857261
transform 1 0 176936 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4024
timestamp 1624857261
transform 1 0 176936 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4023
timestamp 1624857261
transform 1 0 176936 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4022
timestamp 1624857261
transform 1 0 176936 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4021
timestamp 1624857261
transform 1 0 178160 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4020
timestamp 1624857261
transform 1 0 178160 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4019
timestamp 1624857261
transform 1 0 178160 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4018
timestamp 1624857261
transform 1 0 178160 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4017
timestamp 1624857261
transform 1 0 178976 0 1 126621
box 0 0 1 1
use contact_32  contact_32_4016
timestamp 1624857261
transform 1 0 178976 0 1 127029
box 0 0 1 1
use contact_32  contact_32_4015
timestamp 1624857261
transform 1 0 179112 0 1 23669
box 0 0 1 1
use contact_32  contact_32_4014
timestamp 1624857261
transform 1 0 179112 0 1 24349
box 0 0 1 1
use contact_32  contact_32_4013
timestamp 1624857261
transform 1 0 179520 0 1 127165
box 0 0 1 1
use contact_32  contact_32_4012
timestamp 1624857261
transform 1 0 179520 0 1 131789
box 0 0 1 1
use contact_32  contact_32_4011
timestamp 1624857261
transform 1 0 179520 0 1 16325
box 0 0 1 1
use contact_32  contact_32_4010
timestamp 1624857261
transform 1 0 179520 0 1 15509
box 0 0 1 1
use contact_32  contact_32_4009
timestamp 1624857261
transform 1 0 179656 0 1 16461
box 0 0 1 1
use contact_32  contact_32_4008
timestamp 1624857261
transform 1 0 179656 0 1 17957
box 0 0 1 1
use contact_32  contact_32_4007
timestamp 1624857261
transform 1 0 179656 0 1 131925
box 0 0 1 1
use contact_32  contact_32_4006
timestamp 1624857261
transform 1 0 179656 0 1 132605
box 0 0 1 1
use contact_32  contact_32_4005
timestamp 1624857261
transform 1 0 179656 0 1 18773
box 0 0 1 1
use contact_32  contact_32_4004
timestamp 1624857261
transform 1 0 179656 0 1 18093
box 0 0 1 1
use contact_32  contact_32_4003
timestamp 1624857261
transform 1 0 180200 0 1 18909
box 0 0 1 1
use contact_32  contact_32_4002
timestamp 1624857261
transform 1 0 180200 0 1 23533
box 0 0 1 1
use contact_32  contact_32_4001
timestamp 1624857261
transform 1 0 180200 0 1 24213
box 0 0 1 1
use contact_32  contact_32_4000
timestamp 1624857261
transform 1 0 180200 0 1 23669
box 0 0 1 1
use contact_32  contact_32_3999
timestamp 1624857261
transform 1 0 180200 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3998
timestamp 1624857261
transform 1 0 180200 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3997
timestamp 1624857261
transform 1 0 180608 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3996
timestamp 1624857261
transform 1 0 180608 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3995
timestamp 1624857261
transform 1 0 181424 0 1 24213
box 0 0 1 1
use contact_32  contact_32_3994
timestamp 1624857261
transform 1 0 181424 0 1 23669
box 0 0 1 1
use contact_32  contact_32_3993
timestamp 1624857261
transform 1 0 181424 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3992
timestamp 1624857261
transform 1 0 181424 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3991
timestamp 1624857261
transform 1 0 181968 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3990
timestamp 1624857261
transform 1 0 181968 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3989
timestamp 1624857261
transform 1 0 183192 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3988
timestamp 1624857261
transform 1 0 183192 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3987
timestamp 1624857261
transform 1 0 183192 0 1 23669
box 0 0 1 1
use contact_32  contact_32_3986
timestamp 1624857261
transform 1 0 183192 0 1 24213
box 0 0 1 1
use contact_32  contact_32_3985
timestamp 1624857261
transform 1 0 184008 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3984
timestamp 1624857261
transform 1 0 184008 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3983
timestamp 1624857261
transform 1 0 184280 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3982
timestamp 1624857261
transform 1 0 184280 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3981
timestamp 1624857261
transform 1 0 184416 0 1 127165
box 0 0 1 1
use contact_32  contact_32_3980
timestamp 1624857261
transform 1 0 184416 0 1 131789
box 0 0 1 1
use contact_32  contact_32_3979
timestamp 1624857261
transform 1 0 184416 0 1 23533
box 0 0 1 1
use contact_32  contact_32_3978
timestamp 1624857261
transform 1 0 184416 0 1 18909
box 0 0 1 1
use contact_32  contact_32_3977
timestamp 1624857261
transform 1 0 184416 0 1 16325
box 0 0 1 1
use contact_32  contact_32_3976
timestamp 1624857261
transform 1 0 184416 0 1 15509
box 0 0 1 1
use contact_32  contact_32_3975
timestamp 1624857261
transform 1 0 184416 0 1 16461
box 0 0 1 1
use contact_32  contact_32_3974
timestamp 1624857261
transform 1 0 184416 0 1 17957
box 0 0 1 1
use contact_32  contact_32_3973
timestamp 1624857261
transform 1 0 189040 0 1 15509
box 0 0 1 1
use contact_32  contact_32_3972
timestamp 1624857261
transform 1 0 189040 0 1 15101
box 0 0 1 1
use contact_32  contact_32_3971
timestamp 1624857261
transform 1 0 184960 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3970
timestamp 1624857261
transform 1 0 184960 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3969
timestamp 1624857261
transform 1 0 184416 0 1 18773
box 0 0 1 1
use contact_32  contact_32_3968
timestamp 1624857261
transform 1 0 184416 0 1 18093
box 0 0 1 1
use contact_32  contact_32_3967
timestamp 1624857261
transform 1 0 184416 0 1 131925
box 0 0 1 1
use contact_32  contact_32_3966
timestamp 1624857261
transform 1 0 184416 0 1 132605
box 0 0 1 1
use contact_32  contact_32_3965
timestamp 1624857261
transform 1 0 185232 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3964
timestamp 1624857261
transform 1 0 185232 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3963
timestamp 1624857261
transform 1 0 185368 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3962
timestamp 1624857261
transform 1 0 185368 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3961
timestamp 1624857261
transform 1 0 185640 0 1 23669
box 0 0 1 1
use contact_32  contact_32_3960
timestamp 1624857261
transform 1 0 185640 0 1 24213
box 0 0 1 1
use contact_32  contact_32_3959
timestamp 1624857261
transform 1 0 186456 0 1 24213
box 0 0 1 1
use contact_32  contact_32_3958
timestamp 1624857261
transform 1 0 186456 0 1 23669
box 0 0 1 1
use contact_32  contact_32_3957
timestamp 1624857261
transform 1 0 187000 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3956
timestamp 1624857261
transform 1 0 187000 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3955
timestamp 1624857261
transform 1 0 187680 0 1 24213
box 0 0 1 1
use contact_32  contact_32_3954
timestamp 1624857261
transform 1 0 187680 0 1 23669
box 0 0 1 1
use contact_32  contact_32_3953
timestamp 1624857261
transform 1 0 188224 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3952
timestamp 1624857261
transform 1 0 188224 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3951
timestamp 1624857261
transform 1 0 188904 0 1 24213
box 0 0 1 1
use contact_32  contact_32_3950
timestamp 1624857261
transform 1 0 188904 0 1 23669
box 0 0 1 1
use contact_32  contact_32_3949
timestamp 1624857261
transform 1 0 188904 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3948
timestamp 1624857261
transform 1 0 188904 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3947
timestamp 1624857261
transform 1 0 189448 0 1 127029
box 0 0 1 1
use contact_32  contact_32_3946
timestamp 1624857261
transform 1 0 189448 0 1 126621
box 0 0 1 1
use contact_32  contact_32_3945
timestamp 1624857261
transform 1 0 191488 0 1 126485
box 0 0 1 1
use contact_32  contact_32_3944
timestamp 1624857261
transform 1 0 191488 0 1 126213
box 0 0 1 1
use contact_32  contact_32_3943
timestamp 1624857261
transform 1 0 195024 0 1 24349
box 0 0 1 1
use contact_32  contact_32_3942
timestamp 1624857261
transform 1 0 195024 0 1 25165
box 0 0 1 1
use contact_32  contact_32_3941
timestamp 1624857261
transform 1 0 194888 0 1 126077
box 0 0 1 1
use contact_32  contact_32_3940
timestamp 1624857261
transform 1 0 194888 0 1 125669
box 0 0 1 1
use contact_32  contact_32_3939
timestamp 1624857261
transform 1 0 195160 0 1 126077
box 0 0 1 1
use contact_32  contact_32_3938
timestamp 1624857261
transform 1 0 195160 0 1 125669
box 0 0 1 1
use contact_32  contact_32_3937
timestamp 1624857261
transform 1 0 196520 0 1 126213
box 0 0 1 1
use contact_32  contact_32_3936
timestamp 1624857261
transform 1 0 196520 0 1 129749
box 0 0 1 1
use contact_32  contact_32_3935
timestamp 1624857261
transform 1 0 195160 0 1 53997
box 0 0 1 1
use contact_32  contact_32_3934
timestamp 1624857261
transform 1 0 195160 0 1 53725
box 0 0 1 1
use contact_32  contact_32_3933
timestamp 1624857261
transform 1 0 195160 0 1 54133
box 0 0 1 1
use contact_32  contact_32_3932
timestamp 1624857261
transform 1 0 195160 0 1 54405
box 0 0 1 1
use contact_32  contact_32_3931
timestamp 1624857261
transform 1 0 195160 0 1 120365
box 0 0 1 1
use contact_32  contact_32_3930
timestamp 1624857261
transform 1 0 195160 0 1 120093
box 0 0 1 1
use contact_32  contact_32_3929
timestamp 1624857261
transform 1 0 195160 0 1 120501
box 0 0 1 1
use contact_32  contact_32_3928
timestamp 1624857261
transform 1 0 195160 0 1 120773
box 0 0 1 1
use contact_32  contact_32_3927
timestamp 1624857261
transform 1 0 195160 0 1 103093
box 0 0 1 1
use contact_32  contact_32_3926
timestamp 1624857261
transform 1 0 195160 0 1 103365
box 0 0 1 1
use contact_32  contact_32_3925
timestamp 1624857261
transform 1 0 195160 0 1 102957
box 0 0 1 1
use contact_32  contact_32_3924
timestamp 1624857261
transform 1 0 195160 0 1 102685
box 0 0 1 1
use contact_32  contact_32_3923
timestamp 1624857261
transform 1 0 195160 0 1 109349
box 0 0 1 1
use contact_32  contact_32_3922
timestamp 1624857261
transform 1 0 195160 0 1 109621
box 0 0 1 1
use contact_32  contact_32_3921
timestamp 1624857261
transform 1 0 195160 0 1 37949
box 0 0 1 1
use contact_32  contact_32_3920
timestamp 1624857261
transform 1 0 195160 0 1 38221
box 0 0 1 1
use contact_32  contact_32_3919
timestamp 1624857261
transform 1 0 195160 0 1 37813
box 0 0 1 1
use contact_32  contact_32_3918
timestamp 1624857261
transform 1 0 195160 0 1 37541
box 0 0 1 1
use contact_32  contact_32_3917
timestamp 1624857261
transform 1 0 195024 0 1 50189
box 0 0 1 1
use contact_32  contact_32_3916
timestamp 1624857261
transform 1 0 195024 0 1 50461
box 0 0 1 1
use contact_32  contact_32_3915
timestamp 1624857261
transform 1 0 195024 0 1 50053
box 0 0 1 1
use contact_32  contact_32_3914
timestamp 1624857261
transform 1 0 195024 0 1 49781
box 0 0 1 1
use contact_32  contact_32_3913
timestamp 1624857261
transform 1 0 195160 0 1 47741
box 0 0 1 1
use contact_32  contact_32_3912
timestamp 1624857261
transform 1 0 195160 0 1 48013
box 0 0 1 1
use contact_32  contact_32_3911
timestamp 1624857261
transform 1 0 195160 0 1 47605
box 0 0 1 1
use contact_32  contact_32_3910
timestamp 1624857261
transform 1 0 195160 0 1 47333
box 0 0 1 1
use contact_32  contact_32_3909
timestamp 1624857261
transform 1 0 195160 0 1 28021
box 0 0 1 1
use contact_32  contact_32_3908
timestamp 1624857261
transform 1 0 195160 0 1 28293
box 0 0 1 1
use contact_32  contact_32_3907
timestamp 1624857261
transform 1 0 195160 0 1 27885
box 0 0 1 1
use contact_32  contact_32_3906
timestamp 1624857261
transform 1 0 195160 0 1 27613
box 0 0 1 1
use contact_32  contact_32_3905
timestamp 1624857261
transform 1 0 195160 0 1 74669
box 0 0 1 1
use contact_32  contact_32_3904
timestamp 1624857261
transform 1 0 195160 0 1 74941
box 0 0 1 1
use contact_32  contact_32_3903
timestamp 1624857261
transform 1 0 195160 0 1 74533
box 0 0 1 1
use contact_32  contact_32_3902
timestamp 1624857261
transform 1 0 195160 0 1 74261
box 0 0 1 1
use contact_32  contact_32_3901
timestamp 1624857261
transform 1 0 195160 0 1 110845
box 0 0 1 1
use contact_32  contact_32_3900
timestamp 1624857261
transform 1 0 195160 0 1 110573
box 0 0 1 1
use contact_32  contact_32_3899
timestamp 1624857261
transform 1 0 195024 0 1 110981
box 0 0 1 1
use contact_32  contact_32_3898
timestamp 1624857261
transform 1 0 195024 0 1 111253
box 0 0 1 1
use contact_32  contact_32_3897
timestamp 1624857261
transform 1 0 195160 0 1 110437
box 0 0 1 1
use contact_32  contact_32_3896
timestamp 1624857261
transform 1 0 195160 0 1 110165
box 0 0 1 1
use contact_32  contact_32_3895
timestamp 1624857261
transform 1 0 195160 0 1 83373
box 0 0 1 1
use contact_32  contact_32_3894
timestamp 1624857261
transform 1 0 195160 0 1 83645
box 0 0 1 1
use contact_32  contact_32_3893
timestamp 1624857261
transform 1 0 195160 0 1 83237
box 0 0 1 1
use contact_32  contact_32_3892
timestamp 1624857261
transform 1 0 195160 0 1 82965
box 0 0 1 1
use contact_32  contact_32_3891
timestamp 1624857261
transform 1 0 195160 0 1 65829
box 0 0 1 1
use contact_32  contact_32_3890
timestamp 1624857261
transform 1 0 195160 0 1 65557
box 0 0 1 1
use contact_32  contact_32_3889
timestamp 1624857261
transform 1 0 195160 0 1 65965
box 0 0 1 1
use contact_32  contact_32_3888
timestamp 1624857261
transform 1 0 195160 0 1 66237
box 0 0 1 1
use contact_32  contact_32_3887
timestamp 1624857261
transform 1 0 195160 0 1 36725
box 0 0 1 1
use contact_32  contact_32_3886
timestamp 1624857261
transform 1 0 195160 0 1 36997
box 0 0 1 1
use contact_32  contact_32_3885
timestamp 1624857261
transform 1 0 195160 0 1 36589
box 0 0 1 1
use contact_32  contact_32_3884
timestamp 1624857261
transform 1 0 195160 0 1 36317
box 0 0 1 1
use contact_32  contact_32_3883
timestamp 1624857261
transform 1 0 195160 0 1 81197
box 0 0 1 1
use contact_32  contact_32_3882
timestamp 1624857261
transform 1 0 195160 0 1 80925
box 0 0 1 1
use contact_32  contact_32_3881
timestamp 1624857261
transform 1 0 195160 0 1 81333
box 0 0 1 1
use contact_32  contact_32_3880
timestamp 1624857261
transform 1 0 195160 0 1 81605
box 0 0 1 1
use contact_32  contact_32_3879
timestamp 1624857261
transform 1 0 195024 0 1 108125
box 0 0 1 1
use contact_32  contact_32_3878
timestamp 1624857261
transform 1 0 195024 0 1 107853
box 0 0 1 1
use contact_32  contact_32_3877
timestamp 1624857261
transform 1 0 195024 0 1 49237
box 0 0 1 1
use contact_32  contact_32_3876
timestamp 1624857261
transform 1 0 195024 0 1 48965
box 0 0 1 1
use contact_32  contact_32_3875
timestamp 1624857261
transform 1 0 195024 0 1 49373
box 0 0 1 1
use contact_32  contact_32_3874
timestamp 1624857261
transform 1 0 195024 0 1 49645
box 0 0 1 1
use contact_32  contact_32_3873
timestamp 1624857261
transform 1 0 195024 0 1 107037
box 0 0 1 1
use contact_32  contact_32_3872
timestamp 1624857261
transform 1 0 195024 0 1 107309
box 0 0 1 1
use contact_32  contact_32_3871
timestamp 1624857261
transform 1 0 195024 0 1 106901
box 0 0 1 1
use contact_32  contact_32_3870
timestamp 1624857261
transform 1 0 195024 0 1 106629
box 0 0 1 1
use contact_32  contact_32_3869
timestamp 1624857261
transform 1 0 195024 0 1 114381
box 0 0 1 1
use contact_32  contact_32_3868
timestamp 1624857261
transform 1 0 195024 0 1 114109
box 0 0 1 1
use contact_32  contact_32_3867
timestamp 1624857261
transform 1 0 195024 0 1 114517
box 0 0 1 1
use contact_32  contact_32_3866
timestamp 1624857261
transform 1 0 195024 0 1 114789
box 0 0 1 1
use contact_32  contact_32_3865
timestamp 1624857261
transform 1 0 195024 0 1 68549
box 0 0 1 1
use contact_32  contact_32_3864
timestamp 1624857261
transform 1 0 195024 0 1 68277
box 0 0 1 1
use contact_32  contact_32_3863
timestamp 1624857261
transform 1 0 195024 0 1 68685
box 0 0 1 1
use contact_32  contact_32_3862
timestamp 1624857261
transform 1 0 195024 0 1 68957
box 0 0 1 1
use contact_32  contact_32_3861
timestamp 1624857261
transform 1 0 195160 0 1 122405
box 0 0 1 1
use contact_32  contact_32_3860
timestamp 1624857261
transform 1 0 195160 0 1 122677
box 0 0 1 1
use contact_32  contact_32_3859
timestamp 1624857261
transform 1 0 195024 0 1 122269
box 0 0 1 1
use contact_32  contact_32_3858
timestamp 1624857261
transform 1 0 195024 0 1 121997
box 0 0 1 1
use contact_32  contact_32_3857
timestamp 1624857261
transform 1 0 195024 0 1 43661
box 0 0 1 1
use contact_32  contact_32_3856
timestamp 1624857261
transform 1 0 195024 0 1 43389
box 0 0 1 1
use contact_32  contact_32_3855
timestamp 1624857261
transform 1 0 195024 0 1 43797
box 0 0 1 1
use contact_32  contact_32_3854
timestamp 1624857261
transform 1 0 195024 0 1 44069
box 0 0 1 1
use contact_32  contact_32_3853
timestamp 1624857261
transform 1 0 195024 0 1 103501
box 0 0 1 1
use contact_32  contact_32_3852
timestamp 1624857261
transform 1 0 195024 0 1 103773
box 0 0 1 1
use contact_32  contact_32_3851
timestamp 1624857261
transform 1 0 195160 0 1 78885
box 0 0 1 1
use contact_32  contact_32_3850
timestamp 1624857261
transform 1 0 195160 0 1 78613
box 0 0 1 1
use contact_32  contact_32_3849
timestamp 1624857261
transform 1 0 195160 0 1 79021
box 0 0 1 1
use contact_32  contact_32_3848
timestamp 1624857261
transform 1 0 195160 0 1 79293
box 0 0 1 1
use contact_32  contact_32_3847
timestamp 1624857261
transform 1 0 195024 0 1 73037
box 0 0 1 1
use contact_32  contact_32_3846
timestamp 1624857261
transform 1 0 195024 0 1 73309
box 0 0 1 1
use contact_32  contact_32_3845
timestamp 1624857261
transform 1 0 195024 0 1 72901
box 0 0 1 1
use contact_32  contact_32_3844
timestamp 1624857261
transform 1 0 195024 0 1 72629
box 0 0 1 1
use contact_32  contact_32_3843
timestamp 1624857261
transform 1 0 195160 0 1 32373
box 0 0 1 1
use contact_32  contact_32_3842
timestamp 1624857261
transform 1 0 195160 0 1 32645
box 0 0 1 1
use contact_32  contact_32_3841
timestamp 1624857261
transform 1 0 195160 0 1 32237
box 0 0 1 1
use contact_32  contact_32_3840
timestamp 1624857261
transform 1 0 195160 0 1 31965
box 0 0 1 1
use contact_32  contact_32_3839
timestamp 1624857261
transform 1 0 195024 0 1 66645
box 0 0 1 1
use contact_32  contact_32_3838
timestamp 1624857261
transform 1 0 195024 0 1 66373
box 0 0 1 1
use contact_32  contact_32_3837
timestamp 1624857261
transform 1 0 195024 0 1 66781
box 0 0 1 1
use contact_32  contact_32_3836
timestamp 1624857261
transform 1 0 195024 0 1 67053
box 0 0 1 1
use contact_32  contact_32_3835
timestamp 1624857261
transform 1 0 195160 0 1 39037
box 0 0 1 1
use contact_32  contact_32_3834
timestamp 1624857261
transform 1 0 195160 0 1 39309
box 0 0 1 1
use contact_32  contact_32_3833
timestamp 1624857261
transform 1 0 195024 0 1 57941
box 0 0 1 1
use contact_32  contact_32_3832
timestamp 1624857261
transform 1 0 195024 0 1 57669
box 0 0 1 1
use contact_32  contact_32_3831
timestamp 1624857261
transform 1 0 195024 0 1 58077
box 0 0 1 1
use contact_32  contact_32_3830
timestamp 1624857261
transform 1 0 195024 0 1 58349
box 0 0 1 1
use contact_32  contact_32_3829
timestamp 1624857261
transform 1 0 195160 0 1 82149
box 0 0 1 1
use contact_32  contact_32_3828
timestamp 1624857261
transform 1 0 195160 0 1 82421
box 0 0 1 1
use contact_32  contact_32_3827
timestamp 1624857261
transform 1 0 195024 0 1 82013
box 0 0 1 1
use contact_32  contact_32_3826
timestamp 1624857261
transform 1 0 195024 0 1 81741
box 0 0 1 1
use contact_32  contact_32_3825
timestamp 1624857261
transform 1 0 195024 0 1 30741
box 0 0 1 1
use contact_32  contact_32_3824
timestamp 1624857261
transform 1 0 195024 0 1 31013
box 0 0 1 1
use contact_32  contact_32_3823
timestamp 1624857261
transform 1 0 195024 0 1 80789
box 0 0 1 1
use contact_32  contact_32_3822
timestamp 1624857261
transform 1 0 195024 0 1 80517
box 0 0 1 1
use contact_32  contact_32_3821
timestamp 1624857261
transform 1 0 195160 0 1 105405
box 0 0 1 1
use contact_32  contact_32_3820
timestamp 1624857261
transform 1 0 195160 0 1 105677
box 0 0 1 1
use contact_32  contact_32_3819
timestamp 1624857261
transform 1 0 195024 0 1 95885
box 0 0 1 1
use contact_32  contact_32_3818
timestamp 1624857261
transform 1 0 195024 0 1 95613
box 0 0 1 1
use contact_32  contact_32_3817
timestamp 1624857261
transform 1 0 195024 0 1 101325
box 0 0 1 1
use contact_32  contact_32_3816
timestamp 1624857261
transform 1 0 195024 0 1 101053
box 0 0 1 1
use contact_32  contact_32_3815
timestamp 1624857261
transform 1 0 195024 0 1 101461
box 0 0 1 1
use contact_32  contact_32_3814
timestamp 1624857261
transform 1 0 195024 0 1 101733
box 0 0 1 1
use contact_32  contact_32_3813
timestamp 1624857261
transform 1 0 195024 0 1 53589
box 0 0 1 1
use contact_32  contact_32_3812
timestamp 1624857261
transform 1 0 195024 0 1 53317
box 0 0 1 1
use contact_32  contact_32_3811
timestamp 1624857261
transform 1 0 195024 0 1 93845
box 0 0 1 1
use contact_32  contact_32_3810
timestamp 1624857261
transform 1 0 195024 0 1 93573
box 0 0 1 1
use contact_32  contact_32_3809
timestamp 1624857261
transform 1 0 195024 0 1 93981
box 0 0 1 1
use contact_32  contact_32_3808
timestamp 1624857261
transform 1 0 195024 0 1 94253
box 0 0 1 1
use contact_32  contact_32_3807
timestamp 1624857261
transform 1 0 195024 0 1 100237
box 0 0 1 1
use contact_32  contact_32_3806
timestamp 1624857261
transform 1 0 195024 0 1 99965
box 0 0 1 1
use contact_32  contact_32_3805
timestamp 1624857261
transform 1 0 195160 0 1 116149
box 0 0 1 1
use contact_32  contact_32_3804
timestamp 1624857261
transform 1 0 195160 0 1 116421
box 0 0 1 1
use contact_32  contact_32_3803
timestamp 1624857261
transform 1 0 195160 0 1 116013
box 0 0 1 1
use contact_32  contact_32_3802
timestamp 1624857261
transform 1 0 195160 0 1 115741
box 0 0 1 1
use contact_32  contact_32_3801
timestamp 1624857261
transform 1 0 195160 0 1 107445
box 0 0 1 1
use contact_32  contact_32_3800
timestamp 1624857261
transform 1 0 195160 0 1 107717
box 0 0 1 1
use contact_32  contact_32_3799
timestamp 1624857261
transform 1 0 195024 0 1 65421
box 0 0 1 1
use contact_32  contact_32_3798
timestamp 1624857261
transform 1 0 195024 0 1 65149
box 0 0 1 1
use contact_32  contact_32_3797
timestamp 1624857261
transform 1 0 195160 0 1 56037
box 0 0 1 1
use contact_32  contact_32_3796
timestamp 1624857261
transform 1 0 195160 0 1 56309
box 0 0 1 1
use contact_32  contact_32_3795
timestamp 1624857261
transform 1 0 195024 0 1 55901
box 0 0 1 1
use contact_32  contact_32_3794
timestamp 1624857261
transform 1 0 195024 0 1 55629
box 0 0 1 1
use contact_32  contact_32_3793
timestamp 1624857261
transform 1 0 195024 0 1 86093
box 0 0 1 1
use contact_32  contact_32_3792
timestamp 1624857261
transform 1 0 195024 0 1 86365
box 0 0 1 1
use contact_32  contact_32_3791
timestamp 1624857261
transform 1 0 195024 0 1 85957
box 0 0 1 1
use contact_32  contact_32_3790
timestamp 1624857261
transform 1 0 195024 0 1 85685
box 0 0 1 1
use contact_32  contact_32_3789
timestamp 1624857261
transform 1 0 195024 0 1 72221
box 0 0 1 1
use contact_32  contact_32_3788
timestamp 1624857261
transform 1 0 195024 0 1 72493
box 0 0 1 1
use contact_32  contact_32_3787
timestamp 1624857261
transform 1 0 195024 0 1 59981
box 0 0 1 1
use contact_32  contact_32_3786
timestamp 1624857261
transform 1 0 195024 0 1 60253
box 0 0 1 1
use contact_32  contact_32_3785
timestamp 1624857261
transform 1 0 195160 0 1 53181
box 0 0 1 1
use contact_32  contact_32_3784
timestamp 1624857261
transform 1 0 195160 0 1 52909
box 0 0 1 1
use contact_32  contact_32_3783
timestamp 1624857261
transform 1 0 195024 0 1 27205
box 0 0 1 1
use contact_32  contact_32_3782
timestamp 1624857261
transform 1 0 195024 0 1 27477
box 0 0 1 1
use contact_32  contact_32_3781
timestamp 1624857261
transform 1 0 195160 0 1 27069
box 0 0 1 1
use contact_32  contact_32_3780
timestamp 1624857261
transform 1 0 195160 0 1 26797
box 0 0 1 1
use contact_32  contact_32_3779
timestamp 1624857261
transform 1 0 195160 0 1 28837
box 0 0 1 1
use contact_32  contact_32_3778
timestamp 1624857261
transform 1 0 195160 0 1 29109
box 0 0 1 1
use contact_32  contact_32_3777
timestamp 1624857261
transform 1 0 195024 0 1 28701
box 0 0 1 1
use contact_32  contact_32_3776
timestamp 1624857261
transform 1 0 195024 0 1 28429
box 0 0 1 1
use contact_32  contact_32_3775
timestamp 1624857261
transform 1 0 195160 0 1 45429
box 0 0 1 1
use contact_32  contact_32_3774
timestamp 1624857261
transform 1 0 195160 0 1 45701
box 0 0 1 1
use contact_32  contact_32_3773
timestamp 1624857261
transform 1 0 195160 0 1 45293
box 0 0 1 1
use contact_32  contact_32_3772
timestamp 1624857261
transform 1 0 195160 0 1 45021
box 0 0 1 1
use contact_32  contact_32_3771
timestamp 1624857261
transform 1 0 195160 0 1 29245
box 0 0 1 1
use contact_32  contact_32_3770
timestamp 1624857261
transform 1 0 195160 0 1 29517
box 0 0 1 1
use contact_32  contact_32_3769
timestamp 1624857261
transform 1 0 195024 0 1 112477
box 0 0 1 1
use contact_32  contact_32_3768
timestamp 1624857261
transform 1 0 195024 0 1 112205
box 0 0 1 1
use contact_32  contact_32_3767
timestamp 1624857261
transform 1 0 195024 0 1 99421
box 0 0 1 1
use contact_32  contact_32_3766
timestamp 1624857261
transform 1 0 195024 0 1 99149
box 0 0 1 1
use contact_32  contact_32_3765
timestamp 1624857261
transform 1 0 195160 0 1 99557
box 0 0 1 1
use contact_32  contact_32_3764
timestamp 1624857261
transform 1 0 195160 0 1 99829
box 0 0 1 1
use contact_32  contact_32_3763
timestamp 1624857261
transform 1 0 195024 0 1 97109
box 0 0 1 1
use contact_32  contact_32_3762
timestamp 1624857261
transform 1 0 195024 0 1 97381
box 0 0 1 1
use contact_32  contact_32_3761
timestamp 1624857261
transform 1 0 195024 0 1 70997
box 0 0 1 1
use contact_32  contact_32_3760
timestamp 1624857261
transform 1 0 195024 0 1 70725
box 0 0 1 1
use contact_32  contact_32_3759
timestamp 1624857261
transform 1 0 195024 0 1 62021
box 0 0 1 1
use contact_32  contact_32_3758
timestamp 1624857261
transform 1 0 195024 0 1 62293
box 0 0 1 1
use contact_32  contact_32_3757
timestamp 1624857261
transform 1 0 195160 0 1 61885
box 0 0 1 1
use contact_32  contact_32_3756
timestamp 1624857261
transform 1 0 195160 0 1 61613
box 0 0 1 1
use contact_32  contact_32_3755
timestamp 1624857261
transform 1 0 195160 0 1 73717
box 0 0 1 1
use contact_32  contact_32_3754
timestamp 1624857261
transform 1 0 195160 0 1 73445
box 0 0 1 1
use contact_32  contact_32_3753
timestamp 1624857261
transform 1 0 195160 0 1 73853
box 0 0 1 1
use contact_32  contact_32_3752
timestamp 1624857261
transform 1 0 195160 0 1 74125
box 0 0 1 1
use contact_32  contact_32_3751
timestamp 1624857261
transform 1 0 195024 0 1 112069
box 0 0 1 1
use contact_32  contact_32_3750
timestamp 1624857261
transform 1 0 195024 0 1 111797
box 0 0 1 1
use contact_32  contact_32_3749
timestamp 1624857261
transform 1 0 195024 0 1 99013
box 0 0 1 1
use contact_32  contact_32_3748
timestamp 1624857261
transform 1 0 195024 0 1 98741
box 0 0 1 1
use contact_32  contact_32_3747
timestamp 1624857261
transform 1 0 195024 0 1 48149
box 0 0 1 1
use contact_32  contact_32_3746
timestamp 1624857261
transform 1 0 195024 0 1 48421
box 0 0 1 1
use contact_32  contact_32_3745
timestamp 1624857261
transform 1 0 195160 0 1 78069
box 0 0 1 1
use contact_32  contact_32_3744
timestamp 1624857261
transform 1 0 195160 0 1 77797
box 0 0 1 1
use contact_32  contact_32_3743
timestamp 1624857261
transform 1 0 195160 0 1 78205
box 0 0 1 1
use contact_32  contact_32_3742
timestamp 1624857261
transform 1 0 195160 0 1 78477
box 0 0 1 1
use contact_32  contact_32_3741
timestamp 1624857261
transform 1 0 195024 0 1 97925
box 0 0 1 1
use contact_32  contact_32_3740
timestamp 1624857261
transform 1 0 195024 0 1 98197
box 0 0 1 1
use contact_32  contact_32_3739
timestamp 1624857261
transform 1 0 195160 0 1 97789
box 0 0 1 1
use contact_32  contact_32_3738
timestamp 1624857261
transform 1 0 195160 0 1 97517
box 0 0 1 1
use contact_32  contact_32_3737
timestamp 1624857261
transform 1 0 195160 0 1 70589
box 0 0 1 1
use contact_32  contact_32_3736
timestamp 1624857261
transform 1 0 195160 0 1 70317
box 0 0 1 1
use contact_32  contact_32_3735
timestamp 1624857261
transform 1 0 195160 0 1 57533
box 0 0 1 1
use contact_32  contact_32_3734
timestamp 1624857261
transform 1 0 195160 0 1 57261
box 0 0 1 1
use contact_32  contact_32_3733
timestamp 1624857261
transform 1 0 195160 0 1 48829
box 0 0 1 1
use contact_32  contact_32_3732
timestamp 1624857261
transform 1 0 195160 0 1 48557
box 0 0 1 1
use contact_32  contact_32_3731
timestamp 1624857261
transform 1 0 195160 0 1 93437
box 0 0 1 1
use contact_32  contact_32_3730
timestamp 1624857261
transform 1 0 195160 0 1 93165
box 0 0 1 1
use contact_32  contact_32_3729
timestamp 1624857261
transform 1 0 195024 0 1 94661
box 0 0 1 1
use contact_32  contact_32_3728
timestamp 1624857261
transform 1 0 195024 0 1 94389
box 0 0 1 1
use contact_32  contact_32_3727
timestamp 1624857261
transform 1 0 195024 0 1 94797
box 0 0 1 1
use contact_32  contact_32_3726
timestamp 1624857261
transform 1 0 195024 0 1 95069
box 0 0 1 1
use contact_32  contact_32_3725
timestamp 1624857261
transform 1 0 195024 0 1 118733
box 0 0 1 1
use contact_32  contact_32_3724
timestamp 1624857261
transform 1 0 195024 0 1 118461
box 0 0 1 1
use contact_32  contact_32_3723
timestamp 1624857261
transform 1 0 195024 0 1 118869
box 0 0 1 1
use contact_32  contact_32_3722
timestamp 1624857261
transform 1 0 195024 0 1 119141
box 0 0 1 1
use contact_32  contact_32_3721
timestamp 1624857261
transform 1 0 195160 0 1 113973
box 0 0 1 1
use contact_32  contact_32_3720
timestamp 1624857261
transform 1 0 195160 0 1 113701
box 0 0 1 1
use contact_32  contact_32_3719
timestamp 1624857261
transform 1 0 195024 0 1 77661
box 0 0 1 1
use contact_32  contact_32_3718
timestamp 1624857261
transform 1 0 195024 0 1 77389
box 0 0 1 1
use contact_32  contact_32_3717
timestamp 1624857261
transform 1 0 195160 0 1 35501
box 0 0 1 1
use contact_32  contact_32_3716
timestamp 1624857261
transform 1 0 195160 0 1 35773
box 0 0 1 1
use contact_32  contact_32_3715
timestamp 1624857261
transform 1 0 195160 0 1 35365
box 0 0 1 1
use contact_32  contact_32_3714
timestamp 1624857261
transform 1 0 195160 0 1 35093
box 0 0 1 1
use contact_32  contact_32_3713
timestamp 1624857261
transform 1 0 195160 0 1 31421
box 0 0 1 1
use contact_32  contact_32_3712
timestamp 1624857261
transform 1 0 195160 0 1 31149
box 0 0 1 1
use contact_32  contact_32_3711
timestamp 1624857261
transform 1 0 195024 0 1 31557
box 0 0 1 1
use contact_32  contact_32_3710
timestamp 1624857261
transform 1 0 195024 0 1 31829
box 0 0 1 1
use contact_32  contact_32_3709
timestamp 1624857261
transform 1 0 195160 0 1 51685
box 0 0 1 1
use contact_32  contact_32_3708
timestamp 1624857261
transform 1 0 195160 0 1 51957
box 0 0 1 1
use contact_32  contact_32_3707
timestamp 1624857261
transform 1 0 195160 0 1 41077
box 0 0 1 1
use contact_32  contact_32_3706
timestamp 1624857261
transform 1 0 195160 0 1 41349
box 0 0 1 1
use contact_32  contact_32_3705
timestamp 1624857261
transform 1 0 195160 0 1 40941
box 0 0 1 1
use contact_32  contact_32_3704
timestamp 1624857261
transform 1 0 195160 0 1 40669
box 0 0 1 1
use contact_32  contact_32_3703
timestamp 1624857261
transform 1 0 195160 0 1 39853
box 0 0 1 1
use contact_32  contact_32_3702
timestamp 1624857261
transform 1 0 195160 0 1 40125
box 0 0 1 1
use contact_32  contact_32_3701
timestamp 1624857261
transform 1 0 195160 0 1 39717
box 0 0 1 1
use contact_32  contact_32_3700
timestamp 1624857261
transform 1 0 195160 0 1 39445
box 0 0 1 1
use contact_32  contact_32_3699
timestamp 1624857261
transform 1 0 195160 0 1 123901
box 0 0 1 1
use contact_32  contact_32_3698
timestamp 1624857261
transform 1 0 195160 0 1 123629
box 0 0 1 1
use contact_32  contact_32_3697
timestamp 1624857261
transform 1 0 195024 0 1 124037
box 0 0 1 1
use contact_32  contact_32_3696
timestamp 1624857261
transform 1 0 195024 0 1 124309
box 0 0 1 1
use contact_32  contact_32_3695
timestamp 1624857261
transform 1 0 195024 0 1 62429
box 0 0 1 1
use contact_32  contact_32_3694
timestamp 1624857261
transform 1 0 195024 0 1 62701
box 0 0 1 1
use contact_32  contact_32_3693
timestamp 1624857261
transform 1 0 195024 0 1 111389
box 0 0 1 1
use contact_32  contact_32_3692
timestamp 1624857261
transform 1 0 195024 0 1 111661
box 0 0 1 1
use contact_32  contact_32_3691
timestamp 1624857261
transform 1 0 195160 0 1 42165
box 0 0 1 1
use contact_32  contact_32_3690
timestamp 1624857261
transform 1 0 195160 0 1 41893
box 0 0 1 1
use contact_32  contact_32_3689
timestamp 1624857261
transform 1 0 195160 0 1 29925
box 0 0 1 1
use contact_32  contact_32_3688
timestamp 1624857261
transform 1 0 195160 0 1 29653
box 0 0 1 1
use contact_32  contact_32_3687
timestamp 1624857261
transform 1 0 195024 0 1 69909
box 0 0 1 1
use contact_32  contact_32_3686
timestamp 1624857261
transform 1 0 195024 0 1 70181
box 0 0 1 1
use contact_32  contact_32_3685
timestamp 1624857261
transform 1 0 195024 0 1 69773
box 0 0 1 1
use contact_32  contact_32_3684
timestamp 1624857261
transform 1 0 195024 0 1 69501
box 0 0 1 1
use contact_32  contact_32_3683
timestamp 1624857261
transform 1 0 195024 0 1 119957
box 0 0 1 1
use contact_32  contact_32_3682
timestamp 1624857261
transform 1 0 195024 0 1 119685
box 0 0 1 1
use contact_32  contact_32_3681
timestamp 1624857261
transform 1 0 195024 0 1 35909
box 0 0 1 1
use contact_32  contact_32_3680
timestamp 1624857261
transform 1 0 195024 0 1 36181
box 0 0 1 1
use contact_32  contact_32_3679
timestamp 1624857261
transform 1 0 195160 0 1 52093
box 0 0 1 1
use contact_32  contact_32_3678
timestamp 1624857261
transform 1 0 195160 0 1 52365
box 0 0 1 1
use contact_32  contact_32_3677
timestamp 1624857261
transform 1 0 195160 0 1 61477
box 0 0 1 1
use contact_32  contact_32_3676
timestamp 1624857261
transform 1 0 195160 0 1 61205
box 0 0 1 1
use contact_32  contact_32_3675
timestamp 1624857261
transform 1 0 195160 0 1 46517
box 0 0 1 1
use contact_32  contact_32_3674
timestamp 1624857261
transform 1 0 195160 0 1 46245
box 0 0 1 1
use contact_32  contact_32_3673
timestamp 1624857261
transform 1 0 195024 0 1 45837
box 0 0 1 1
use contact_32  contact_32_3672
timestamp 1624857261
transform 1 0 195024 0 1 46109
box 0 0 1 1
use contact_32  contact_32_3671
timestamp 1624857261
transform 1 0 195024 0 1 32781
box 0 0 1 1
use contact_32  contact_32_3670
timestamp 1624857261
transform 1 0 195024 0 1 33053
box 0 0 1 1
use contact_32  contact_32_3669
timestamp 1624857261
transform 1 0 195024 0 1 37133
box 0 0 1 1
use contact_32  contact_32_3668
timestamp 1624857261
transform 1 0 195024 0 1 37405
box 0 0 1 1
use contact_32  contact_32_3667
timestamp 1624857261
transform 1 0 195160 0 1 118053
box 0 0 1 1
use contact_32  contact_32_3666
timestamp 1624857261
transform 1 0 195160 0 1 118325
box 0 0 1 1
use contact_32  contact_32_3665
timestamp 1624857261
transform 1 0 195024 0 1 117917
box 0 0 1 1
use contact_32  contact_32_3664
timestamp 1624857261
transform 1 0 195024 0 1 117645
box 0 0 1 1
use contact_32  contact_32_3663
timestamp 1624857261
transform 1 0 195024 0 1 75349
box 0 0 1 1
use contact_32  contact_32_3662
timestamp 1624857261
transform 1 0 195024 0 1 75077
box 0 0 1 1
use contact_32  contact_32_3661
timestamp 1624857261
transform 1 0 195024 0 1 90717
box 0 0 1 1
use contact_32  contact_32_3660
timestamp 1624857261
transform 1 0 195024 0 1 90445
box 0 0 1 1
use contact_32  contact_32_3659
timestamp 1624857261
transform 1 0 195160 0 1 90853
box 0 0 1 1
use contact_32  contact_32_3658
timestamp 1624857261
transform 1 0 195160 0 1 91125
box 0 0 1 1
use contact_32  contact_32_3657
timestamp 1624857261
transform 1 0 195160 0 1 123493
box 0 0 1 1
use contact_32  contact_32_3656
timestamp 1624857261
transform 1 0 195160 0 1 123221
box 0 0 1 1
use contact_32  contact_32_3655
timestamp 1624857261
transform 1 0 195024 0 1 41485
box 0 0 1 1
use contact_32  contact_32_3654
timestamp 1624857261
transform 1 0 195024 0 1 41757
box 0 0 1 1
use contact_32  contact_32_3653
timestamp 1624857261
transform 1 0 195024 0 1 90309
box 0 0 1 1
use contact_32  contact_32_3652
timestamp 1624857261
transform 1 0 195024 0 1 90037
box 0 0 1 1
use contact_32  contact_32_3651
timestamp 1624857261
transform 1 0 195024 0 1 40261
box 0 0 1 1
use contact_32  contact_32_3650
timestamp 1624857261
transform 1 0 195024 0 1 40533
box 0 0 1 1
use contact_32  contact_32_3649
timestamp 1624857261
transform 1 0 195160 0 1 102141
box 0 0 1 1
use contact_32  contact_32_3648
timestamp 1624857261
transform 1 0 195160 0 1 101869
box 0 0 1 1
use contact_32  contact_32_3647
timestamp 1624857261
transform 1 0 195024 0 1 102277
box 0 0 1 1
use contact_32  contact_32_3646
timestamp 1624857261
transform 1 0 195024 0 1 102549
box 0 0 1 1
use contact_32  contact_32_3645
timestamp 1624857261
transform 1 0 195160 0 1 57125
box 0 0 1 1
use contact_32  contact_32_3644
timestamp 1624857261
transform 1 0 195160 0 1 56853
box 0 0 1 1
use contact_32  contact_32_3643
timestamp 1624857261
transform 1 0 195024 0 1 92757
box 0 0 1 1
use contact_32  contact_32_3642
timestamp 1624857261
transform 1 0 195024 0 1 93029
box 0 0 1 1
use contact_32  contact_32_3641
timestamp 1624857261
transform 1 0 195160 0 1 33597
box 0 0 1 1
use contact_32  contact_32_3640
timestamp 1624857261
transform 1 0 195160 0 1 33869
box 0 0 1 1
use contact_32  contact_32_3639
timestamp 1624857261
transform 1 0 195160 0 1 33461
box 0 0 1 1
use contact_32  contact_32_3638
timestamp 1624857261
transform 1 0 195160 0 1 33189
box 0 0 1 1
use contact_32  contact_32_3637
timestamp 1624857261
transform 1 0 195024 0 1 44613
box 0 0 1 1
use contact_32  contact_32_3636
timestamp 1624857261
transform 1 0 195024 0 1 44885
box 0 0 1 1
use contact_32  contact_32_3635
timestamp 1624857261
transform 1 0 195160 0 1 44477
box 0 0 1 1
use contact_32  contact_32_3634
timestamp 1624857261
transform 1 0 195160 0 1 44205
box 0 0 1 1
use contact_32  contact_32_3633
timestamp 1624857261
transform 1 0 195160 0 1 76981
box 0 0 1 1
use contact_32  contact_32_3632
timestamp 1624857261
transform 1 0 195160 0 1 77253
box 0 0 1 1
use contact_32  contact_32_3631
timestamp 1624857261
transform 1 0 195160 0 1 76845
box 0 0 1 1
use contact_32  contact_32_3630
timestamp 1624857261
transform 1 0 195160 0 1 76573
box 0 0 1 1
use contact_32  contact_32_3629
timestamp 1624857261
transform 1 0 195160 0 1 52773
box 0 0 1 1
use contact_32  contact_32_3628
timestamp 1624857261
transform 1 0 195160 0 1 52501
box 0 0 1 1
use contact_32  contact_32_3627
timestamp 1624857261
transform 1 0 195160 0 1 114925
box 0 0 1 1
use contact_32  contact_32_3626
timestamp 1624857261
transform 1 0 195160 0 1 115197
box 0 0 1 1
use contact_32  contact_32_3625
timestamp 1624857261
transform 1 0 195160 0 1 86501
box 0 0 1 1
use contact_32  contact_32_3624
timestamp 1624857261
transform 1 0 195160 0 1 86773
box 0 0 1 1
use contact_32  contact_32_3623
timestamp 1624857261
transform 1 0 195160 0 1 58485
box 0 0 1 1
use contact_32  contact_32_3622
timestamp 1624857261
transform 1 0 195160 0 1 58757
box 0 0 1 1
use contact_32  contact_32_3621
timestamp 1624857261
transform 1 0 195160 0 1 91941
box 0 0 1 1
use contact_32  contact_32_3620
timestamp 1624857261
transform 1 0 195160 0 1 91669
box 0 0 1 1
use contact_32  contact_32_3619
timestamp 1624857261
transform 1 0 195024 0 1 91533
box 0 0 1 1
use contact_32  contact_32_3618
timestamp 1624857261
transform 1 0 195024 0 1 91261
box 0 0 1 1
use contact_32  contact_32_3617
timestamp 1624857261
transform 1 0 195024 0 1 110029
box 0 0 1 1
use contact_32  contact_32_3616
timestamp 1624857261
transform 1 0 195024 0 1 109757
box 0 0 1 1
use contact_32  contact_32_3615
timestamp 1624857261
transform 1 0 195160 0 1 82557
box 0 0 1 1
use contact_32  contact_32_3614
timestamp 1624857261
transform 1 0 195160 0 1 82829
box 0 0 1 1
use contact_32  contact_32_3613
timestamp 1624857261
transform 1 0 195160 0 1 95477
box 0 0 1 1
use contact_32  contact_32_3612
timestamp 1624857261
transform 1 0 195160 0 1 95205
box 0 0 1 1
use contact_32  contact_32_3611
timestamp 1624857261
transform 1 0 195024 0 1 89221
box 0 0 1 1
use contact_32  contact_32_3610
timestamp 1624857261
transform 1 0 195024 0 1 89493
box 0 0 1 1
use contact_32  contact_32_3609
timestamp 1624857261
transform 1 0 195160 0 1 89085
box 0 0 1 1
use contact_32  contact_32_3608
timestamp 1624857261
transform 1 0 195160 0 1 88813
box 0 0 1 1
use contact_32  contact_32_3607
timestamp 1624857261
transform 1 0 195024 0 1 61069
box 0 0 1 1
use contact_32  contact_32_3606
timestamp 1624857261
transform 1 0 195024 0 1 60797
box 0 0 1 1
use contact_32  contact_32_3605
timestamp 1624857261
transform 1 0 195024 0 1 25301
box 0 0 1 1
use contact_32  contact_32_3604
timestamp 1624857261
transform 1 0 195024 0 1 25573
box 0 0 1 1
use contact_32  contact_32_3603
timestamp 1624857261
transform 1 0 195024 0 1 89629
box 0 0 1 1
use contact_32  contact_32_3602
timestamp 1624857261
transform 1 0 195024 0 1 89901
box 0 0 1 1
use contact_32  contact_32_3601
timestamp 1624857261
transform 1 0 195160 0 1 122813
box 0 0 1 1
use contact_32  contact_32_3600
timestamp 1624857261
transform 1 0 195160 0 1 123085
box 0 0 1 1
use contact_32  contact_32_3599
timestamp 1624857261
transform 1 0 195160 0 1 60661
box 0 0 1 1
use contact_32  contact_32_3598
timestamp 1624857261
transform 1 0 195160 0 1 60389
box 0 0 1 1
use contact_32  contact_32_3597
timestamp 1624857261
transform 1 0 195160 0 1 56445
box 0 0 1 1
use contact_32  contact_32_3596
timestamp 1624857261
transform 1 0 195160 0 1 56717
box 0 0 1 1
use contact_32  contact_32_3595
timestamp 1624857261
transform 1 0 195024 0 1 98333
box 0 0 1 1
use contact_32  contact_32_3594
timestamp 1624857261
transform 1 0 195024 0 1 98605
box 0 0 1 1
use contact_32  contact_32_3593
timestamp 1624857261
transform 1 0 195024 0 1 85141
box 0 0 1 1
use contact_32  contact_32_3592
timestamp 1624857261
transform 1 0 195024 0 1 84869
box 0 0 1 1
use contact_32  contact_32_3591
timestamp 1624857261
transform 1 0 195024 0 1 85277
box 0 0 1 1
use contact_32  contact_32_3590
timestamp 1624857261
transform 1 0 195024 0 1 85549
box 0 0 1 1
use contact_32  contact_32_3589
timestamp 1624857261
transform 1 0 195024 0 1 87317
box 0 0 1 1
use contact_32  contact_32_3588
timestamp 1624857261
transform 1 0 195024 0 1 87589
box 0 0 1 1
use contact_32  contact_32_3587
timestamp 1624857261
transform 1 0 195024 0 1 87181
box 0 0 1 1
use contact_32  contact_32_3586
timestamp 1624857261
transform 1 0 195024 0 1 86909
box 0 0 1 1
use contact_32  contact_32_3585
timestamp 1624857261
transform 1 0 195160 0 1 65013
box 0 0 1 1
use contact_32  contact_32_3584
timestamp 1624857261
transform 1 0 195160 0 1 64741
box 0 0 1 1
use contact_32  contact_32_3583
timestamp 1624857261
transform 1 0 195160 0 1 69093
box 0 0 1 1
use contact_32  contact_32_3582
timestamp 1624857261
transform 1 0 195160 0 1 69365
box 0 0 1 1
use contact_32  contact_32_3581
timestamp 1624857261
transform 1 0 195160 0 1 106221
box 0 0 1 1
use contact_32  contact_32_3580
timestamp 1624857261
transform 1 0 195160 0 1 106493
box 0 0 1 1
use contact_32  contact_32_3579
timestamp 1624857261
transform 1 0 195160 0 1 106085
box 0 0 1 1
use contact_32  contact_32_3578
timestamp 1624857261
transform 1 0 195160 0 1 105813
box 0 0 1 1
use contact_32  contact_32_3577
timestamp 1624857261
transform 1 0 195160 0 1 63925
box 0 0 1 1
use contact_32  contact_32_3576
timestamp 1624857261
transform 1 0 195160 0 1 64197
box 0 0 1 1
use contact_32  contact_32_3575
timestamp 1624857261
transform 1 0 195160 0 1 84733
box 0 0 1 1
use contact_32  contact_32_3574
timestamp 1624857261
transform 1 0 195160 0 1 84461
box 0 0 1 1
use contact_32  contact_32_3573
timestamp 1624857261
transform 1 0 195024 0 1 115605
box 0 0 1 1
use contact_32  contact_32_3572
timestamp 1624857261
transform 1 0 195024 0 1 115333
box 0 0 1 1
use contact_32  contact_32_3571
timestamp 1624857261
transform 1 0 195024 0 1 64333
box 0 0 1 1
use contact_32  contact_32_3570
timestamp 1624857261
transform 1 0 195024 0 1 64605
box 0 0 1 1
use contact_32  contact_32_3569
timestamp 1624857261
transform 1 0 195160 0 1 119277
box 0 0 1 1
use contact_32  contact_32_3568
timestamp 1624857261
transform 1 0 195160 0 1 119549
box 0 0 1 1
use contact_32  contact_32_3567
timestamp 1624857261
transform 1 0 195160 0 1 104181
box 0 0 1 1
use contact_32  contact_32_3566
timestamp 1624857261
transform 1 0 195160 0 1 103909
box 0 0 1 1
use contact_32  contact_32_3565
timestamp 1624857261
transform 1 0 195160 0 1 124717
box 0 0 1 1
use contact_32  contact_32_3564
timestamp 1624857261
transform 1 0 195160 0 1 124445
box 0 0 1 1
use contact_32  contact_32_3563
timestamp 1624857261
transform 1 0 195840 0 1 82149
box 0 0 1 1
use contact_32  contact_32_3562
timestamp 1624857261
transform 1 0 195840 0 1 82421
box 0 0 1 1
use contact_32  contact_32_3561
timestamp 1624857261
transform 1 0 195976 0 1 82013
box 0 0 1 1
use contact_32  contact_32_3560
timestamp 1624857261
transform 1 0 195976 0 1 81741
box 0 0 1 1
use contact_32  contact_32_3559
timestamp 1624857261
transform 1 0 195840 0 1 104181
box 0 0 1 1
use contact_32  contact_32_3558
timestamp 1624857261
transform 1 0 195840 0 1 103909
box 0 0 1 1
use contact_32  contact_32_3557
timestamp 1624857261
transform 1 0 195840 0 1 86773
box 0 0 1 1
use contact_32  contact_32_3556
timestamp 1624857261
transform 1 0 195840 0 1 86501
box 0 0 1 1
use contact_32  contact_32_3555
timestamp 1624857261
transform 1 0 195840 0 1 29925
box 0 0 1 1
use contact_32  contact_32_3554
timestamp 1624857261
transform 1 0 195840 0 1 29653
box 0 0 1 1
use contact_32  contact_32_3553
timestamp 1624857261
transform 1 0 195840 0 1 60661
box 0 0 1 1
use contact_32  contact_32_3552
timestamp 1624857261
transform 1 0 195840 0 1 60389
box 0 0 1 1
use contact_32  contact_32_3551
timestamp 1624857261
transform 1 0 195840 0 1 48829
box 0 0 1 1
use contact_32  contact_32_3550
timestamp 1624857261
transform 1 0 195840 0 1 48557
box 0 0 1 1
use contact_32  contact_32_3549
timestamp 1624857261
transform 1 0 195840 0 1 31421
box 0 0 1 1
use contact_32  contact_32_3548
timestamp 1624857261
transform 1 0 195840 0 1 31149
box 0 0 1 1
use contact_32  contact_32_3547
timestamp 1624857261
transform 1 0 195976 0 1 86365
box 0 0 1 1
use contact_32  contact_32_3546
timestamp 1624857261
transform 1 0 195976 0 1 86093
box 0 0 1 1
use contact_32  contact_32_3545
timestamp 1624857261
transform 1 0 196112 0 1 86365
box 0 0 1 1
use contact_32  contact_32_3544
timestamp 1624857261
transform 1 0 196112 0 1 86093
box 0 0 1 1
use contact_32  contact_32_3543
timestamp 1624857261
transform 1 0 196112 0 1 86501
box 0 0 1 1
use contact_32  contact_32_3542
timestamp 1624857261
transform 1 0 196112 0 1 86773
box 0 0 1 1
use contact_32  contact_32_3541
timestamp 1624857261
transform 1 0 195840 0 1 97789
box 0 0 1 1
use contact_32  contact_32_3540
timestamp 1624857261
transform 1 0 195840 0 1 97517
box 0 0 1 1
use contact_32  contact_32_3539
timestamp 1624857261
transform 1 0 195976 0 1 119685
box 0 0 1 1
use contact_32  contact_32_3538
timestamp 1624857261
transform 1 0 195976 0 1 119957
box 0 0 1 1
use contact_32  contact_32_3537
timestamp 1624857261
transform 1 0 195840 0 1 119549
box 0 0 1 1
use contact_32  contact_32_3536
timestamp 1624857261
transform 1 0 195840 0 1 119277
box 0 0 1 1
use contact_32  contact_32_3535
timestamp 1624857261
transform 1 0 195976 0 1 123221
box 0 0 1 1
use contact_32  contact_32_3534
timestamp 1624857261
transform 1 0 195976 0 1 123493
box 0 0 1 1
use contact_32  contact_32_3533
timestamp 1624857261
transform 1 0 196112 0 1 123221
box 0 0 1 1
use contact_32  contact_32_3532
timestamp 1624857261
transform 1 0 196112 0 1 123493
box 0 0 1 1
use contact_32  contact_32_3531
timestamp 1624857261
transform 1 0 195976 0 1 114517
box 0 0 1 1
use contact_32  contact_32_3530
timestamp 1624857261
transform 1 0 195976 0 1 114789
box 0 0 1 1
use contact_32  contact_32_3529
timestamp 1624857261
transform 1 0 195976 0 1 120093
box 0 0 1 1
use contact_32  contact_32_3528
timestamp 1624857261
transform 1 0 195976 0 1 120365
box 0 0 1 1
use contact_32  contact_32_3527
timestamp 1624857261
transform 1 0 195976 0 1 32645
box 0 0 1 1
use contact_32  contact_32_3526
timestamp 1624857261
transform 1 0 195976 0 1 32373
box 0 0 1 1
use contact_32  contact_32_3525
timestamp 1624857261
transform 1 0 195976 0 1 32781
box 0 0 1 1
use contact_32  contact_32_3524
timestamp 1624857261
transform 1 0 195976 0 1 33053
box 0 0 1 1
use contact_32  contact_32_3523
timestamp 1624857261
transform 1 0 196112 0 1 32781
box 0 0 1 1
use contact_32  contact_32_3522
timestamp 1624857261
transform 1 0 196112 0 1 33053
box 0 0 1 1
use contact_32  contact_32_3521
timestamp 1624857261
transform 1 0 195976 0 1 58077
box 0 0 1 1
use contact_32  contact_32_3520
timestamp 1624857261
transform 1 0 195976 0 1 58349
box 0 0 1 1
use contact_32  contact_32_3519
timestamp 1624857261
transform 1 0 196112 0 1 58077
box 0 0 1 1
use contact_32  contact_32_3518
timestamp 1624857261
transform 1 0 196112 0 1 58349
box 0 0 1 1
use contact_32  contact_32_3517
timestamp 1624857261
transform 1 0 195976 0 1 115741
box 0 0 1 1
use contact_32  contact_32_3516
timestamp 1624857261
transform 1 0 195976 0 1 116013
box 0 0 1 1
use contact_32  contact_32_3515
timestamp 1624857261
transform 1 0 196112 0 1 115741
box 0 0 1 1
use contact_32  contact_32_3514
timestamp 1624857261
transform 1 0 196112 0 1 116013
box 0 0 1 1
use contact_32  contact_32_3513
timestamp 1624857261
transform 1 0 195976 0 1 80925
box 0 0 1 1
use contact_32  contact_32_3512
timestamp 1624857261
transform 1 0 195976 0 1 81197
box 0 0 1 1
use contact_32  contact_32_3511
timestamp 1624857261
transform 1 0 196112 0 1 80925
box 0 0 1 1
use contact_32  contact_32_3510
timestamp 1624857261
transform 1 0 196112 0 1 81197
box 0 0 1 1
use contact_32  contact_32_3509
timestamp 1624857261
transform 1 0 195840 0 1 120501
box 0 0 1 1
use contact_32  contact_32_3508
timestamp 1624857261
transform 1 0 195840 0 1 120773
box 0 0 1 1
use contact_32  contact_32_3507
timestamp 1624857261
transform 1 0 195840 0 1 83645
box 0 0 1 1
use contact_32  contact_32_3506
timestamp 1624857261
transform 1 0 195840 0 1 83373
box 0 0 1 1
use contact_32  contact_32_3505
timestamp 1624857261
transform 1 0 195976 0 1 52501
box 0 0 1 1
use contact_32  contact_32_3504
timestamp 1624857261
transform 1 0 195976 0 1 52773
box 0 0 1 1
use contact_32  contact_32_3503
timestamp 1624857261
transform 1 0 196112 0 1 52501
box 0 0 1 1
use contact_32  contact_32_3502
timestamp 1624857261
transform 1 0 196112 0 1 52773
box 0 0 1 1
use contact_32  contact_32_3501
timestamp 1624857261
transform 1 0 195976 0 1 89085
box 0 0 1 1
use contact_32  contact_32_3500
timestamp 1624857261
transform 1 0 195976 0 1 88813
box 0 0 1 1
use contact_32  contact_32_3499
timestamp 1624857261
transform 1 0 195840 0 1 53181
box 0 0 1 1
use contact_32  contact_32_3498
timestamp 1624857261
transform 1 0 195840 0 1 52909
box 0 0 1 1
use contact_32  contact_32_3497
timestamp 1624857261
transform 1 0 195840 0 1 57125
box 0 0 1 1
use contact_32  contact_32_3496
timestamp 1624857261
transform 1 0 195840 0 1 56853
box 0 0 1 1
use contact_32  contact_32_3495
timestamp 1624857261
transform 1 0 195840 0 1 119141
box 0 0 1 1
use contact_32  contact_32_3494
timestamp 1624857261
transform 1 0 195840 0 1 118869
box 0 0 1 1
use contact_32  contact_32_3493
timestamp 1624857261
transform 1 0 195976 0 1 113293
box 0 0 1 1
use contact_32  contact_32_3492
timestamp 1624857261
transform 1 0 195976 0 1 113565
box 0 0 1 1
use contact_32  contact_32_3491
timestamp 1624857261
transform 1 0 196112 0 1 113293
box 0 0 1 1
use contact_32  contact_32_3490
timestamp 1624857261
transform 1 0 196112 0 1 113565
box 0 0 1 1
use contact_32  contact_32_3489
timestamp 1624857261
transform 1 0 195840 0 1 29109
box 0 0 1 1
use contact_32  contact_32_3488
timestamp 1624857261
transform 1 0 195840 0 1 28837
box 0 0 1 1
use contact_32  contact_32_3487
timestamp 1624857261
transform 1 0 195840 0 1 29245
box 0 0 1 1
use contact_32  contact_32_3486
timestamp 1624857261
transform 1 0 195840 0 1 29517
box 0 0 1 1
use contact_32  contact_32_3485
timestamp 1624857261
transform 1 0 195976 0 1 107037
box 0 0 1 1
use contact_32  contact_32_3484
timestamp 1624857261
transform 1 0 195976 0 1 107309
box 0 0 1 1
use contact_32  contact_32_3483
timestamp 1624857261
transform 1 0 196112 0 1 106901
box 0 0 1 1
use contact_32  contact_32_3482
timestamp 1624857261
transform 1 0 196112 0 1 106629
box 0 0 1 1
use contact_32  contact_32_3481
timestamp 1624857261
transform 1 0 195976 0 1 89629
box 0 0 1 1
use contact_32  contact_32_3480
timestamp 1624857261
transform 1 0 195976 0 1 89901
box 0 0 1 1
use contact_32  contact_32_3479
timestamp 1624857261
transform 1 0 196112 0 1 89629
box 0 0 1 1
use contact_32  contact_32_3478
timestamp 1624857261
transform 1 0 196112 0 1 89901
box 0 0 1 1
use contact_32  contact_32_3477
timestamp 1624857261
transform 1 0 195976 0 1 124445
box 0 0 1 1
use contact_32  contact_32_3476
timestamp 1624857261
transform 1 0 195976 0 1 124717
box 0 0 1 1
use contact_32  contact_32_3475
timestamp 1624857261
transform 1 0 195976 0 1 124309
box 0 0 1 1
use contact_32  contact_32_3474
timestamp 1624857261
transform 1 0 195976 0 1 124037
box 0 0 1 1
use contact_32  contact_32_3473
timestamp 1624857261
transform 1 0 196112 0 1 124309
box 0 0 1 1
use contact_32  contact_32_3472
timestamp 1624857261
transform 1 0 196112 0 1 124037
box 0 0 1 1
use contact_32  contact_32_3471
timestamp 1624857261
transform 1 0 196112 0 1 124445
box 0 0 1 1
use contact_32  contact_32_3470
timestamp 1624857261
transform 1 0 196112 0 1 124717
box 0 0 1 1
use contact_32  contact_32_3469
timestamp 1624857261
transform 1 0 195976 0 1 63517
box 0 0 1 1
use contact_32  contact_32_3468
timestamp 1624857261
transform 1 0 195976 0 1 63789
box 0 0 1 1
use contact_32  contact_32_3467
timestamp 1624857261
transform 1 0 195840 0 1 106221
box 0 0 1 1
use contact_32  contact_32_3466
timestamp 1624857261
transform 1 0 195840 0 1 106493
box 0 0 1 1
use contact_32  contact_32_3465
timestamp 1624857261
transform 1 0 196112 0 1 121997
box 0 0 1 1
use contact_32  contact_32_3464
timestamp 1624857261
transform 1 0 196112 0 1 122269
box 0 0 1 1
use contact_32  contact_32_3463
timestamp 1624857261
transform 1 0 195976 0 1 61205
box 0 0 1 1
use contact_32  contact_32_3462
timestamp 1624857261
transform 1 0 195976 0 1 61477
box 0 0 1 1
use contact_32  contact_32_3461
timestamp 1624857261
transform 1 0 196112 0 1 61069
box 0 0 1 1
use contact_32  contact_32_3460
timestamp 1624857261
transform 1 0 196112 0 1 60797
box 0 0 1 1
use contact_32  contact_32_3459
timestamp 1624857261
transform 1 0 195976 0 1 94797
box 0 0 1 1
use contact_32  contact_32_3458
timestamp 1624857261
transform 1 0 195976 0 1 95069
box 0 0 1 1
use contact_32  contact_32_3457
timestamp 1624857261
transform 1 0 196112 0 1 94661
box 0 0 1 1
use contact_32  contact_32_3456
timestamp 1624857261
transform 1 0 196112 0 1 94389
box 0 0 1 1
use contact_32  contact_32_3455
timestamp 1624857261
transform 1 0 195840 0 1 103093
box 0 0 1 1
use contact_32  contact_32_3454
timestamp 1624857261
transform 1 0 195840 0 1 103365
box 0 0 1 1
use contact_32  contact_32_3453
timestamp 1624857261
transform 1 0 196112 0 1 109621
box 0 0 1 1
use contact_32  contact_32_3452
timestamp 1624857261
transform 1 0 196112 0 1 109349
box 0 0 1 1
use contact_32  contact_32_3451
timestamp 1624857261
transform 1 0 195840 0 1 84325
box 0 0 1 1
use contact_32  contact_32_3450
timestamp 1624857261
transform 1 0 195840 0 1 84053
box 0 0 1 1
use contact_32  contact_32_3449
timestamp 1624857261
transform 1 0 195840 0 1 41077
box 0 0 1 1
use contact_32  contact_32_3448
timestamp 1624857261
transform 1 0 195840 0 1 41349
box 0 0 1 1
use contact_32  contact_32_3447
timestamp 1624857261
transform 1 0 195840 0 1 91125
box 0 0 1 1
use contact_32  contact_32_3446
timestamp 1624857261
transform 1 0 195840 0 1 90853
box 0 0 1 1
use contact_32  contact_32_3445
timestamp 1624857261
transform 1 0 195840 0 1 51957
box 0 0 1 1
use contact_32  contact_32_3444
timestamp 1624857261
transform 1 0 195840 0 1 51685
box 0 0 1 1
use contact_32  contact_32_3443
timestamp 1624857261
transform 1 0 195840 0 1 78069
box 0 0 1 1
use contact_32  contact_32_3442
timestamp 1624857261
transform 1 0 195840 0 1 77797
box 0 0 1 1
use contact_32  contact_32_3441
timestamp 1624857261
transform 1 0 195840 0 1 78205
box 0 0 1 1
use contact_32  contact_32_3440
timestamp 1624857261
transform 1 0 195840 0 1 78477
box 0 0 1 1
use contact_32  contact_32_3439
timestamp 1624857261
transform 1 0 196112 0 1 31965
box 0 0 1 1
use contact_32  contact_32_3438
timestamp 1624857261
transform 1 0 196112 0 1 32237
box 0 0 1 1
use contact_32  contact_32_3437
timestamp 1624857261
transform 1 0 195840 0 1 69365
box 0 0 1 1
use contact_32  contact_32_3436
timestamp 1624857261
transform 1 0 195840 0 1 69093
box 0 0 1 1
use contact_32  contact_32_3435
timestamp 1624857261
transform 1 0 195976 0 1 85277
box 0 0 1 1
use contact_32  contact_32_3434
timestamp 1624857261
transform 1 0 195976 0 1 85549
box 0 0 1 1
use contact_32  contact_32_3433
timestamp 1624857261
transform 1 0 195840 0 1 73445
box 0 0 1 1
use contact_32  contact_32_3432
timestamp 1624857261
transform 1 0 195840 0 1 73717
box 0 0 1 1
use contact_32  contact_32_3431
timestamp 1624857261
transform 1 0 195976 0 1 73309
box 0 0 1 1
use contact_32  contact_32_3430
timestamp 1624857261
transform 1 0 195976 0 1 73037
box 0 0 1 1
use contact_32  contact_32_3429
timestamp 1624857261
transform 1 0 195840 0 1 122677
box 0 0 1 1
use contact_32  contact_32_3428
timestamp 1624857261
transform 1 0 195840 0 1 122405
box 0 0 1 1
use contact_32  contact_32_3427
timestamp 1624857261
transform 1 0 196112 0 1 63109
box 0 0 1 1
use contact_32  contact_32_3426
timestamp 1624857261
transform 1 0 196112 0 1 62837
box 0 0 1 1
use contact_32  contact_32_3425
timestamp 1624857261
transform 1 0 195976 0 1 59165
box 0 0 1 1
use contact_32  contact_32_3424
timestamp 1624857261
transform 1 0 195976 0 1 58893
box 0 0 1 1
use contact_32  contact_32_3423
timestamp 1624857261
transform 1 0 195976 0 1 55901
box 0 0 1 1
use contact_32  contact_32_3422
timestamp 1624857261
transform 1 0 195976 0 1 55629
box 0 0 1 1
use contact_32  contact_32_3421
timestamp 1624857261
transform 1 0 196112 0 1 55901
box 0 0 1 1
use contact_32  contact_32_3420
timestamp 1624857261
transform 1 0 196112 0 1 55629
box 0 0 1 1
use contact_32  contact_32_3419
timestamp 1624857261
transform 1 0 195976 0 1 93845
box 0 0 1 1
use contact_32  contact_32_3418
timestamp 1624857261
transform 1 0 195976 0 1 93573
box 0 0 1 1
use contact_32  contact_32_3417
timestamp 1624857261
transform 1 0 195976 0 1 93981
box 0 0 1 1
use contact_32  contact_32_3416
timestamp 1624857261
transform 1 0 195976 0 1 94253
box 0 0 1 1
use contact_32  contact_32_3415
timestamp 1624857261
transform 1 0 196112 0 1 93981
box 0 0 1 1
use contact_32  contact_32_3414
timestamp 1624857261
transform 1 0 196112 0 1 94253
box 0 0 1 1
use contact_32  contact_32_3413
timestamp 1624857261
transform 1 0 195840 0 1 101733
box 0 0 1 1
use contact_32  contact_32_3412
timestamp 1624857261
transform 1 0 195840 0 1 101461
box 0 0 1 1
use contact_32  contact_32_3411
timestamp 1624857261
transform 1 0 195976 0 1 27613
box 0 0 1 1
use contact_32  contact_32_3410
timestamp 1624857261
transform 1 0 195976 0 1 27885
box 0 0 1 1
use contact_32  contact_32_3409
timestamp 1624857261
transform 1 0 195976 0 1 69909
box 0 0 1 1
use contact_32  contact_32_3408
timestamp 1624857261
transform 1 0 195976 0 1 70181
box 0 0 1 1
use contact_32  contact_32_3407
timestamp 1624857261
transform 1 0 196112 0 1 69909
box 0 0 1 1
use contact_32  contact_32_3406
timestamp 1624857261
transform 1 0 196112 0 1 70181
box 0 0 1 1
use contact_32  contact_32_3405
timestamp 1624857261
transform 1 0 196112 0 1 69093
box 0 0 1 1
use contact_32  contact_32_3404
timestamp 1624857261
transform 1 0 196112 0 1 69365
box 0 0 1 1
use contact_32  contact_32_3403
timestamp 1624857261
transform 1 0 195840 0 1 76437
box 0 0 1 1
use contact_32  contact_32_3402
timestamp 1624857261
transform 1 0 195840 0 1 76165
box 0 0 1 1
use contact_32  contact_32_3401
timestamp 1624857261
transform 1 0 196112 0 1 76437
box 0 0 1 1
use contact_32  contact_32_3400
timestamp 1624857261
transform 1 0 196112 0 1 76165
box 0 0 1 1
use contact_32  contact_32_3399
timestamp 1624857261
transform 1 0 195840 0 1 78885
box 0 0 1 1
use contact_32  contact_32_3398
timestamp 1624857261
transform 1 0 195840 0 1 78613
box 0 0 1 1
use contact_32  contact_32_3397
timestamp 1624857261
transform 1 0 195840 0 1 48421
box 0 0 1 1
use contact_32  contact_32_3396
timestamp 1624857261
transform 1 0 195840 0 1 48149
box 0 0 1 1
use contact_32  contact_32_3395
timestamp 1624857261
transform 1 0 196112 0 1 84053
box 0 0 1 1
use contact_32  contact_32_3394
timestamp 1624857261
transform 1 0 196112 0 1 84325
box 0 0 1 1
use contact_32  contact_32_3393
timestamp 1624857261
transform 1 0 195840 0 1 118325
box 0 0 1 1
use contact_32  contact_32_3392
timestamp 1624857261
transform 1 0 195840 0 1 118053
box 0 0 1 1
use contact_32  contact_32_3391
timestamp 1624857261
transform 1 0 195840 0 1 118461
box 0 0 1 1
use contact_32  contact_32_3390
timestamp 1624857261
transform 1 0 195840 0 1 118733
box 0 0 1 1
use contact_32  contact_32_3389
timestamp 1624857261
transform 1 0 195976 0 1 64333
box 0 0 1 1
use contact_32  contact_32_3388
timestamp 1624857261
transform 1 0 195976 0 1 64605
box 0 0 1 1
use contact_32  contact_32_3387
timestamp 1624857261
transform 1 0 195840 0 1 104997
box 0 0 1 1
use contact_32  contact_32_3386
timestamp 1624857261
transform 1 0 195840 0 1 104725
box 0 0 1 1
use contact_32  contact_32_3385
timestamp 1624857261
transform 1 0 195840 0 1 85685
box 0 0 1 1
use contact_32  contact_32_3384
timestamp 1624857261
transform 1 0 195840 0 1 85957
box 0 0 1 1
use contact_32  contact_32_3383
timestamp 1624857261
transform 1 0 195976 0 1 35093
box 0 0 1 1
use contact_32  contact_32_3382
timestamp 1624857261
transform 1 0 195976 0 1 35365
box 0 0 1 1
use contact_32  contact_32_3381
timestamp 1624857261
transform 1 0 196112 0 1 35093
box 0 0 1 1
use contact_32  contact_32_3380
timestamp 1624857261
transform 1 0 196112 0 1 35365
box 0 0 1 1
use contact_32  contact_32_3379
timestamp 1624857261
transform 1 0 195976 0 1 50189
box 0 0 1 1
use contact_32  contact_32_3378
timestamp 1624857261
transform 1 0 195976 0 1 50461
box 0 0 1 1
use contact_32  contact_32_3377
timestamp 1624857261
transform 1 0 195840 0 1 38629
box 0 0 1 1
use contact_32  contact_32_3376
timestamp 1624857261
transform 1 0 195840 0 1 38357
box 0 0 1 1
use contact_32  contact_32_3375
timestamp 1624857261
transform 1 0 195840 0 1 90037
box 0 0 1 1
use contact_32  contact_32_3374
timestamp 1624857261
transform 1 0 195840 0 1 90309
box 0 0 1 1
use contact_32  contact_32_3373
timestamp 1624857261
transform 1 0 196112 0 1 48149
box 0 0 1 1
use contact_32  contact_32_3372
timestamp 1624857261
transform 1 0 196112 0 1 48421
box 0 0 1 1
use contact_32  contact_32_3371
timestamp 1624857261
transform 1 0 196112 0 1 121589
box 0 0 1 1
use contact_32  contact_32_3370
timestamp 1624857261
transform 1 0 196112 0 1 121317
box 0 0 1 1
use contact_32  contact_32_3369
timestamp 1624857261
transform 1 0 195840 0 1 39853
box 0 0 1 1
use contact_32  contact_32_3368
timestamp 1624857261
transform 1 0 195840 0 1 40125
box 0 0 1 1
use contact_32  contact_32_3367
timestamp 1624857261
transform 1 0 195840 0 1 64741
box 0 0 1 1
use contact_32  contact_32_3366
timestamp 1624857261
transform 1 0 195840 0 1 65013
box 0 0 1 1
use contact_32  contact_32_3365
timestamp 1624857261
transform 1 0 196112 0 1 64741
box 0 0 1 1
use contact_32  contact_32_3364
timestamp 1624857261
transform 1 0 196112 0 1 65013
box 0 0 1 1
use contact_32  contact_32_3363
timestamp 1624857261
transform 1 0 195976 0 1 112613
box 0 0 1 1
use contact_32  contact_32_3362
timestamp 1624857261
transform 1 0 195976 0 1 112885
box 0 0 1 1
use contact_32  contact_32_3361
timestamp 1624857261
transform 1 0 196112 0 1 57533
box 0 0 1 1
use contact_32  contact_32_3360
timestamp 1624857261
transform 1 0 196112 0 1 57261
box 0 0 1 1
use contact_32  contact_32_3359
timestamp 1624857261
transform 1 0 195840 0 1 49645
box 0 0 1 1
use contact_32  contact_32_3358
timestamp 1624857261
transform 1 0 195840 0 1 49373
box 0 0 1 1
use contact_32  contact_32_3357
timestamp 1624857261
transform 1 0 195976 0 1 43797
box 0 0 1 1
use contact_32  contact_32_3356
timestamp 1624857261
transform 1 0 195976 0 1 44069
box 0 0 1 1
use contact_32  contact_32_3355
timestamp 1624857261
transform 1 0 195840 0 1 45293
box 0 0 1 1
use contact_32  contact_32_3354
timestamp 1624857261
transform 1 0 195840 0 1 45021
box 0 0 1 1
use contact_32  contact_32_3353
timestamp 1624857261
transform 1 0 195840 0 1 45429
box 0 0 1 1
use contact_32  contact_32_3352
timestamp 1624857261
transform 1 0 195840 0 1 45701
box 0 0 1 1
use contact_32  contact_32_3351
timestamp 1624857261
transform 1 0 195976 0 1 77661
box 0 0 1 1
use contact_32  contact_32_3350
timestamp 1624857261
transform 1 0 195976 0 1 77389
box 0 0 1 1
use contact_32  contact_32_3349
timestamp 1624857261
transform 1 0 195976 0 1 96021
box 0 0 1 1
use contact_32  contact_32_3348
timestamp 1624857261
transform 1 0 195976 0 1 96293
box 0 0 1 1
use contact_32  contact_32_3347
timestamp 1624857261
transform 1 0 196112 0 1 96021
box 0 0 1 1
use contact_32  contact_32_3346
timestamp 1624857261
transform 1 0 196112 0 1 96293
box 0 0 1 1
use contact_32  contact_32_3345
timestamp 1624857261
transform 1 0 195976 0 1 111389
box 0 0 1 1
use contact_32  contact_32_3344
timestamp 1624857261
transform 1 0 195976 0 1 111661
box 0 0 1 1
use contact_32  contact_32_3343
timestamp 1624857261
transform 1 0 195840 0 1 100917
box 0 0 1 1
use contact_32  contact_32_3342
timestamp 1624857261
transform 1 0 195840 0 1 100645
box 0 0 1 1
use contact_32  contact_32_3341
timestamp 1624857261
transform 1 0 196112 0 1 90445
box 0 0 1 1
use contact_32  contact_32_3340
timestamp 1624857261
transform 1 0 196112 0 1 90717
box 0 0 1 1
use contact_32  contact_32_3339
timestamp 1624857261
transform 1 0 195976 0 1 87317
box 0 0 1 1
use contact_32  contact_32_3338
timestamp 1624857261
transform 1 0 195976 0 1 87589
box 0 0 1 1
use contact_32  contact_32_3337
timestamp 1624857261
transform 1 0 195976 0 1 80381
box 0 0 1 1
use contact_32  contact_32_3336
timestamp 1624857261
transform 1 0 195976 0 1 80109
box 0 0 1 1
use contact_32  contact_32_3335
timestamp 1624857261
transform 1 0 195840 0 1 99965
box 0 0 1 1
use contact_32  contact_32_3334
timestamp 1624857261
transform 1 0 195840 0 1 100237
box 0 0 1 1
use contact_32  contact_32_3333
timestamp 1624857261
transform 1 0 196112 0 1 92349
box 0 0 1 1
use contact_32  contact_32_3332
timestamp 1624857261
transform 1 0 196112 0 1 92077
box 0 0 1 1
use contact_32  contact_32_3331
timestamp 1624857261
transform 1 0 195840 0 1 116557
box 0 0 1 1
use contact_32  contact_32_3330
timestamp 1624857261
transform 1 0 195840 0 1 116829
box 0 0 1 1
use contact_32  contact_32_3329
timestamp 1624857261
transform 1 0 196112 0 1 116557
box 0 0 1 1
use contact_32  contact_32_3328
timestamp 1624857261
transform 1 0 196112 0 1 116829
box 0 0 1 1
use contact_32  contact_32_3327
timestamp 1624857261
transform 1 0 195840 0 1 115197
box 0 0 1 1
use contact_32  contact_32_3326
timestamp 1624857261
transform 1 0 195840 0 1 114925
box 0 0 1 1
use contact_32  contact_32_3325
timestamp 1624857261
transform 1 0 195976 0 1 102549
box 0 0 1 1
use contact_32  contact_32_3324
timestamp 1624857261
transform 1 0 195976 0 1 102277
box 0 0 1 1
use contact_32  contact_32_3323
timestamp 1624857261
transform 1 0 195840 0 1 74533
box 0 0 1 1
use contact_32  contact_32_3322
timestamp 1624857261
transform 1 0 195840 0 1 74261
box 0 0 1 1
use contact_32  contact_32_3321
timestamp 1624857261
transform 1 0 196112 0 1 107853
box 0 0 1 1
use contact_32  contact_32_3320
timestamp 1624857261
transform 1 0 196112 0 1 108125
box 0 0 1 1
use contact_32  contact_32_3319
timestamp 1624857261
transform 1 0 196112 0 1 33461
box 0 0 1 1
use contact_32  contact_32_3318
timestamp 1624857261
transform 1 0 196112 0 1 33189
box 0 0 1 1
use contact_32  contact_32_3317
timestamp 1624857261
transform 1 0 195840 0 1 76981
box 0 0 1 1
use contact_32  contact_32_3316
timestamp 1624857261
transform 1 0 195840 0 1 77253
box 0 0 1 1
use contact_32  contact_32_3315
timestamp 1624857261
transform 1 0 195840 0 1 34685
box 0 0 1 1
use contact_32  contact_32_3314
timestamp 1624857261
transform 1 0 195840 0 1 34413
box 0 0 1 1
use contact_32  contact_32_3313
timestamp 1624857261
transform 1 0 195840 0 1 54133
box 0 0 1 1
use contact_32  contact_32_3312
timestamp 1624857261
transform 1 0 195840 0 1 54405
box 0 0 1 1
use contact_32  contact_32_3311
timestamp 1624857261
transform 1 0 196112 0 1 72221
box 0 0 1 1
use contact_32  contact_32_3310
timestamp 1624857261
transform 1 0 196112 0 1 72493
box 0 0 1 1
use contact_32  contact_32_3309
timestamp 1624857261
transform 1 0 196112 0 1 102141
box 0 0 1 1
use contact_32  contact_32_3308
timestamp 1624857261
transform 1 0 196112 0 1 101869
box 0 0 1 1
use contact_32  contact_32_3307
timestamp 1624857261
transform 1 0 195840 0 1 66237
box 0 0 1 1
use contact_32  contact_32_3306
timestamp 1624857261
transform 1 0 195840 0 1 65965
box 0 0 1 1
use contact_32  contact_32_3305
timestamp 1624857261
transform 1 0 196112 0 1 99013
box 0 0 1 1
use contact_32  contact_32_3304
timestamp 1624857261
transform 1 0 196112 0 1 98741
box 0 0 1 1
use contact_32  contact_32_3303
timestamp 1624857261
transform 1 0 196112 0 1 56853
box 0 0 1 1
use contact_32  contact_32_3302
timestamp 1624857261
transform 1 0 196112 0 1 57125
box 0 0 1 1
use contact_32  contact_32_3301
timestamp 1624857261
transform 1 0 196112 0 1 70589
box 0 0 1 1
use contact_32  contact_32_3300
timestamp 1624857261
transform 1 0 196112 0 1 70317
box 0 0 1 1
use contact_32  contact_32_3299
timestamp 1624857261
transform 1 0 196112 0 1 104725
box 0 0 1 1
use contact_32  contact_32_3298
timestamp 1624857261
transform 1 0 196112 0 1 104997
box 0 0 1 1
use contact_32  contact_32_3297
timestamp 1624857261
transform 1 0 195840 0 1 110437
box 0 0 1 1
use contact_32  contact_32_3296
timestamp 1624857261
transform 1 0 195840 0 1 110165
box 0 0 1 1
use contact_32  contact_32_3295
timestamp 1624857261
transform 1 0 195840 0 1 117237
box 0 0 1 1
use contact_32  contact_32_3294
timestamp 1624857261
transform 1 0 195840 0 1 117509
box 0 0 1 1
use contact_32  contact_32_3293
timestamp 1624857261
transform 1 0 195976 0 1 98333
box 0 0 1 1
use contact_32  contact_32_3292
timestamp 1624857261
transform 1 0 195976 0 1 98605
box 0 0 1 1
use contact_32  contact_32_3291
timestamp 1624857261
transform 1 0 196112 0 1 78613
box 0 0 1 1
use contact_32  contact_32_3290
timestamp 1624857261
transform 1 0 196112 0 1 78885
box 0 0 1 1
use contact_32  contact_32_3289
timestamp 1624857261
transform 1 0 196112 0 1 108669
box 0 0 1 1
use contact_32  contact_32_3288
timestamp 1624857261
transform 1 0 196112 0 1 108941
box 0 0 1 1
use contact_32  contact_32_3287
timestamp 1624857261
transform 1 0 196112 0 1 118053
box 0 0 1 1
use contact_32  contact_32_3286
timestamp 1624857261
transform 1 0 196112 0 1 118325
box 0 0 1 1
use contact_32  contact_32_3285
timestamp 1624857261
transform 1 0 195976 0 1 82965
box 0 0 1 1
use contact_32  contact_32_3284
timestamp 1624857261
transform 1 0 195976 0 1 83237
box 0 0 1 1
use contact_32  contact_32_3283
timestamp 1624857261
transform 1 0 195976 0 1 62021
box 0 0 1 1
use contact_32  contact_32_3282
timestamp 1624857261
transform 1 0 195976 0 1 62293
box 0 0 1 1
use contact_32  contact_32_3281
timestamp 1624857261
transform 1 0 196112 0 1 61885
box 0 0 1 1
use contact_32  contact_32_3280
timestamp 1624857261
transform 1 0 196112 0 1 61613
box 0 0 1 1
use contact_32  contact_32_3279
timestamp 1624857261
transform 1 0 196112 0 1 45021
box 0 0 1 1
use contact_32  contact_32_3278
timestamp 1624857261
transform 1 0 196112 0 1 45293
box 0 0 1 1
use contact_32  contact_32_3277
timestamp 1624857261
transform 1 0 195976 0 1 51277
box 0 0 1 1
use contact_32  contact_32_3276
timestamp 1624857261
transform 1 0 195976 0 1 51005
box 0 0 1 1
use contact_32  contact_32_3275
timestamp 1624857261
transform 1 0 196112 0 1 118869
box 0 0 1 1
use contact_32  contact_32_3274
timestamp 1624857261
transform 1 0 196112 0 1 119141
box 0 0 1 1
use contact_32  contact_32_3273
timestamp 1624857261
transform 1 0 196112 0 1 75485
box 0 0 1 1
use contact_32  contact_32_3272
timestamp 1624857261
transform 1 0 196112 0 1 75757
box 0 0 1 1
use contact_32  contact_32_3271
timestamp 1624857261
transform 1 0 196112 0 1 81605
box 0 0 1 1
use contact_32  contact_32_3270
timestamp 1624857261
transform 1 0 196112 0 1 81333
box 0 0 1 1
use contact_32  contact_32_3269
timestamp 1624857261
transform 1 0 195976 0 1 65557
box 0 0 1 1
use contact_32  contact_32_3268
timestamp 1624857261
transform 1 0 195976 0 1 65829
box 0 0 1 1
use contact_32  contact_32_3267
timestamp 1624857261
transform 1 0 196112 0 1 65557
box 0 0 1 1
use contact_32  contact_32_3266
timestamp 1624857261
transform 1 0 196112 0 1 65829
box 0 0 1 1
use contact_32  contact_32_3265
timestamp 1624857261
transform 1 0 196112 0 1 73037
box 0 0 1 1
use contact_32  contact_32_3264
timestamp 1624857261
transform 1 0 196112 0 1 73309
box 0 0 1 1
use contact_32  contact_32_3263
timestamp 1624857261
transform 1 0 196112 0 1 88405
box 0 0 1 1
use contact_32  contact_32_3262
timestamp 1624857261
transform 1 0 196112 0 1 88133
box 0 0 1 1
use contact_32  contact_32_3261
timestamp 1624857261
transform 1 0 196112 0 1 55221
box 0 0 1 1
use contact_32  contact_32_3260
timestamp 1624857261
transform 1 0 196112 0 1 54949
box 0 0 1 1
use contact_32  contact_32_3259
timestamp 1624857261
transform 1 0 196112 0 1 74125
box 0 0 1 1
use contact_32  contact_32_3258
timestamp 1624857261
transform 1 0 196112 0 1 73853
box 0 0 1 1
use contact_32  contact_32_3257
timestamp 1624857261
transform 1 0 196112 0 1 95477
box 0 0 1 1
use contact_32  contact_32_3256
timestamp 1624857261
transform 1 0 196112 0 1 95205
box 0 0 1 1
use contact_32  contact_32_3255
timestamp 1624857261
transform 1 0 196112 0 1 95613
box 0 0 1 1
use contact_32  contact_32_3254
timestamp 1624857261
transform 1 0 196248 0 1 95749
box 0 0 1 1
use contact_32  contact_32_3253
timestamp 1624857261
transform 1 0 196112 0 1 108261
box 0 0 1 1
use contact_32  contact_32_3252
timestamp 1624857261
transform 1 0 196248 0 1 108397
box 0 0 1 1
use contact_32  contact_32_3251
timestamp 1624857261
transform 1 0 195840 0 1 68277
box 0 0 1 1
use contact_32  contact_32_3250
timestamp 1624857261
transform 1 0 195840 0 1 68549
box 0 0 1 1
use contact_32  contact_32_3249
timestamp 1624857261
transform 1 0 196384 0 1 28293
box 0 0 1 1
use contact_32  contact_32_3248
timestamp 1624857261
transform 1 0 196384 0 1 28021
box 0 0 1 1
use contact_32  contact_32_3247
timestamp 1624857261
transform 1 0 196384 0 1 33189
box 0 0 1 1
use contact_32  contact_32_3246
timestamp 1624857261
transform 1 0 196384 0 1 33461
box 0 0 1 1
use contact_32  contact_32_3245
timestamp 1624857261
transform 1 0 196384 0 1 79701
box 0 0 1 1
use contact_32  contact_32_3244
timestamp 1624857261
transform 1 0 196384 0 1 79429
box 0 0 1 1
use contact_32  contact_32_3243
timestamp 1624857261
transform 1 0 196248 0 1 82557
box 0 0 1 1
use contact_32  contact_32_3242
timestamp 1624857261
transform 1 0 196248 0 1 82829
box 0 0 1 1
use contact_32  contact_32_3241
timestamp 1624857261
transform 1 0 196248 0 1 82421
box 0 0 1 1
use contact_32  contact_32_3240
timestamp 1624857261
transform 1 0 196248 0 1 82149
box 0 0 1 1
use contact_32  contact_32_3239
timestamp 1624857261
transform 1 0 196384 0 1 40533
box 0 0 1 1
use contact_32  contact_32_3238
timestamp 1624857261
transform 1 0 196384 0 1 40261
box 0 0 1 1
use contact_32  contact_32_3237
timestamp 1624857261
transform 1 0 196384 0 1 54405
box 0 0 1 1
use contact_32  contact_32_3236
timestamp 1624857261
transform 1 0 196384 0 1 54133
box 0 0 1 1
use contact_32  contact_32_3235
timestamp 1624857261
transform 1 0 196248 0 1 48557
box 0 0 1 1
use contact_32  contact_32_3234
timestamp 1624857261
transform 1 0 196248 0 1 48829
box 0 0 1 1
use contact_32  contact_32_3233
timestamp 1624857261
transform 1 0 196384 0 1 42301
box 0 0 1 1
use contact_32  contact_32_3232
timestamp 1624857261
transform 1 0 196384 0 1 42573
box 0 0 1 1
use contact_32  contact_32_3231
timestamp 1624857261
transform 1 0 196248 0 1 115197
box 0 0 1 1
use contact_32  contact_32_3230
timestamp 1624857261
transform 1 0 196248 0 1 114925
box 0 0 1 1
use contact_32  contact_32_3229
timestamp 1624857261
transform 1 0 196384 0 1 115333
box 0 0 1 1
use contact_32  contact_32_3228
timestamp 1624857261
transform 1 0 196384 0 1 115605
box 0 0 1 1
use contact_32  contact_32_3227
timestamp 1624857261
transform 1 0 196248 0 1 123629
box 0 0 1 1
use contact_32  contact_32_3226
timestamp 1624857261
transform 1 0 196248 0 1 123901
box 0 0 1 1
use contact_32  contact_32_3225
timestamp 1624857261
transform 1 0 196248 0 1 25981
box 0 0 1 1
use contact_32  contact_32_3224
timestamp 1624857261
transform 1 0 196248 0 1 25709
box 0 0 1 1
use contact_32  contact_32_3223
timestamp 1624857261
transform 1 0 196384 0 1 53589
box 0 0 1 1
use contact_32  contact_32_3222
timestamp 1624857261
transform 1 0 196384 0 1 53317
box 0 0 1 1
use contact_32  contact_32_3221
timestamp 1624857261
transform 1 0 196248 0 1 119277
box 0 0 1 1
use contact_32  contact_32_3220
timestamp 1624857261
transform 1 0 196248 0 1 119549
box 0 0 1 1
use contact_32  contact_32_3219
timestamp 1624857261
transform 1 0 196248 0 1 46517
box 0 0 1 1
use contact_32  contact_32_3218
timestamp 1624857261
transform 1 0 196248 0 1 46245
box 0 0 1 1
use contact_32  contact_32_3217
timestamp 1624857261
transform 1 0 196384 0 1 33869
box 0 0 1 1
use contact_32  contact_32_3216
timestamp 1624857261
transform 1 0 196384 0 1 33597
box 0 0 1 1
use contact_32  contact_32_3215
timestamp 1624857261
transform 1 0 196384 0 1 98197
box 0 0 1 1
use contact_32  contact_32_3214
timestamp 1624857261
transform 1 0 196384 0 1 97925
box 0 0 1 1
use contact_32  contact_32_3213
timestamp 1624857261
transform 1 0 196384 0 1 43253
box 0 0 1 1
use contact_32  contact_32_3212
timestamp 1624857261
transform 1 0 196384 0 1 42981
box 0 0 1 1
use contact_32  contact_32_3211
timestamp 1624857261
transform 1 0 196384 0 1 50053
box 0 0 1 1
use contact_32  contact_32_3210
timestamp 1624857261
transform 1 0 196384 0 1 49781
box 0 0 1 1
use contact_32  contact_32_3209
timestamp 1624857261
transform 1 0 196384 0 1 114381
box 0 0 1 1
use contact_32  contact_32_3208
timestamp 1624857261
transform 1 0 196384 0 1 114109
box 0 0 1 1
use contact_32  contact_32_3207
timestamp 1624857261
transform 1 0 196248 0 1 28837
box 0 0 1 1
use contact_32  contact_32_3206
timestamp 1624857261
transform 1 0 196248 0 1 29109
box 0 0 1 1
use contact_32  contact_32_3205
timestamp 1624857261
transform 1 0 196384 0 1 52501
box 0 0 1 1
use contact_32  contact_32_3204
timestamp 1624857261
transform 1 0 196384 0 1 52773
box 0 0 1 1
use contact_32  contact_32_3203
timestamp 1624857261
transform 1 0 196248 0 1 37541
box 0 0 1 1
use contact_32  contact_32_3202
timestamp 1624857261
transform 1 0 196248 0 1 37813
box 0 0 1 1
use contact_32  contact_32_3201
timestamp 1624857261
transform 1 0 196248 0 1 69501
box 0 0 1 1
use contact_32  contact_32_3200
timestamp 1624857261
transform 1 0 196248 0 1 69773
box 0 0 1 1
use contact_32  contact_32_3199
timestamp 1624857261
transform 1 0 196248 0 1 86909
box 0 0 1 1
use contact_32  contact_32_3198
timestamp 1624857261
transform 1 0 196248 0 1 87181
box 0 0 1 1
use contact_32  contact_32_3197
timestamp 1624857261
transform 1 0 196384 0 1 66645
box 0 0 1 1
use contact_32  contact_32_3196
timestamp 1624857261
transform 1 0 196384 0 1 66373
box 0 0 1 1
use contact_32  contact_32_3195
timestamp 1624857261
transform 1 0 196248 0 1 31149
box 0 0 1 1
use contact_32  contact_32_3194
timestamp 1624857261
transform 1 0 196248 0 1 31421
box 0 0 1 1
use contact_32  contact_32_3193
timestamp 1624857261
transform 1 0 196248 0 1 105405
box 0 0 1 1
use contact_32  contact_32_3192
timestamp 1624857261
transform 1 0 196248 0 1 105677
box 0 0 1 1
use contact_32  contact_32_3191
timestamp 1624857261
transform 1 0 196248 0 1 94253
box 0 0 1 1
use contact_32  contact_32_3190
timestamp 1624857261
transform 1 0 196248 0 1 93981
box 0 0 1 1
use contact_32  contact_32_3189
timestamp 1624857261
transform 1 0 196384 0 1 107717
box 0 0 1 1
use contact_32  contact_32_3188
timestamp 1624857261
transform 1 0 196384 0 1 107445
box 0 0 1 1
use contact_32  contact_32_3187
timestamp 1624857261
transform 1 0 196248 0 1 96701
box 0 0 1 1
use contact_32  contact_32_3186
timestamp 1624857261
transform 1 0 196248 0 1 96973
box 0 0 1 1
use contact_32  contact_32_3185
timestamp 1624857261
transform 1 0 196384 0 1 70997
box 0 0 1 1
use contact_32  contact_32_3184
timestamp 1624857261
transform 1 0 196384 0 1 70725
box 0 0 1 1
use contact_32  contact_32_3183
timestamp 1624857261
transform 1 0 196248 0 1 107309
box 0 0 1 1
use contact_32  contact_32_3182
timestamp 1624857261
transform 1 0 196248 0 1 107037
box 0 0 1 1
use contact_32  contact_32_3181
timestamp 1624857261
transform 1 0 196384 0 1 43797
box 0 0 1 1
use contact_32  contact_32_3180
timestamp 1624857261
transform 1 0 196384 0 1 44069
box 0 0 1 1
use contact_32  contact_32_3179
timestamp 1624857261
transform 1 0 196384 0 1 36181
box 0 0 1 1
use contact_32  contact_32_3178
timestamp 1624857261
transform 1 0 196384 0 1 35909
box 0 0 1 1
use contact_32  contact_32_3177
timestamp 1624857261
transform 1 0 196248 0 1 65149
box 0 0 1 1
use contact_32  contact_32_3176
timestamp 1624857261
transform 1 0 196248 0 1 65421
box 0 0 1 1
use contact_32  contact_32_3175
timestamp 1624857261
transform 1 0 196384 0 1 82965
box 0 0 1 1
use contact_32  contact_32_3174
timestamp 1624857261
transform 1 0 196384 0 1 83237
box 0 0 1 1
use contact_32  contact_32_3173
timestamp 1624857261
transform 1 0 196248 0 1 70317
box 0 0 1 1
use contact_32  contact_32_3172
timestamp 1624857261
transform 1 0 196248 0 1 70589
box 0 0 1 1
use contact_32  contact_32_3171
timestamp 1624857261
transform 1 0 196248 0 1 39037
box 0 0 1 1
use contact_32  contact_32_3170
timestamp 1624857261
transform 1 0 196248 0 1 39309
box 0 0 1 1
use contact_32  contact_32_3169
timestamp 1624857261
transform 1 0 196248 0 1 110573
box 0 0 1 1
use contact_32  contact_32_3168
timestamp 1624857261
transform 1 0 196248 0 1 110845
box 0 0 1 1
use contact_32  contact_32_3167
timestamp 1624857261
transform 1 0 196384 0 1 75485
box 0 0 1 1
use contact_32  contact_32_3166
timestamp 1624857261
transform 1 0 196384 0 1 75757
box 0 0 1 1
use contact_32  contact_32_3165
timestamp 1624857261
transform 1 0 196248 0 1 65965
box 0 0 1 1
use contact_32  contact_32_3164
timestamp 1624857261
transform 1 0 196248 0 1 66237
box 0 0 1 1
use contact_32  contact_32_3163
timestamp 1624857261
transform 1 0 196384 0 1 111253
box 0 0 1 1
use contact_32  contact_32_3162
timestamp 1624857261
transform 1 0 196384 0 1 110981
box 0 0 1 1
use contact_32  contact_32_3161
timestamp 1624857261
transform 1 0 196384 0 1 77661
box 0 0 1 1
use contact_32  contact_32_3160
timestamp 1624857261
transform 1 0 196384 0 1 77389
box 0 0 1 1
use contact_32  contact_32_3159
timestamp 1624857261
transform 1 0 196248 0 1 97517
box 0 0 1 1
use contact_32  contact_32_3158
timestamp 1624857261
transform 1 0 196248 0 1 97789
box 0 0 1 1
use contact_32  contact_32_3157
timestamp 1624857261
transform 1 0 196384 0 1 87317
box 0 0 1 1
use contact_32  contact_32_3156
timestamp 1624857261
transform 1 0 196384 0 1 87589
box 0 0 1 1
use contact_32  contact_32_3155
timestamp 1624857261
transform 1 0 196248 0 1 60389
box 0 0 1 1
use contact_32  contact_32_3154
timestamp 1624857261
transform 1 0 196248 0 1 60661
box 0 0 1 1
use contact_32  contact_32_3153
timestamp 1624857261
transform 1 0 196248 0 1 40125
box 0 0 1 1
use contact_32  contact_32_3152
timestamp 1624857261
transform 1 0 196248 0 1 39853
box 0 0 1 1
use contact_32  contact_32_3151
timestamp 1624857261
transform 1 0 196384 0 1 102549
box 0 0 1 1
use contact_32  contact_32_3150
timestamp 1624857261
transform 1 0 196384 0 1 102277
box 0 0 1 1
use contact_32  contact_32_3149
timestamp 1624857261
transform 1 0 196248 0 1 30333
box 0 0 1 1
use contact_32  contact_32_3148
timestamp 1624857261
transform 1 0 196248 0 1 30605
box 0 0 1 1
use contact_32  contact_32_3147
timestamp 1624857261
transform 1 0 196248 0 1 91261
box 0 0 1 1
use contact_32  contact_32_3146
timestamp 1624857261
transform 1 0 196248 0 1 91533
box 0 0 1 1
use contact_32  contact_32_3145
timestamp 1624857261
transform 1 0 196384 0 1 85141
box 0 0 1 1
use contact_32  contact_32_3144
timestamp 1624857261
transform 1 0 196384 0 1 84869
box 0 0 1 1
use contact_32  contact_32_3143
timestamp 1624857261
transform 1 0 198832 0 1 31013
box 0 0 1 1
use contact_32  contact_32_3142
timestamp 1624857261
transform 1 0 198832 0 1 31421
box 0 0 1 1
use contact_32  contact_32_3141
timestamp 1624857261
transform 1 0 196248 0 1 61885
box 0 0 1 1
use contact_32  contact_32_3140
timestamp 1624857261
transform 1 0 196248 0 1 61613
box 0 0 1 1
use contact_32  contact_32_3139
timestamp 1624857261
transform 1 0 196248 0 1 47741
box 0 0 1 1
use contact_32  contact_32_3138
timestamp 1624857261
transform 1 0 196248 0 1 48013
box 0 0 1 1
use contact_32  contact_32_3137
timestamp 1624857261
transform 1 0 196248 0 1 122813
box 0 0 1 1
use contact_32  contact_32_3136
timestamp 1624857261
transform 1 0 196248 0 1 123085
box 0 0 1 1
use contact_32  contact_32_3135
timestamp 1624857261
transform 1 0 196384 0 1 74261
box 0 0 1 1
use contact_32  contact_32_3134
timestamp 1624857261
transform 1 0 196384 0 1 74533
box 0 0 1 1
use contact_32  contact_32_3133
timestamp 1624857261
transform 1 0 196248 0 1 44205
box 0 0 1 1
use contact_32  contact_32_3132
timestamp 1624857261
transform 1 0 196248 0 1 44477
box 0 0 1 1
use contact_32  contact_32_3131
timestamp 1624857261
transform 1 0 196248 0 1 74669
box 0 0 1 1
use contact_32  contact_32_3130
timestamp 1624857261
transform 1 0 196248 0 1 74941
box 0 0 1 1
use contact_32  contact_32_3129
timestamp 1624857261
transform 1 0 196248 0 1 73445
box 0 0 1 1
use contact_32  contact_32_3128
timestamp 1624857261
transform 1 0 196248 0 1 73717
box 0 0 1 1
use contact_32  contact_32_3127
timestamp 1624857261
transform 1 0 196384 0 1 77253
box 0 0 1 1
use contact_32  contact_32_3126
timestamp 1624857261
transform 1 0 196384 0 1 76981
box 0 0 1 1
use contact_32  contact_32_3125
timestamp 1624857261
transform 1 0 196384 0 1 41349
box 0 0 1 1
use contact_32  contact_32_3124
timestamp 1624857261
transform 1 0 196384 0 1 41077
box 0 0 1 1
use contact_32  contact_32_3123
timestamp 1624857261
transform 1 0 196384 0 1 26389
box 0 0 1 1
use contact_32  contact_32_3122
timestamp 1624857261
transform 1 0 196384 0 1 26661
box 0 0 1 1
use contact_32  contact_32_3121
timestamp 1624857261
transform 1 0 196248 0 1 88813
box 0 0 1 1
use contact_32  contact_32_3120
timestamp 1624857261
transform 1 0 196248 0 1 89085
box 0 0 1 1
use contact_32  contact_32_3119
timestamp 1624857261
transform 1 0 196248 0 1 106221
box 0 0 1 1
use contact_32  contact_32_3118
timestamp 1624857261
transform 1 0 196248 0 1 106493
box 0 0 1 1
use contact_32  contact_32_3117
timestamp 1624857261
transform 1 0 196248 0 1 100645
box 0 0 1 1
use contact_32  contact_32_3116
timestamp 1624857261
transform 1 0 196248 0 1 100917
box 0 0 1 1
use contact_32  contact_32_3115
timestamp 1624857261
transform 1 0 196384 0 1 53181
box 0 0 1 1
use contact_32  contact_32_3114
timestamp 1624857261
transform 1 0 196384 0 1 52909
box 0 0 1 1
use contact_32  contact_32_3113
timestamp 1624857261
transform 1 0 196384 0 1 71813
box 0 0 1 1
use contact_32  contact_32_3112
timestamp 1624857261
transform 1 0 196384 0 1 71541
box 0 0 1 1
use contact_32  contact_32_3111
timestamp 1624857261
transform 1 0 196384 0 1 32645
box 0 0 1 1
use contact_32  contact_32_3110
timestamp 1624857261
transform 1 0 196384 0 1 32373
box 0 0 1 1
use contact_32  contact_32_3109
timestamp 1624857261
transform 1 0 196384 0 1 48965
box 0 0 1 1
use contact_32  contact_32_3108
timestamp 1624857261
transform 1 0 196384 0 1 49237
box 0 0 1 1
use contact_32  contact_32_3107
timestamp 1624857261
transform 1 0 196384 0 1 44885
box 0 0 1 1
use contact_32  contact_32_3106
timestamp 1624857261
transform 1 0 196384 0 1 44613
box 0 0 1 1
use contact_32  contact_32_3105
timestamp 1624857261
transform 1 0 196248 0 1 56445
box 0 0 1 1
use contact_32  contact_32_3104
timestamp 1624857261
transform 1 0 196248 0 1 56717
box 0 0 1 1
use contact_32  contact_32_3103
timestamp 1624857261
transform 1 0 196384 0 1 27477
box 0 0 1 1
use contact_32  contact_32_3102
timestamp 1624857261
transform 1 0 196384 0 1 27205
box 0 0 1 1
use contact_32  contact_32_3101
timestamp 1624857261
transform 1 0 196384 0 1 57941
box 0 0 1 1
use contact_32  contact_32_3100
timestamp 1624857261
transform 1 0 196384 0 1 57669
box 0 0 1 1
use contact_32  contact_32_3099
timestamp 1624857261
transform 1 0 196384 0 1 31557
box 0 0 1 1
use contact_32  contact_32_3098
timestamp 1624857261
transform 1 0 196384 0 1 31829
box 0 0 1 1
use contact_32  contact_32_3097
timestamp 1624857261
transform 1 0 196248 0 1 57261
box 0 0 1 1
use contact_32  contact_32_3096
timestamp 1624857261
transform 1 0 196248 0 1 57533
box 0 0 1 1
use contact_32  contact_32_3095
timestamp 1624857261
transform 1 0 196656 0 1 138317
box 0 0 1 1
use contact_32  contact_32_3094
timestamp 1624857261
transform 1 0 196656 0 1 135597
box 0 0 1 1
use contact_32  contact_32_3093
timestamp 1624857261
transform 1 0 196520 0 1 132605
box 0 0 1 1
use contact_32  contact_32_3092
timestamp 1624857261
transform 1 0 196520 0 1 130021
box 0 0 1 1
use contact_32  contact_32_3091
timestamp 1624857261
transform 1 0 198016 0 1 135461
box 0 0 1 1
use contact_32  contact_32_3090
timestamp 1624857261
transform 1 0 198016 0 1 132741
box 0 0 1 1
use contact_32  contact_32_3089
timestamp 1624857261
transform 1 0 198152 0 1 138453
box 0 0 1 1
use contact_32  contact_32_3088
timestamp 1624857261
transform 1 0 198152 0 1 140493
box 0 0 1 1
use contact_32  contact_32_3087
timestamp 1624857261
transform 1 0 203456 0 1 132741
box 0 0 1 1
use contact_32  contact_32_3086
timestamp 1624857261
transform 1 0 203456 0 1 133829
box 0 0 1 1
use contact_32  contact_32_3085
timestamp 1624857261
transform 1 0 198152 0 1 140629
box 0 0 1 1
use contact_32  contact_32_3084
timestamp 1624857261
transform 1 0 198152 0 1 143485
box 0 0 1 1
use contact_32  contact_32_3083
timestamp 1624857261
transform 1 0 198832 0 1 33189
box 0 0 1 1
use contact_32  contact_32_3082
timestamp 1624857261
transform 1 0 198832 0 1 33869
box 0 0 1 1
use contact_32  contact_32_3081
timestamp 1624857261
transform 1 0 198832 0 1 29109
box 0 0 1 1
use contact_32  contact_32_3080
timestamp 1624857261
transform 1 0 198832 0 1 28429
box 0 0 1 1
use contact_32  contact_32_3079
timestamp 1624857261
transform 1 0 198968 0 1 27613
box 0 0 1 1
use contact_32  contact_32_3078
timestamp 1624857261
transform 1 0 198968 0 1 28293
box 0 0 1 1
use contact_32  contact_32_3077
timestamp 1624857261
transform 1 0 198968 0 1 26117
box 0 0 1 1
use contact_32  contact_32_3076
timestamp 1624857261
transform 1 0 198968 0 1 27341
box 0 0 1 1
use contact_32  contact_32_3075
timestamp 1624857261
transform 1 0 198968 0 1 31557
box 0 0 1 1
use contact_32  contact_32_3074
timestamp 1624857261
transform 1 0 198968 0 1 32237
box 0 0 1 1
use contact_32  contact_32_3073
timestamp 1624857261
transform 1 0 199648 0 1 25301
box 0 0 1 1
use contact_32  contact_32_3072
timestamp 1624857261
transform 1 0 199648 0 1 25981
box 0 0 1 1
use contact_32  contact_32_3071
timestamp 1624857261
transform 1 0 199784 0 1 30061
box 0 0 1 1
use contact_32  contact_32_3070
timestamp 1624857261
transform 1 0 199784 0 1 31421
box 0 0 1 1
use contact_32  contact_32_3069
timestamp 1624857261
transform 1 0 199784 0 1 29245
box 0 0 1 1
use contact_32  contact_32_3068
timestamp 1624857261
transform 1 0 199920 0 1 29925
box 0 0 1 1
use contact_32  contact_32_3067
timestamp 1624857261
transform 1 0 199784 0 1 33053
box 0 0 1 1
use contact_32  contact_32_3066
timestamp 1624857261
transform 1 0 199920 0 1 32373
box 0 0 1 1
use contact_32  contact_32_3065
timestamp 1624857261
transform 1 0 201144 0 1 25165
box 0 0 1 1
use contact_32  contact_32_3064
timestamp 1624857261
transform 1 0 201144 0 1 23533
box 0 0 1 1
use contact_32  contact_32_3063
timestamp 1624857261
transform 1 0 203592 0 1 133829
box 0 0 1 1
use contact_32  contact_32_3062
timestamp 1624857261
transform 1 0 203592 0 1 131109
box 0 0 1 1
use contact_32  contact_32_3061
timestamp 1624857261
transform 1 0 203592 0 1 130973
box 0 0 1 1
use contact_32  contact_32_3060
timestamp 1624857261
transform 1 0 203592 0 1 128389
box 0 0 1 1
use contact_32  contact_32_3059
timestamp 1624857261
transform 1 0 204136 0 1 14965
box 0 0 1 1
use contact_32  contact_32_3058
timestamp 1624857261
transform 1 0 204136 0 1 17685
box 0 0 1 1
use contact_32  contact_32_3057
timestamp 1624857261
transform 1 0 204000 0 1 23261
box 0 0 1 1
use contact_32  contact_32_3056
timestamp 1624857261
transform 1 0 204000 0 1 20677
box 0 0 1 1
use contact_32  contact_32_3055
timestamp 1624857261
transform 1 0 204000 0 1 17821
box 0 0 1 1
use contact_32  contact_32_3054
timestamp 1624857261
transform 1 0 204000 0 1 20541
box 0 0 1 1
use contact_32  contact_32_3053
timestamp 1624857261
transform 1 0 218144 0 1 129613
box 0 0 1 1
use contact_32  contact_32_3052
timestamp 1624857261
transform 1 0 218144 0 1 123901
box 0 0 1 1
use contact_32  contact_32_3051
timestamp 1624857261
transform 1 0 218144 0 1 118461
box 0 0 1 1
use contact_32  contact_32_3050
timestamp 1624857261
transform 1 0 218144 0 1 126893
box 0 0 1 1
use contact_32  contact_32_3049
timestamp 1624857261
transform 1 0 218144 0 1 121045
box 0 0 1 1
use contact_32  contact_32_3048
timestamp 1624857261
transform 1 0 218144 0 1 133829
box 0 0 1 1
use contact_32  contact_32_3047
timestamp 1624857261
transform 1 0 1224 0 1 54133
box 0 0 1 1
use contact_32  contact_32_3046
timestamp 1624857261
transform 1 0 1224 0 1 126485
box 0 0 1 1
use contact_32  contact_32_3045
timestamp 1624857261
transform 1 0 1224 0 1 104725
box 0 0 1 1
use contact_32  contact_32_3044
timestamp 1624857261
transform 1 0 1224 0 1 123221
box 0 0 1 1
use contact_32  contact_32_3043
timestamp 1624857261
transform 1 0 1224 0 1 128117
box 0 0 1 1
use contact_32  contact_32_3042
timestamp 1624857261
transform 1 0 1224 0 1 13877
box 0 0 1 1
use contact_32  contact_32_3041
timestamp 1624857261
transform 1 0 1224 0 1 15509
box 0 0 1 1
use contact_32  contact_32_3040
timestamp 1624857261
transform 1 0 1224 0 1 49237
box 0 0 1 1
use contact_32  contact_32_3039
timestamp 1624857261
transform 1 0 1224 0 1 47605
box 0 0 1 1
use contact_32  contact_32_3038
timestamp 1624857261
transform 1 0 1224 0 1 2181
box 0 0 1 1
use contact_32  contact_32_3037
timestamp 1624857261
transform 1 0 1224 0 1 60933
box 0 0 1 1
use contact_32  contact_32_3036
timestamp 1624857261
transform 1 0 1224 0 1 114653
box 0 0 1 1
use contact_32  contact_32_3035
timestamp 1624857261
transform 1 0 1904 0 1 27477
box 0 0 1 1
use contact_32  contact_32_3034
timestamp 1624857261
transform 1 0 1904 0 1 28021
box 0 0 1 1
use contact_32  contact_32_3033
timestamp 1624857261
transform 1 0 1224 0 1 27477
box 0 0 1 1
use contact_32  contact_32_3032
timestamp 1624857261
transform 1 0 1224 0 1 10613
box 0 0 1 1
use contact_32  contact_32_3031
timestamp 1624857261
transform 1 0 1224 0 1 82693
box 0 0 1 1
use contact_32  contact_32_3030
timestamp 1624857261
transform 1 0 1224 0 1 72629
box 0 0 1 1
use contact_32  contact_32_3029
timestamp 1624857261
transform 1 0 1224 0 1 76165
box 0 0 1 1
use contact_32  contact_32_3028
timestamp 1624857261
transform 1 0 1224 0 1 57669
box 0 0 1 1
use contact_32  contact_32_3027
timestamp 1624857261
transform 1 0 1224 0 1 141717
box 0 0 1 1
use contact_32  contact_32_3026
timestamp 1624857261
transform 1 0 1224 0 1 79565
box 0 0 1 1
use contact_32  contact_32_3025
timestamp 1624857261
transform 1 0 1224 0 1 55901
box 0 0 1 1
use contact_32  contact_32_3024
timestamp 1624857261
transform 1 0 1224 0 1 111253
box 0 0 1 1
use contact_32  contact_32_3023
timestamp 1624857261
transform 1 0 1224 0 1 94661
box 0 0 1 1
use contact_32  contact_32_3022
timestamp 1624857261
transform 1 0 1224 0 1 84461
box 0 0 1 1
use contact_32  contact_32_3021
timestamp 1624857261
transform 1 0 1224 0 1 3813
box 0 0 1 1
use contact_32  contact_32_3020
timestamp 1624857261
transform 1 0 1224 0 1 44069
box 0 0 1 1
use contact_32  contact_32_3019
timestamp 1624857261
transform 1 0 1224 0 1 129749
box 0 0 1 1
use contact_32  contact_32_3018
timestamp 1624857261
transform 1 0 1224 0 1 131517
box 0 0 1 1
use contact_32  contact_32_3017
timestamp 1624857261
transform 1 0 1224 0 1 18909
box 0 0 1 1
use contact_32  contact_32_3016
timestamp 1624857261
transform 1 0 1224 0 1 121317
box 0 0 1 1
use contact_32  contact_32_3015
timestamp 1624857261
transform 1 0 1224 0 1 70997
box 0 0 1 1
use contact_32  contact_32_3014
timestamp 1624857261
transform 1 0 1224 0 1 92757
box 0 0 1 1
use contact_32  contact_32_3013
timestamp 1624857261
transform 1 0 1224 0 1 86229
box 0 0 1 1
use contact_32  contact_32_3012
timestamp 1624857261
transform 1 0 1224 0 1 66101
box 0 0 1 1
use contact_32  contact_32_3011
timestamp 1624857261
transform 1 0 1224 0 1 96157
box 0 0 1 1
use contact_32  contact_32_3010
timestamp 1624857261
transform 1 0 1224 0 1 116421
box 0 0 1 1
use contact_32  contact_32_3009
timestamp 1624857261
transform 1 0 1224 0 1 74533
box 0 0 1 1
use contact_32  contact_32_3008
timestamp 1624857261
transform 1 0 1224 0 1 138181
box 0 0 1 1
use contact_32  contact_32_3007
timestamp 1624857261
transform 1 0 1224 0 1 134917
box 0 0 1 1
use contact_32  contact_32_3006
timestamp 1624857261
transform 1 0 1224 0 1 45973
box 0 0 1 1
use contact_32  contact_32_3005
timestamp 1624857261
transform 1 0 1224 0 1 77661
box 0 0 1 1
use contact_32  contact_32_3004
timestamp 1624857261
transform 1 0 1224 0 1 8981
box 0 0 1 1
use contact_32  contact_32_3003
timestamp 1624857261
transform 1 0 1224 0 1 40805
box 0 0 1 1
use contact_32  contact_32_3002
timestamp 1624857261
transform 1 0 1224 0 1 133149
box 0 0 1 1
use contact_32  contact_32_3001
timestamp 1624857261
transform 1 0 1224 0 1 109621
box 0 0 1 1
use contact_32  contact_32_3000
timestamp 1624857261
transform 1 0 1224 0 1 64197
box 0 0 1 1
use contact_32  contact_32_2999
timestamp 1624857261
transform 1 0 1224 0 1 118053
box 0 0 1 1
use contact_32  contact_32_2998
timestamp 1624857261
transform 1 0 1224 0 1 91125
box 0 0 1 1
use contact_32  contact_32_2997
timestamp 1624857261
transform 1 0 1224 0 1 29109
box 0 0 1 1
use contact_32  contact_32_2996
timestamp 1624857261
transform 1 0 1224 0 1 50869
box 0 0 1 1
use contact_32  contact_32_2995
timestamp 1624857261
transform 1 0 1224 0 1 101189
box 0 0 1 1
use contact_32  contact_32_2994
timestamp 1624857261
transform 1 0 1224 0 1 124853
box 0 0 1 1
use contact_32  contact_32_2993
timestamp 1624857261
transform 1 0 1224 0 1 106357
box 0 0 1 1
use contact_32  contact_32_2992
timestamp 1624857261
transform 1 0 1224 0 1 32373
box 0 0 1 1
use contact_32  contact_32_2991
timestamp 1624857261
transform 1 0 1224 0 1 39173
box 0 0 1 1
use contact_32  contact_32_2990
timestamp 1624857261
transform 1 0 1224 0 1 139813
box 0 0 1 1
use contact_32  contact_32_2989
timestamp 1624857261
transform 1 0 1224 0 1 30741
box 0 0 1 1
use contact_32  contact_32_2988
timestamp 1624857261
transform 1 0 1224 0 1 62565
box 0 0 1 1
use contact_32  contact_32_2987
timestamp 1624857261
transform 1 0 1224 0 1 136685
box 0 0 1 1
use contact_32  contact_32_2986
timestamp 1624857261
transform 1 0 2040 0 1 12245
box 0 0 1 1
use contact_32  contact_32_2985
timestamp 1624857261
transform 1 0 2040 0 1 12517
box 0 0 1 1
use contact_32  contact_32_2984
timestamp 1624857261
transform 1 0 1224 0 1 12245
box 0 0 1 1
use contact_32  contact_32_2983
timestamp 1624857261
transform 1 0 1224 0 1 67733
box 0 0 1 1
use contact_32  contact_32_2982
timestamp 1624857261
transform 1 0 1224 0 1 119685
box 0 0 1 1
use contact_32  contact_32_2981
timestamp 1624857261
transform 1 0 1224 0 1 113021
box 0 0 1 1
use contact_32  contact_32_2980
timestamp 1624857261
transform 1 0 1224 0 1 37405
box 0 0 1 1
use contact_32  contact_32_2979
timestamp 1624857261
transform 1 0 1224 0 1 89493
box 0 0 1 1
use contact_32  contact_32_2978
timestamp 1624857261
transform 1 0 1224 0 1 87861
box 0 0 1 1
use contact_32  contact_32_2977
timestamp 1624857261
transform 1 0 1224 0 1 34005
box 0 0 1 1
use contact_32  contact_32_2976
timestamp 1624857261
transform 1 0 1224 0 1 81061
box 0 0 1 1
use contact_32  contact_32_2975
timestamp 1624857261
transform 1 0 1224 0 1 99557
box 0 0 1 1
use contact_32  contact_32_2974
timestamp 1624857261
transform 1 0 1224 0 1 35637
box 0 0 1 1
use contact_32  contact_32_2973
timestamp 1624857261
transform 1 0 1224 0 1 7077
box 0 0 1 1
use contact_32  contact_32_2972
timestamp 1624857261
transform 1 0 1224 0 1 97925
box 0 0 1 1
use contact_32  contact_32_2971
timestamp 1624857261
transform 1 0 1224 0 1 69365
box 0 0 1 1
use contact_32  contact_32_2970
timestamp 1624857261
transform 1 0 1224 0 1 59165
box 0 0 1 1
use contact_32  contact_32_2969
timestamp 1624857261
transform 1 0 1224 0 1 108125
box 0 0 1 1
use contact_32  contact_32_2968
timestamp 1624857261
transform 1 0 1224 0 1 103093
box 0 0 1 1
use contact_32  contact_32_2967
timestamp 1624857261
transform 1 0 1224 0 1 52501
box 0 0 1 1
use contact_32  contact_32_2966
timestamp 1624857261
transform 1 0 1224 0 1 5445
box 0 0 1 1
use contact_32  contact_32_2965
timestamp 1624857261
transform 1 0 1224 0 1 17277
box 0 0 1 1
use contact_32  contact_32_2964
timestamp 1624857261
transform 1 0 1224 0 1 25573
box 0 0 1 1
use contact_32  contact_32_2963
timestamp 1624857261
transform 1 0 1224 0 1 22309
box 0 0 1 1
use contact_32  contact_32_2962
timestamp 1624857261
transform 1 0 1224 0 1 42437
box 0 0 1 1
use contact_32  contact_32_2961
timestamp 1624857261
transform 1 0 1224 0 1 23941
box 0 0 1 1
use contact_32  contact_32_2960
timestamp 1624857261
transform 1 0 2720 0 1 20541
box 0 0 1 1
use contact_32  contact_32_2959
timestamp 1624857261
transform 1 0 2720 0 1 19725
box 0 0 1 1
use contact_32  contact_32_2958
timestamp 1624857261
transform 1 0 1224 0 1 20677
box 0 0 1 1
use contact_32  contact_32_2957
timestamp 1624857261
transform 1 0 1904 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2956
timestamp 1624857261
transform 1 0 1904 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2955
timestamp 1624857261
transform 1 0 3672 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2954
timestamp 1624857261
transform 1 0 3672 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2953
timestamp 1624857261
transform 1 0 3672 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2952
timestamp 1624857261
transform 1 0 3672 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2951
timestamp 1624857261
transform 1 0 5440 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2950
timestamp 1624857261
transform 1 0 5440 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2949
timestamp 1624857261
transform 1 0 5440 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2948
timestamp 1624857261
transform 1 0 5440 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2947
timestamp 1624857261
transform 1 0 6936 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2946
timestamp 1624857261
transform 1 0 6936 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2945
timestamp 1624857261
transform 1 0 7208 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2944
timestamp 1624857261
transform 1 0 7208 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2943
timestamp 1624857261
transform 1 0 8704 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2942
timestamp 1624857261
transform 1 0 8704 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2941
timestamp 1624857261
transform 1 0 8704 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2940
timestamp 1624857261
transform 1 0 8704 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2939
timestamp 1624857261
transform 1 0 10472 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2938
timestamp 1624857261
transform 1 0 10472 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2937
timestamp 1624857261
transform 1 0 10472 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2936
timestamp 1624857261
transform 1 0 10472 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2935
timestamp 1624857261
transform 1 0 12240 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2934
timestamp 1624857261
transform 1 0 12240 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2933
timestamp 1624857261
transform 1 0 12104 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2932
timestamp 1624857261
transform 1 0 12104 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2931
timestamp 1624857261
transform 1 0 13736 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2930
timestamp 1624857261
transform 1 0 13736 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2929
timestamp 1624857261
transform 1 0 13736 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2928
timestamp 1624857261
transform 1 0 13736 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2927
timestamp 1624857261
transform 1 0 14688 0 1 36997
box 0 0 1 1
use contact_32  contact_32_2926
timestamp 1624857261
transform 1 0 14688 0 1 34413
box 0 0 1 1
use contact_32  contact_32_2925
timestamp 1624857261
transform 1 0 14688 0 1 37133
box 0 0 1 1
use contact_32  contact_32_2924
timestamp 1624857261
transform 1 0 14688 0 1 39853
box 0 0 1 1
use contact_32  contact_32_2923
timestamp 1624857261
transform 1 0 16592 0 1 34141
box 0 0 1 1
use contact_32  contact_32_2922
timestamp 1624857261
transform 1 0 16592 0 1 31557
box 0 0 1 1
use contact_32  contact_32_2921
timestamp 1624857261
transform 1 0 14688 0 1 45565
box 0 0 1 1
use contact_32  contact_32_2920
timestamp 1624857261
transform 1 0 14688 0 1 42845
box 0 0 1 1
use contact_32  contact_32_2919
timestamp 1624857261
transform 1 0 14688 0 1 39989
box 0 0 1 1
use contact_32  contact_32_2918
timestamp 1624857261
transform 1 0 14688 0 1 42709
box 0 0 1 1
use contact_32  contact_32_2917
timestamp 1624857261
transform 1 0 15232 0 1 23805
box 0 0 1 1
use contact_32  contact_32_2916
timestamp 1624857261
transform 1 0 15232 0 1 21085
box 0 0 1 1
use contact_32  contact_32_2915
timestamp 1624857261
transform 1 0 17136 0 1 23941
box 0 0 1 1
use contact_32  contact_32_2914
timestamp 1624857261
transform 1 0 17136 0 1 25165
box 0 0 1 1
use contact_32  contact_32_2913
timestamp 1624857261
transform 1 0 15232 0 1 20949
box 0 0 1 1
use contact_32  contact_32_2912
timestamp 1624857261
transform 1 0 15232 0 1 18365
box 0 0 1 1
use contact_32  contact_32_2911
timestamp 1624857261
transform 1 0 15232 0 1 12653
box 0 0 1 1
use contact_32  contact_32_2910
timestamp 1624857261
transform 1 0 15232 0 1 15373
box 0 0 1 1
use contact_32  contact_32_2909
timestamp 1624857261
transform 1 0 15232 0 1 18093
box 0 0 1 1
use contact_32  contact_32_2908
timestamp 1624857261
transform 1 0 15232 0 1 15509
box 0 0 1 1
use contact_32  contact_32_2907
timestamp 1624857261
transform 1 0 15368 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2906
timestamp 1624857261
transform 1 0 15368 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2905
timestamp 1624857261
transform 1 0 15504 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2904
timestamp 1624857261
transform 1 0 15504 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2903
timestamp 1624857261
transform 1 0 17136 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2902
timestamp 1624857261
transform 1 0 17136 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2901
timestamp 1624857261
transform 1 0 17136 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2900
timestamp 1624857261
transform 1 0 17136 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2899
timestamp 1624857261
transform 1 0 18088 0 1 27613
box 0 0 1 1
use contact_32  contact_32_2898
timestamp 1624857261
transform 1 0 18088 0 1 28293
box 0 0 1 1
use contact_32  contact_32_2897
timestamp 1624857261
transform 1 0 18224 0 1 29925
box 0 0 1 1
use contact_32  contact_32_2896
timestamp 1624857261
transform 1 0 18224 0 1 29245
box 0 0 1 1
use contact_32  contact_32_2895
timestamp 1624857261
transform 1 0 18224 0 1 28429
box 0 0 1 1
use contact_32  contact_32_2894
timestamp 1624857261
transform 1 0 18224 0 1 29109
box 0 0 1 1
use contact_32  contact_32_2893
timestamp 1624857261
transform 1 0 18360 0 1 28293
box 0 0 1 1
use contact_32  contact_32_2892
timestamp 1624857261
transform 1 0 18360 0 1 28021
box 0 0 1 1
use contact_32  contact_32_2891
timestamp 1624857261
transform 1 0 19312 0 1 28021
box 0 0 1 1
use contact_32  contact_32_2890
timestamp 1624857261
transform 1 0 19312 0 1 28293
box 0 0 1 1
use contact_32  contact_32_2889
timestamp 1624857261
transform 1 0 18088 0 1 33053
box 0 0 1 1
use contact_32  contact_32_2888
timestamp 1624857261
transform 1 0 18088 0 1 32373
box 0 0 1 1
use contact_32  contact_32_2887
timestamp 1624857261
transform 1 0 18224 0 1 33189
box 0 0 1 1
use contact_32  contact_32_2886
timestamp 1624857261
transform 1 0 18224 0 1 33869
box 0 0 1 1
use contact_32  contact_32_2885
timestamp 1624857261
transform 1 0 18088 0 1 32237
box 0 0 1 1
use contact_32  contact_32_2884
timestamp 1624857261
transform 1 0 18088 0 1 31557
box 0 0 1 1
use contact_32  contact_32_2883
timestamp 1624857261
transform 1 0 18632 0 1 25301
box 0 0 1 1
use contact_32  contact_32_2882
timestamp 1624857261
transform 1 0 18632 0 1 25981
box 0 0 1 1
use contact_32  contact_32_2881
timestamp 1624857261
transform 1 0 18768 0 1 25301
box 0 0 1 1
use contact_32  contact_32_2880
timestamp 1624857261
transform 1 0 18768 0 1 25573
box 0 0 1 1
use contact_32  contact_32_2879
timestamp 1624857261
transform 1 0 19312 0 1 25573
box 0 0 1 1
use contact_32  contact_32_2878
timestamp 1624857261
transform 1 0 19312 0 1 25301
box 0 0 1 1
use contact_32  contact_32_2877
timestamp 1624857261
transform 1 0 19040 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2876
timestamp 1624857261
transform 1 0 19040 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2875
timestamp 1624857261
transform 1 0 18904 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2874
timestamp 1624857261
transform 1 0 18904 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2873
timestamp 1624857261
transform 1 0 19448 0 1 31557
box 0 0 1 1
use contact_32  contact_32_2872
timestamp 1624857261
transform 1 0 19448 0 1 32237
box 0 0 1 1
use contact_32  contact_32_2871
timestamp 1624857261
transform 1 0 19312 0 1 31421
box 0 0 1 1
use contact_32  contact_32_2870
timestamp 1624857261
transform 1 0 19312 0 1 30061
box 0 0 1 1
use contact_32  contact_32_2869
timestamp 1624857261
transform 1 0 19448 0 1 27613
box 0 0 1 1
use contact_32  contact_32_2868
timestamp 1624857261
transform 1 0 19448 0 1 28293
box 0 0 1 1
use contact_32  contact_32_2867
timestamp 1624857261
transform 1 0 19448 0 1 27477
box 0 0 1 1
use contact_32  contact_32_2866
timestamp 1624857261
transform 1 0 19448 0 1 26117
box 0 0 1 1
use contact_32  contact_32_2865
timestamp 1624857261
transform 1 0 19312 0 1 33189
box 0 0 1 1
use contact_32  contact_32_2864
timestamp 1624857261
transform 1 0 19312 0 1 33869
box 0 0 1 1
use contact_32  contact_32_2863
timestamp 1624857261
transform 1 0 19448 0 1 33053
box 0 0 1 1
use contact_32  contact_32_2862
timestamp 1624857261
transform 1 0 19448 0 1 32373
box 0 0 1 1
use contact_32  contact_32_2861
timestamp 1624857261
transform 1 0 19448 0 1 28429
box 0 0 1 1
use contact_32  contact_32_2860
timestamp 1624857261
transform 1 0 19448 0 1 29109
box 0 0 1 1
use contact_32  contact_32_2859
timestamp 1624857261
transform 1 0 19312 0 1 29245
box 0 0 1 1
use contact_32  contact_32_2858
timestamp 1624857261
transform 1 0 19312 0 1 29925
box 0 0 1 1
use contact_32  contact_32_2857
timestamp 1624857261
transform 1 0 19448 0 1 25301
box 0 0 1 1
use contact_32  contact_32_2856
timestamp 1624857261
transform 1 0 19448 0 1 25845
box 0 0 1 1
use contact_32  contact_32_2855
timestamp 1624857261
transform 1 0 20400 0 1 13741
box 0 0 1 1
use contact_32  contact_32_2854
timestamp 1624857261
transform 1 0 20400 0 1 11021
box 0 0 1 1
use contact_32  contact_32_2853
timestamp 1624857261
transform 1 0 20400 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2852
timestamp 1624857261
transform 1 0 20400 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2851
timestamp 1624857261
transform 1 0 20400 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2850
timestamp 1624857261
transform 1 0 20400 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2849
timestamp 1624857261
transform 1 0 21896 0 1 79429
box 0 0 1 1
use contact_32  contact_32_2848
timestamp 1624857261
transform 1 0 21896 0 1 79701
box 0 0 1 1
use contact_32  contact_32_2847
timestamp 1624857261
transform 1 0 21760 0 1 79293
box 0 0 1 1
use contact_32  contact_32_2846
timestamp 1624857261
transform 1 0 21760 0 1 79021
box 0 0 1 1
use contact_32  contact_32_2845
timestamp 1624857261
transform 1 0 21896 0 1 61205
box 0 0 1 1
use contact_32  contact_32_2844
timestamp 1624857261
transform 1 0 21896 0 1 61477
box 0 0 1 1
use contact_32  contact_32_2843
timestamp 1624857261
transform 1 0 21896 0 1 61069
box 0 0 1 1
use contact_32  contact_32_2842
timestamp 1624857261
transform 1 0 21896 0 1 60797
box 0 0 1 1
use contact_32  contact_32_2841
timestamp 1624857261
transform 1 0 21896 0 1 68685
box 0 0 1 1
use contact_32  contact_32_2840
timestamp 1624857261
transform 1 0 21896 0 1 68957
box 0 0 1 1
use contact_32  contact_32_2839
timestamp 1624857261
transform 1 0 21896 0 1 92757
box 0 0 1 1
use contact_32  contact_32_2838
timestamp 1624857261
transform 1 0 21896 0 1 92485
box 0 0 1 1
use contact_32  contact_32_2837
timestamp 1624857261
transform 1 0 21760 0 1 73717
box 0 0 1 1
use contact_32  contact_32_2836
timestamp 1624857261
transform 1 0 21760 0 1 73445
box 0 0 1 1
use contact_32  contact_32_2835
timestamp 1624857261
transform 1 0 21760 0 1 73853
box 0 0 1 1
use contact_32  contact_32_2834
timestamp 1624857261
transform 1 0 21760 0 1 74125
box 0 0 1 1
use contact_32  contact_32_2833
timestamp 1624857261
transform 1 0 21760 0 1 49645
box 0 0 1 1
use contact_32  contact_32_2832
timestamp 1624857261
transform 1 0 21760 0 1 49373
box 0 0 1 1
use contact_32  contact_32_2831
timestamp 1624857261
transform 1 0 21760 0 1 49781
box 0 0 1 1
use contact_32  contact_32_2830
timestamp 1624857261
transform 1 0 21760 0 1 50053
box 0 0 1 1
use contact_32  contact_32_2829
timestamp 1624857261
transform 1 0 21760 0 1 30333
box 0 0 1 1
use contact_32  contact_32_2828
timestamp 1624857261
transform 1 0 21760 0 1 30061
box 0 0 1 1
use contact_32  contact_32_2827
timestamp 1624857261
transform 1 0 21760 0 1 91941
box 0 0 1 1
use contact_32  contact_32_2826
timestamp 1624857261
transform 1 0 21760 0 1 91669
box 0 0 1 1
use contact_32  contact_32_2825
timestamp 1624857261
transform 1 0 21760 0 1 92077
box 0 0 1 1
use contact_32  contact_32_2824
timestamp 1624857261
transform 1 0 21760 0 1 92349
box 0 0 1 1
use contact_32  contact_32_2823
timestamp 1624857261
transform 1 0 21760 0 1 103909
box 0 0 1 1
use contact_32  contact_32_2822
timestamp 1624857261
transform 1 0 21760 0 1 104181
box 0 0 1 1
use contact_32  contact_32_2821
timestamp 1624857261
transform 1 0 21896 0 1 103773
box 0 0 1 1
use contact_32  contact_32_2820
timestamp 1624857261
transform 1 0 21896 0 1 103501
box 0 0 1 1
use contact_32  contact_32_2819
timestamp 1624857261
transform 1 0 21760 0 1 42981
box 0 0 1 1
use contact_32  contact_32_2818
timestamp 1624857261
transform 1 0 21760 0 1 42709
box 0 0 1 1
use contact_32  contact_32_2817
timestamp 1624857261
transform 1 0 21760 0 1 105133
box 0 0 1 1
use contact_32  contact_32_2816
timestamp 1624857261
transform 1 0 21760 0 1 105405
box 0 0 1 1
use contact_32  contact_32_2815
timestamp 1624857261
transform 1 0 21760 0 1 104997
box 0 0 1 1
use contact_32  contact_32_2814
timestamp 1624857261
transform 1 0 21760 0 1 104725
box 0 0 1 1
use contact_32  contact_32_2813
timestamp 1624857261
transform 1 0 21896 0 1 28293
box 0 0 1 1
use contact_32  contact_32_2812
timestamp 1624857261
transform 1 0 21896 0 1 28021
box 0 0 1 1
use contact_32  contact_32_2811
timestamp 1624857261
transform 1 0 21896 0 1 28429
box 0 0 1 1
use contact_32  contact_32_2810
timestamp 1624857261
transform 1 0 21896 0 1 28701
box 0 0 1 1
use contact_32  contact_32_2809
timestamp 1624857261
transform 1 0 21896 0 1 107853
box 0 0 1 1
use contact_32  contact_32_2808
timestamp 1624857261
transform 1 0 21896 0 1 108125
box 0 0 1 1
use contact_32  contact_32_2807
timestamp 1624857261
transform 1 0 21896 0 1 107717
box 0 0 1 1
use contact_32  contact_32_2806
timestamp 1624857261
transform 1 0 21896 0 1 107445
box 0 0 1 1
use contact_32  contact_32_2805
timestamp 1624857261
transform 1 0 21760 0 1 65013
box 0 0 1 1
use contact_32  contact_32_2804
timestamp 1624857261
transform 1 0 21760 0 1 64741
box 0 0 1 1
use contact_32  contact_32_2803
timestamp 1624857261
transform 1 0 21896 0 1 36317
box 0 0 1 1
use contact_32  contact_32_2802
timestamp 1624857261
transform 1 0 21896 0 1 36589
box 0 0 1 1
use contact_32  contact_32_2801
timestamp 1624857261
transform 1 0 21760 0 1 109349
box 0 0 1 1
use contact_32  contact_32_2800
timestamp 1624857261
transform 1 0 21760 0 1 109077
box 0 0 1 1
use contact_32  contact_32_2799
timestamp 1624857261
transform 1 0 21896 0 1 25301
box 0 0 1 1
use contact_32  contact_32_2798
timestamp 1624857261
transform 1 0 21896 0 1 25573
box 0 0 1 1
use contact_32  contact_32_2797
timestamp 1624857261
transform 1 0 21896 0 1 25165
box 0 0 1 1
use contact_32  contact_32_2796
timestamp 1624857261
transform 1 0 21896 0 1 22309
box 0 0 1 1
use contact_32  contact_32_2795
timestamp 1624857261
transform 1 0 21760 0 1 112613
box 0 0 1 1
use contact_32  contact_32_2794
timestamp 1624857261
transform 1 0 21760 0 1 112885
box 0 0 1 1
use contact_32  contact_32_2793
timestamp 1624857261
transform 1 0 21896 0 1 112477
box 0 0 1 1
use contact_32  contact_32_2792
timestamp 1624857261
transform 1 0 21896 0 1 112205
box 0 0 1 1
use contact_32  contact_32_2791
timestamp 1624857261
transform 1 0 21760 0 1 81333
box 0 0 1 1
use contact_32  contact_32_2790
timestamp 1624857261
transform 1 0 21760 0 1 81605
box 0 0 1 1
use contact_32  contact_32_2789
timestamp 1624857261
transform 1 0 21896 0 1 64333
box 0 0 1 1
use contact_32  contact_32_2788
timestamp 1624857261
transform 1 0 21896 0 1 64061
box 0 0 1 1
use contact_32  contact_32_2787
timestamp 1624857261
transform 1 0 21760 0 1 82557
box 0 0 1 1
use contact_32  contact_32_2786
timestamp 1624857261
transform 1 0 21760 0 1 82829
box 0 0 1 1
use contact_32  contact_32_2785
timestamp 1624857261
transform 1 0 21760 0 1 82421
box 0 0 1 1
use contact_32  contact_32_2784
timestamp 1624857261
transform 1 0 21760 0 1 82149
box 0 0 1 1
use contact_32  contact_32_2783
timestamp 1624857261
transform 1 0 21896 0 1 48149
box 0 0 1 1
use contact_32  contact_32_2782
timestamp 1624857261
transform 1 0 21896 0 1 48421
box 0 0 1 1
use contact_32  contact_32_2781
timestamp 1624857261
transform 1 0 21760 0 1 52909
box 0 0 1 1
use contact_32  contact_32_2780
timestamp 1624857261
transform 1 0 21760 0 1 53181
box 0 0 1 1
use contact_32  contact_32_2779
timestamp 1624857261
transform 1 0 21896 0 1 91533
box 0 0 1 1
use contact_32  contact_32_2778
timestamp 1624857261
transform 1 0 21896 0 1 91261
box 0 0 1 1
use contact_32  contact_32_2777
timestamp 1624857261
transform 1 0 21896 0 1 80925
box 0 0 1 1
use contact_32  contact_32_2776
timestamp 1624857261
transform 1 0 21896 0 1 80653
box 0 0 1 1
use contact_32  contact_32_2775
timestamp 1624857261
transform 1 0 21760 0 1 121317
box 0 0 1 1
use contact_32  contact_32_2774
timestamp 1624857261
transform 1 0 21760 0 1 121589
box 0 0 1 1
use contact_32  contact_32_2773
timestamp 1624857261
transform 1 0 21896 0 1 121181
box 0 0 1 1
use contact_32  contact_32_2772
timestamp 1624857261
transform 1 0 21896 0 1 120909
box 0 0 1 1
use contact_32  contact_32_2771
timestamp 1624857261
transform 1 0 21896 0 1 36997
box 0 0 1 1
use contact_32  contact_32_2770
timestamp 1624857261
transform 1 0 21896 0 1 36725
box 0 0 1 1
use contact_32  contact_32_2769
timestamp 1624857261
transform 1 0 21896 0 1 37133
box 0 0 1 1
use contact_32  contact_32_2768
timestamp 1624857261
transform 1 0 21896 0 1 37405
box 0 0 1 1
use contact_32  contact_32_2767
timestamp 1624857261
transform 1 0 21896 0 1 32781
box 0 0 1 1
use contact_32  contact_32_2766
timestamp 1624857261
transform 1 0 21896 0 1 33053
box 0 0 1 1
use contact_32  contact_32_2765
timestamp 1624857261
transform 1 0 21896 0 1 32645
box 0 0 1 1
use contact_32  contact_32_2764
timestamp 1624857261
transform 1 0 21896 0 1 32373
box 0 0 1 1
use contact_32  contact_32_2763
timestamp 1624857261
transform 1 0 21760 0 1 95477
box 0 0 1 1
use contact_32  contact_32_2762
timestamp 1624857261
transform 1 0 21760 0 1 95205
box 0 0 1 1
use contact_32  contact_32_2761
timestamp 1624857261
transform 1 0 21760 0 1 95613
box 0 0 1 1
use contact_32  contact_32_2760
timestamp 1624857261
transform 1 0 21760 0 1 95885
box 0 0 1 1
use contact_32  contact_32_2759
timestamp 1624857261
transform 1 0 21760 0 1 83373
box 0 0 1 1
use contact_32  contact_32_2758
timestamp 1624857261
transform 1 0 21760 0 1 83645
box 0 0 1 1
use contact_32  contact_32_2757
timestamp 1624857261
transform 1 0 21760 0 1 83237
box 0 0 1 1
use contact_32  contact_32_2756
timestamp 1624857261
transform 1 0 21760 0 1 82965
box 0 0 1 1
use contact_32  contact_32_2755
timestamp 1624857261
transform 1 0 21760 0 1 98605
box 0 0 1 1
use contact_32  contact_32_2754
timestamp 1624857261
transform 1 0 21760 0 1 98333
box 0 0 1 1
use contact_32  contact_32_2753
timestamp 1624857261
transform 1 0 21760 0 1 98741
box 0 0 1 1
use contact_32  contact_32_2752
timestamp 1624857261
transform 1 0 21760 0 1 99013
box 0 0 1 1
use contact_32  contact_32_2751
timestamp 1624857261
transform 1 0 21896 0 1 38221
box 0 0 1 1
use contact_32  contact_32_2750
timestamp 1624857261
transform 1 0 21896 0 1 37949
box 0 0 1 1
use contact_32  contact_32_2749
timestamp 1624857261
transform 1 0 21896 0 1 38357
box 0 0 1 1
use contact_32  contact_32_2748
timestamp 1624857261
transform 1 0 21896 0 1 38629
box 0 0 1 1
use contact_32  contact_32_2747
timestamp 1624857261
transform 1 0 21896 0 1 83781
box 0 0 1 1
use contact_32  contact_32_2746
timestamp 1624857261
transform 1 0 21896 0 1 84053
box 0 0 1 1
use contact_32  contact_32_2745
timestamp 1624857261
transform 1 0 21896 0 1 35093
box 0 0 1 1
use contact_32  contact_32_2744
timestamp 1624857261
transform 1 0 21896 0 1 34821
box 0 0 1 1
use contact_32  contact_32_2743
timestamp 1624857261
transform 1 0 21896 0 1 58077
box 0 0 1 1
use contact_32  contact_32_2742
timestamp 1624857261
transform 1 0 21896 0 1 58349
box 0 0 1 1
use contact_32  contact_32_2741
timestamp 1624857261
transform 1 0 21896 0 1 57941
box 0 0 1 1
use contact_32  contact_32_2740
timestamp 1624857261
transform 1 0 21896 0 1 57669
box 0 0 1 1
use contact_32  contact_32_2739
timestamp 1624857261
transform 1 0 21896 0 1 106629
box 0 0 1 1
use contact_32  contact_32_2738
timestamp 1624857261
transform 1 0 21896 0 1 106901
box 0 0 1 1
use contact_32  contact_32_2737
timestamp 1624857261
transform 1 0 21760 0 1 58485
box 0 0 1 1
use contact_32  contact_32_2736
timestamp 1624857261
transform 1 0 21760 0 1 58757
box 0 0 1 1
use contact_32  contact_32_2735
timestamp 1624857261
transform 1 0 21760 0 1 42165
box 0 0 1 1
use contact_32  contact_32_2734
timestamp 1624857261
transform 1 0 21760 0 1 41893
box 0 0 1 1
use contact_32  contact_32_2733
timestamp 1624857261
transform 1 0 21760 0 1 42301
box 0 0 1 1
use contact_32  contact_32_2732
timestamp 1624857261
transform 1 0 21760 0 1 42573
box 0 0 1 1
use contact_32  contact_32_2731
timestamp 1624857261
transform 1 0 21896 0 1 70997
box 0 0 1 1
use contact_32  contact_32_2730
timestamp 1624857261
transform 1 0 21896 0 1 70725
box 0 0 1 1
use contact_32  contact_32_2729
timestamp 1624857261
transform 1 0 21896 0 1 71133
box 0 0 1 1
use contact_32  contact_32_2728
timestamp 1624857261
transform 1 0 21896 0 1 71405
box 0 0 1 1
use contact_32  contact_32_2727
timestamp 1624857261
transform 1 0 21760 0 1 68277
box 0 0 1 1
use contact_32  contact_32_2726
timestamp 1624857261
transform 1 0 21760 0 1 68005
box 0 0 1 1
use contact_32  contact_32_2725
timestamp 1624857261
transform 1 0 21760 0 1 114925
box 0 0 1 1
use contact_32  contact_32_2724
timestamp 1624857261
transform 1 0 21760 0 1 115197
box 0 0 1 1
use contact_32  contact_32_2723
timestamp 1624857261
transform 1 0 21760 0 1 114789
box 0 0 1 1
use contact_32  contact_32_2722
timestamp 1624857261
transform 1 0 21760 0 1 114517
box 0 0 1 1
use contact_32  contact_32_2721
timestamp 1624857261
transform 1 0 21760 0 1 27885
box 0 0 1 1
use contact_32  contact_32_2720
timestamp 1624857261
transform 1 0 21760 0 1 27613
box 0 0 1 1
use contact_32  contact_32_2719
timestamp 1624857261
transform 1 0 21896 0 1 63109
box 0 0 1 1
use contact_32  contact_32_2718
timestamp 1624857261
transform 1 0 21896 0 1 62837
box 0 0 1 1
use contact_32  contact_32_2717
timestamp 1624857261
transform 1 0 21896 0 1 63245
box 0 0 1 1
use contact_32  contact_32_2716
timestamp 1624857261
transform 1 0 21896 0 1 63517
box 0 0 1 1
use contact_32  contact_32_2715
timestamp 1624857261
transform 1 0 21896 0 1 102685
box 0 0 1 1
use contact_32  contact_32_2714
timestamp 1624857261
transform 1 0 21896 0 1 102957
box 0 0 1 1
use contact_32  contact_32_2713
timestamp 1624857261
transform 1 0 21896 0 1 95069
box 0 0 1 1
use contact_32  contact_32_2712
timestamp 1624857261
transform 1 0 21896 0 1 94797
box 0 0 1 1
use contact_32  contact_32_2711
timestamp 1624857261
transform 1 0 21760 0 1 80109
box 0 0 1 1
use contact_32  contact_32_2710
timestamp 1624857261
transform 1 0 21760 0 1 79837
box 0 0 1 1
use contact_32  contact_32_2709
timestamp 1624857261
transform 1 0 21760 0 1 120365
box 0 0 1 1
use contact_32  contact_32_2708
timestamp 1624857261
transform 1 0 21760 0 1 120093
box 0 0 1 1
use contact_32  contact_32_2707
timestamp 1624857261
transform 1 0 21760 0 1 120501
box 0 0 1 1
use contact_32  contact_32_2706
timestamp 1624857261
transform 1 0 21760 0 1 120773
box 0 0 1 1
use contact_32  contact_32_2705
timestamp 1624857261
transform 1 0 21896 0 1 49237
box 0 0 1 1
use contact_32  contact_32_2704
timestamp 1624857261
transform 1 0 21896 0 1 48965
box 0 0 1 1
use contact_32  contact_32_2703
timestamp 1624857261
transform 1 0 21760 0 1 121725
box 0 0 1 1
use contact_32  contact_32_2702
timestamp 1624857261
transform 1 0 21760 0 1 121997
box 0 0 1 1
use contact_32  contact_32_2701
timestamp 1624857261
transform 1 0 21896 0 1 98197
box 0 0 1 1
use contact_32  contact_32_2700
timestamp 1624857261
transform 1 0 21896 0 1 97925
box 0 0 1 1
use contact_32  contact_32_2699
timestamp 1624857261
transform 1 0 21896 0 1 125533
box 0 0 1 1
use contact_32  contact_32_2698
timestamp 1624857261
transform 1 0 21896 0 1 125261
box 0 0 1 1
use contact_32  contact_32_2697
timestamp 1624857261
transform 1 0 21760 0 1 113021
box 0 0 1 1
use contact_32  contact_32_2696
timestamp 1624857261
transform 1 0 21760 0 1 113293
box 0 0 1 1
use contact_32  contact_32_2695
timestamp 1624857261
transform 1 0 21760 0 1 59573
box 0 0 1 1
use contact_32  contact_32_2694
timestamp 1624857261
transform 1 0 21760 0 1 59301
box 0 0 1 1
use contact_32  contact_32_2693
timestamp 1624857261
transform 1 0 21896 0 1 115333
box 0 0 1 1
use contact_32  contact_32_2692
timestamp 1624857261
transform 1 0 21896 0 1 115605
box 0 0 1 1
use contact_32  contact_32_2691
timestamp 1624857261
transform 1 0 21760 0 1 55357
box 0 0 1 1
use contact_32  contact_32_2690
timestamp 1624857261
transform 1 0 21760 0 1 55629
box 0 0 1 1
use contact_32  contact_32_2689
timestamp 1624857261
transform 1 0 21760 0 1 55221
box 0 0 1 1
use contact_32  contact_32_2688
timestamp 1624857261
transform 1 0 21760 0 1 54949
box 0 0 1 1
use contact_32  contact_32_2687
timestamp 1624857261
transform 1 0 21760 0 1 31149
box 0 0 1 1
use contact_32  contact_32_2686
timestamp 1624857261
transform 1 0 21760 0 1 30877
box 0 0 1 1
use contact_32  contact_32_2685
timestamp 1624857261
transform 1 0 21896 0 1 81741
box 0 0 1 1
use contact_32  contact_32_2684
timestamp 1624857261
transform 1 0 21896 0 1 82013
box 0 0 1 1
use contact_32  contact_32_2683
timestamp 1624857261
transform 1 0 21760 0 1 122405
box 0 0 1 1
use contact_32  contact_32_2682
timestamp 1624857261
transform 1 0 21760 0 1 122677
box 0 0 1 1
use contact_32  contact_32_2681
timestamp 1624857261
transform 1 0 21760 0 1 74669
box 0 0 1 1
use contact_32  contact_32_2680
timestamp 1624857261
transform 1 0 21760 0 1 74941
box 0 0 1 1
use contact_32  contact_32_2679
timestamp 1624857261
transform 1 0 21760 0 1 74533
box 0 0 1 1
use contact_32  contact_32_2678
timestamp 1624857261
transform 1 0 21760 0 1 74261
box 0 0 1 1
use contact_32  contact_32_2677
timestamp 1624857261
transform 1 0 21896 0 1 58893
box 0 0 1 1
use contact_32  contact_32_2676
timestamp 1624857261
transform 1 0 21896 0 1 59165
box 0 0 1 1
use contact_32  contact_32_2675
timestamp 1624857261
transform 1 0 21760 0 1 33461
box 0 0 1 1
use contact_32  contact_32_2674
timestamp 1624857261
transform 1 0 21760 0 1 33189
box 0 0 1 1
use contact_32  contact_32_2673
timestamp 1624857261
transform 1 0 21760 0 1 33597
box 0 0 1 1
use contact_32  contact_32_2672
timestamp 1624857261
transform 1 0 21760 0 1 33869
box 0 0 1 1
use contact_32  contact_32_2671
timestamp 1624857261
transform 1 0 21896 0 1 78613
box 0 0 1 1
use contact_32  contact_32_2670
timestamp 1624857261
transform 1 0 21896 0 1 78885
box 0 0 1 1
use contact_32  contact_32_2669
timestamp 1624857261
transform 1 0 21896 0 1 78477
box 0 0 1 1
use contact_32  contact_32_2668
timestamp 1624857261
transform 1 0 21896 0 1 78205
box 0 0 1 1
use contact_32  contact_32_2667
timestamp 1624857261
transform 1 0 21896 0 1 46109
box 0 0 1 1
use contact_32  contact_32_2666
timestamp 1624857261
transform 1 0 21896 0 1 45837
box 0 0 1 1
use contact_32  contact_32_2665
timestamp 1624857261
transform 1 0 21760 0 1 46245
box 0 0 1 1
use contact_32  contact_32_2664
timestamp 1624857261
transform 1 0 21760 0 1 46517
box 0 0 1 1
use contact_32  contact_32_2663
timestamp 1624857261
transform 1 0 21896 0 1 47469
box 0 0 1 1
use contact_32  contact_32_2662
timestamp 1624857261
transform 1 0 21896 0 1 47741
box 0 0 1 1
use contact_32  contact_32_2661
timestamp 1624857261
transform 1 0 21760 0 1 104317
box 0 0 1 1
use contact_32  contact_32_2660
timestamp 1624857261
transform 1 0 21760 0 1 104589
box 0 0 1 1
use contact_32  contact_32_2659
timestamp 1624857261
transform 1 0 21896 0 1 90445
box 0 0 1 1
use contact_32  contact_32_2658
timestamp 1624857261
transform 1 0 21896 0 1 90717
box 0 0 1 1
use contact_32  contact_32_2657
timestamp 1624857261
transform 1 0 21896 0 1 90309
box 0 0 1 1
use contact_32  contact_32_2656
timestamp 1624857261
transform 1 0 21896 0 1 90037
box 0 0 1 1
use contact_32  contact_32_2655
timestamp 1624857261
transform 1 0 21760 0 1 57261
box 0 0 1 1
use contact_32  contact_32_2654
timestamp 1624857261
transform 1 0 21760 0 1 57533
box 0 0 1 1
use contact_32  contact_32_2653
timestamp 1624857261
transform 1 0 21760 0 1 57125
box 0 0 1 1
use contact_32  contact_32_2652
timestamp 1624857261
transform 1 0 21760 0 1 56853
box 0 0 1 1
use contact_32  contact_32_2651
timestamp 1624857261
transform 1 0 21760 0 1 124853
box 0 0 1 1
use contact_32  contact_32_2650
timestamp 1624857261
transform 1 0 21760 0 1 125125
box 0 0 1 1
use contact_32  contact_32_2649
timestamp 1624857261
transform 1 0 21760 0 1 124717
box 0 0 1 1
use contact_32  contact_32_2648
timestamp 1624857261
transform 1 0 21760 0 1 124445
box 0 0 1 1
use contact_32  contact_32_2647
timestamp 1624857261
transform 1 0 21896 0 1 53725
box 0 0 1 1
use contact_32  contact_32_2646
timestamp 1624857261
transform 1 0 21896 0 1 53997
box 0 0 1 1
use contact_32  contact_32_2645
timestamp 1624857261
transform 1 0 21896 0 1 53589
box 0 0 1 1
use contact_32  contact_32_2644
timestamp 1624857261
transform 1 0 21896 0 1 53317
box 0 0 1 1
use contact_32  contact_32_2643
timestamp 1624857261
transform 1 0 21896 0 1 88541
box 0 0 1 1
use contact_32  contact_32_2642
timestamp 1624857261
transform 1 0 21896 0 1 88813
box 0 0 1 1
use contact_32  contact_32_2641
timestamp 1624857261
transform 1 0 21896 0 1 88405
box 0 0 1 1
use contact_32  contact_32_2640
timestamp 1624857261
transform 1 0 21896 0 1 88133
box 0 0 1 1
use contact_32  contact_32_2639
timestamp 1624857261
transform 1 0 21760 0 1 108261
box 0 0 1 1
use contact_32  contact_32_2638
timestamp 1624857261
transform 1 0 21760 0 1 108533
box 0 0 1 1
use contact_32  contact_32_2637
timestamp 1624857261
transform 1 0 21896 0 1 124037
box 0 0 1 1
use contact_32  contact_32_2636
timestamp 1624857261
transform 1 0 21896 0 1 124309
box 0 0 1 1
use contact_32  contact_32_2635
timestamp 1624857261
transform 1 0 21760 0 1 123901
box 0 0 1 1
use contact_32  contact_32_2634
timestamp 1624857261
transform 1 0 21760 0 1 123629
box 0 0 1 1
use contact_32  contact_32_2633
timestamp 1624857261
transform 1 0 21760 0 1 61613
box 0 0 1 1
use contact_32  contact_32_2632
timestamp 1624857261
transform 1 0 21760 0 1 61885
box 0 0 1 1
use contact_32  contact_32_2631
timestamp 1624857261
transform 1 0 21760 0 1 28837
box 0 0 1 1
use contact_32  contact_32_2630
timestamp 1624857261
transform 1 0 21760 0 1 29109
box 0 0 1 1
use contact_32  contact_32_2629
timestamp 1624857261
transform 1 0 21760 0 1 50597
box 0 0 1 1
use contact_32  contact_32_2628
timestamp 1624857261
transform 1 0 21760 0 1 50869
box 0 0 1 1
use contact_32  contact_32_2627
timestamp 1624857261
transform 1 0 21896 0 1 50461
box 0 0 1 1
use contact_32  contact_32_2626
timestamp 1624857261
transform 1 0 21896 0 1 50189
box 0 0 1 1
use contact_32  contact_32_2625
timestamp 1624857261
transform 1 0 21896 0 1 115741
box 0 0 1 1
use contact_32  contact_32_2624
timestamp 1624857261
transform 1 0 21896 0 1 116013
box 0 0 1 1
use contact_32  contact_32_2623
timestamp 1624857261
transform 1 0 21896 0 1 40533
box 0 0 1 1
use contact_32  contact_32_2622
timestamp 1624857261
transform 1 0 21896 0 1 40261
box 0 0 1 1
use contact_32  contact_32_2621
timestamp 1624857261
transform 1 0 21896 0 1 40669
box 0 0 1 1
use contact_32  contact_32_2620
timestamp 1624857261
transform 1 0 21896 0 1 40941
box 0 0 1 1
use contact_32  contact_32_2619
timestamp 1624857261
transform 1 0 21896 0 1 84869
box 0 0 1 1
use contact_32  contact_32_2618
timestamp 1624857261
transform 1 0 21896 0 1 84597
box 0 0 1 1
use contact_32  contact_32_2617
timestamp 1624857261
transform 1 0 21760 0 1 117237
box 0 0 1 1
use contact_32  contact_32_2616
timestamp 1624857261
transform 1 0 21760 0 1 116965
box 0 0 1 1
use contact_32  contact_32_2615
timestamp 1624857261
transform 1 0 21760 0 1 75893
box 0 0 1 1
use contact_32  contact_32_2614
timestamp 1624857261
transform 1 0 21760 0 1 76165
box 0 0 1 1
use contact_32  contact_32_2613
timestamp 1624857261
transform 1 0 21760 0 1 75757
box 0 0 1 1
use contact_32  contact_32_2612
timestamp 1624857261
transform 1 0 21760 0 1 75485
box 0 0 1 1
use contact_32  contact_32_2611
timestamp 1624857261
transform 1 0 21760 0 1 65829
box 0 0 1 1
use contact_32  contact_32_2610
timestamp 1624857261
transform 1 0 21760 0 1 65557
box 0 0 1 1
use contact_32  contact_32_2609
timestamp 1624857261
transform 1 0 21760 0 1 65965
box 0 0 1 1
use contact_32  contact_32_2608
timestamp 1624857261
transform 1 0 21760 0 1 66237
box 0 0 1 1
use contact_32  contact_32_2607
timestamp 1624857261
transform 1 0 21896 0 1 77661
box 0 0 1 1
use contact_32  contact_32_2606
timestamp 1624857261
transform 1 0 21896 0 1 77389
box 0 0 1 1
use contact_32  contact_32_2605
timestamp 1624857261
transform 1 0 21760 0 1 77797
box 0 0 1 1
use contact_32  contact_32_2604
timestamp 1624857261
transform 1 0 21760 0 1 78069
box 0 0 1 1
use contact_32  contact_32_2603
timestamp 1624857261
transform 1 0 21760 0 1 103093
box 0 0 1 1
use contact_32  contact_32_2602
timestamp 1624857261
transform 1 0 21760 0 1 103365
box 0 0 1 1
use contact_32  contact_32_2601
timestamp 1624857261
transform 1 0 21896 0 1 27205
box 0 0 1 1
use contact_32  contact_32_2600
timestamp 1624857261
transform 1 0 21896 0 1 26933
box 0 0 1 1
use contact_32  contact_32_2599
timestamp 1624857261
transform 1 0 21760 0 1 69501
box 0 0 1 1
use contact_32  contact_32_2598
timestamp 1624857261
transform 1 0 21760 0 1 69773
box 0 0 1 1
use contact_32  contact_32_2597
timestamp 1624857261
transform 1 0 21760 0 1 62701
box 0 0 1 1
use contact_32  contact_32_2596
timestamp 1624857261
transform 1 0 21760 0 1 62429
box 0 0 1 1
use contact_32  contact_32_2595
timestamp 1624857261
transform 1 0 21896 0 1 26117
box 0 0 1 1
use contact_32  contact_32_2594
timestamp 1624857261
transform 1 0 21896 0 1 26389
box 0 0 1 1
use contact_32  contact_32_2593
timestamp 1624857261
transform 1 0 21760 0 1 25981
box 0 0 1 1
use contact_32  contact_32_2592
timestamp 1624857261
transform 1 0 21760 0 1 25709
box 0 0 1 1
use contact_32  contact_32_2591
timestamp 1624857261
transform 1 0 21760 0 1 87725
box 0 0 1 1
use contact_32  contact_32_2590
timestamp 1624857261
transform 1 0 21760 0 1 87997
box 0 0 1 1
use contact_32  contact_32_2589
timestamp 1624857261
transform 1 0 21760 0 1 87589
box 0 0 1 1
use contact_32  contact_32_2588
timestamp 1624857261
transform 1 0 21760 0 1 87317
box 0 0 1 1
use contact_32  contact_32_2587
timestamp 1624857261
transform 1 0 21896 0 1 86093
box 0 0 1 1
use contact_32  contact_32_2586
timestamp 1624857261
transform 1 0 21896 0 1 86365
box 0 0 1 1
use contact_32  contact_32_2585
timestamp 1624857261
transform 1 0 21896 0 1 111253
box 0 0 1 1
use contact_32  contact_32_2584
timestamp 1624857261
transform 1 0 21896 0 1 110981
box 0 0 1 1
use contact_32  contact_32_2583
timestamp 1624857261
transform 1 0 21896 0 1 111389
box 0 0 1 1
use contact_32  contact_32_2582
timestamp 1624857261
transform 1 0 21896 0 1 111661
box 0 0 1 1
use contact_32  contact_32_2581
timestamp 1624857261
transform 1 0 21760 0 1 34277
box 0 0 1 1
use contact_32  contact_32_2580
timestamp 1624857261
transform 1 0 21760 0 1 34005
box 0 0 1 1
use contact_32  contact_32_2579
timestamp 1624857261
transform 1 0 21760 0 1 34413
box 0 0 1 1
use contact_32  contact_32_2578
timestamp 1624857261
transform 1 0 21760 0 1 34685
box 0 0 1 1
use contact_32  contact_32_2577
timestamp 1624857261
transform 1 0 21760 0 1 123493
box 0 0 1 1
use contact_32  contact_32_2576
timestamp 1624857261
transform 1 0 21760 0 1 123221
box 0 0 1 1
use contact_32  contact_32_2575
timestamp 1624857261
transform 1 0 21896 0 1 66781
box 0 0 1 1
use contact_32  contact_32_2574
timestamp 1624857261
transform 1 0 21896 0 1 67053
box 0 0 1 1
use contact_32  contact_32_2573
timestamp 1624857261
transform 1 0 21896 0 1 66645
box 0 0 1 1
use contact_32  contact_32_2572
timestamp 1624857261
transform 1 0 21896 0 1 66373
box 0 0 1 1
use contact_32  contact_32_2571
timestamp 1624857261
transform 1 0 21896 0 1 62293
box 0 0 1 1
use contact_32  contact_32_2570
timestamp 1624857261
transform 1 0 21896 0 1 62021
box 0 0 1 1
use contact_32  contact_32_2569
timestamp 1624857261
transform 1 0 21896 0 1 72221
box 0 0 1 1
use contact_32  contact_32_2568
timestamp 1624857261
transform 1 0 21896 0 1 71949
box 0 0 1 1
use contact_32  contact_32_2567
timestamp 1624857261
transform 1 0 21896 0 1 112069
box 0 0 1 1
use contact_32  contact_32_2566
timestamp 1624857261
transform 1 0 21896 0 1 111797
box 0 0 1 1
use contact_32  contact_32_2565
timestamp 1624857261
transform 1 0 21760 0 1 70589
box 0 0 1 1
use contact_32  contact_32_2564
timestamp 1624857261
transform 1 0 21760 0 1 70317
box 0 0 1 1
use contact_32  contact_32_2563
timestamp 1624857261
transform 1 0 21760 0 1 37541
box 0 0 1 1
use contact_32  contact_32_2562
timestamp 1624857261
transform 1 0 21760 0 1 37813
box 0 0 1 1
use contact_32  contact_32_2561
timestamp 1624857261
transform 1 0 21760 0 1 51005
box 0 0 1 1
use contact_32  contact_32_2560
timestamp 1624857261
transform 1 0 21760 0 1 51277
box 0 0 1 1
use contact_32  contact_32_2559
timestamp 1624857261
transform 1 0 21896 0 1 118733
box 0 0 1 1
use contact_32  contact_32_2558
timestamp 1624857261
transform 1 0 21896 0 1 118461
box 0 0 1 1
use contact_32  contact_32_2557
timestamp 1624857261
transform 1 0 21896 0 1 69909
box 0 0 1 1
use contact_32  contact_32_2556
timestamp 1624857261
transform 1 0 21896 0 1 70181
box 0 0 1 1
use contact_32  contact_32_2555
timestamp 1624857261
transform 1 0 21896 0 1 41757
box 0 0 1 1
use contact_32  contact_32_2554
timestamp 1624857261
transform 1 0 21896 0 1 41485
box 0 0 1 1
use contact_32  contact_32_2553
timestamp 1624857261
transform 1 0 21760 0 1 90853
box 0 0 1 1
use contact_32  contact_32_2552
timestamp 1624857261
transform 1 0 21760 0 1 91125
box 0 0 1 1
use contact_32  contact_32_2551
timestamp 1624857261
transform 1 0 21896 0 1 67869
box 0 0 1 1
use contact_32  contact_32_2550
timestamp 1624857261
transform 1 0 21896 0 1 67597
box 0 0 1 1
use contact_32  contact_32_2549
timestamp 1624857261
transform 1 0 21896 0 1 101461
box 0 0 1 1
use contact_32  contact_32_2548
timestamp 1624857261
transform 1 0 21896 0 1 101189
box 0 0 1 1
use contact_32  contact_32_2547
timestamp 1624857261
transform 1 0 21760 0 1 54133
box 0 0 1 1
use contact_32  contact_32_2546
timestamp 1624857261
transform 1 0 21760 0 1 54405
box 0 0 1 1
use contact_32  contact_32_2545
timestamp 1624857261
transform 1 0 21896 0 1 41349
box 0 0 1 1
use contact_32  contact_32_2544
timestamp 1624857261
transform 1 0 21896 0 1 41077
box 0 0 1 1
use contact_32  contact_32_2543
timestamp 1624857261
transform 1 0 21896 0 1 54813
box 0 0 1 1
use contact_32  contact_32_2542
timestamp 1624857261
transform 1 0 21896 0 1 54541
box 0 0 1 1
use contact_32  contact_32_2541
timestamp 1624857261
transform 1 0 21760 0 1 44205
box 0 0 1 1
use contact_32  contact_32_2540
timestamp 1624857261
transform 1 0 21760 0 1 44477
box 0 0 1 1
use contact_32  contact_32_2539
timestamp 1624857261
transform 1 0 21760 0 1 99965
box 0 0 1 1
use contact_32  contact_32_2538
timestamp 1624857261
transform 1 0 21760 0 1 100237
box 0 0 1 1
use contact_32  contact_32_2537
timestamp 1624857261
transform 1 0 21760 0 1 99829
box 0 0 1 1
use contact_32  contact_32_2536
timestamp 1624857261
transform 1 0 21760 0 1 99557
box 0 0 1 1
use contact_32  contact_32_2535
timestamp 1624857261
transform 1 0 21896 0 1 75349
box 0 0 1 1
use contact_32  contact_32_2534
timestamp 1624857261
transform 1 0 21896 0 1 75077
box 0 0 1 1
use contact_32  contact_32_2533
timestamp 1624857261
transform 1 0 21896 0 1 44613
box 0 0 1 1
use contact_32  contact_32_2532
timestamp 1624857261
transform 1 0 21896 0 1 44885
box 0 0 1 1
use contact_32  contact_32_2531
timestamp 1624857261
transform 1 0 21896 0 1 116829
box 0 0 1 1
use contact_32  contact_32_2530
timestamp 1624857261
transform 1 0 21896 0 1 116557
box 0 0 1 1
use contact_32  contact_32_2529
timestamp 1624857261
transform 1 0 21896 0 1 45021
box 0 0 1 1
use contact_32  contact_32_2528
timestamp 1624857261
transform 1 0 21896 0 1 45293
box 0 0 1 1
use contact_32  contact_32_2527
timestamp 1624857261
transform 1 0 21896 0 1 116421
box 0 0 1 1
use contact_32  contact_32_2526
timestamp 1624857261
transform 1 0 21896 0 1 116149
box 0 0 1 1
use contact_32  contact_32_2525
timestamp 1624857261
transform 1 0 21760 0 1 118053
box 0 0 1 1
use contact_32  contact_32_2524
timestamp 1624857261
transform 1 0 21760 0 1 117781
box 0 0 1 1
use contact_32  contact_32_2523
timestamp 1624857261
transform 1 0 21760 0 1 110573
box 0 0 1 1
use contact_32  contact_32_2522
timestamp 1624857261
transform 1 0 21760 0 1 110845
box 0 0 1 1
use contact_32  contact_32_2521
timestamp 1624857261
transform 1 0 21760 0 1 39037
box 0 0 1 1
use contact_32  contact_32_2520
timestamp 1624857261
transform 1 0 21760 0 1 38765
box 0 0 1 1
use contact_32  contact_32_2519
timestamp 1624857261
transform 1 0 21896 0 1 102141
box 0 0 1 1
use contact_32  contact_32_2518
timestamp 1624857261
transform 1 0 21896 0 1 101869
box 0 0 1 1
use contact_32  contact_32_2517
timestamp 1624857261
transform 1 0 21896 0 1 107037
box 0 0 1 1
use contact_32  contact_32_2516
timestamp 1624857261
transform 1 0 21896 0 1 107309
box 0 0 1 1
use contact_32  contact_32_2515
timestamp 1624857261
transform 1 0 21896 0 1 51413
box 0 0 1 1
use contact_32  contact_32_2514
timestamp 1624857261
transform 1 0 21896 0 1 51685
box 0 0 1 1
use contact_32  contact_32_2513
timestamp 1624857261
transform 1 0 21896 0 1 85277
box 0 0 1 1
use contact_32  contact_32_2512
timestamp 1624857261
transform 1 0 21896 0 1 85549
box 0 0 1 1
use contact_32  contact_32_2511
timestamp 1624857261
transform 1 0 21760 0 1 94389
box 0 0 1 1
use contact_32  contact_32_2510
timestamp 1624857261
transform 1 0 21760 0 1 94661
box 0 0 1 1
use contact_32  contact_32_2509
timestamp 1624857261
transform 1 0 21760 0 1 94253
box 0 0 1 1
use contact_32  contact_32_2508
timestamp 1624857261
transform 1 0 21760 0 1 93981
box 0 0 1 1
use contact_32  contact_32_2507
timestamp 1624857261
transform 1 0 21760 0 1 96293
box 0 0 1 1
use contact_32  contact_32_2506
timestamp 1624857261
transform 1 0 21760 0 1 96021
box 0 0 1 1
use contact_32  contact_32_2505
timestamp 1624857261
transform 1 0 21760 0 1 96429
box 0 0 1 1
use contact_32  contact_32_2504
timestamp 1624857261
transform 1 0 21760 0 1 96701
box 0 0 1 1
use contact_32  contact_32_2503
timestamp 1624857261
transform 1 0 21760 0 1 119277
box 0 0 1 1
use contact_32  contact_32_2502
timestamp 1624857261
transform 1 0 21760 0 1 119549
box 0 0 1 1
use contact_32  contact_32_2501
timestamp 1624857261
transform 1 0 21896 0 1 46925
box 0 0 1 1
use contact_32  contact_32_2500
timestamp 1624857261
transform 1 0 21896 0 1 46653
box 0 0 1 1
use contact_32  contact_32_2499
timestamp 1624857261
transform 1 0 21760 0 1 86501
box 0 0 1 1
use contact_32  contact_32_2498
timestamp 1624857261
transform 1 0 21760 0 1 86773
box 0 0 1 1
use contact_32  contact_32_2497
timestamp 1624857261
transform 1 0 21896 0 1 71813
box 0 0 1 1
use contact_32  contact_32_2496
timestamp 1624857261
transform 1 0 21896 0 1 71541
box 0 0 1 1
use contact_32  contact_32_2495
timestamp 1624857261
transform 1 0 21896 0 1 31557
box 0 0 1 1
use contact_32  contact_32_2494
timestamp 1624857261
transform 1 0 21896 0 1 31829
box 0 0 1 1
use contact_32  contact_32_2493
timestamp 1624857261
transform 1 0 21896 0 1 67461
box 0 0 1 1
use contact_32  contact_32_2492
timestamp 1624857261
transform 1 0 21896 0 1 67189
box 0 0 1 1
use contact_32  contact_32_2491
timestamp 1624857261
transform 1 0 21896 0 1 45701
box 0 0 1 1
use contact_32  contact_32_2490
timestamp 1624857261
transform 1 0 21896 0 1 45429
box 0 0 1 1
use contact_32  contact_32_2489
timestamp 1624857261
transform 1 0 21896 0 1 29517
box 0 0 1 1
use contact_32  contact_32_2488
timestamp 1624857261
transform 1 0 21896 0 1 29245
box 0 0 1 1
use contact_32  contact_32_2487
timestamp 1624857261
transform 1 0 21896 0 1 29653
box 0 0 1 1
use contact_32  contact_32_2486
timestamp 1624857261
transform 1 0 21896 0 1 29925
box 0 0 1 1
use contact_32  contact_32_2485
timestamp 1624857261
transform 1 0 21760 0 1 86909
box 0 0 1 1
use contact_32  contact_32_2484
timestamp 1624857261
transform 1 0 21760 0 1 87181
box 0 0 1 1
use contact_32  contact_32_2483
timestamp 1624857261
transform 1 0 21896 0 1 119957
box 0 0 1 1
use contact_32  contact_32_2482
timestamp 1624857261
transform 1 0 21896 0 1 119685
box 0 0 1 1
use contact_32  contact_32_2481
timestamp 1624857261
transform 1 0 21760 0 1 100645
box 0 0 1 1
use contact_32  contact_32_2480
timestamp 1624857261
transform 1 0 21760 0 1 100373
box 0 0 1 1
use contact_32  contact_32_2479
timestamp 1624857261
transform 1 0 21760 0 1 108669
box 0 0 1 1
use contact_32  contact_32_2478
timestamp 1624857261
transform 1 0 21760 0 1 108941
box 0 0 1 1
use contact_32  contact_32_2477
timestamp 1624857261
transform 1 0 21896 0 1 99149
box 0 0 1 1
use contact_32  contact_32_2476
timestamp 1624857261
transform 1 0 21896 0 1 99421
box 0 0 1 1
use contact_32  contact_32_2475
timestamp 1624857261
transform 1 0 21760 0 1 13877
box 0 0 1 1
use contact_32  contact_32_2474
timestamp 1624857261
transform 1 0 21760 0 1 16461
box 0 0 1 1
use contact_32  contact_32_2473
timestamp 1624857261
transform 1 0 21760 0 1 19453
box 0 0 1 1
use contact_32  contact_32_2472
timestamp 1624857261
transform 1 0 21760 0 1 22173
box 0 0 1 1
use contact_32  contact_32_2471
timestamp 1624857261
transform 1 0 21760 0 1 19317
box 0 0 1 1
use contact_32  contact_32_2470
timestamp 1624857261
transform 1 0 21760 0 1 16733
box 0 0 1 1
use contact_32  contact_32_2469
timestamp 1624857261
transform 1 0 22168 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2468
timestamp 1624857261
transform 1 0 22168 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2467
timestamp 1624857261
transform 1 0 22168 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2466
timestamp 1624857261
transform 1 0 22168 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2465
timestamp 1624857261
transform 1 0 23256 0 1 75621
box 0 0 1 1
use contact_32  contact_32_2464
timestamp 1624857261
transform 1 0 23256 0 1 75213
box 0 0 1 1
use contact_32  contact_32_2463
timestamp 1624857261
transform 1 0 22984 0 1 93845
box 0 0 1 1
use contact_32  contact_32_2462
timestamp 1624857261
transform 1 0 22984 0 1 93573
box 0 0 1 1
use contact_32  contact_32_2461
timestamp 1624857261
transform 1 0 22984 0 1 93981
box 0 0 1 1
use contact_32  contact_32_2460
timestamp 1624857261
transform 1 0 22984 0 1 94253
box 0 0 1 1
use contact_32  contact_32_2459
timestamp 1624857261
transform 1 0 23120 0 1 83373
box 0 0 1 1
use contact_32  contact_32_2458
timestamp 1624857261
transform 1 0 23120 0 1 83645
box 0 0 1 1
use contact_32  contact_32_2457
timestamp 1624857261
transform 1 0 23120 0 1 83237
box 0 0 1 1
use contact_32  contact_32_2456
timestamp 1624857261
transform 1 0 23120 0 1 82965
box 0 0 1 1
use contact_32  contact_32_2455
timestamp 1624857261
transform 1 0 23120 0 1 97925
box 0 0 1 1
use contact_32  contact_32_2454
timestamp 1624857261
transform 1 0 23120 0 1 98197
box 0 0 1 1
use contact_32  contact_32_2453
timestamp 1624857261
transform 1 0 22984 0 1 97789
box 0 0 1 1
use contact_32  contact_32_2452
timestamp 1624857261
transform 1 0 22984 0 1 97517
box 0 0 1 1
use contact_32  contact_32_2451
timestamp 1624857261
transform 1 0 22984 0 1 30741
box 0 0 1 1
use contact_32  contact_32_2450
timestamp 1624857261
transform 1 0 22984 0 1 31013
box 0 0 1 1
use contact_32  contact_32_2449
timestamp 1624857261
transform 1 0 22984 0 1 56445
box 0 0 1 1
use contact_32  contact_32_2448
timestamp 1624857261
transform 1 0 22984 0 1 56717
box 0 0 1 1
use contact_32  contact_32_2447
timestamp 1624857261
transform 1 0 22984 0 1 56309
box 0 0 1 1
use contact_32  contact_32_2446
timestamp 1624857261
transform 1 0 22984 0 1 56037
box 0 0 1 1
use contact_32  contact_32_2445
timestamp 1624857261
transform 1 0 23120 0 1 81741
box 0 0 1 1
use contact_32  contact_32_2444
timestamp 1624857261
transform 1 0 23120 0 1 82013
box 0 0 1 1
use contact_32  contact_32_2443
timestamp 1624857261
transform 1 0 23120 0 1 81605
box 0 0 1 1
use contact_32  contact_32_2442
timestamp 1624857261
transform 1 0 23120 0 1 81333
box 0 0 1 1
use contact_32  contact_32_2441
timestamp 1624857261
transform 1 0 22984 0 1 53181
box 0 0 1 1
use contact_32  contact_32_2440
timestamp 1624857261
transform 1 0 22984 0 1 52909
box 0 0 1 1
use contact_32  contact_32_2439
timestamp 1624857261
transform 1 0 23120 0 1 53317
box 0 0 1 1
use contact_32  contact_32_2438
timestamp 1624857261
transform 1 0 23120 0 1 53589
box 0 0 1 1
use contact_32  contact_32_2437
timestamp 1624857261
transform 1 0 23120 0 1 48965
box 0 0 1 1
use contact_32  contact_32_2436
timestamp 1624857261
transform 1 0 23120 0 1 49237
box 0 0 1 1
use contact_32  contact_32_2435
timestamp 1624857261
transform 1 0 22984 0 1 48829
box 0 0 1 1
use contact_32  contact_32_2434
timestamp 1624857261
transform 1 0 22984 0 1 48557
box 0 0 1 1
use contact_32  contact_32_2433
timestamp 1624857261
transform 1 0 23120 0 1 31557
box 0 0 1 1
use contact_32  contact_32_2432
timestamp 1624857261
transform 1 0 23120 0 1 31829
box 0 0 1 1
use contact_32  contact_32_2431
timestamp 1624857261
transform 1 0 22984 0 1 31421
box 0 0 1 1
use contact_32  contact_32_2430
timestamp 1624857261
transform 1 0 22984 0 1 31149
box 0 0 1 1
use contact_32  contact_32_2429
timestamp 1624857261
transform 1 0 22984 0 1 123901
box 0 0 1 1
use contact_32  contact_32_2428
timestamp 1624857261
transform 1 0 22984 0 1 123629
box 0 0 1 1
use contact_32  contact_32_2427
timestamp 1624857261
transform 1 0 23120 0 1 124037
box 0 0 1 1
use contact_32  contact_32_2426
timestamp 1624857261
transform 1 0 23120 0 1 124309
box 0 0 1 1
use contact_32  contact_32_2425
timestamp 1624857261
transform 1 0 22984 0 1 52501
box 0 0 1 1
use contact_32  contact_32_2424
timestamp 1624857261
transform 1 0 22984 0 1 52773
box 0 0 1 1
use contact_32  contact_32_2423
timestamp 1624857261
transform 1 0 22984 0 1 52365
box 0 0 1 1
use contact_32  contact_32_2422
timestamp 1624857261
transform 1 0 22984 0 1 52093
box 0 0 1 1
use contact_32  contact_32_2421
timestamp 1624857261
transform 1 0 23120 0 1 123493
box 0 0 1 1
use contact_32  contact_32_2420
timestamp 1624857261
transform 1 0 23120 0 1 123221
box 0 0 1 1
use contact_32  contact_32_2419
timestamp 1624857261
transform 1 0 22984 0 1 33053
box 0 0 1 1
use contact_32  contact_32_2418
timestamp 1624857261
transform 1 0 22984 0 1 32781
box 0 0 1 1
use contact_32  contact_32_2417
timestamp 1624857261
transform 1 0 23120 0 1 33189
box 0 0 1 1
use contact_32  contact_32_2416
timestamp 1624857261
transform 1 0 23120 0 1 33461
box 0 0 1 1
use contact_32  contact_32_2415
timestamp 1624857261
transform 1 0 23120 0 1 120773
box 0 0 1 1
use contact_32  contact_32_2414
timestamp 1624857261
transform 1 0 23120 0 1 120501
box 0 0 1 1
use contact_32  contact_32_2413
timestamp 1624857261
transform 1 0 22984 0 1 58349
box 0 0 1 1
use contact_32  contact_32_2412
timestamp 1624857261
transform 1 0 22984 0 1 58077
box 0 0 1 1
use contact_32  contact_32_2411
timestamp 1624857261
transform 1 0 22984 0 1 58485
box 0 0 1 1
use contact_32  contact_32_2410
timestamp 1624857261
transform 1 0 22984 0 1 58757
box 0 0 1 1
use contact_32  contact_32_2409
timestamp 1624857261
transform 1 0 22984 0 1 107445
box 0 0 1 1
use contact_32  contact_32_2408
timestamp 1624857261
transform 1 0 22984 0 1 107717
box 0 0 1 1
use contact_32  contact_32_2407
timestamp 1624857261
transform 1 0 22984 0 1 107309
box 0 0 1 1
use contact_32  contact_32_2406
timestamp 1624857261
transform 1 0 22984 0 1 107037
box 0 0 1 1
use contact_32  contact_32_2405
timestamp 1624857261
transform 1 0 23120 0 1 121997
box 0 0 1 1
use contact_32  contact_32_2404
timestamp 1624857261
transform 1 0 23120 0 1 122269
box 0 0 1 1
use contact_32  contact_32_2403
timestamp 1624857261
transform 1 0 22984 0 1 111797
box 0 0 1 1
use contact_32  contact_32_2402
timestamp 1624857261
transform 1 0 22984 0 1 112069
box 0 0 1 1
use contact_32  contact_32_2401
timestamp 1624857261
transform 1 0 23120 0 1 111661
box 0 0 1 1
use contact_32  contact_32_2400
timestamp 1624857261
transform 1 0 23120 0 1 111389
box 0 0 1 1
use contact_32  contact_32_2399
timestamp 1624857261
transform 1 0 23120 0 1 62021
box 0 0 1 1
use contact_32  contact_32_2398
timestamp 1624857261
transform 1 0 23120 0 1 62293
box 0 0 1 1
use contact_32  contact_32_2397
timestamp 1624857261
transform 1 0 22984 0 1 61885
box 0 0 1 1
use contact_32  contact_32_2396
timestamp 1624857261
transform 1 0 22984 0 1 61613
box 0 0 1 1
use contact_32  contact_32_2395
timestamp 1624857261
transform 1 0 23120 0 1 110437
box 0 0 1 1
use contact_32  contact_32_2394
timestamp 1624857261
transform 1 0 23120 0 1 110165
box 0 0 1 1
use contact_32  contact_32_2393
timestamp 1624857261
transform 1 0 23120 0 1 110573
box 0 0 1 1
use contact_32  contact_32_2392
timestamp 1624857261
transform 1 0 23120 0 1 110845
box 0 0 1 1
use contact_32  contact_32_2391
timestamp 1624857261
transform 1 0 23120 0 1 86093
box 0 0 1 1
use contact_32  contact_32_2390
timestamp 1624857261
transform 1 0 23120 0 1 86365
box 0 0 1 1
use contact_32  contact_32_2389
timestamp 1624857261
transform 1 0 23120 0 1 85957
box 0 0 1 1
use contact_32  contact_32_2388
timestamp 1624857261
transform 1 0 23120 0 1 85685
box 0 0 1 1
use contact_32  contact_32_2387
timestamp 1624857261
transform 1 0 23120 0 1 84461
box 0 0 1 1
use contact_32  contact_32_2386
timestamp 1624857261
transform 1 0 23120 0 1 84733
box 0 0 1 1
use contact_32  contact_32_2385
timestamp 1624857261
transform 1 0 23120 0 1 29925
box 0 0 1 1
use contact_32  contact_32_2384
timestamp 1624857261
transform 1 0 23120 0 1 29653
box 0 0 1 1
use contact_32  contact_32_2383
timestamp 1624857261
transform 1 0 23120 0 1 99013
box 0 0 1 1
use contact_32  contact_32_2382
timestamp 1624857261
transform 1 0 23120 0 1 98741
box 0 0 1 1
use contact_32  contact_32_2381
timestamp 1624857261
transform 1 0 23120 0 1 99149
box 0 0 1 1
use contact_32  contact_32_2380
timestamp 1624857261
transform 1 0 23120 0 1 99421
box 0 0 1 1
use contact_32  contact_32_2379
timestamp 1624857261
transform 1 0 22984 0 1 124445
box 0 0 1 1
use contact_32  contact_32_2378
timestamp 1624857261
transform 1 0 22984 0 1 124717
box 0 0 1 1
use contact_32  contact_32_2377
timestamp 1624857261
transform 1 0 22984 0 1 72221
box 0 0 1 1
use contact_32  contact_32_2376
timestamp 1624857261
transform 1 0 22984 0 1 72493
box 0 0 1 1
use contact_32  contact_32_2375
timestamp 1624857261
transform 1 0 23120 0 1 112205
box 0 0 1 1
use contact_32  contact_32_2374
timestamp 1624857261
transform 1 0 23120 0 1 112477
box 0 0 1 1
use contact_32  contact_32_2373
timestamp 1624857261
transform 1 0 23120 0 1 101733
box 0 0 1 1
use contact_32  contact_32_2372
timestamp 1624857261
transform 1 0 23120 0 1 101461
box 0 0 1 1
use contact_32  contact_32_2371
timestamp 1624857261
transform 1 0 23120 0 1 101869
box 0 0 1 1
use contact_32  contact_32_2370
timestamp 1624857261
transform 1 0 23120 0 1 102141
box 0 0 1 1
use contact_32  contact_32_2369
timestamp 1624857261
transform 1 0 22984 0 1 91669
box 0 0 1 1
use contact_32  contact_32_2368
timestamp 1624857261
transform 1 0 22984 0 1 91941
box 0 0 1 1
use contact_32  contact_32_2367
timestamp 1624857261
transform 1 0 23120 0 1 91533
box 0 0 1 1
use contact_32  contact_32_2366
timestamp 1624857261
transform 1 0 23120 0 1 91261
box 0 0 1 1
use contact_32  contact_32_2365
timestamp 1624857261
transform 1 0 23120 0 1 65965
box 0 0 1 1
use contact_32  contact_32_2364
timestamp 1624857261
transform 1 0 23120 0 1 66237
box 0 0 1 1
use contact_32  contact_32_2363
timestamp 1624857261
transform 1 0 23120 0 1 65829
box 0 0 1 1
use contact_32  contact_32_2362
timestamp 1624857261
transform 1 0 23120 0 1 65557
box 0 0 1 1
use contact_32  contact_32_2361
timestamp 1624857261
transform 1 0 22984 0 1 93437
box 0 0 1 1
use contact_32  contact_32_2360
timestamp 1624857261
transform 1 0 22984 0 1 93165
box 0 0 1 1
use contact_32  contact_32_2359
timestamp 1624857261
transform 1 0 22984 0 1 44477
box 0 0 1 1
use contact_32  contact_32_2358
timestamp 1624857261
transform 1 0 22984 0 1 44205
box 0 0 1 1
use contact_32  contact_32_2357
timestamp 1624857261
transform 1 0 23120 0 1 44613
box 0 0 1 1
use contact_32  contact_32_2356
timestamp 1624857261
transform 1 0 23120 0 1 44885
box 0 0 1 1
use contact_32  contact_32_2355
timestamp 1624857261
transform 1 0 23120 0 1 86501
box 0 0 1 1
use contact_32  contact_32_2354
timestamp 1624857261
transform 1 0 23120 0 1 86773
box 0 0 1 1
use contact_32  contact_32_2353
timestamp 1624857261
transform 1 0 22984 0 1 104181
box 0 0 1 1
use contact_32  contact_32_2352
timestamp 1624857261
transform 1 0 22984 0 1 103909
box 0 0 1 1
use contact_32  contact_32_2351
timestamp 1624857261
transform 1 0 22984 0 1 90037
box 0 0 1 1
use contact_32  contact_32_2350
timestamp 1624857261
transform 1 0 22984 0 1 90309
box 0 0 1 1
use contact_32  contact_32_2349
timestamp 1624857261
transform 1 0 22984 0 1 89901
box 0 0 1 1
use contact_32  contact_32_2348
timestamp 1624857261
transform 1 0 22984 0 1 89629
box 0 0 1 1
use contact_32  contact_32_2347
timestamp 1624857261
transform 1 0 23120 0 1 105813
box 0 0 1 1
use contact_32  contact_32_2346
timestamp 1624857261
transform 1 0 23120 0 1 106085
box 0 0 1 1
use contact_32  contact_32_2345
timestamp 1624857261
transform 1 0 23120 0 1 105677
box 0 0 1 1
use contact_32  contact_32_2344
timestamp 1624857261
transform 1 0 23120 0 1 105405
box 0 0 1 1
use contact_32  contact_32_2343
timestamp 1624857261
transform 1 0 23120 0 1 41893
box 0 0 1 1
use contact_32  contact_32_2342
timestamp 1624857261
transform 1 0 23120 0 1 42165
box 0 0 1 1
use contact_32  contact_32_2341
timestamp 1624857261
transform 1 0 22984 0 1 41757
box 0 0 1 1
use contact_32  contact_32_2340
timestamp 1624857261
transform 1 0 22984 0 1 41485
box 0 0 1 1
use contact_32  contact_32_2339
timestamp 1624857261
transform 1 0 23120 0 1 85549
box 0 0 1 1
use contact_32  contact_32_2338
timestamp 1624857261
transform 1 0 23120 0 1 85277
box 0 0 1 1
use contact_32  contact_32_2337
timestamp 1624857261
transform 1 0 23120 0 1 113701
box 0 0 1 1
use contact_32  contact_32_2336
timestamp 1624857261
transform 1 0 23120 0 1 113973
box 0 0 1 1
use contact_32  contact_32_2335
timestamp 1624857261
transform 1 0 23120 0 1 67053
box 0 0 1 1
use contact_32  contact_32_2334
timestamp 1624857261
transform 1 0 23120 0 1 66781
box 0 0 1 1
use contact_32  contact_32_2333
timestamp 1624857261
transform 1 0 23120 0 1 114789
box 0 0 1 1
use contact_32  contact_32_2332
timestamp 1624857261
transform 1 0 23120 0 1 114517
box 0 0 1 1
use contact_32  contact_32_2331
timestamp 1624857261
transform 1 0 23120 0 1 114925
box 0 0 1 1
use contact_32  contact_32_2330
timestamp 1624857261
transform 1 0 23120 0 1 115197
box 0 0 1 1
use contact_32  contact_32_2329
timestamp 1624857261
transform 1 0 23120 0 1 106221
box 0 0 1 1
use contact_32  contact_32_2328
timestamp 1624857261
transform 1 0 23120 0 1 106493
box 0 0 1 1
use contact_32  contact_32_2327
timestamp 1624857261
transform 1 0 22984 0 1 101053
box 0 0 1 1
use contact_32  contact_32_2326
timestamp 1624857261
transform 1 0 22984 0 1 101325
box 0 0 1 1
use contact_32  contact_32_2325
timestamp 1624857261
transform 1 0 22984 0 1 57941
box 0 0 1 1
use contact_32  contact_32_2324
timestamp 1624857261
transform 1 0 22984 0 1 57669
box 0 0 1 1
use contact_32  contact_32_2323
timestamp 1624857261
transform 1 0 22984 0 1 37949
box 0 0 1 1
use contact_32  contact_32_2322
timestamp 1624857261
transform 1 0 22984 0 1 38221
box 0 0 1 1
use contact_32  contact_32_2321
timestamp 1624857261
transform 1 0 22984 0 1 37813
box 0 0 1 1
use contact_32  contact_32_2320
timestamp 1624857261
transform 1 0 22984 0 1 37541
box 0 0 1 1
use contact_32  contact_32_2319
timestamp 1624857261
transform 1 0 22984 0 1 46517
box 0 0 1 1
use contact_32  contact_32_2318
timestamp 1624857261
transform 1 0 22984 0 1 46245
box 0 0 1 1
use contact_32  contact_32_2317
timestamp 1624857261
transform 1 0 22984 0 1 86909
box 0 0 1 1
use contact_32  contact_32_2316
timestamp 1624857261
transform 1 0 22984 0 1 87181
box 0 0 1 1
use contact_32  contact_32_2315
timestamp 1624857261
transform 1 0 23120 0 1 84869
box 0 0 1 1
use contact_32  contact_32_2314
timestamp 1624857261
transform 1 0 23120 0 1 85141
box 0 0 1 1
use contact_32  contact_32_2313
timestamp 1624857261
transform 1 0 23120 0 1 51685
box 0 0 1 1
use contact_32  contact_32_2312
timestamp 1624857261
transform 1 0 23120 0 1 51957
box 0 0 1 1
use contact_32  contact_32_2311
timestamp 1624857261
transform 1 0 23120 0 1 64333
box 0 0 1 1
use contact_32  contact_32_2310
timestamp 1624857261
transform 1 0 23120 0 1 64605
box 0 0 1 1
use contact_32  contact_32_2309
timestamp 1624857261
transform 1 0 23120 0 1 64197
box 0 0 1 1
use contact_32  contact_32_2308
timestamp 1624857261
transform 1 0 23120 0 1 63925
box 0 0 1 1
use contact_32  contact_32_2307
timestamp 1624857261
transform 1 0 22984 0 1 49645
box 0 0 1 1
use contact_32  contact_32_2306
timestamp 1624857261
transform 1 0 22984 0 1 49373
box 0 0 1 1
use contact_32  contact_32_2305
timestamp 1624857261
transform 1 0 22984 0 1 49781
box 0 0 1 1
use contact_32  contact_32_2304
timestamp 1624857261
transform 1 0 22984 0 1 50053
box 0 0 1 1
use contact_32  contact_32_2303
timestamp 1624857261
transform 1 0 22984 0 1 114381
box 0 0 1 1
use contact_32  contact_32_2302
timestamp 1624857261
transform 1 0 22984 0 1 114109
box 0 0 1 1
use contact_32  contact_32_2301
timestamp 1624857261
transform 1 0 22984 0 1 109757
box 0 0 1 1
use contact_32  contact_32_2300
timestamp 1624857261
transform 1 0 22984 0 1 110029
box 0 0 1 1
use contact_32  contact_32_2299
timestamp 1624857261
transform 1 0 22984 0 1 109621
box 0 0 1 1
use contact_32  contact_32_2298
timestamp 1624857261
transform 1 0 22984 0 1 109349
box 0 0 1 1
use contact_32  contact_32_2297
timestamp 1624857261
transform 1 0 23120 0 1 44069
box 0 0 1 1
use contact_32  contact_32_2296
timestamp 1624857261
transform 1 0 23120 0 1 43797
box 0 0 1 1
use contact_32  contact_32_2295
timestamp 1624857261
transform 1 0 22984 0 1 102685
box 0 0 1 1
use contact_32  contact_32_2294
timestamp 1624857261
transform 1 0 22984 0 1 102957
box 0 0 1 1
use contact_32  contact_32_2293
timestamp 1624857261
transform 1 0 22984 0 1 102549
box 0 0 1 1
use contact_32  contact_32_2292
timestamp 1624857261
transform 1 0 22984 0 1 102277
box 0 0 1 1
use contact_32  contact_32_2291
timestamp 1624857261
transform 1 0 23120 0 1 88813
box 0 0 1 1
use contact_32  contact_32_2290
timestamp 1624857261
transform 1 0 23120 0 1 89085
box 0 0 1 1
use contact_32  contact_32_2289
timestamp 1624857261
transform 1 0 22984 0 1 66645
box 0 0 1 1
use contact_32  contact_32_2288
timestamp 1624857261
transform 1 0 22984 0 1 66373
box 0 0 1 1
use contact_32  contact_32_2287
timestamp 1624857261
transform 1 0 22984 0 1 80789
box 0 0 1 1
use contact_32  contact_32_2286
timestamp 1624857261
transform 1 0 22984 0 1 80517
box 0 0 1 1
use contact_32  contact_32_2285
timestamp 1624857261
transform 1 0 22984 0 1 80925
box 0 0 1 1
use contact_32  contact_32_2284
timestamp 1624857261
transform 1 0 22984 0 1 81197
box 0 0 1 1
use contact_32  contact_32_2283
timestamp 1624857261
transform 1 0 22984 0 1 122677
box 0 0 1 1
use contact_32  contact_32_2282
timestamp 1624857261
transform 1 0 22984 0 1 122405
box 0 0 1 1
use contact_32  contact_32_2281
timestamp 1624857261
transform 1 0 22984 0 1 122813
box 0 0 1 1
use contact_32  contact_32_2280
timestamp 1624857261
transform 1 0 22984 0 1 123085
box 0 0 1 1
use contact_32  contact_32_2279
timestamp 1624857261
transform 1 0 23120 0 1 64741
box 0 0 1 1
use contact_32  contact_32_2278
timestamp 1624857261
transform 1 0 23120 0 1 65013
box 0 0 1 1
use contact_32  contact_32_2277
timestamp 1624857261
transform 1 0 22984 0 1 28701
box 0 0 1 1
use contact_32  contact_32_2276
timestamp 1624857261
transform 1 0 22984 0 1 28429
box 0 0 1 1
use contact_32  contact_32_2275
timestamp 1624857261
transform 1 0 23120 0 1 28837
box 0 0 1 1
use contact_32  contact_32_2274
timestamp 1624857261
transform 1 0 23120 0 1 29109
box 0 0 1 1
use contact_32  contact_32_2273
timestamp 1624857261
transform 1 0 23120 0 1 93029
box 0 0 1 1
use contact_32  contact_32_2272
timestamp 1624857261
transform 1 0 23120 0 1 92757
box 0 0 1 1
use contact_32  contact_32_2271
timestamp 1624857261
transform 1 0 22984 0 1 94389
box 0 0 1 1
use contact_32  contact_32_2270
timestamp 1624857261
transform 1 0 22984 0 1 94661
box 0 0 1 1
use contact_32  contact_32_2269
timestamp 1624857261
transform 1 0 23120 0 1 110981
box 0 0 1 1
use contact_32  contact_32_2268
timestamp 1624857261
transform 1 0 23120 0 1 111253
box 0 0 1 1
use contact_32  contact_32_2267
timestamp 1624857261
transform 1 0 23120 0 1 82149
box 0 0 1 1
use contact_32  contact_32_2266
timestamp 1624857261
transform 1 0 23120 0 1 82421
box 0 0 1 1
use contact_32  contact_32_2265
timestamp 1624857261
transform 1 0 22984 0 1 69773
box 0 0 1 1
use contact_32  contact_32_2264
timestamp 1624857261
transform 1 0 22984 0 1 69501
box 0 0 1 1
use contact_32  contact_32_2263
timestamp 1624857261
transform 1 0 22984 0 1 69909
box 0 0 1 1
use contact_32  contact_32_2262
timestamp 1624857261
transform 1 0 22984 0 1 70181
box 0 0 1 1
use contact_32  contact_32_2261
timestamp 1624857261
transform 1 0 23120 0 1 117645
box 0 0 1 1
use contact_32  contact_32_2260
timestamp 1624857261
transform 1 0 23120 0 1 117917
box 0 0 1 1
use contact_32  contact_32_2259
timestamp 1624857261
transform 1 0 23120 0 1 82829
box 0 0 1 1
use contact_32  contact_32_2258
timestamp 1624857261
transform 1 0 23120 0 1 82557
box 0 0 1 1
use contact_32  contact_32_2257
timestamp 1624857261
transform 1 0 22984 0 1 70997
box 0 0 1 1
use contact_32  contact_32_2256
timestamp 1624857261
transform 1 0 22984 0 1 70725
box 0 0 1 1
use contact_32  contact_32_2255
timestamp 1624857261
transform 1 0 22984 0 1 57533
box 0 0 1 1
use contact_32  contact_32_2254
timestamp 1624857261
transform 1 0 22984 0 1 57261
box 0 0 1 1
use contact_32  contact_32_2253
timestamp 1624857261
transform 1 0 23120 0 1 100237
box 0 0 1 1
use contact_32  contact_32_2252
timestamp 1624857261
transform 1 0 23120 0 1 99965
box 0 0 1 1
use contact_32  contact_32_2251
timestamp 1624857261
transform 1 0 23120 0 1 25573
box 0 0 1 1
use contact_32  contact_32_2250
timestamp 1624857261
transform 1 0 23120 0 1 25301
box 0 0 1 1
use contact_32  contact_32_2249
timestamp 1624857261
transform 1 0 23120 0 1 45837
box 0 0 1 1
use contact_32  contact_32_2248
timestamp 1624857261
transform 1 0 23120 0 1 46109
box 0 0 1 1
use contact_32  contact_32_2247
timestamp 1624857261
transform 1 0 23120 0 1 45701
box 0 0 1 1
use contact_32  contact_32_2246
timestamp 1624857261
transform 1 0 23120 0 1 45429
box 0 0 1 1
use contact_32  contact_32_2245
timestamp 1624857261
transform 1 0 22984 0 1 69365
box 0 0 1 1
use contact_32  contact_32_2244
timestamp 1624857261
transform 1 0 22984 0 1 69093
box 0 0 1 1
use contact_32  contact_32_2243
timestamp 1624857261
transform 1 0 22984 0 1 78477
box 0 0 1 1
use contact_32  contact_32_2242
timestamp 1624857261
transform 1 0 22984 0 1 78205
box 0 0 1 1
use contact_32  contact_32_2241
timestamp 1624857261
transform 1 0 22984 0 1 78613
box 0 0 1 1
use contact_32  contact_32_2240
timestamp 1624857261
transform 1 0 22984 0 1 78885
box 0 0 1 1
use contact_32  contact_32_2239
timestamp 1624857261
transform 1 0 23120 0 1 106629
box 0 0 1 1
use contact_32  contact_32_2238
timestamp 1624857261
transform 1 0 23120 0 1 106901
box 0 0 1 1
use contact_32  contact_32_2237
timestamp 1624857261
transform 1 0 22984 0 1 70589
box 0 0 1 1
use contact_32  contact_32_2236
timestamp 1624857261
transform 1 0 22984 0 1 70317
box 0 0 1 1
use contact_32  contact_32_2235
timestamp 1624857261
transform 1 0 22984 0 1 78069
box 0 0 1 1
use contact_32  contact_32_2234
timestamp 1624857261
transform 1 0 22984 0 1 77797
box 0 0 1 1
use contact_32  contact_32_2233
timestamp 1624857261
transform 1 0 23120 0 1 119277
box 0 0 1 1
use contact_32  contact_32_2232
timestamp 1624857261
transform 1 0 23120 0 1 119549
box 0 0 1 1
use contact_32  contact_32_2231
timestamp 1624857261
transform 1 0 23120 0 1 119141
box 0 0 1 1
use contact_32  contact_32_2230
timestamp 1624857261
transform 1 0 23120 0 1 118869
box 0 0 1 1
use contact_32  contact_32_2229
timestamp 1624857261
transform 1 0 23120 0 1 73037
box 0 0 1 1
use contact_32  contact_32_2228
timestamp 1624857261
transform 1 0 23120 0 1 73309
box 0 0 1 1
use contact_32  contact_32_2227
timestamp 1624857261
transform 1 0 23120 0 1 72901
box 0 0 1 1
use contact_32  contact_32_2226
timestamp 1624857261
transform 1 0 23120 0 1 72629
box 0 0 1 1
use contact_32  contact_32_2225
timestamp 1624857261
transform 1 0 23120 0 1 87589
box 0 0 1 1
use contact_32  contact_32_2224
timestamp 1624857261
transform 1 0 23120 0 1 87317
box 0 0 1 1
use contact_32  contact_32_2223
timestamp 1624857261
transform 1 0 23120 0 1 26797
box 0 0 1 1
use contact_32  contact_32_2222
timestamp 1624857261
transform 1 0 23120 0 1 27069
box 0 0 1 1
use contact_32  contact_32_2221
timestamp 1624857261
transform 1 0 23120 0 1 89221
box 0 0 1 1
use contact_32  contact_32_2220
timestamp 1624857261
transform 1 0 23120 0 1 89493
box 0 0 1 1
use contact_32  contact_32_2219
timestamp 1624857261
transform 1 0 22984 0 1 98605
box 0 0 1 1
use contact_32  contact_32_2218
timestamp 1624857261
transform 1 0 22984 0 1 98333
box 0 0 1 1
use contact_32  contact_32_2217
timestamp 1624857261
transform 1 0 22984 0 1 40125
box 0 0 1 1
use contact_32  contact_32_2216
timestamp 1624857261
transform 1 0 22984 0 1 39853
box 0 0 1 1
use contact_32  contact_32_2215
timestamp 1624857261
transform 1 0 23120 0 1 40261
box 0 0 1 1
use contact_32  contact_32_2214
timestamp 1624857261
transform 1 0 23120 0 1 40533
box 0 0 1 1
use contact_32  contact_32_2213
timestamp 1624857261
transform 1 0 22984 0 1 60661
box 0 0 1 1
use contact_32  contact_32_2212
timestamp 1624857261
transform 1 0 22984 0 1 60389
box 0 0 1 1
use contact_32  contact_32_2211
timestamp 1624857261
transform 1 0 22984 0 1 60797
box 0 0 1 1
use contact_32  contact_32_2210
timestamp 1624857261
transform 1 0 22984 0 1 61069
box 0 0 1 1
use contact_32  contact_32_2209
timestamp 1624857261
transform 1 0 22984 0 1 91125
box 0 0 1 1
use contact_32  contact_32_2208
timestamp 1624857261
transform 1 0 22984 0 1 90853
box 0 0 1 1
use contact_32  contact_32_2207
timestamp 1624857261
transform 1 0 22984 0 1 68277
box 0 0 1 1
use contact_32  contact_32_2206
timestamp 1624857261
transform 1 0 22984 0 1 68549
box 0 0 1 1
use contact_32  contact_32_2205
timestamp 1624857261
transform 1 0 22984 0 1 76573
box 0 0 1 1
use contact_32  contact_32_2204
timestamp 1624857261
transform 1 0 22984 0 1 76845
box 0 0 1 1
use contact_32  contact_32_2203
timestamp 1624857261
transform 1 0 22984 0 1 103773
box 0 0 1 1
use contact_32  contact_32_2202
timestamp 1624857261
transform 1 0 22984 0 1 103501
box 0 0 1 1
use contact_32  contact_32_2201
timestamp 1624857261
transform 1 0 23120 0 1 90445
box 0 0 1 1
use contact_32  contact_32_2200
timestamp 1624857261
transform 1 0 23120 0 1 90717
box 0 0 1 1
use contact_32  contact_32_2199
timestamp 1624857261
transform 1 0 23120 0 1 94797
box 0 0 1 1
use contact_32  contact_32_2198
timestamp 1624857261
transform 1 0 23120 0 1 95069
box 0 0 1 1
use contact_32  contact_32_2197
timestamp 1624857261
transform 1 0 23120 0 1 107853
box 0 0 1 1
use contact_32  contact_32_2196
timestamp 1624857261
transform 1 0 23120 0 1 108125
box 0 0 1 1
use contact_32  contact_32_2195
timestamp 1624857261
transform 1 0 23120 0 1 59981
box 0 0 1 1
use contact_32  contact_32_2194
timestamp 1624857261
transform 1 0 23120 0 1 60253
box 0 0 1 1
use contact_32  contact_32_2193
timestamp 1624857261
transform 1 0 22984 0 1 76981
box 0 0 1 1
use contact_32  contact_32_2192
timestamp 1624857261
transform 1 0 22984 0 1 77253
box 0 0 1 1
use contact_32  contact_32_2191
timestamp 1624857261
transform 1 0 23120 0 1 57125
box 0 0 1 1
use contact_32  contact_32_2190
timestamp 1624857261
transform 1 0 23120 0 1 56853
box 0 0 1 1
use contact_32  contact_32_2189
timestamp 1624857261
transform 1 0 23120 0 1 68685
box 0 0 1 1
use contact_32  contact_32_2188
timestamp 1624857261
transform 1 0 23120 0 1 68957
box 0 0 1 1
use contact_32  contact_32_2187
timestamp 1624857261
transform 1 0 23120 0 1 116421
box 0 0 1 1
use contact_32  contact_32_2186
timestamp 1624857261
transform 1 0 23120 0 1 116149
box 0 0 1 1
use contact_32  contact_32_2185
timestamp 1624857261
transform 1 0 22984 0 1 28021
box 0 0 1 1
use contact_32  contact_32_2184
timestamp 1624857261
transform 1 0 22984 0 1 28293
box 0 0 1 1
use contact_32  contact_32_2183
timestamp 1624857261
transform 1 0 23120 0 1 27885
box 0 0 1 1
use contact_32  contact_32_2182
timestamp 1624857261
transform 1 0 23120 0 1 27613
box 0 0 1 1
use contact_32  contact_32_2181
timestamp 1624857261
transform 1 0 22984 0 1 47605
box 0 0 1 1
use contact_32  contact_32_2180
timestamp 1624857261
transform 1 0 22984 0 1 47333
box 0 0 1 1
use contact_32  contact_32_2179
timestamp 1624857261
transform 1 0 22984 0 1 47741
box 0 0 1 1
use contact_32  contact_32_2178
timestamp 1624857261
transform 1 0 22984 0 1 48013
box 0 0 1 1
use contact_32  contact_32_2177
timestamp 1624857261
transform 1 0 22984 0 1 31965
box 0 0 1 1
use contact_32  contact_32_2176
timestamp 1624857261
transform 1 0 22984 0 1 32237
box 0 0 1 1
use contact_32  contact_32_2175
timestamp 1624857261
transform 1 0 23120 0 1 79021
box 0 0 1 1
use contact_32  contact_32_2174
timestamp 1624857261
transform 1 0 23120 0 1 79293
box 0 0 1 1
use contact_32  contact_32_2173
timestamp 1624857261
transform 1 0 22984 0 1 29517
box 0 0 1 1
use contact_32  contact_32_2172
timestamp 1624857261
transform 1 0 22984 0 1 29245
box 0 0 1 1
use contact_32  contact_32_2171
timestamp 1624857261
transform 1 0 22984 0 1 95477
box 0 0 1 1
use contact_32  contact_32_2170
timestamp 1624857261
transform 1 0 22984 0 1 95205
box 0 0 1 1
use contact_32  contact_32_2169
timestamp 1624857261
transform 1 0 22984 0 1 95613
box 0 0 1 1
use contact_32  contact_32_2168
timestamp 1624857261
transform 1 0 22984 0 1 95885
box 0 0 1 1
use contact_32  contact_32_2167
timestamp 1624857261
transform 1 0 22984 0 1 65149
box 0 0 1 1
use contact_32  contact_32_2166
timestamp 1624857261
transform 1 0 22984 0 1 65421
box 0 0 1 1
use contact_32  contact_32_2165
timestamp 1624857261
transform 1 0 22984 0 1 43661
box 0 0 1 1
use contact_32  contact_32_2164
timestamp 1624857261
transform 1 0 22984 0 1 43389
box 0 0 1 1
use contact_32  contact_32_2163
timestamp 1624857261
transform 1 0 23120 0 1 48421
box 0 0 1 1
use contact_32  contact_32_2162
timestamp 1624857261
transform 1 0 23120 0 1 48149
box 0 0 1 1
use contact_32  contact_32_2161
timestamp 1624857261
transform 1 0 22984 0 1 50461
box 0 0 1 1
use contact_32  contact_32_2160
timestamp 1624857261
transform 1 0 22984 0 1 50189
box 0 0 1 1
use contact_32  contact_32_2159
timestamp 1624857261
transform 1 0 23120 0 1 103093
box 0 0 1 1
use contact_32  contact_32_2158
timestamp 1624857261
transform 1 0 23120 0 1 103365
box 0 0 1 1
use contact_32  contact_32_2157
timestamp 1624857261
transform 1 0 22984 0 1 115741
box 0 0 1 1
use contact_32  contact_32_2156
timestamp 1624857261
transform 1 0 22984 0 1 116013
box 0 0 1 1
use contact_32  contact_32_2155
timestamp 1624857261
transform 1 0 22984 0 1 115605
box 0 0 1 1
use contact_32  contact_32_2154
timestamp 1624857261
transform 1 0 22984 0 1 115333
box 0 0 1 1
use contact_32  contact_32_2153
timestamp 1624857261
transform 1 0 23120 0 1 119685
box 0 0 1 1
use contact_32  contact_32_2152
timestamp 1624857261
transform 1 0 23120 0 1 119957
box 0 0 1 1
use contact_32  contact_32_2151
timestamp 1624857261
transform 1 0 22984 0 1 53725
box 0 0 1 1
use contact_32  contact_32_2150
timestamp 1624857261
transform 1 0 22984 0 1 53997
box 0 0 1 1
use contact_32  contact_32_2149
timestamp 1624857261
transform 1 0 23120 0 1 118053
box 0 0 1 1
use contact_32  contact_32_2148
timestamp 1624857261
transform 1 0 23120 0 1 118325
box 0 0 1 1
use contact_32  contact_32_2147
timestamp 1624857261
transform 1 0 22984 0 1 39309
box 0 0 1 1
use contact_32  contact_32_2146
timestamp 1624857261
transform 1 0 22984 0 1 39037
box 0 0 1 1
use contact_32  contact_32_2145
timestamp 1624857261
transform 1 0 22984 0 1 39445
box 0 0 1 1
use contact_32  contact_32_2144
timestamp 1624857261
transform 1 0 22984 0 1 39717
box 0 0 1 1
use contact_32  contact_32_2143
timestamp 1624857261
transform 1 0 22984 0 1 45293
box 0 0 1 1
use contact_32  contact_32_2142
timestamp 1624857261
transform 1 0 22984 0 1 45021
box 0 0 1 1
use contact_32  contact_32_2141
timestamp 1624857261
transform 1 0 22984 0 1 97109
box 0 0 1 1
use contact_32  contact_32_2140
timestamp 1624857261
transform 1 0 22984 0 1 97381
box 0 0 1 1
use contact_32  contact_32_2139
timestamp 1624857261
transform 1 0 23120 0 1 99557
box 0 0 1 1
use contact_32  contact_32_2138
timestamp 1624857261
transform 1 0 23120 0 1 99829
box 0 0 1 1
use contact_32  contact_32_2137
timestamp 1624857261
transform 1 0 22984 0 1 77661
box 0 0 1 1
use contact_32  contact_32_2136
timestamp 1624857261
transform 1 0 22984 0 1 77389
box 0 0 1 1
use contact_32  contact_32_2135
timestamp 1624857261
transform 1 0 22984 0 1 62429
box 0 0 1 1
use contact_32  contact_32_2134
timestamp 1624857261
transform 1 0 22984 0 1 62701
box 0 0 1 1
use contact_32  contact_32_2133
timestamp 1624857261
transform 1 0 23120 0 1 27205
box 0 0 1 1
use contact_32  contact_32_2132
timestamp 1624857261
transform 1 0 23120 0 1 27477
box 0 0 1 1
use contact_32  contact_32_2131
timestamp 1624857261
transform 1 0 23120 0 1 120365
box 0 0 1 1
use contact_32  contact_32_2130
timestamp 1624857261
transform 1 0 23120 0 1 120093
box 0 0 1 1
use contact_32  contact_32_2129
timestamp 1624857261
transform 1 0 23120 0 1 32645
box 0 0 1 1
use contact_32  contact_32_2128
timestamp 1624857261
transform 1 0 23120 0 1 32373
box 0 0 1 1
use contact_32  contact_32_2127
timestamp 1624857261
transform 1 0 23120 0 1 35909
box 0 0 1 1
use contact_32  contact_32_2126
timestamp 1624857261
transform 1 0 23120 0 1 36181
box 0 0 1 1
use contact_32  contact_32_2125
timestamp 1624857261
transform 1 0 22984 0 1 35773
box 0 0 1 1
use contact_32  contact_32_2124
timestamp 1624857261
transform 1 0 22984 0 1 35501
box 0 0 1 1
use contact_32  contact_32_2123
timestamp 1624857261
transform 1 0 23120 0 1 54133
box 0 0 1 1
use contact_32  contact_32_2122
timestamp 1624857261
transform 1 0 23120 0 1 54405
box 0 0 1 1
use contact_32  contact_32_2121
timestamp 1624857261
transform 1 0 22984 0 1 55901
box 0 0 1 1
use contact_32  contact_32_2120
timestamp 1624857261
transform 1 0 22984 0 1 55629
box 0 0 1 1
use contact_32  contact_32_2119
timestamp 1624857261
transform 1 0 22984 0 1 37405
box 0 0 1 1
use contact_32  contact_32_2118
timestamp 1624857261
transform 1 0 22984 0 1 37133
box 0 0 1 1
use contact_32  contact_32_2117
timestamp 1624857261
transform 1 0 22984 0 1 33597
box 0 0 1 1
use contact_32  contact_32_2116
timestamp 1624857261
transform 1 0 22984 0 1 33869
box 0 0 1 1
use contact_32  contact_32_2115
timestamp 1624857261
transform 1 0 23120 0 1 41349
box 0 0 1 1
use contact_32  contact_32_2114
timestamp 1624857261
transform 1 0 23120 0 1 41077
box 0 0 1 1
use contact_32  contact_32_2113
timestamp 1624857261
transform 1 0 22984 0 1 118461
box 0 0 1 1
use contact_32  contact_32_2112
timestamp 1624857261
transform 1 0 22984 0 1 118733
box 0 0 1 1
use contact_32  contact_32_2111
timestamp 1624857261
transform 1 0 23120 0 1 73445
box 0 0 1 1
use contact_32  contact_32_2110
timestamp 1624857261
transform 1 0 23120 0 1 73717
box 0 0 1 1
use contact_32  contact_32_2109
timestamp 1624857261
transform 1 0 23120 0 1 75077
box 0 0 1 1
use contact_32  contact_32_2108
timestamp 1624857261
transform 1 0 23120 0 1 75349
box 0 0 1 1
use contact_32  contact_32_2107
timestamp 1624857261
transform 1 0 22984 0 1 74941
box 0 0 1 1
use contact_32  contact_32_2106
timestamp 1624857261
transform 1 0 22984 0 1 74669
box 0 0 1 1
use contact_32  contact_32_2105
timestamp 1624857261
transform 1 0 22984 0 1 36317
box 0 0 1 1
use contact_32  contact_32_2104
timestamp 1624857261
transform 1 0 22984 0 1 36589
box 0 0 1 1
use contact_32  contact_32_2103
timestamp 1624857261
transform 1 0 22984 0 1 74125
box 0 0 1 1
use contact_32  contact_32_2102
timestamp 1624857261
transform 1 0 22984 0 1 73853
box 0 0 1 1
use contact_32  contact_32_2101
timestamp 1624857261
transform 1 0 22984 0 1 74261
box 0 0 1 1
use contact_32  contact_32_2100
timestamp 1624857261
transform 1 0 22984 0 1 74533
box 0 0 1 1
use contact_32  contact_32_2099
timestamp 1624857261
transform 1 0 22984 0 1 36725
box 0 0 1 1
use contact_32  contact_32_2098
timestamp 1624857261
transform 1 0 22984 0 1 36997
box 0 0 1 1
use contact_32  contact_32_2097
timestamp 1624857261
transform 1 0 22984 0 1 40941
box 0 0 1 1
use contact_32  contact_32_2096
timestamp 1624857261
transform 1 0 22984 0 1 40669
box 0 0 1 1
use contact_32  contact_32_2095
timestamp 1624857261
transform 1 0 23120 0 1 61477
box 0 0 1 1
use contact_32  contact_32_2094
timestamp 1624857261
transform 1 0 23120 0 1 61205
box 0 0 1 1
use contact_32  contact_32_2093
timestamp 1624857261
transform 1 0 22984 0 1 35093
box 0 0 1 1
use contact_32  contact_32_2092
timestamp 1624857261
transform 1 0 22984 0 1 35365
box 0 0 1 1
use contact_32  contact_32_2091
timestamp 1624857261
transform 1 0 23936 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2090
timestamp 1624857261
transform 1 0 23936 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2089
timestamp 1624857261
transform 1 0 23936 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2088
timestamp 1624857261
transform 1 0 23936 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2087
timestamp 1624857261
transform 1 0 25296 0 1 75077
box 0 0 1 1
use contact_32  contact_32_2086
timestamp 1624857261
transform 1 0 25296 0 1 75349
box 0 0 1 1
use contact_32  contact_32_2085
timestamp 1624857261
transform 1 0 25432 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2084
timestamp 1624857261
transform 1 0 25432 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2083
timestamp 1624857261
transform 1 0 25432 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2082
timestamp 1624857261
transform 1 0 25432 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2081
timestamp 1624857261
transform 1 0 27200 0 1 142397
box 0 0 1 1
use contact_32  contact_32_2080
timestamp 1624857261
transform 1 0 27200 0 1 142805
box 0 0 1 1
use contact_32  contact_32_2079
timestamp 1624857261
transform 1 0 27200 0 1 1773
box 0 0 1 1
use contact_32  contact_32_2078
timestamp 1624857261
transform 1 0 27200 0 1 1229
box 0 0 1 1
use contact_32  contact_32_2077
timestamp 1624857261
transform 1 0 29920 0 1 24621
box 0 0 1 1
use contact_32  contact_32_2076
timestamp 1624857261
transform 1 0 29920 0 1 22173
box 0 0 1 1
use contact_32  contact_32_2075
timestamp 1624857261
transform 1 0 29240 0 1 14013
box 0 0 1 1
use contact_32  contact_32_2074
timestamp 1624857261
transform 1 0 29240 0 1 15781
box 0 0 1 1
use contact_32  contact_32_2073
timestamp 1624857261
transform 1 0 28288 0 1 126213
box 0 0 1 1
use contact_32  contact_32_2072
timestamp 1624857261
transform 1 0 28288 0 1 125941
box 0 0 1 1
use contact_32  contact_32_2071
timestamp 1624857261
transform 1 0 28832 0 1 126349
box 0 0 1 1
use contact_32  contact_32_2070
timestamp 1624857261
transform 1 0 28832 0 1 128525
box 0 0 1 1
use contact_32  contact_32_2069
timestamp 1624857261
transform 1 0 28560 0 1 92485
box 0 0 1 1
use contact_32  contact_32_2068
timestamp 1624857261
transform 1 0 28560 0 1 92213
box 0 0 1 1
use contact_32  contact_32_2067
timestamp 1624857261
transform 1 0 28424 0 1 71269
box 0 0 1 1
use contact_32  contact_32_2066
timestamp 1624857261
transform 1 0 28424 0 1 70997
box 0 0 1 1
use contact_32  contact_32_2065
timestamp 1624857261
transform 1 0 28288 0 1 121453
box 0 0 1 1
use contact_32  contact_32_2064
timestamp 1624857261
transform 1 0 28288 0 1 121725
box 0 0 1 1
use contact_32  contact_32_2063
timestamp 1624857261
transform 1 0 28288 0 1 121317
box 0 0 1 1
use contact_32  contact_32_2062
timestamp 1624857261
transform 1 0 28288 0 1 121045
box 0 0 1 1
use contact_32  contact_32_2061
timestamp 1624857261
transform 1 0 28424 0 1 107581
box 0 0 1 1
use contact_32  contact_32_2060
timestamp 1624857261
transform 1 0 28424 0 1 107853
box 0 0 1 1
use contact_32  contact_32_2059
timestamp 1624857261
transform 1 0 28424 0 1 75485
box 0 0 1 1
use contact_32  contact_32_2058
timestamp 1624857261
transform 1 0 28424 0 1 75213
box 0 0 1 1
use contact_32  contact_32_2057
timestamp 1624857261
transform 1 0 28424 0 1 75621
box 0 0 1 1
use contact_32  contact_32_2056
timestamp 1624857261
transform 1 0 28424 0 1 75893
box 0 0 1 1
use contact_32  contact_32_2055
timestamp 1624857261
transform 1 0 28288 0 1 72901
box 0 0 1 1
use contact_32  contact_32_2054
timestamp 1624857261
transform 1 0 28288 0 1 72493
box 0 0 1 1
use contact_32  contact_32_2053
timestamp 1624857261
transform 1 0 28424 0 1 117373
box 0 0 1 1
use contact_32  contact_32_2052
timestamp 1624857261
transform 1 0 28424 0 1 117101
box 0 0 1 1
use contact_32  contact_32_2051
timestamp 1624857261
transform 1 0 28288 0 1 60253
box 0 0 1 1
use contact_32  contact_32_2050
timestamp 1624857261
transform 1 0 28288 0 1 59845
box 0 0 1 1
use contact_32  contact_32_2049
timestamp 1624857261
transform 1 0 28288 0 1 55085
box 0 0 1 1
use contact_32  contact_32_2048
timestamp 1624857261
transform 1 0 28288 0 1 55357
box 0 0 1 1
use contact_32  contact_32_2047
timestamp 1624857261
transform 1 0 28560 0 1 54949
box 0 0 1 1
use contact_32  contact_32_2046
timestamp 1624857261
transform 1 0 28560 0 1 54677
box 0 0 1 1
use contact_32  contact_32_2045
timestamp 1624857261
transform 1 0 28424 0 1 101597
box 0 0 1 1
use contact_32  contact_32_2044
timestamp 1624857261
transform 1 0 28424 0 1 101325
box 0 0 1 1
use contact_32  contact_32_2043
timestamp 1624857261
transform 1 0 28288 0 1 41213
box 0 0 1 1
use contact_32  contact_32_2042
timestamp 1624857261
transform 1 0 28288 0 1 41485
box 0 0 1 1
use contact_32  contact_32_2041
timestamp 1624857261
transform 1 0 28560 0 1 26525
box 0 0 1 1
use contact_32  contact_32_2040
timestamp 1624857261
transform 1 0 28560 0 1 26253
box 0 0 1 1
use contact_32  contact_32_2039
timestamp 1624857261
transform 1 0 28288 0 1 38493
box 0 0 1 1
use contact_32  contact_32_2038
timestamp 1624857261
transform 1 0 28288 0 1 38765
box 0 0 1 1
use contact_32  contact_32_2037
timestamp 1624857261
transform 1 0 28288 0 1 55493
box 0 0 1 1
use contact_32  contact_32_2036
timestamp 1624857261
transform 1 0 28288 0 1 55765
box 0 0 1 1
use contact_32  contact_32_2035
timestamp 1624857261
transform 1 0 28288 0 1 54405
box 0 0 1 1
use contact_32  contact_32_2034
timestamp 1624857261
transform 1 0 28288 0 1 54677
box 0 0 1 1
use contact_32  contact_32_2033
timestamp 1624857261
transform 1 0 28288 0 1 34141
box 0 0 1 1
use contact_32  contact_32_2032
timestamp 1624857261
transform 1 0 28288 0 1 34413
box 0 0 1 1
use contact_32  contact_32_2031
timestamp 1624857261
transform 1 0 28424 0 1 113021
box 0 0 1 1
use contact_32  contact_32_2030
timestamp 1624857261
transform 1 0 28424 0 1 112749
box 0 0 1 1
use contact_32  contact_32_2029
timestamp 1624857261
transform 1 0 28424 0 1 83373
box 0 0 1 1
use contact_32  contact_32_2028
timestamp 1624857261
transform 1 0 28424 0 1 83101
box 0 0 1 1
use contact_32  contact_32_2027
timestamp 1624857261
transform 1 0 28288 0 1 93437
box 0 0 1 1
use contact_32  contact_32_2026
timestamp 1624857261
transform 1 0 28288 0 1 93709
box 0 0 1 1
use contact_32  contact_32_2025
timestamp 1624857261
transform 1 0 28288 0 1 51141
box 0 0 1 1
use contact_32  contact_32_2024
timestamp 1624857261
transform 1 0 28288 0 1 51413
box 0 0 1 1
use contact_32  contact_32_2023
timestamp 1624857261
transform 1 0 28560 0 1 76301
box 0 0 1 1
use contact_32  contact_32_2022
timestamp 1624857261
transform 1 0 28560 0 1 76029
box 0 0 1 1
use contact_32  contact_32_2021
timestamp 1624857261
transform 1 0 28288 0 1 67325
box 0 0 1 1
use contact_32  contact_32_2020
timestamp 1624857261
transform 1 0 28288 0 1 67597
box 0 0 1 1
use contact_32  contact_32_2019
timestamp 1624857261
transform 1 0 28424 0 1 88541
box 0 0 1 1
use contact_32  contact_32_2018
timestamp 1624857261
transform 1 0 28424 0 1 88269
box 0 0 1 1
use contact_32  contact_32_2017
timestamp 1624857261
transform 1 0 28560 0 1 70725
box 0 0 1 1
use contact_32  contact_32_2016
timestamp 1624857261
transform 1 0 28560 0 1 70453
box 0 0 1 1
use contact_32  contact_32_2015
timestamp 1624857261
transform 1 0 28288 0 1 46789
box 0 0 1 1
use contact_32  contact_32_2014
timestamp 1624857261
transform 1 0 28288 0 1 47061
box 0 0 1 1
use contact_32  contact_32_2013
timestamp 1624857261
transform 1 0 28424 0 1 80789
box 0 0 1 1
use contact_32  contact_32_2012
timestamp 1624857261
transform 1 0 28424 0 1 80381
box 0 0 1 1
use contact_32  contact_32_2011
timestamp 1624857261
transform 1 0 28288 0 1 120501
box 0 0 1 1
use contact_32  contact_32_2010
timestamp 1624857261
transform 1 0 28288 0 1 120229
box 0 0 1 1
use contact_32  contact_32_2009
timestamp 1624857261
transform 1 0 28424 0 1 67733
box 0 0 1 1
use contact_32  contact_32_2008
timestamp 1624857261
transform 1 0 28424 0 1 68005
box 0 0 1 1
use contact_32  contact_32_2007
timestamp 1624857261
transform 1 0 28560 0 1 116693
box 0 0 1 1
use contact_32  contact_32_2006
timestamp 1624857261
transform 1 0 28560 0 1 116965
box 0 0 1 1
use contact_32  contact_32_2005
timestamp 1624857261
transform 1 0 28424 0 1 116557
box 0 0 1 1
use contact_32  contact_32_2004
timestamp 1624857261
transform 1 0 28424 0 1 116285
box 0 0 1 1
use contact_32  contact_32_2003
timestamp 1624857261
transform 1 0 28424 0 1 58077
box 0 0 1 1
use contact_32  contact_32_2002
timestamp 1624857261
transform 1 0 28424 0 1 57805
box 0 0 1 1
use contact_32  contact_32_2001
timestamp 1624857261
transform 1 0 28424 0 1 63381
box 0 0 1 1
use contact_32  contact_32_2000
timestamp 1624857261
transform 1 0 28424 0 1 63653
box 0 0 1 1
use contact_32  contact_32_1999
timestamp 1624857261
transform 1 0 28560 0 1 80789
box 0 0 1 1
use contact_32  contact_32_1998
timestamp 1624857261
transform 1 0 28560 0 1 81061
box 0 0 1 1
use contact_32  contact_32_1997
timestamp 1624857261
transform 1 0 28424 0 1 34549
box 0 0 1 1
use contact_32  contact_32_1996
timestamp 1624857261
transform 1 0 28424 0 1 34821
box 0 0 1 1
use contact_32  contact_32_1995
timestamp 1624857261
transform 1 0 28560 0 1 31285
box 0 0 1 1
use contact_32  contact_32_1994
timestamp 1624857261
transform 1 0 28560 0 1 31013
box 0 0 1 1
use contact_32  contact_32_1993
timestamp 1624857261
transform 1 0 28288 0 1 125805
box 0 0 1 1
use contact_32  contact_32_1992
timestamp 1624857261
transform 1 0 28288 0 1 125397
box 0 0 1 1
use contact_32  contact_32_1991
timestamp 1624857261
transform 1 0 28288 0 1 108397
box 0 0 1 1
use contact_32  contact_32_1990
timestamp 1624857261
transform 1 0 28288 0 1 108669
box 0 0 1 1
use contact_32  contact_32_1989
timestamp 1624857261
transform 1 0 28424 0 1 84189
box 0 0 1 1
use contact_32  contact_32_1988
timestamp 1624857261
transform 1 0 28424 0 1 84461
box 0 0 1 1
use contact_32  contact_32_1987
timestamp 1624857261
transform 1 0 28288 0 1 36045
box 0 0 1 1
use contact_32  contact_32_1986
timestamp 1624857261
transform 1 0 28288 0 1 35773
box 0 0 1 1
use contact_32  contact_32_1985
timestamp 1624857261
transform 1 0 28288 0 1 80245
box 0 0 1 1
use contact_32  contact_32_1984
timestamp 1624857261
transform 1 0 28288 0 1 79973
box 0 0 1 1
use contact_32  contact_32_1983
timestamp 1624857261
transform 1 0 28288 0 1 25437
box 0 0 1 1
use contact_32  contact_32_1982
timestamp 1624857261
transform 1 0 28288 0 1 25709
box 0 0 1 1
use contact_32  contact_32_1981
timestamp 1624857261
transform 1 0 28424 0 1 25845
box 0 0 1 1
use contact_32  contact_32_1980
timestamp 1624857261
transform 1 0 28424 0 1 26117
box 0 0 1 1
use contact_32  contact_32_1979
timestamp 1624857261
transform 1 0 28424 0 1 79973
box 0 0 1 1
use contact_32  contact_32_1978
timestamp 1624857261
transform 1 0 28424 0 1 79565
box 0 0 1 1
use contact_32  contact_32_1977
timestamp 1624857261
transform 1 0 28560 0 1 89765
box 0 0 1 1
use contact_32  contact_32_1976
timestamp 1624857261
transform 1 0 28560 0 1 89493
box 0 0 1 1
use contact_32  contact_32_1975
timestamp 1624857261
transform 1 0 28560 0 1 105541
box 0 0 1 1
use contact_32  contact_32_1974
timestamp 1624857261
transform 1 0 28560 0 1 105269
box 0 0 1 1
use contact_32  contact_32_1973
timestamp 1624857261
transform 1 0 28560 0 1 72357
box 0 0 1 1
use contact_32  contact_32_1972
timestamp 1624857261
transform 1 0 28560 0 1 72085
box 0 0 1 1
use contact_32  contact_32_1971
timestamp 1624857261
transform 1 0 28560 0 1 59301
box 0 0 1 1
use contact_32  contact_32_1970
timestamp 1624857261
transform 1 0 28560 0 1 59029
box 0 0 1 1
use contact_32  contact_32_1969
timestamp 1624857261
transform 1 0 28424 0 1 120909
box 0 0 1 1
use contact_32  contact_32_1968
timestamp 1624857261
transform 1 0 28424 0 1 120501
box 0 0 1 1
use contact_32  contact_32_1967
timestamp 1624857261
transform 1 0 28288 0 1 111797
box 0 0 1 1
use contact_32  contact_32_1966
timestamp 1624857261
transform 1 0 28288 0 1 111525
box 0 0 1 1
use contact_32  contact_32_1965
timestamp 1624857261
transform 1 0 28288 0 1 66509
box 0 0 1 1
use contact_32  contact_32_1964
timestamp 1624857261
transform 1 0 28288 0 1 66781
box 0 0 1 1
use contact_32  contact_32_1963
timestamp 1624857261
transform 1 0 28424 0 1 87045
box 0 0 1 1
use contact_32  contact_32_1962
timestamp 1624857261
transform 1 0 28424 0 1 87317
box 0 0 1 1
use contact_32  contact_32_1961
timestamp 1624857261
transform 1 0 28560 0 1 96837
box 0 0 1 1
use contact_32  contact_32_1960
timestamp 1624857261
transform 1 0 28560 0 1 96565
box 0 0 1 1
use contact_32  contact_32_1959
timestamp 1624857261
transform 1 0 28288 0 1 49917
box 0 0 1 1
use contact_32  contact_32_1958
timestamp 1624857261
transform 1 0 28288 0 1 50189
box 0 0 1 1
use contact_32  contact_32_1957
timestamp 1624857261
transform 1 0 28424 0 1 108805
box 0 0 1 1
use contact_32  contact_32_1956
timestamp 1624857261
transform 1 0 28424 0 1 109077
box 0 0 1 1
use contact_32  contact_32_1955
timestamp 1624857261
transform 1 0 28560 0 1 84189
box 0 0 1 1
use contact_32  contact_32_1954
timestamp 1624857261
transform 1 0 28560 0 1 83917
box 0 0 1 1
use contact_32  contact_32_1953
timestamp 1624857261
transform 1 0 28560 0 1 79157
box 0 0 1 1
use contact_32  contact_32_1952
timestamp 1624857261
transform 1 0 28560 0 1 79429
box 0 0 1 1
use contact_32  contact_32_1951
timestamp 1624857261
transform 1 0 28560 0 1 114245
box 0 0 1 1
use contact_32  contact_32_1950
timestamp 1624857261
transform 1 0 28560 0 1 113973
box 0 0 1 1
use contact_32  contact_32_1949
timestamp 1624857261
transform 1 0 28560 0 1 71949
box 0 0 1 1
use contact_32  contact_32_1948
timestamp 1624857261
transform 1 0 28560 0 1 71677
box 0 0 1 1
use contact_32  contact_32_1947
timestamp 1624857261
transform 1 0 28288 0 1 39717
box 0 0 1 1
use contact_32  contact_32_1946
timestamp 1624857261
transform 1 0 28288 0 1 39989
box 0 0 1 1
use contact_32  contact_32_1945
timestamp 1624857261
transform 1 0 28288 0 1 43117
box 0 0 1 1
use contact_32  contact_32_1944
timestamp 1624857261
transform 1 0 28288 0 1 42845
box 0 0 1 1
use contact_32  contact_32_1943
timestamp 1624857261
transform 1 0 28288 0 1 62973
box 0 0 1 1
use contact_32  contact_32_1942
timestamp 1624857261
transform 1 0 28288 0 1 63381
box 0 0 1 1
use contact_32  contact_32_1941
timestamp 1624857261
transform 1 0 28424 0 1 124989
box 0 0 1 1
use contact_32  contact_32_1940
timestamp 1624857261
transform 1 0 28424 0 1 125261
box 0 0 1 1
use contact_32  contact_32_1939
timestamp 1624857261
transform 1 0 28288 0 1 117373
box 0 0 1 1
use contact_32  contact_32_1938
timestamp 1624857261
transform 1 0 28288 0 1 117645
box 0 0 1 1
use contact_32  contact_32_1937
timestamp 1624857261
transform 1 0 28560 0 1 83781
box 0 0 1 1
use contact_32  contact_32_1936
timestamp 1624857261
transform 1 0 28560 0 1 83373
box 0 0 1 1
use contact_32  contact_32_1935
timestamp 1624857261
transform 1 0 28288 0 1 84733
box 0 0 1 1
use contact_32  contact_32_1934
timestamp 1624857261
transform 1 0 28288 0 1 85005
box 0 0 1 1
use contact_32  contact_32_1933
timestamp 1624857261
transform 1 0 28288 0 1 42437
box 0 0 1 1
use contact_32  contact_32_1932
timestamp 1624857261
transform 1 0 28288 0 1 42709
box 0 0 1 1
use contact_32  contact_32_1931
timestamp 1624857261
transform 1 0 28560 0 1 42437
box 0 0 1 1
use contact_32  contact_32_1930
timestamp 1624857261
transform 1 0 28560 0 1 42845
box 0 0 1 1
use contact_32  contact_32_1929
timestamp 1624857261
transform 1 0 28424 0 1 105133
box 0 0 1 1
use contact_32  contact_32_1928
timestamp 1624857261
transform 1 0 28424 0 1 104861
box 0 0 1 1
use contact_32  contact_32_1927
timestamp 1624857261
transform 1 0 28424 0 1 96429
box 0 0 1 1
use contact_32  contact_32_1926
timestamp 1624857261
transform 1 0 28424 0 1 96157
box 0 0 1 1
use contact_32  contact_32_1925
timestamp 1624857261
transform 1 0 28560 0 1 88133
box 0 0 1 1
use contact_32  contact_32_1924
timestamp 1624857261
transform 1 0 28560 0 1 87861
box 0 0 1 1
use contact_32  contact_32_1923
timestamp 1624857261
transform 1 0 28424 0 1 95749
box 0 0 1 1
use contact_32  contact_32_1922
timestamp 1624857261
transform 1 0 28424 0 1 96021
box 0 0 1 1
use contact_32  contact_32_1921
timestamp 1624857261
transform 1 0 28560 0 1 125669
box 0 0 1 1
use contact_32  contact_32_1920
timestamp 1624857261
transform 1 0 28560 0 1 125397
box 0 0 1 1
use contact_32  contact_32_1919
timestamp 1624857261
transform 1 0 28560 0 1 58893
box 0 0 1 1
use contact_32  contact_32_1918
timestamp 1624857261
transform 1 0 28560 0 1 58621
box 0 0 1 1
use contact_32  contact_32_1917
timestamp 1624857261
transform 1 0 28288 0 1 51549
box 0 0 1 1
use contact_32  contact_32_1916
timestamp 1624857261
transform 1 0 28288 0 1 51821
box 0 0 1 1
use contact_32  contact_32_1915
timestamp 1624857261
transform 1 0 28288 0 1 70725
box 0 0 1 1
use contact_32  contact_32_1914
timestamp 1624857261
transform 1 0 28288 0 1 71133
box 0 0 1 1
use contact_32  contact_32_1913
timestamp 1624857261
transform 1 0 28288 0 1 113701
box 0 0 1 1
use contact_32  contact_32_1912
timestamp 1624857261
transform 1 0 28288 0 1 113429
box 0 0 1 1
use contact_32  contact_32_1911
timestamp 1624857261
transform 1 0 28424 0 1 33869
box 0 0 1 1
use contact_32  contact_32_1910
timestamp 1624857261
transform 1 0 28424 0 1 34141
box 0 0 1 1
use contact_32  contact_32_1909
timestamp 1624857261
transform 1 0 28560 0 1 64469
box 0 0 1 1
use contact_32  contact_32_1908
timestamp 1624857261
transform 1 0 28560 0 1 64197
box 0 0 1 1
use contact_32  contact_32_1907
timestamp 1624857261
transform 1 0 28832 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1906
timestamp 1624857261
transform 1 0 28832 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1905
timestamp 1624857261
transform 1 0 28968 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1904
timestamp 1624857261
transform 1 0 28968 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1903
timestamp 1624857261
transform 1 0 29784 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1902
timestamp 1624857261
transform 1 0 29784 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1901
timestamp 1624857261
transform 1 0 29784 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1900
timestamp 1624857261
transform 1 0 29784 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1899
timestamp 1624857261
transform 1 0 30056 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1898
timestamp 1624857261
transform 1 0 30056 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1897
timestamp 1624857261
transform 1 0 29920 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1896
timestamp 1624857261
transform 1 0 29920 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1895
timestamp 1624857261
transform 1 0 29920 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1894
timestamp 1624857261
transform 1 0 29920 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1893
timestamp 1624857261
transform 1 0 29920 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1892
timestamp 1624857261
transform 1 0 29920 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1891
timestamp 1624857261
transform 1 0 30464 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1890
timestamp 1624857261
transform 1 0 30464 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1889
timestamp 1624857261
transform 1 0 30464 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1888
timestamp 1624857261
transform 1 0 30464 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1887
timestamp 1624857261
transform 1 0 32368 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1886
timestamp 1624857261
transform 1 0 32368 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1885
timestamp 1624857261
transform 1 0 32232 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1884
timestamp 1624857261
transform 1 0 32232 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1883
timestamp 1624857261
transform 1 0 33864 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1882
timestamp 1624857261
transform 1 0 33864 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1881
timestamp 1624857261
transform 1 0 33864 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1880
timestamp 1624857261
transform 1 0 33864 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1879
timestamp 1624857261
transform 1 0 34952 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1878
timestamp 1624857261
transform 1 0 34952 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1877
timestamp 1624857261
transform 1 0 34952 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1876
timestamp 1624857261
transform 1 0 34952 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1875
timestamp 1624857261
transform 1 0 34816 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1874
timestamp 1624857261
transform 1 0 34816 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1873
timestamp 1624857261
transform 1 0 34952 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1872
timestamp 1624857261
transform 1 0 34952 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1871
timestamp 1624857261
transform 1 0 35088 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1870
timestamp 1624857261
transform 1 0 35088 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1869
timestamp 1624857261
transform 1 0 34952 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1868
timestamp 1624857261
transform 1 0 34952 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1867
timestamp 1624857261
transform 1 0 35496 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1866
timestamp 1624857261
transform 1 0 35496 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1865
timestamp 1624857261
transform 1 0 35496 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1864
timestamp 1624857261
transform 1 0 35496 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1863
timestamp 1624857261
transform 1 0 37400 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1862
timestamp 1624857261
transform 1 0 37400 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1861
timestamp 1624857261
transform 1 0 37264 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1860
timestamp 1624857261
transform 1 0 37264 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1859
timestamp 1624857261
transform 1 0 38896 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1858
timestamp 1624857261
transform 1 0 38896 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1857
timestamp 1624857261
transform 1 0 38896 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1856
timestamp 1624857261
transform 1 0 38896 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1855
timestamp 1624857261
transform 1 0 39848 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1854
timestamp 1624857261
transform 1 0 39848 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1853
timestamp 1624857261
transform 1 0 39848 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1852
timestamp 1624857261
transform 1 0 39848 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1851
timestamp 1624857261
transform 1 0 39848 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1850
timestamp 1624857261
transform 1 0 39848 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1849
timestamp 1624857261
transform 1 0 39848 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1848
timestamp 1624857261
transform 1 0 39848 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1847
timestamp 1624857261
transform 1 0 39984 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1846
timestamp 1624857261
transform 1 0 39984 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1845
timestamp 1624857261
transform 1 0 39984 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1844
timestamp 1624857261
transform 1 0 39984 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1843
timestamp 1624857261
transform 1 0 40664 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1842
timestamp 1624857261
transform 1 0 40664 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1841
timestamp 1624857261
transform 1 0 40800 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1840
timestamp 1624857261
transform 1 0 40800 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1839
timestamp 1624857261
transform 1 0 42432 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1838
timestamp 1624857261
transform 1 0 42432 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1837
timestamp 1624857261
transform 1 0 42432 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1836
timestamp 1624857261
transform 1 0 42432 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1835
timestamp 1624857261
transform 1 0 43928 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1834
timestamp 1624857261
transform 1 0 43928 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1833
timestamp 1624857261
transform 1 0 43928 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1832
timestamp 1624857261
transform 1 0 43928 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1831
timestamp 1624857261
transform 1 0 44608 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1830
timestamp 1624857261
transform 1 0 44608 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1829
timestamp 1624857261
transform 1 0 44744 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1828
timestamp 1624857261
transform 1 0 44744 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1827
timestamp 1624857261
transform 1 0 44880 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1826
timestamp 1624857261
transform 1 0 44880 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1825
timestamp 1624857261
transform 1 0 45016 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1824
timestamp 1624857261
transform 1 0 45016 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1823
timestamp 1624857261
transform 1 0 44880 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1822
timestamp 1624857261
transform 1 0 44880 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1821
timestamp 1624857261
transform 1 0 44880 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1820
timestamp 1624857261
transform 1 0 44880 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1819
timestamp 1624857261
transform 1 0 45696 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1818
timestamp 1624857261
transform 1 0 45696 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1817
timestamp 1624857261
transform 1 0 45696 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1816
timestamp 1624857261
transform 1 0 45696 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1815
timestamp 1624857261
transform 1 0 47464 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1814
timestamp 1624857261
transform 1 0 47464 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1813
timestamp 1624857261
transform 1 0 47464 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1812
timestamp 1624857261
transform 1 0 47464 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1811
timestamp 1624857261
transform 1 0 48960 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1810
timestamp 1624857261
transform 1 0 48960 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1809
timestamp 1624857261
transform 1 0 48960 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1808
timestamp 1624857261
transform 1 0 48960 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1807
timestamp 1624857261
transform 1 0 49912 0 1 15917
box 0 0 1 1
use contact_32  contact_32_1806
timestamp 1624857261
transform 1 0 49912 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1805
timestamp 1624857261
transform 1 0 50048 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1804
timestamp 1624857261
transform 1 0 50048 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1803
timestamp 1624857261
transform 1 0 49912 0 1 17141
box 0 0 1 1
use contact_32  contact_32_1802
timestamp 1624857261
transform 1 0 49912 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1801
timestamp 1624857261
transform 1 0 49912 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1800
timestamp 1624857261
transform 1 0 49912 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1799
timestamp 1624857261
transform 1 0 49912 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1798
timestamp 1624857261
transform 1 0 49912 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1797
timestamp 1624857261
transform 1 0 49912 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1796
timestamp 1624857261
transform 1 0 49912 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1795
timestamp 1624857261
transform 1 0 50048 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1794
timestamp 1624857261
transform 1 0 50048 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1793
timestamp 1624857261
transform 1 0 50728 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1792
timestamp 1624857261
transform 1 0 50728 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1791
timestamp 1624857261
transform 1 0 50728 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1790
timestamp 1624857261
transform 1 0 50728 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1789
timestamp 1624857261
transform 1 0 52360 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1788
timestamp 1624857261
transform 1 0 52360 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1787
timestamp 1624857261
transform 1 0 52360 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1786
timestamp 1624857261
transform 1 0 52360 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1785
timestamp 1624857261
transform 1 0 54808 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1784
timestamp 1624857261
transform 1 0 54808 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1783
timestamp 1624857261
transform 1 0 53992 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1782
timestamp 1624857261
transform 1 0 53992 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1781
timestamp 1624857261
transform 1 0 54128 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1780
timestamp 1624857261
transform 1 0 54128 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1779
timestamp 1624857261
transform 1 0 54944 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1778
timestamp 1624857261
transform 1 0 54944 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1777
timestamp 1624857261
transform 1 0 54944 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1776
timestamp 1624857261
transform 1 0 54944 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1775
timestamp 1624857261
transform 1 0 54808 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1774
timestamp 1624857261
transform 1 0 54808 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1773
timestamp 1624857261
transform 1 0 54944 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1772
timestamp 1624857261
transform 1 0 54944 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1771
timestamp 1624857261
transform 1 0 55080 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1770
timestamp 1624857261
transform 1 0 55080 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1769
timestamp 1624857261
transform 1 0 55896 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1768
timestamp 1624857261
transform 1 0 55896 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1767
timestamp 1624857261
transform 1 0 55896 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1766
timestamp 1624857261
transform 1 0 55896 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1765
timestamp 1624857261
transform 1 0 57392 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1764
timestamp 1624857261
transform 1 0 57392 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1763
timestamp 1624857261
transform 1 0 57664 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1762
timestamp 1624857261
transform 1 0 57664 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1761
timestamp 1624857261
transform 1 0 59704 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1760
timestamp 1624857261
transform 1 0 59704 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1759
timestamp 1624857261
transform 1 0 59160 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1758
timestamp 1624857261
transform 1 0 59160 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1757
timestamp 1624857261
transform 1 0 59160 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1756
timestamp 1624857261
transform 1 0 59160 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1755
timestamp 1624857261
transform 1 0 59568 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1754
timestamp 1624857261
transform 1 0 59568 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1753
timestamp 1624857261
transform 1 0 59704 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1752
timestamp 1624857261
transform 1 0 59704 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1751
timestamp 1624857261
transform 1 0 59976 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1750
timestamp 1624857261
transform 1 0 59976 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1749
timestamp 1624857261
transform 1 0 59840 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1748
timestamp 1624857261
transform 1 0 59840 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1747
timestamp 1624857261
transform 1 0 59976 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1746
timestamp 1624857261
transform 1 0 59976 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1745
timestamp 1624857261
transform 1 0 61064 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1744
timestamp 1624857261
transform 1 0 61064 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1743
timestamp 1624857261
transform 1 0 60928 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1742
timestamp 1624857261
transform 1 0 60928 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1741
timestamp 1624857261
transform 1 0 62424 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1740
timestamp 1624857261
transform 1 0 62424 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1739
timestamp 1624857261
transform 1 0 62424 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1738
timestamp 1624857261
transform 1 0 62424 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1737
timestamp 1624857261
transform 1 0 64056 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1736
timestamp 1624857261
transform 1 0 64056 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1735
timestamp 1624857261
transform 1 0 64056 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1734
timestamp 1624857261
transform 1 0 64056 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1733
timestamp 1624857261
transform 1 0 64872 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1732
timestamp 1624857261
transform 1 0 64872 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1731
timestamp 1624857261
transform 1 0 64872 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1730
timestamp 1624857261
transform 1 0 64872 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1729
timestamp 1624857261
transform 1 0 65008 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1728
timestamp 1624857261
transform 1 0 65008 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1727
timestamp 1624857261
transform 1 0 64736 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1726
timestamp 1624857261
transform 1 0 64736 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1725
timestamp 1624857261
transform 1 0 64872 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1724
timestamp 1624857261
transform 1 0 64872 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1723
timestamp 1624857261
transform 1 0 64872 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1722
timestamp 1624857261
transform 1 0 64872 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1721
timestamp 1624857261
transform 1 0 65960 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1720
timestamp 1624857261
transform 1 0 65960 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1719
timestamp 1624857261
transform 1 0 65960 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1718
timestamp 1624857261
transform 1 0 65960 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1717
timestamp 1624857261
transform 1 0 67456 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1716
timestamp 1624857261
transform 1 0 67456 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1715
timestamp 1624857261
transform 1 0 67456 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1714
timestamp 1624857261
transform 1 0 67456 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1713
timestamp 1624857261
transform 1 0 69360 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1712
timestamp 1624857261
transform 1 0 69360 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1711
timestamp 1624857261
transform 1 0 69224 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1710
timestamp 1624857261
transform 1 0 69224 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1709
timestamp 1624857261
transform 1 0 69904 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1708
timestamp 1624857261
transform 1 0 69904 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1707
timestamp 1624857261
transform 1 0 69904 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1706
timestamp 1624857261
transform 1 0 69904 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1705
timestamp 1624857261
transform 1 0 69904 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1704
timestamp 1624857261
transform 1 0 69904 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1703
timestamp 1624857261
transform 1 0 69904 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1702
timestamp 1624857261
transform 1 0 69904 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1701
timestamp 1624857261
transform 1 0 69904 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1700
timestamp 1624857261
transform 1 0 69904 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1699
timestamp 1624857261
transform 1 0 70040 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1698
timestamp 1624857261
transform 1 0 70040 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1697
timestamp 1624857261
transform 1 0 70856 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1696
timestamp 1624857261
transform 1 0 70856 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1695
timestamp 1624857261
transform 1 0 70856 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1694
timestamp 1624857261
transform 1 0 70856 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1693
timestamp 1624857261
transform 1 0 72488 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1692
timestamp 1624857261
transform 1 0 72488 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1691
timestamp 1624857261
transform 1 0 72488 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1690
timestamp 1624857261
transform 1 0 72488 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1689
timestamp 1624857261
transform 1 0 74256 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1688
timestamp 1624857261
transform 1 0 74256 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1687
timestamp 1624857261
transform 1 0 74256 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1686
timestamp 1624857261
transform 1 0 74256 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1685
timestamp 1624857261
transform 1 0 74664 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1684
timestamp 1624857261
transform 1 0 74664 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1683
timestamp 1624857261
transform 1 0 74664 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1682
timestamp 1624857261
transform 1 0 74664 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1681
timestamp 1624857261
transform 1 0 74800 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1680
timestamp 1624857261
transform 1 0 74800 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1679
timestamp 1624857261
transform 1 0 74936 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1678
timestamp 1624857261
transform 1 0 74936 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1677
timestamp 1624857261
transform 1 0 75072 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1676
timestamp 1624857261
transform 1 0 75072 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1675
timestamp 1624857261
transform 1 0 74936 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1674
timestamp 1624857261
transform 1 0 74936 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1673
timestamp 1624857261
transform 1 0 75888 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1672
timestamp 1624857261
transform 1 0 75888 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1671
timestamp 1624857261
transform 1 0 75888 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1670
timestamp 1624857261
transform 1 0 75888 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1669
timestamp 1624857261
transform 1 0 77656 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1668
timestamp 1624857261
transform 1 0 77656 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1667
timestamp 1624857261
transform 1 0 77656 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1666
timestamp 1624857261
transform 1 0 77656 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1665
timestamp 1624857261
transform 1 0 79424 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1664
timestamp 1624857261
transform 1 0 79424 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1663
timestamp 1624857261
transform 1 0 79288 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1662
timestamp 1624857261
transform 1 0 79288 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1661
timestamp 1624857261
transform 1 0 79288 0 1 16053
box 0 0 1 1
use contact_32  contact_32_1660
timestamp 1624857261
transform 1 0 79288 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1659
timestamp 1624857261
transform 1 0 79968 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1658
timestamp 1624857261
transform 1 0 79968 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1657
timestamp 1624857261
transform 1 0 79696 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1656
timestamp 1624857261
transform 1 0 79696 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1655
timestamp 1624857261
transform 1 0 79968 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1654
timestamp 1624857261
transform 1 0 79968 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1653
timestamp 1624857261
transform 1 0 79832 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1652
timestamp 1624857261
transform 1 0 79832 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1651
timestamp 1624857261
transform 1 0 79832 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1650
timestamp 1624857261
transform 1 0 79832 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1649
timestamp 1624857261
transform 1 0 79832 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1648
timestamp 1624857261
transform 1 0 79832 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1647
timestamp 1624857261
transform 1 0 80920 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1646
timestamp 1624857261
transform 1 0 80920 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1645
timestamp 1624857261
transform 1 0 80920 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1644
timestamp 1624857261
transform 1 0 80920 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1643
timestamp 1624857261
transform 1 0 82688 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1642
timestamp 1624857261
transform 1 0 82688 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1641
timestamp 1624857261
transform 1 0 82688 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1640
timestamp 1624857261
transform 1 0 82688 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1639
timestamp 1624857261
transform 1 0 84592 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1638
timestamp 1624857261
transform 1 0 84592 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1637
timestamp 1624857261
transform 1 0 84592 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1636
timestamp 1624857261
transform 1 0 84592 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1635
timestamp 1624857261
transform 1 0 84864 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1634
timestamp 1624857261
transform 1 0 84864 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1633
timestamp 1624857261
transform 1 0 84864 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1632
timestamp 1624857261
transform 1 0 84864 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1631
timestamp 1624857261
transform 1 0 84864 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1630
timestamp 1624857261
transform 1 0 84864 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1629
timestamp 1624857261
transform 1 0 84864 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1628
timestamp 1624857261
transform 1 0 84864 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1627
timestamp 1624857261
transform 1 0 84864 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1626
timestamp 1624857261
transform 1 0 84864 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1625
timestamp 1624857261
transform 1 0 85000 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1624
timestamp 1624857261
transform 1 0 85000 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1623
timestamp 1624857261
transform 1 0 85952 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1622
timestamp 1624857261
transform 1 0 85952 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1621
timestamp 1624857261
transform 1 0 85952 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1620
timestamp 1624857261
transform 1 0 85952 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1619
timestamp 1624857261
transform 1 0 87720 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1618
timestamp 1624857261
transform 1 0 87720 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1617
timestamp 1624857261
transform 1 0 87720 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1616
timestamp 1624857261
transform 1 0 87720 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1615
timestamp 1624857261
transform 1 0 89488 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1614
timestamp 1624857261
transform 1 0 89488 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1613
timestamp 1624857261
transform 1 0 89488 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1612
timestamp 1624857261
transform 1 0 89488 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1611
timestamp 1624857261
transform 1 0 89624 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1610
timestamp 1624857261
transform 1 0 89624 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1609
timestamp 1624857261
transform 1 0 89624 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1608
timestamp 1624857261
transform 1 0 89624 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1607
timestamp 1624857261
transform 1 0 89896 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1606
timestamp 1624857261
transform 1 0 89896 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1605
timestamp 1624857261
transform 1 0 89896 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1604
timestamp 1624857261
transform 1 0 89896 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1603
timestamp 1624857261
transform 1 0 89896 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1602
timestamp 1624857261
transform 1 0 89896 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1601
timestamp 1624857261
transform 1 0 90032 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1600
timestamp 1624857261
transform 1 0 90032 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1599
timestamp 1624857261
transform 1 0 91120 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1598
timestamp 1624857261
transform 1 0 91120 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1597
timestamp 1624857261
transform 1 0 90984 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1596
timestamp 1624857261
transform 1 0 90984 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1595
timestamp 1624857261
transform 1 0 92616 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1594
timestamp 1624857261
transform 1 0 92616 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1593
timestamp 1624857261
transform 1 0 92888 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1592
timestamp 1624857261
transform 1 0 92888 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1591
timestamp 1624857261
transform 1 0 94384 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1590
timestamp 1624857261
transform 1 0 94384 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1589
timestamp 1624857261
transform 1 0 94656 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1588
timestamp 1624857261
transform 1 0 94656 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1587
timestamp 1624857261
transform 1 0 94928 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1586
timestamp 1624857261
transform 1 0 94928 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1585
timestamp 1624857261
transform 1 0 94656 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1584
timestamp 1624857261
transform 1 0 94656 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1583
timestamp 1624857261
transform 1 0 94928 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1582
timestamp 1624857261
transform 1 0 94928 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1581
timestamp 1624857261
transform 1 0 94928 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1580
timestamp 1624857261
transform 1 0 94928 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1579
timestamp 1624857261
transform 1 0 94792 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1578
timestamp 1624857261
transform 1 0 94792 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1577
timestamp 1624857261
transform 1 0 94928 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1576
timestamp 1624857261
transform 1 0 94928 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1575
timestamp 1624857261
transform 1 0 96152 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1574
timestamp 1624857261
transform 1 0 96152 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1573
timestamp 1624857261
transform 1 0 96152 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1572
timestamp 1624857261
transform 1 0 96152 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1571
timestamp 1624857261
transform 1 0 97784 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1570
timestamp 1624857261
transform 1 0 97784 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1569
timestamp 1624857261
transform 1 0 97784 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1568
timestamp 1624857261
transform 1 0 97784 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1567
timestamp 1624857261
transform 1 0 99552 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1566
timestamp 1624857261
transform 1 0 99552 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1565
timestamp 1624857261
transform 1 0 99552 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1564
timestamp 1624857261
transform 1 0 99552 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1563
timestamp 1624857261
transform 1 0 99688 0 1 16053
box 0 0 1 1
use contact_32  contact_32_1562
timestamp 1624857261
transform 1 0 99688 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1561
timestamp 1624857261
transform 1 0 99824 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1560
timestamp 1624857261
transform 1 0 99824 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1559
timestamp 1624857261
transform 1 0 99688 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1558
timestamp 1624857261
transform 1 0 99688 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1557
timestamp 1624857261
transform 1 0 99824 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1556
timestamp 1624857261
transform 1 0 99824 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1555
timestamp 1624857261
transform 1 0 99824 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1554
timestamp 1624857261
transform 1 0 99824 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1553
timestamp 1624857261
transform 1 0 99960 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1552
timestamp 1624857261
transform 1 0 99960 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1551
timestamp 1624857261
transform 1 0 99824 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1550
timestamp 1624857261
transform 1 0 99824 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1549
timestamp 1624857261
transform 1 0 101184 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1548
timestamp 1624857261
transform 1 0 101184 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1547
timestamp 1624857261
transform 1 0 101184 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1546
timestamp 1624857261
transform 1 0 101184 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1545
timestamp 1624857261
transform 1 0 102952 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1544
timestamp 1624857261
transform 1 0 102952 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1543
timestamp 1624857261
transform 1 0 102952 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1542
timestamp 1624857261
transform 1 0 102952 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1541
timestamp 1624857261
transform 1 0 104448 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1540
timestamp 1624857261
transform 1 0 104448 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1539
timestamp 1624857261
transform 1 0 104448 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1538
timestamp 1624857261
transform 1 0 104448 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1537
timestamp 1624857261
transform 1 0 104448 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1536
timestamp 1624857261
transform 1 0 104448 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1535
timestamp 1624857261
transform 1 0 104584 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1534
timestamp 1624857261
transform 1 0 104584 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1533
timestamp 1624857261
transform 1 0 104856 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1532
timestamp 1624857261
transform 1 0 104856 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1531
timestamp 1624857261
transform 1 0 104720 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1530
timestamp 1624857261
transform 1 0 104720 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1529
timestamp 1624857261
transform 1 0 104856 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1528
timestamp 1624857261
transform 1 0 104856 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1527
timestamp 1624857261
transform 1 0 104992 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1526
timestamp 1624857261
transform 1 0 104992 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1525
timestamp 1624857261
transform 1 0 106216 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1524
timestamp 1624857261
transform 1 0 106216 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1523
timestamp 1624857261
transform 1 0 106216 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1522
timestamp 1624857261
transform 1 0 106216 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1521
timestamp 1624857261
transform 1 0 107848 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1520
timestamp 1624857261
transform 1 0 107848 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1519
timestamp 1624857261
transform 1 0 107848 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1518
timestamp 1624857261
transform 1 0 107848 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1517
timestamp 1624857261
transform 1 0 109616 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1516
timestamp 1624857261
transform 1 0 109616 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1515
timestamp 1624857261
transform 1 0 109480 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1514
timestamp 1624857261
transform 1 0 109480 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1513
timestamp 1624857261
transform 1 0 109480 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1512
timestamp 1624857261
transform 1 0 109480 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1511
timestamp 1624857261
transform 1 0 109616 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1510
timestamp 1624857261
transform 1 0 109616 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1509
timestamp 1624857261
transform 1 0 109888 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1508
timestamp 1624857261
transform 1 0 109888 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1507
timestamp 1624857261
transform 1 0 109888 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1506
timestamp 1624857261
transform 1 0 109888 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1505
timestamp 1624857261
transform 1 0 110024 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1504
timestamp 1624857261
transform 1 0 110024 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1503
timestamp 1624857261
transform 1 0 109888 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1502
timestamp 1624857261
transform 1 0 109888 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1501
timestamp 1624857261
transform 1 0 111112 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1500
timestamp 1624857261
transform 1 0 111112 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1499
timestamp 1624857261
transform 1 0 111112 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1498
timestamp 1624857261
transform 1 0 111112 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1497
timestamp 1624857261
transform 1 0 112880 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1496
timestamp 1624857261
transform 1 0 112880 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1495
timestamp 1624857261
transform 1 0 112880 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1494
timestamp 1624857261
transform 1 0 112880 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1493
timestamp 1624857261
transform 1 0 114648 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1492
timestamp 1624857261
transform 1 0 114648 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1491
timestamp 1624857261
transform 1 0 114648 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1490
timestamp 1624857261
transform 1 0 114648 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1489
timestamp 1624857261
transform 1 0 114648 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1488
timestamp 1624857261
transform 1 0 114648 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1487
timestamp 1624857261
transform 1 0 114648 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1486
timestamp 1624857261
transform 1 0 114648 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1485
timestamp 1624857261
transform 1 0 114648 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1484
timestamp 1624857261
transform 1 0 114648 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1483
timestamp 1624857261
transform 1 0 114784 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1482
timestamp 1624857261
transform 1 0 114648 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1481
timestamp 1624857261
transform 1 0 114920 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1480
timestamp 1624857261
transform 1 0 114920 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1479
timestamp 1624857261
transform 1 0 114784 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1478
timestamp 1624857261
transform 1 0 114784 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1477
timestamp 1624857261
transform 1 0 116144 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1476
timestamp 1624857261
transform 1 0 116144 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1475
timestamp 1624857261
transform 1 0 116144 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1474
timestamp 1624857261
transform 1 0 116144 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1473
timestamp 1624857261
transform 1 0 117912 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1472
timestamp 1624857261
transform 1 0 117912 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1471
timestamp 1624857261
transform 1 0 117912 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1470
timestamp 1624857261
transform 1 0 117912 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1469
timestamp 1624857261
transform 1 0 119544 0 1 16053
box 0 0 1 1
use contact_32  contact_32_1468
timestamp 1624857261
transform 1 0 119544 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1467
timestamp 1624857261
transform 1 0 119816 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1466
timestamp 1624857261
transform 1 0 119816 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1465
timestamp 1624857261
transform 1 0 119816 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1464
timestamp 1624857261
transform 1 0 119816 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1463
timestamp 1624857261
transform 1 0 119680 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1462
timestamp 1624857261
transform 1 0 119680 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1461
timestamp 1624857261
transform 1 0 119680 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1460
timestamp 1624857261
transform 1 0 119680 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1459
timestamp 1624857261
transform 1 0 119680 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1458
timestamp 1624857261
transform 1 0 119680 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1457
timestamp 1624857261
transform 1 0 119816 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1456
timestamp 1624857261
transform 1 0 119816 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1455
timestamp 1624857261
transform 1 0 119816 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1454
timestamp 1624857261
transform 1 0 119816 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1453
timestamp 1624857261
transform 1 0 119952 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1452
timestamp 1624857261
transform 1 0 119952 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1451
timestamp 1624857261
transform 1 0 121448 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1450
timestamp 1624857261
transform 1 0 121448 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1449
timestamp 1624857261
transform 1 0 121312 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1448
timestamp 1624857261
transform 1 0 121312 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1447
timestamp 1624857261
transform 1 0 122944 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1446
timestamp 1624857261
transform 1 0 122944 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1445
timestamp 1624857261
transform 1 0 122944 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1444
timestamp 1624857261
transform 1 0 122944 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1443
timestamp 1624857261
transform 1 0 124848 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1442
timestamp 1624857261
transform 1 0 124848 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1441
timestamp 1624857261
transform 1 0 124576 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1440
timestamp 1624857261
transform 1 0 124576 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1439
timestamp 1624857261
transform 1 0 124848 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1438
timestamp 1624857261
transform 1 0 124848 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1437
timestamp 1624857261
transform 1 0 124712 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1436
timestamp 1624857261
transform 1 0 124712 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1435
timestamp 1624857261
transform 1 0 124712 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1434
timestamp 1624857261
transform 1 0 124712 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1433
timestamp 1624857261
transform 1 0 124712 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1432
timestamp 1624857261
transform 1 0 124712 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1431
timestamp 1624857261
transform 1 0 124984 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1430
timestamp 1624857261
transform 1 0 124984 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1429
timestamp 1624857261
transform 1 0 124848 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1428
timestamp 1624857261
transform 1 0 124848 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1427
timestamp 1624857261
transform 1 0 126208 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1426
timestamp 1624857261
transform 1 0 126208 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1425
timestamp 1624857261
transform 1 0 126208 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1424
timestamp 1624857261
transform 1 0 126208 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1423
timestamp 1624857261
transform 1 0 127976 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1422
timestamp 1624857261
transform 1 0 127976 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1421
timestamp 1624857261
transform 1 0 127976 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1420
timestamp 1624857261
transform 1 0 127976 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1419
timestamp 1624857261
transform 1 0 129880 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1418
timestamp 1624857261
transform 1 0 129880 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1417
timestamp 1624857261
transform 1 0 129608 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1416
timestamp 1624857261
transform 1 0 129608 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1415
timestamp 1624857261
transform 1 0 129744 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1414
timestamp 1624857261
transform 1 0 129744 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1413
timestamp 1624857261
transform 1 0 129880 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1412
timestamp 1624857261
transform 1 0 129880 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1411
timestamp 1624857261
transform 1 0 129608 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1410
timestamp 1624857261
transform 1 0 129608 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1409
timestamp 1624857261
transform 1 0 129608 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1408
timestamp 1624857261
transform 1 0 129608 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1407
timestamp 1624857261
transform 1 0 129744 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1406
timestamp 1624857261
transform 1 0 129744 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1405
timestamp 1624857261
transform 1 0 129744 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1404
timestamp 1624857261
transform 1 0 129744 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1403
timestamp 1624857261
transform 1 0 131376 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1402
timestamp 1624857261
transform 1 0 131376 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1401
timestamp 1624857261
transform 1 0 131376 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1400
timestamp 1624857261
transform 1 0 131376 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1399
timestamp 1624857261
transform 1 0 133144 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1398
timestamp 1624857261
transform 1 0 133144 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1397
timestamp 1624857261
transform 1 0 133144 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1396
timestamp 1624857261
transform 1 0 133144 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1395
timestamp 1624857261
transform 1 0 134776 0 1 15917
box 0 0 1 1
use contact_32  contact_32_1394
timestamp 1624857261
transform 1 0 134776 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1393
timestamp 1624857261
transform 1 0 134912 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1392
timestamp 1624857261
transform 1 0 134912 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1391
timestamp 1624857261
transform 1 0 134776 0 1 17141
box 0 0 1 1
use contact_32  contact_32_1390
timestamp 1624857261
transform 1 0 134776 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1389
timestamp 1624857261
transform 1 0 134776 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1388
timestamp 1624857261
transform 1 0 134776 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1387
timestamp 1624857261
transform 1 0 134776 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1386
timestamp 1624857261
transform 1 0 134776 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1385
timestamp 1624857261
transform 1 0 134912 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1384
timestamp 1624857261
transform 1 0 134912 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1383
timestamp 1624857261
transform 1 0 134776 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1382
timestamp 1624857261
transform 1 0 134776 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1381
timestamp 1624857261
transform 1 0 134640 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1380
timestamp 1624857261
transform 1 0 134640 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1379
timestamp 1624857261
transform 1 0 134640 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1378
timestamp 1624857261
transform 1 0 134640 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1377
timestamp 1624857261
transform 1 0 136408 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1376
timestamp 1624857261
transform 1 0 136408 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1375
timestamp 1624857261
transform 1 0 136408 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1374
timestamp 1624857261
transform 1 0 136408 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1373
timestamp 1624857261
transform 1 0 138176 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1372
timestamp 1624857261
transform 1 0 138176 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1371
timestamp 1624857261
transform 1 0 138176 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1370
timestamp 1624857261
transform 1 0 138176 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1369
timestamp 1624857261
transform 1 0 139808 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1368
timestamp 1624857261
transform 1 0 139808 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1367
timestamp 1624857261
transform 1 0 139536 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1366
timestamp 1624857261
transform 1 0 139536 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1365
timestamp 1624857261
transform 1 0 139808 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1364
timestamp 1624857261
transform 1 0 139808 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1363
timestamp 1624857261
transform 1 0 139672 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1362
timestamp 1624857261
transform 1 0 139672 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1361
timestamp 1624857261
transform 1 0 139944 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1360
timestamp 1624857261
transform 1 0 139944 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1359
timestamp 1624857261
transform 1 0 139808 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1358
timestamp 1624857261
transform 1 0 139808 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1357
timestamp 1624857261
transform 1 0 139672 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1356
timestamp 1624857261
transform 1 0 139672 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1355
timestamp 1624857261
transform 1 0 139672 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1354
timestamp 1624857261
transform 1 0 139672 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1353
timestamp 1624857261
transform 1 0 141440 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1352
timestamp 1624857261
transform 1 0 141440 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1351
timestamp 1624857261
transform 1 0 141440 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1350
timestamp 1624857261
transform 1 0 141440 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1349
timestamp 1624857261
transform 1 0 143208 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1348
timestamp 1624857261
transform 1 0 143208 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1347
timestamp 1624857261
transform 1 0 143208 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1346
timestamp 1624857261
transform 1 0 143208 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1345
timestamp 1624857261
transform 1 0 144840 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1344
timestamp 1624857261
transform 1 0 144840 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1343
timestamp 1624857261
transform 1 0 144568 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1342
timestamp 1624857261
transform 1 0 144568 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1341
timestamp 1624857261
transform 1 0 144704 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1340
timestamp 1624857261
transform 1 0 144704 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1339
timestamp 1624857261
transform 1 0 144840 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1338
timestamp 1624857261
transform 1 0 144840 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1337
timestamp 1624857261
transform 1 0 144840 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1336
timestamp 1624857261
transform 1 0 144840 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1335
timestamp 1624857261
transform 1 0 144704 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1334
timestamp 1624857261
transform 1 0 144840 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1333
timestamp 1624857261
transform 1 0 144704 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1332
timestamp 1624857261
transform 1 0 144704 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1331
timestamp 1624857261
transform 1 0 144704 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1330
timestamp 1624857261
transform 1 0 144704 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1329
timestamp 1624857261
transform 1 0 146472 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1328
timestamp 1624857261
transform 1 0 146472 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1327
timestamp 1624857261
transform 1 0 146472 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1326
timestamp 1624857261
transform 1 0 146472 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1325
timestamp 1624857261
transform 1 0 148104 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1324
timestamp 1624857261
transform 1 0 148104 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1323
timestamp 1624857261
transform 1 0 148104 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1322
timestamp 1624857261
transform 1 0 148104 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1321
timestamp 1624857261
transform 1 0 149600 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1320
timestamp 1624857261
transform 1 0 149600 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1319
timestamp 1624857261
transform 1 0 149464 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1318
timestamp 1624857261
transform 1 0 149464 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1317
timestamp 1624857261
transform 1 0 149600 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1316
timestamp 1624857261
transform 1 0 149600 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1315
timestamp 1624857261
transform 1 0 149736 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1314
timestamp 1624857261
transform 1 0 149736 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1313
timestamp 1624857261
transform 1 0 149872 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1312
timestamp 1624857261
transform 1 0 149872 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1311
timestamp 1624857261
transform 1 0 149736 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1310
timestamp 1624857261
transform 1 0 149736 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1309
timestamp 1624857261
transform 1 0 150008 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1308
timestamp 1624857261
transform 1 0 150008 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1307
timestamp 1624857261
transform 1 0 149736 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1306
timestamp 1624857261
transform 1 0 149736 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1305
timestamp 1624857261
transform 1 0 151640 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1304
timestamp 1624857261
transform 1 0 151640 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1303
timestamp 1624857261
transform 1 0 151640 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1302
timestamp 1624857261
transform 1 0 151640 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1301
timestamp 1624857261
transform 1 0 153136 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1300
timestamp 1624857261
transform 1 0 153136 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1299
timestamp 1624857261
transform 1 0 153136 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1298
timestamp 1624857261
transform 1 0 153136 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1297
timestamp 1624857261
transform 1 0 154768 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1296
timestamp 1624857261
transform 1 0 154768 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1295
timestamp 1624857261
transform 1 0 154768 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1294
timestamp 1624857261
transform 1 0 154768 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1293
timestamp 1624857261
transform 1 0 154768 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1292
timestamp 1624857261
transform 1 0 154768 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1291
timestamp 1624857261
transform 1 0 154768 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1290
timestamp 1624857261
transform 1 0 154768 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1289
timestamp 1624857261
transform 1 0 154768 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1288
timestamp 1624857261
transform 1 0 154768 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1287
timestamp 1624857261
transform 1 0 154904 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1286
timestamp 1624857261
transform 1 0 154904 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1285
timestamp 1624857261
transform 1 0 154904 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1284
timestamp 1624857261
transform 1 0 154904 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1283
timestamp 1624857261
transform 1 0 154768 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1282
timestamp 1624857261
transform 1 0 154768 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1281
timestamp 1624857261
transform 1 0 156672 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1280
timestamp 1624857261
transform 1 0 156672 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1279
timestamp 1624857261
transform 1 0 156672 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1278
timestamp 1624857261
transform 1 0 156672 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1277
timestamp 1624857261
transform 1 0 158168 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1276
timestamp 1624857261
transform 1 0 158168 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1275
timestamp 1624857261
transform 1 0 158168 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1274
timestamp 1624857261
transform 1 0 158168 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1273
timestamp 1624857261
transform 1 0 159528 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1272
timestamp 1624857261
transform 1 0 159528 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1271
timestamp 1624857261
transform 1 0 159528 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1270
timestamp 1624857261
transform 1 0 159528 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1269
timestamp 1624857261
transform 1 0 159800 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1268
timestamp 1624857261
transform 1 0 159800 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1267
timestamp 1624857261
transform 1 0 159800 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1266
timestamp 1624857261
transform 1 0 159800 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1265
timestamp 1624857261
transform 1 0 159936 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1264
timestamp 1624857261
transform 1 0 159936 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1263
timestamp 1624857261
transform 1 0 159800 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1262
timestamp 1624857261
transform 1 0 159800 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1261
timestamp 1624857261
transform 1 0 159936 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1260
timestamp 1624857261
transform 1 0 159936 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1259
timestamp 1624857261
transform 1 0 159936 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1258
timestamp 1624857261
transform 1 0 159936 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1257
timestamp 1624857261
transform 1 0 161704 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1256
timestamp 1624857261
transform 1 0 161704 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1255
timestamp 1624857261
transform 1 0 161704 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1254
timestamp 1624857261
transform 1 0 161704 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1253
timestamp 1624857261
transform 1 0 163200 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1252
timestamp 1624857261
transform 1 0 163200 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1251
timestamp 1624857261
transform 1 0 163200 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1250
timestamp 1624857261
transform 1 0 163200 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1249
timestamp 1624857261
transform 1 0 164696 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1248
timestamp 1624857261
transform 1 0 164696 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1247
timestamp 1624857261
transform 1 0 164696 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1246
timestamp 1624857261
transform 1 0 164696 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1245
timestamp 1624857261
transform 1 0 164696 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1244
timestamp 1624857261
transform 1 0 164696 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1243
timestamp 1624857261
transform 1 0 164696 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1242
timestamp 1624857261
transform 1 0 164696 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1241
timestamp 1624857261
transform 1 0 164832 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1240
timestamp 1624857261
transform 1 0 164832 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1239
timestamp 1624857261
transform 1 0 164696 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1238
timestamp 1624857261
transform 1 0 164696 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1237
timestamp 1624857261
transform 1 0 164968 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1236
timestamp 1624857261
transform 1 0 164968 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1235
timestamp 1624857261
transform 1 0 164968 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1234
timestamp 1624857261
transform 1 0 164968 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1233
timestamp 1624857261
transform 1 0 166600 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1232
timestamp 1624857261
transform 1 0 166600 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1231
timestamp 1624857261
transform 1 0 166600 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1230
timestamp 1624857261
transform 1 0 166600 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1229
timestamp 1624857261
transform 1 0 168232 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1228
timestamp 1624857261
transform 1 0 168232 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1227
timestamp 1624857261
transform 1 0 168368 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1226
timestamp 1624857261
transform 1 0 168368 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1225
timestamp 1624857261
transform 1 0 169456 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1224
timestamp 1624857261
transform 1 0 169456 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1223
timestamp 1624857261
transform 1 0 169728 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1222
timestamp 1624857261
transform 1 0 169728 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1221
timestamp 1624857261
transform 1 0 169728 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1220
timestamp 1624857261
transform 1 0 169728 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1219
timestamp 1624857261
transform 1 0 169728 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1218
timestamp 1624857261
transform 1 0 169728 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1217
timestamp 1624857261
transform 1 0 169728 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1216
timestamp 1624857261
transform 1 0 169728 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1215
timestamp 1624857261
transform 1 0 169864 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1214
timestamp 1624857261
transform 1 0 169864 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1213
timestamp 1624857261
transform 1 0 170136 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1212
timestamp 1624857261
transform 1 0 170136 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1211
timestamp 1624857261
transform 1 0 170136 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1210
timestamp 1624857261
transform 1 0 170136 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1209
timestamp 1624857261
transform 1 0 171632 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1208
timestamp 1624857261
transform 1 0 171632 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1207
timestamp 1624857261
transform 1 0 171632 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1206
timestamp 1624857261
transform 1 0 171632 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1205
timestamp 1624857261
transform 1 0 173400 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1204
timestamp 1624857261
transform 1 0 173400 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1203
timestamp 1624857261
transform 1 0 173400 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1202
timestamp 1624857261
transform 1 0 173400 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1201
timestamp 1624857261
transform 1 0 174624 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1200
timestamp 1624857261
transform 1 0 174624 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1199
timestamp 1624857261
transform 1 0 174760 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1198
timestamp 1624857261
transform 1 0 174760 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1197
timestamp 1624857261
transform 1 0 174488 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1196
timestamp 1624857261
transform 1 0 174488 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1195
timestamp 1624857261
transform 1 0 174760 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1194
timestamp 1624857261
transform 1 0 174760 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1193
timestamp 1624857261
transform 1 0 174760 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1192
timestamp 1624857261
transform 1 0 174760 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1191
timestamp 1624857261
transform 1 0 174896 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1190
timestamp 1624857261
transform 1 0 174896 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1189
timestamp 1624857261
transform 1 0 175168 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1188
timestamp 1624857261
transform 1 0 175168 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1187
timestamp 1624857261
transform 1 0 175168 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1186
timestamp 1624857261
transform 1 0 175168 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1185
timestamp 1624857261
transform 1 0 176664 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1184
timestamp 1624857261
transform 1 0 176664 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1183
timestamp 1624857261
transform 1 0 176664 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1182
timestamp 1624857261
transform 1 0 176664 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1181
timestamp 1624857261
transform 1 0 178432 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1180
timestamp 1624857261
transform 1 0 178432 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1179
timestamp 1624857261
transform 1 0 178432 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1178
timestamp 1624857261
transform 1 0 178432 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1177
timestamp 1624857261
transform 1 0 179792 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1176
timestamp 1624857261
transform 1 0 179792 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1175
timestamp 1624857261
transform 1 0 179520 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1174
timestamp 1624857261
transform 1 0 179520 0 1 17413
box 0 0 1 1
use contact_32  contact_32_1173
timestamp 1624857261
transform 1 0 179792 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1172
timestamp 1624857261
transform 1 0 179792 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1171
timestamp 1624857261
transform 1 0 179792 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1170
timestamp 1624857261
transform 1 0 179792 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1169
timestamp 1624857261
transform 1 0 179792 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1168
timestamp 1624857261
transform 1 0 179792 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1167
timestamp 1624857261
transform 1 0 179656 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1166
timestamp 1624857261
transform 1 0 179656 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1165
timestamp 1624857261
transform 1 0 180200 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1164
timestamp 1624857261
transform 1 0 180200 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1163
timestamp 1624857261
transform 1 0 180200 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1162
timestamp 1624857261
transform 1 0 180200 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1161
timestamp 1624857261
transform 1 0 181696 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1160
timestamp 1624857261
transform 1 0 181696 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1159
timestamp 1624857261
transform 1 0 181696 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1158
timestamp 1624857261
transform 1 0 181696 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1157
timestamp 1624857261
transform 1 0 183464 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1156
timestamp 1624857261
transform 1 0 183464 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1155
timestamp 1624857261
transform 1 0 183328 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1154
timestamp 1624857261
transform 1 0 183328 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1153
timestamp 1624857261
transform 1 0 184552 0 1 16053
box 0 0 1 1
use contact_32  contact_32_1152
timestamp 1624857261
transform 1 0 184552 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1151
timestamp 1624857261
transform 1 0 189176 0 1 15781
box 0 0 1 1
use contact_32  contact_32_1150
timestamp 1624857261
transform 1 0 189176 0 1 14013
box 0 0 1 1
use contact_32  contact_32_1149
timestamp 1624857261
transform 1 0 184688 0 1 16869
box 0 0 1 1
use contact_32  contact_32_1148
timestamp 1624857261
transform 1 0 184688 0 1 16189
box 0 0 1 1
use contact_32  contact_32_1147
timestamp 1624857261
transform 1 0 184552 0 1 17005
box 0 0 1 1
use contact_32  contact_32_1146
timestamp 1624857261
transform 1 0 184552 0 1 17549
box 0 0 1 1
use contact_32  contact_32_1145
timestamp 1624857261
transform 1 0 184552 0 1 133013
box 0 0 1 1
use contact_32  contact_32_1144
timestamp 1624857261
transform 1 0 184552 0 1 131245
box 0 0 1 1
use contact_32  contact_32_1143
timestamp 1624857261
transform 1 0 184552 0 1 17821
box 0 0 1 1
use contact_32  contact_32_1142
timestamp 1624857261
transform 1 0 184552 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1141
timestamp 1624857261
transform 1 0 184688 0 1 131109
box 0 0 1 1
use contact_32  contact_32_1140
timestamp 1624857261
transform 1 0 184688 0 1 128661
box 0 0 1 1
use contact_32  contact_32_1139
timestamp 1624857261
transform 1 0 184688 0 1 19589
box 0 0 1 1
use contact_32  contact_32_1138
timestamp 1624857261
transform 1 0 184688 0 1 22037
box 0 0 1 1
use contact_32  contact_32_1137
timestamp 1624857261
transform 1 0 185096 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1136
timestamp 1624857261
transform 1 0 185096 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1135
timestamp 1624857261
transform 1 0 185096 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1134
timestamp 1624857261
transform 1 0 185096 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1133
timestamp 1624857261
transform 1 0 186728 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1132
timestamp 1624857261
transform 1 0 186728 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1131
timestamp 1624857261
transform 1 0 186864 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1130
timestamp 1624857261
transform 1 0 186864 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1129
timestamp 1624857261
transform 1 0 188632 0 1 142397
box 0 0 1 1
use contact_32  contact_32_1128
timestamp 1624857261
transform 1 0 188632 0 1 142805
box 0 0 1 1
use contact_32  contact_32_1127
timestamp 1624857261
transform 1 0 188632 0 1 1773
box 0 0 1 1
use contact_32  contact_32_1126
timestamp 1624857261
transform 1 0 188632 0 1 1229
box 0 0 1 1
use contact_32  contact_32_1125
timestamp 1624857261
transform 1 0 190400 0 1 128525
box 0 0 1 1
use contact_32  contact_32_1124
timestamp 1624857261
transform 1 0 190400 0 1 126349
box 0 0 1 1
use contact_32  contact_32_1123
timestamp 1624857261
transform 1 0 190264 0 1 66509
box 0 0 1 1
use contact_32  contact_32_1122
timestamp 1624857261
transform 1 0 190264 0 1 66781
box 0 0 1 1
use contact_32  contact_32_1121
timestamp 1624857261
transform 1 0 190128 0 1 39989
box 0 0 1 1
use contact_32  contact_32_1120
timestamp 1624857261
transform 1 0 190128 0 1 39717
box 0 0 1 1
use contact_32  contact_32_1119
timestamp 1624857261
transform 1 0 190264 0 1 79837
box 0 0 1 1
use contact_32  contact_32_1118
timestamp 1624857261
transform 1 0 190264 0 1 79565
box 0 0 1 1
use contact_32  contact_32_1117
timestamp 1624857261
transform 1 0 190128 0 1 79973
box 0 0 1 1
use contact_32  contact_32_1116
timestamp 1624857261
transform 1 0 190128 0 1 80245
box 0 0 1 1
use contact_32  contact_32_1115
timestamp 1624857261
transform 1 0 190264 0 1 87045
box 0 0 1 1
use contact_32  contact_32_1114
timestamp 1624857261
transform 1 0 190264 0 1 87317
box 0 0 1 1
use contact_32  contact_32_1113
timestamp 1624857261
transform 1 0 190128 0 1 41213
box 0 0 1 1
use contact_32  contact_32_1112
timestamp 1624857261
transform 1 0 190128 0 1 41485
box 0 0 1 1
use contact_32  contact_32_1111
timestamp 1624857261
transform 1 0 190128 0 1 68413
box 0 0 1 1
use contact_32  contact_32_1110
timestamp 1624857261
transform 1 0 190128 0 1 68141
box 0 0 1 1
use contact_32  contact_32_1109
timestamp 1624857261
transform 1 0 190128 0 1 38901
box 0 0 1 1
use contact_32  contact_32_1108
timestamp 1624857261
transform 1 0 190128 0 1 38493
box 0 0 1 1
use contact_32  contact_32_1107
timestamp 1624857261
transform 1 0 190264 0 1 101325
box 0 0 1 1
use contact_32  contact_32_1106
timestamp 1624857261
transform 1 0 190264 0 1 100917
box 0 0 1 1
use contact_32  contact_32_1105
timestamp 1624857261
transform 1 0 190264 0 1 26117
box 0 0 1 1
use contact_32  contact_32_1104
timestamp 1624857261
transform 1 0 190264 0 1 25845
box 0 0 1 1
use contact_32  contact_32_1103
timestamp 1624857261
transform 1 0 190264 0 1 26253
box 0 0 1 1
use contact_32  contact_32_1102
timestamp 1624857261
transform 1 0 190264 0 1 26525
box 0 0 1 1
use contact_32  contact_32_1101
timestamp 1624857261
transform 1 0 190264 0 1 42845
box 0 0 1 1
use contact_32  contact_32_1100
timestamp 1624857261
transform 1 0 190264 0 1 43117
box 0 0 1 1
use contact_32  contact_32_1099
timestamp 1624857261
transform 1 0 190264 0 1 42709
box 0 0 1 1
use contact_32  contact_32_1098
timestamp 1624857261
transform 1 0 190264 0 1 42437
box 0 0 1 1
use contact_32  contact_32_1097
timestamp 1624857261
transform 1 0 190128 0 1 34413
box 0 0 1 1
use contact_32  contact_32_1096
timestamp 1624857261
transform 1 0 190128 0 1 34141
box 0 0 1 1
use contact_32  contact_32_1095
timestamp 1624857261
transform 1 0 190128 0 1 34549
box 0 0 1 1
use contact_32  contact_32_1094
timestamp 1624857261
transform 1 0 190128 0 1 34821
box 0 0 1 1
use contact_32  contact_32_1093
timestamp 1624857261
transform 1 0 190128 0 1 58621
box 0 0 1 1
use contact_32  contact_32_1092
timestamp 1624857261
transform 1 0 190128 0 1 58893
box 0 0 1 1
use contact_32  contact_32_1091
timestamp 1624857261
transform 1 0 190128 0 1 63653
box 0 0 1 1
use contact_32  contact_32_1090
timestamp 1624857261
transform 1 0 190128 0 1 63381
box 0 0 1 1
use contact_32  contact_32_1089
timestamp 1624857261
transform 1 0 190128 0 1 88677
box 0 0 1 1
use contact_32  contact_32_1088
timestamp 1624857261
transform 1 0 190128 0 1 88949
box 0 0 1 1
use contact_32  contact_32_1087
timestamp 1624857261
transform 1 0 190264 0 1 104453
box 0 0 1 1
use contact_32  contact_32_1086
timestamp 1624857261
transform 1 0 190264 0 1 104181
box 0 0 1 1
use contact_32  contact_32_1085
timestamp 1624857261
transform 1 0 190264 0 1 125261
box 0 0 1 1
use contact_32  contact_32_1084
timestamp 1624857261
transform 1 0 190264 0 1 124989
box 0 0 1 1
use contact_32  contact_32_1083
timestamp 1624857261
transform 1 0 190128 0 1 112613
box 0 0 1 1
use contact_32  contact_32_1082
timestamp 1624857261
transform 1 0 190128 0 1 113021
box 0 0 1 1
use contact_32  contact_32_1081
timestamp 1624857261
transform 1 0 190264 0 1 113157
box 0 0 1 1
use contact_32  contact_32_1080
timestamp 1624857261
transform 1 0 190264 0 1 112749
box 0 0 1 1
use contact_32  contact_32_1079
timestamp 1624857261
transform 1 0 190128 0 1 30197
box 0 0 1 1
use contact_32  contact_32_1078
timestamp 1624857261
transform 1 0 190128 0 1 30469
box 0 0 1 1
use contact_32  contact_32_1077
timestamp 1624857261
transform 1 0 190128 0 1 125261
box 0 0 1 1
use contact_32  contact_32_1076
timestamp 1624857261
transform 1 0 190128 0 1 125669
box 0 0 1 1
use contact_32  contact_32_1075
timestamp 1624857261
transform 1 0 190128 0 1 113429
box 0 0 1 1
use contact_32  contact_32_1074
timestamp 1624857261
transform 1 0 190128 0 1 113157
box 0 0 1 1
use contact_32  contact_32_1073
timestamp 1624857261
transform 1 0 190264 0 1 116557
box 0 0 1 1
use contact_32  contact_32_1072
timestamp 1624857261
transform 1 0 190264 0 1 116285
box 0 0 1 1
use contact_32  contact_32_1071
timestamp 1624857261
transform 1 0 190264 0 1 116693
box 0 0 1 1
use contact_32  contact_32_1070
timestamp 1624857261
transform 1 0 190264 0 1 116965
box 0 0 1 1
use contact_32  contact_32_1069
timestamp 1624857261
transform 1 0 190128 0 1 31285
box 0 0 1 1
use contact_32  contact_32_1068
timestamp 1624857261
transform 1 0 190128 0 1 31013
box 0 0 1 1
use contact_32  contact_32_1067
timestamp 1624857261
transform 1 0 190128 0 1 87589
box 0 0 1 1
use contact_32  contact_32_1066
timestamp 1624857261
transform 1 0 190128 0 1 87861
box 0 0 1 1
use contact_32  contact_32_1065
timestamp 1624857261
transform 1 0 190128 0 1 62837
box 0 0 1 1
use contact_32  contact_32_1064
timestamp 1624857261
transform 1 0 190128 0 1 62565
box 0 0 1 1
use contact_32  contact_32_1063
timestamp 1624857261
transform 1 0 190128 0 1 62973
box 0 0 1 1
use contact_32  contact_32_1062
timestamp 1624857261
transform 1 0 190128 0 1 63245
box 0 0 1 1
use contact_32  contact_32_1061
timestamp 1624857261
transform 1 0 190264 0 1 76301
box 0 0 1 1
use contact_32  contact_32_1060
timestamp 1624857261
transform 1 0 190264 0 1 76029
box 0 0 1 1
use contact_32  contact_32_1059
timestamp 1624857261
transform 1 0 190128 0 1 71269
box 0 0 1 1
use contact_32  contact_32_1058
timestamp 1624857261
transform 1 0 190128 0 1 71541
box 0 0 1 1
use contact_32  contact_32_1057
timestamp 1624857261
transform 1 0 190264 0 1 104861
box 0 0 1 1
use contact_32  contact_32_1056
timestamp 1624857261
transform 1 0 190264 0 1 105133
box 0 0 1 1
use contact_32  contact_32_1055
timestamp 1624857261
transform 1 0 190128 0 1 70453
box 0 0 1 1
use contact_32  contact_32_1054
timestamp 1624857261
transform 1 0 190128 0 1 70725
box 0 0 1 1
use contact_32  contact_32_1053
timestamp 1624857261
transform 1 0 190264 0 1 110029
box 0 0 1 1
use contact_32  contact_32_1052
timestamp 1624857261
transform 1 0 190264 0 1 110301
box 0 0 1 1
use contact_32  contact_32_1051
timestamp 1624857261
transform 1 0 190128 0 1 96429
box 0 0 1 1
use contact_32  contact_32_1050
timestamp 1624857261
transform 1 0 190128 0 1 96157
box 0 0 1 1
use contact_32  contact_32_1049
timestamp 1624857261
transform 1 0 190264 0 1 114245
box 0 0 1 1
use contact_32  contact_32_1048
timestamp 1624857261
transform 1 0 190264 0 1 113973
box 0 0 1 1
use contact_32  contact_32_1047
timestamp 1624857261
transform 1 0 190264 0 1 35229
box 0 0 1 1
use contact_32  contact_32_1046
timestamp 1624857261
transform 1 0 190264 0 1 34957
box 0 0 1 1
use contact_32  contact_32_1045
timestamp 1624857261
transform 1 0 190128 0 1 55357
box 0 0 1 1
use contact_32  contact_32_1044
timestamp 1624857261
transform 1 0 190128 0 1 55085
box 0 0 1 1
use contact_32  contact_32_1043
timestamp 1624857261
transform 1 0 190264 0 1 83917
box 0 0 1 1
use contact_32  contact_32_1042
timestamp 1624857261
transform 1 0 190264 0 1 84189
box 0 0 1 1
use contact_32  contact_32_1041
timestamp 1624857261
transform 1 0 190128 0 1 92213
box 0 0 1 1
use contact_32  contact_32_1040
timestamp 1624857261
transform 1 0 190128 0 1 92485
box 0 0 1 1
use contact_32  contact_32_1039
timestamp 1624857261
transform 1 0 190264 0 1 54677
box 0 0 1 1
use contact_32  contact_32_1038
timestamp 1624857261
transform 1 0 190264 0 1 54949
box 0 0 1 1
use contact_32  contact_32_1037
timestamp 1624857261
transform 1 0 190128 0 1 121725
box 0 0 1 1
use contact_32  contact_32_1036
timestamp 1624857261
transform 1 0 190128 0 1 121453
box 0 0 1 1
use contact_32  contact_32_1035
timestamp 1624857261
transform 1 0 190264 0 1 70997
box 0 0 1 1
use contact_32  contact_32_1034
timestamp 1624857261
transform 1 0 190264 0 1 71269
box 0 0 1 1
use contact_32  contact_32_1033
timestamp 1624857261
transform 1 0 190264 0 1 107853
box 0 0 1 1
use contact_32  contact_32_1032
timestamp 1624857261
transform 1 0 190264 0 1 107581
box 0 0 1 1
use contact_32  contact_32_1031
timestamp 1624857261
transform 1 0 190264 0 1 109213
box 0 0 1 1
use contact_32  contact_32_1030
timestamp 1624857261
transform 1 0 190264 0 1 109485
box 0 0 1 1
use contact_32  contact_32_1029
timestamp 1624857261
transform 1 0 190264 0 1 109077
box 0 0 1 1
use contact_32  contact_32_1028
timestamp 1624857261
transform 1 0 190264 0 1 108805
box 0 0 1 1
use contact_32  contact_32_1027
timestamp 1624857261
transform 1 0 190128 0 1 43389
box 0 0 1 1
use contact_32  contact_32_1026
timestamp 1624857261
transform 1 0 190128 0 1 43117
box 0 0 1 1
use contact_32  contact_32_1025
timestamp 1624857261
transform 1 0 190264 0 1 88677
box 0 0 1 1
use contact_32  contact_32_1024
timestamp 1624857261
transform 1 0 190264 0 1 88269
box 0 0 1 1
use contact_32  contact_32_1023
timestamp 1624857261
transform 1 0 190128 0 1 46245
box 0 0 1 1
use contact_32  contact_32_1022
timestamp 1624857261
transform 1 0 190128 0 1 45973
box 0 0 1 1
use contact_32  contact_32_1021
timestamp 1624857261
transform 1 0 190128 0 1 37541
box 0 0 1 1
use contact_32  contact_32_1020
timestamp 1624857261
transform 1 0 190128 0 1 37269
box 0 0 1 1
use contact_32  contact_32_1019
timestamp 1624857261
transform 1 0 190128 0 1 120501
box 0 0 1 1
use contact_32  contact_32_1018
timestamp 1624857261
transform 1 0 190128 0 1 120229
box 0 0 1 1
use contact_32  contact_32_1017
timestamp 1624857261
transform 1 0 190400 0 1 125941
box 0 0 1 1
use contact_32  contact_32_1016
timestamp 1624857261
transform 1 0 190400 0 1 126213
box 0 0 1 1
use contact_32  contact_32_1015
timestamp 1624857261
transform 1 0 190264 0 1 38765
box 0 0 1 1
use contact_32  contact_32_1014
timestamp 1624857261
transform 1 0 190264 0 1 38493
box 0 0 1 1
use contact_32  contact_32_1013
timestamp 1624857261
transform 1 0 190264 0 1 79429
box 0 0 1 1
use contact_32  contact_32_1012
timestamp 1624857261
transform 1 0 190264 0 1 79157
box 0 0 1 1
use contact_32  contact_32_1011
timestamp 1624857261
transform 1 0 190264 0 1 120909
box 0 0 1 1
use contact_32  contact_32_1010
timestamp 1624857261
transform 1 0 190264 0 1 120501
box 0 0 1 1
use contact_32  contact_32_1009
timestamp 1624857261
transform 1 0 190264 0 1 121045
box 0 0 1 1
use contact_32  contact_32_1008
timestamp 1624857261
transform 1 0 190264 0 1 121317
box 0 0 1 1
use contact_32  contact_32_1007
timestamp 1624857261
transform 1 0 190264 0 1 95205
box 0 0 1 1
use contact_32  contact_32_1006
timestamp 1624857261
transform 1 0 190264 0 1 94933
box 0 0 1 1
use contact_32  contact_32_1005
timestamp 1624857261
transform 1 0 190264 0 1 56581
box 0 0 1 1
use contact_32  contact_32_1004
timestamp 1624857261
transform 1 0 190264 0 1 56309
box 0 0 1 1
use contact_32  contact_32_1003
timestamp 1624857261
transform 1 0 190264 0 1 51141
box 0 0 1 1
use contact_32  contact_32_1002
timestamp 1624857261
transform 1 0 190264 0 1 51413
box 0 0 1 1
use contact_32  contact_32_1001
timestamp 1624857261
transform 1 0 190264 0 1 75213
box 0 0 1 1
use contact_32  contact_32_1000
timestamp 1624857261
transform 1 0 190264 0 1 75485
box 0 0 1 1
use contact_32  contact_32_999
timestamp 1624857261
transform 1 0 193120 0 1 75077
box 0 0 1 1
use contact_32  contact_32_998
timestamp 1624857261
transform 1 0 193120 0 1 75349
box 0 0 1 1
use contact_32  contact_32_997
timestamp 1624857261
transform 1 0 190128 0 1 71677
box 0 0 1 1
use contact_32  contact_32_996
timestamp 1624857261
transform 1 0 190128 0 1 71949
box 0 0 1 1
use contact_32  contact_32_995
timestamp 1624857261
transform 1 0 190264 0 1 92893
box 0 0 1 1
use contact_32  contact_32_994
timestamp 1624857261
transform 1 0 190264 0 1 92621
box 0 0 1 1
use contact_32  contact_32_993
timestamp 1624857261
transform 1 0 190128 0 1 110029
box 0 0 1 1
use contact_32  contact_32_992
timestamp 1624857261
transform 1 0 190128 0 1 109621
box 0 0 1 1
use contact_32  contact_32_991
timestamp 1624857261
transform 1 0 190264 0 1 59029
box 0 0 1 1
use contact_32  contact_32_990
timestamp 1624857261
transform 1 0 190264 0 1 59301
box 0 0 1 1
use contact_32  contact_32_989
timestamp 1624857261
transform 1 0 190128 0 1 117101
box 0 0 1 1
use contact_32  contact_32_988
timestamp 1624857261
transform 1 0 190128 0 1 117373
box 0 0 1 1
use contact_32  contact_32_987
timestamp 1624857261
transform 1 0 190264 0 1 105541
box 0 0 1 1
use contact_32  contact_32_986
timestamp 1624857261
transform 1 0 190264 0 1 105269
box 0 0 1 1
use contact_32  contact_32_985
timestamp 1624857261
transform 1 0 190128 0 1 68005
box 0 0 1 1
use contact_32  contact_32_984
timestamp 1624857261
transform 1 0 190128 0 1 67733
box 0 0 1 1
use contact_32  contact_32_983
timestamp 1624857261
transform 1 0 190128 0 1 107853
box 0 0 1 1
use contact_32  contact_32_982
timestamp 1624857261
transform 1 0 190128 0 1 108261
box 0 0 1 1
use contact_32  contact_32_981
timestamp 1624857261
transform 1 0 190128 0 1 75893
box 0 0 1 1
use contact_32  contact_32_980
timestamp 1624857261
transform 1 0 190128 0 1 75621
box 0 0 1 1
use contact_32  contact_32_979
timestamp 1624857261
transform 1 0 190128 0 1 108397
box 0 0 1 1
use contact_32  contact_32_978
timestamp 1624857261
transform 1 0 190128 0 1 108669
box 0 0 1 1
use contact_32  contact_32_977
timestamp 1624857261
transform 1 0 190128 0 1 77117
box 0 0 1 1
use contact_32  contact_32_976
timestamp 1624857261
transform 1 0 190128 0 1 76845
box 0 0 1 1
use contact_32  contact_32_975
timestamp 1624857261
transform 1 0 190128 0 1 1773
box 0 0 1 1
use contact_32  contact_32_974
timestamp 1624857261
transform 1 0 190128 0 1 1229
box 0 0 1 1
use contact_32  contact_32_973
timestamp 1624857261
transform 1 0 190128 0 1 142397
box 0 0 1 1
use contact_32  contact_32_972
timestamp 1624857261
transform 1 0 190128 0 1 142805
box 0 0 1 1
use contact_32  contact_32_971
timestamp 1624857261
transform 1 0 191896 0 1 142397
box 0 0 1 1
use contact_32  contact_32_970
timestamp 1624857261
transform 1 0 191896 0 1 142805
box 0 0 1 1
use contact_32  contact_32_969
timestamp 1624857261
transform 1 0 191896 0 1 1773
box 0 0 1 1
use contact_32  contact_32_968
timestamp 1624857261
transform 1 0 191896 0 1 1229
box 0 0 1 1
use contact_32  contact_32_967
timestamp 1624857261
transform 1 0 193664 0 1 1773
box 0 0 1 1
use contact_32  contact_32_966
timestamp 1624857261
transform 1 0 193664 0 1 1229
box 0 0 1 1
use contact_32  contact_32_965
timestamp 1624857261
transform 1 0 193664 0 1 142397
box 0 0 1 1
use contact_32  contact_32_964
timestamp 1624857261
transform 1 0 193664 0 1 142805
box 0 0 1 1
use contact_32  contact_32_963
timestamp 1624857261
transform 1 0 195160 0 1 1773
box 0 0 1 1
use contact_32  contact_32_962
timestamp 1624857261
transform 1 0 195160 0 1 1229
box 0 0 1 1
use contact_32  contact_32_961
timestamp 1624857261
transform 1 0 195160 0 1 142397
box 0 0 1 1
use contact_32  contact_32_960
timestamp 1624857261
transform 1 0 195160 0 1 142805
box 0 0 1 1
use contact_32  contact_32_959
timestamp 1624857261
transform 1 0 195568 0 1 124037
box 0 0 1 1
use contact_32  contact_32_958
timestamp 1624857261
transform 1 0 195568 0 1 124309
box 0 0 1 1
use contact_32  contact_32_957
timestamp 1624857261
transform 1 0 195432 0 1 123901
box 0 0 1 1
use contact_32  contact_32_956
timestamp 1624857261
transform 1 0 195432 0 1 123629
box 0 0 1 1
use contact_32  contact_32_955
timestamp 1624857261
transform 1 0 195568 0 1 99149
box 0 0 1 1
use contact_32  contact_32_954
timestamp 1624857261
transform 1 0 195568 0 1 99421
box 0 0 1 1
use contact_32  contact_32_953
timestamp 1624857261
transform 1 0 195568 0 1 99013
box 0 0 1 1
use contact_32  contact_32_952
timestamp 1624857261
transform 1 0 195568 0 1 98741
box 0 0 1 1
use contact_32  contact_32_951
timestamp 1624857261
transform 1 0 195432 0 1 45021
box 0 0 1 1
use contact_32  contact_32_950
timestamp 1624857261
transform 1 0 195432 0 1 45293
box 0 0 1 1
use contact_32  contact_32_949
timestamp 1624857261
transform 1 0 195432 0 1 44885
box 0 0 1 1
use contact_32  contact_32_948
timestamp 1624857261
transform 1 0 195432 0 1 44613
box 0 0 1 1
use contact_32  contact_32_947
timestamp 1624857261
transform 1 0 195568 0 1 100237
box 0 0 1 1
use contact_32  contact_32_946
timestamp 1624857261
transform 1 0 195568 0 1 99965
box 0 0 1 1
use contact_32  contact_32_945
timestamp 1624857261
transform 1 0 195568 0 1 45701
box 0 0 1 1
use contact_32  contact_32_944
timestamp 1624857261
transform 1 0 195568 0 1 45429
box 0 0 1 1
use contact_32  contact_32_943
timestamp 1624857261
transform 1 0 195568 0 1 45837
box 0 0 1 1
use contact_32  contact_32_942
timestamp 1624857261
transform 1 0 195568 0 1 46109
box 0 0 1 1
use contact_32  contact_32_941
timestamp 1624857261
transform 1 0 195568 0 1 122405
box 0 0 1 1
use contact_32  contact_32_940
timestamp 1624857261
transform 1 0 195568 0 1 122677
box 0 0 1 1
use contact_32  contact_32_939
timestamp 1624857261
transform 1 0 195432 0 1 122269
box 0 0 1 1
use contact_32  contact_32_938
timestamp 1624857261
transform 1 0 195432 0 1 121997
box 0 0 1 1
use contact_32  contact_32_937
timestamp 1624857261
transform 1 0 195432 0 1 108125
box 0 0 1 1
use contact_32  contact_32_936
timestamp 1624857261
transform 1 0 195432 0 1 107853
box 0 0 1 1
use contact_32  contact_32_935
timestamp 1624857261
transform 1 0 195568 0 1 111661
box 0 0 1 1
use contact_32  contact_32_934
timestamp 1624857261
transform 1 0 195568 0 1 111389
box 0 0 1 1
use contact_32  contact_32_933
timestamp 1624857261
transform 1 0 195432 0 1 111797
box 0 0 1 1
use contact_32  contact_32_932
timestamp 1624857261
transform 1 0 195432 0 1 112069
box 0 0 1 1
use contact_32  contact_32_931
timestamp 1624857261
transform 1 0 195432 0 1 35093
box 0 0 1 1
use contact_32  contact_32_930
timestamp 1624857261
transform 1 0 195432 0 1 35365
box 0 0 1 1
use contact_32  contact_32_929
timestamp 1624857261
transform 1 0 195432 0 1 29245
box 0 0 1 1
use contact_32  contact_32_928
timestamp 1624857261
transform 1 0 195432 0 1 29517
box 0 0 1 1
use contact_32  contact_32_927
timestamp 1624857261
transform 1 0 195432 0 1 29109
box 0 0 1 1
use contact_32  contact_32_926
timestamp 1624857261
transform 1 0 195432 0 1 28837
box 0 0 1 1
use contact_32  contact_32_925
timestamp 1624857261
transform 1 0 195432 0 1 107037
box 0 0 1 1
use contact_32  contact_32_924
timestamp 1624857261
transform 1 0 195432 0 1 107309
box 0 0 1 1
use contact_32  contact_32_923
timestamp 1624857261
transform 1 0 195432 0 1 106901
box 0 0 1 1
use contact_32  contact_32_922
timestamp 1624857261
transform 1 0 195432 0 1 106629
box 0 0 1 1
use contact_32  contact_32_921
timestamp 1624857261
transform 1 0 195568 0 1 54405
box 0 0 1 1
use contact_32  contact_32_920
timestamp 1624857261
transform 1 0 195568 0 1 54133
box 0 0 1 1
use contact_32  contact_32_919
timestamp 1624857261
transform 1 0 195432 0 1 116013
box 0 0 1 1
use contact_32  contact_32_918
timestamp 1624857261
transform 1 0 195432 0 1 115741
box 0 0 1 1
use contact_32  contact_32_917
timestamp 1624857261
transform 1 0 195432 0 1 116149
box 0 0 1 1
use contact_32  contact_32_916
timestamp 1624857261
transform 1 0 195432 0 1 116421
box 0 0 1 1
use contact_32  contact_32_915
timestamp 1624857261
transform 1 0 195432 0 1 32237
box 0 0 1 1
use contact_32  contact_32_914
timestamp 1624857261
transform 1 0 195432 0 1 31965
box 0 0 1 1
use contact_32  contact_32_913
timestamp 1624857261
transform 1 0 195432 0 1 32373
box 0 0 1 1
use contact_32  contact_32_912
timestamp 1624857261
transform 1 0 195432 0 1 32645
box 0 0 1 1
use contact_32  contact_32_911
timestamp 1624857261
transform 1 0 195568 0 1 61613
box 0 0 1 1
use contact_32  contact_32_910
timestamp 1624857261
transform 1 0 195568 0 1 61885
box 0 0 1 1
use contact_32  contact_32_909
timestamp 1624857261
transform 1 0 195568 0 1 61477
box 0 0 1 1
use contact_32  contact_32_908
timestamp 1624857261
transform 1 0 195568 0 1 61205
box 0 0 1 1
use contact_32  contact_32_907
timestamp 1624857261
transform 1 0 195432 0 1 56717
box 0 0 1 1
use contact_32  contact_32_906
timestamp 1624857261
transform 1 0 195432 0 1 56445
box 0 0 1 1
use contact_32  contact_32_905
timestamp 1624857261
transform 1 0 195432 0 1 56853
box 0 0 1 1
use contact_32  contact_32_904
timestamp 1624857261
transform 1 0 195432 0 1 57125
box 0 0 1 1
use contact_32  contact_32_903
timestamp 1624857261
transform 1 0 195568 0 1 57669
box 0 0 1 1
use contact_32  contact_32_902
timestamp 1624857261
transform 1 0 195568 0 1 57941
box 0 0 1 1
use contact_32  contact_32_901
timestamp 1624857261
transform 1 0 195432 0 1 57533
box 0 0 1 1
use contact_32  contact_32_900
timestamp 1624857261
transform 1 0 195432 0 1 57261
box 0 0 1 1
use contact_32  contact_32_899
timestamp 1624857261
transform 1 0 195432 0 1 33869
box 0 0 1 1
use contact_32  contact_32_898
timestamp 1624857261
transform 1 0 195432 0 1 33597
box 0 0 1 1
use contact_32  contact_32_897
timestamp 1624857261
transform 1 0 195432 0 1 36181
box 0 0 1 1
use contact_32  contact_32_896
timestamp 1624857261
transform 1 0 195432 0 1 35909
box 0 0 1 1
use contact_32  contact_32_895
timestamp 1624857261
transform 1 0 195432 0 1 36317
box 0 0 1 1
use contact_32  contact_32_894
timestamp 1624857261
transform 1 0 195432 0 1 36589
box 0 0 1 1
use contact_32  contact_32_893
timestamp 1624857261
transform 1 0 195432 0 1 31829
box 0 0 1 1
use contact_32  contact_32_892
timestamp 1624857261
transform 1 0 195432 0 1 31557
box 0 0 1 1
use contact_32  contact_32_891
timestamp 1624857261
transform 1 0 195432 0 1 91669
box 0 0 1 1
use contact_32  contact_32_890
timestamp 1624857261
transform 1 0 195432 0 1 91941
box 0 0 1 1
use contact_32  contact_32_889
timestamp 1624857261
transform 1 0 195432 0 1 91533
box 0 0 1 1
use contact_32  contact_32_888
timestamp 1624857261
transform 1 0 195432 0 1 91261
box 0 0 1 1
use contact_32  contact_32_887
timestamp 1624857261
transform 1 0 195432 0 1 97789
box 0 0 1 1
use contact_32  contact_32_886
timestamp 1624857261
transform 1 0 195432 0 1 97517
box 0 0 1 1
use contact_32  contact_32_885
timestamp 1624857261
transform 1 0 195568 0 1 97925
box 0 0 1 1
use contact_32  contact_32_884
timestamp 1624857261
transform 1 0 195568 0 1 98197
box 0 0 1 1
use contact_32  contact_32_883
timestamp 1624857261
transform 1 0 195432 0 1 86365
box 0 0 1 1
use contact_32  contact_32_882
timestamp 1624857261
transform 1 0 195432 0 1 86093
box 0 0 1 1
use contact_32  contact_32_881
timestamp 1624857261
transform 1 0 195568 0 1 86501
box 0 0 1 1
use contact_32  contact_32_880
timestamp 1624857261
transform 1 0 195568 0 1 86773
box 0 0 1 1
use contact_32  contact_32_879
timestamp 1624857261
transform 1 0 195432 0 1 58485
box 0 0 1 1
use contact_32  contact_32_878
timestamp 1624857261
transform 1 0 195432 0 1 58757
box 0 0 1 1
use contact_32  contact_32_877
timestamp 1624857261
transform 1 0 195432 0 1 58349
box 0 0 1 1
use contact_32  contact_32_876
timestamp 1624857261
transform 1 0 195432 0 1 58077
box 0 0 1 1
use contact_32  contact_32_875
timestamp 1624857261
transform 1 0 195568 0 1 99557
box 0 0 1 1
use contact_32  contact_32_874
timestamp 1624857261
transform 1 0 195568 0 1 99829
box 0 0 1 1
use contact_32  contact_32_873
timestamp 1624857261
transform 1 0 195568 0 1 73445
box 0 0 1 1
use contact_32  contact_32_872
timestamp 1624857261
transform 1 0 195568 0 1 73717
box 0 0 1 1
use contact_32  contact_32_871
timestamp 1624857261
transform 1 0 195432 0 1 73309
box 0 0 1 1
use contact_32  contact_32_870
timestamp 1624857261
transform 1 0 195432 0 1 73037
box 0 0 1 1
use contact_32  contact_32_869
timestamp 1624857261
transform 1 0 195568 0 1 93165
box 0 0 1 1
use contact_32  contact_32_868
timestamp 1624857261
transform 1 0 195568 0 1 93437
box 0 0 1 1
use contact_32  contact_32_867
timestamp 1624857261
transform 1 0 195568 0 1 93029
box 0 0 1 1
use contact_32  contact_32_866
timestamp 1624857261
transform 1 0 195568 0 1 92757
box 0 0 1 1
use contact_32  contact_32_865
timestamp 1624857261
transform 1 0 195568 0 1 120365
box 0 0 1 1
use contact_32  contact_32_864
timestamp 1624857261
transform 1 0 195568 0 1 120093
box 0 0 1 1
use contact_32  contact_32_863
timestamp 1624857261
transform 1 0 195432 0 1 120501
box 0 0 1 1
use contact_32  contact_32_862
timestamp 1624857261
transform 1 0 195432 0 1 120773
box 0 0 1 1
use contact_32  contact_32_861
timestamp 1624857261
transform 1 0 195568 0 1 30741
box 0 0 1 1
use contact_32  contact_32_860
timestamp 1624857261
transform 1 0 195568 0 1 31013
box 0 0 1 1
use contact_32  contact_32_859
timestamp 1624857261
transform 1 0 195432 0 1 40533
box 0 0 1 1
use contact_32  contact_32_858
timestamp 1624857261
transform 1 0 195432 0 1 40261
box 0 0 1 1
use contact_32  contact_32_857
timestamp 1624857261
transform 1 0 195432 0 1 40669
box 0 0 1 1
use contact_32  contact_32_856
timestamp 1624857261
transform 1 0 195432 0 1 40941
box 0 0 1 1
use contact_32  contact_32_855
timestamp 1624857261
transform 1 0 195432 0 1 89493
box 0 0 1 1
use contact_32  contact_32_854
timestamp 1624857261
transform 1 0 195432 0 1 89221
box 0 0 1 1
use contact_32  contact_32_853
timestamp 1624857261
transform 1 0 195432 0 1 89629
box 0 0 1 1
use contact_32  contact_32_852
timestamp 1624857261
transform 1 0 195432 0 1 89901
box 0 0 1 1
use contact_32  contact_32_851
timestamp 1624857261
transform 1 0 195568 0 1 94797
box 0 0 1 1
use contact_32  contact_32_850
timestamp 1624857261
transform 1 0 195568 0 1 95069
box 0 0 1 1
use contact_32  contact_32_849
timestamp 1624857261
transform 1 0 195568 0 1 94661
box 0 0 1 1
use contact_32  contact_32_848
timestamp 1624857261
transform 1 0 195568 0 1 94389
box 0 0 1 1
use contact_32  contact_32_847
timestamp 1624857261
transform 1 0 195432 0 1 46517
box 0 0 1 1
use contact_32  contact_32_846
timestamp 1624857261
transform 1 0 195432 0 1 46245
box 0 0 1 1
use contact_32  contact_32_845
timestamp 1624857261
transform 1 0 195568 0 1 84869
box 0 0 1 1
use contact_32  contact_32_844
timestamp 1624857261
transform 1 0 195568 0 1 85141
box 0 0 1 1
use contact_32  contact_32_843
timestamp 1624857261
transform 1 0 195432 0 1 84733
box 0 0 1 1
use contact_32  contact_32_842
timestamp 1624857261
transform 1 0 195432 0 1 84461
box 0 0 1 1
use contact_32  contact_32_841
timestamp 1624857261
transform 1 0 195568 0 1 53997
box 0 0 1 1
use contact_32  contact_32_840
timestamp 1624857261
transform 1 0 195568 0 1 53725
box 0 0 1 1
use contact_32  contact_32_839
timestamp 1624857261
transform 1 0 195432 0 1 55901
box 0 0 1 1
use contact_32  contact_32_838
timestamp 1624857261
transform 1 0 195432 0 1 55629
box 0 0 1 1
use contact_32  contact_32_837
timestamp 1624857261
transform 1 0 195568 0 1 56037
box 0 0 1 1
use contact_32  contact_32_836
timestamp 1624857261
transform 1 0 195568 0 1 56309
box 0 0 1 1
use contact_32  contact_32_835
timestamp 1624857261
transform 1 0 195568 0 1 44205
box 0 0 1 1
use contact_32  contact_32_834
timestamp 1624857261
transform 1 0 195568 0 1 44477
box 0 0 1 1
use contact_32  contact_32_833
timestamp 1624857261
transform 1 0 195568 0 1 44069
box 0 0 1 1
use contact_32  contact_32_832
timestamp 1624857261
transform 1 0 195568 0 1 43797
box 0 0 1 1
use contact_32  contact_32_831
timestamp 1624857261
transform 1 0 195568 0 1 87589
box 0 0 1 1
use contact_32  contact_32_830
timestamp 1624857261
transform 1 0 195568 0 1 87317
box 0 0 1 1
use contact_32  contact_32_829
timestamp 1624857261
transform 1 0 195568 0 1 41893
box 0 0 1 1
use contact_32  contact_32_828
timestamp 1624857261
transform 1 0 195568 0 1 42165
box 0 0 1 1
use contact_32  contact_32_827
timestamp 1624857261
transform 1 0 195432 0 1 41757
box 0 0 1 1
use contact_32  contact_32_826
timestamp 1624857261
transform 1 0 195432 0 1 41485
box 0 0 1 1
use contact_32  contact_32_825
timestamp 1624857261
transform 1 0 195432 0 1 73853
box 0 0 1 1
use contact_32  contact_32_824
timestamp 1624857261
transform 1 0 195432 0 1 74125
box 0 0 1 1
use contact_32  contact_32_823
timestamp 1624857261
transform 1 0 195568 0 1 70725
box 0 0 1 1
use contact_32  contact_32_822
timestamp 1624857261
transform 1 0 195568 0 1 70997
box 0 0 1 1
use contact_32  contact_32_821
timestamp 1624857261
transform 1 0 195432 0 1 70589
box 0 0 1 1
use contact_32  contact_32_820
timestamp 1624857261
transform 1 0 195432 0 1 70317
box 0 0 1 1
use contact_32  contact_32_819
timestamp 1624857261
transform 1 0 195432 0 1 47605
box 0 0 1 1
use contact_32  contact_32_818
timestamp 1624857261
transform 1 0 195432 0 1 47333
box 0 0 1 1
use contact_32  contact_32_817
timestamp 1624857261
transform 1 0 195432 0 1 47741
box 0 0 1 1
use contact_32  contact_32_816
timestamp 1624857261
transform 1 0 195432 0 1 48013
box 0 0 1 1
use contact_32  contact_32_815
timestamp 1624857261
transform 1 0 195432 0 1 78613
box 0 0 1 1
use contact_32  contact_32_814
timestamp 1624857261
transform 1 0 195432 0 1 78885
box 0 0 1 1
use contact_32  contact_32_813
timestamp 1624857261
transform 1 0 195568 0 1 78477
box 0 0 1 1
use contact_32  contact_32_812
timestamp 1624857261
transform 1 0 195568 0 1 78205
box 0 0 1 1
use contact_32  contact_32_811
timestamp 1624857261
transform 1 0 195432 0 1 93845
box 0 0 1 1
use contact_32  contact_32_810
timestamp 1624857261
transform 1 0 195432 0 1 93573
box 0 0 1 1
use contact_32  contact_32_809
timestamp 1624857261
transform 1 0 195432 0 1 93981
box 0 0 1 1
use contact_32  contact_32_808
timestamp 1624857261
transform 1 0 195432 0 1 94253
box 0 0 1 1
use contact_32  contact_32_807
timestamp 1624857261
transform 1 0 195432 0 1 118325
box 0 0 1 1
use contact_32  contact_32_806
timestamp 1624857261
transform 1 0 195432 0 1 118053
box 0 0 1 1
use contact_32  contact_32_805
timestamp 1624857261
transform 1 0 195432 0 1 118461
box 0 0 1 1
use contact_32  contact_32_804
timestamp 1624857261
transform 1 0 195432 0 1 118733
box 0 0 1 1
use contact_32  contact_32_803
timestamp 1624857261
transform 1 0 195432 0 1 111253
box 0 0 1 1
use contact_32  contact_32_802
timestamp 1624857261
transform 1 0 195432 0 1 110981
box 0 0 1 1
use contact_32  contact_32_801
timestamp 1624857261
transform 1 0 195568 0 1 119685
box 0 0 1 1
use contact_32  contact_32_800
timestamp 1624857261
transform 1 0 195568 0 1 119957
box 0 0 1 1
use contact_32  contact_32_799
timestamp 1624857261
transform 1 0 195432 0 1 119549
box 0 0 1 1
use contact_32  contact_32_798
timestamp 1624857261
transform 1 0 195432 0 1 119277
box 0 0 1 1
use contact_32  contact_32_797
timestamp 1624857261
transform 1 0 195568 0 1 97381
box 0 0 1 1
use contact_32  contact_32_796
timestamp 1624857261
transform 1 0 195568 0 1 97109
box 0 0 1 1
use contact_32  contact_32_795
timestamp 1624857261
transform 1 0 195568 0 1 112205
box 0 0 1 1
use contact_32  contact_32_794
timestamp 1624857261
transform 1 0 195568 0 1 112477
box 0 0 1 1
use contact_32  contact_32_793
timestamp 1624857261
transform 1 0 195432 0 1 27613
box 0 0 1 1
use contact_32  contact_32_792
timestamp 1624857261
transform 1 0 195432 0 1 27885
box 0 0 1 1
use contact_32  contact_32_791
timestamp 1624857261
transform 1 0 195432 0 1 27477
box 0 0 1 1
use contact_32  contact_32_790
timestamp 1624857261
transform 1 0 195432 0 1 27205
box 0 0 1 1
use contact_32  contact_32_789
timestamp 1624857261
transform 1 0 195432 0 1 28021
box 0 0 1 1
use contact_32  contact_32_788
timestamp 1624857261
transform 1 0 195432 0 1 28293
box 0 0 1 1
use contact_32  contact_32_787
timestamp 1624857261
transform 1 0 195432 0 1 117917
box 0 0 1 1
use contact_32  contact_32_786
timestamp 1624857261
transform 1 0 195432 0 1 117645
box 0 0 1 1
use contact_32  contact_32_785
timestamp 1624857261
transform 1 0 195568 0 1 79021
box 0 0 1 1
use contact_32  contact_32_784
timestamp 1624857261
transform 1 0 195568 0 1 79293
box 0 0 1 1
use contact_32  contact_32_783
timestamp 1624857261
transform 1 0 195568 0 1 95205
box 0 0 1 1
use contact_32  contact_32_782
timestamp 1624857261
transform 1 0 195568 0 1 95477
box 0 0 1 1
use contact_32  contact_32_781
timestamp 1624857261
transform 1 0 195432 0 1 81197
box 0 0 1 1
use contact_32  contact_32_780
timestamp 1624857261
transform 1 0 195432 0 1 80925
box 0 0 1 1
use contact_32  contact_32_779
timestamp 1624857261
transform 1 0 195432 0 1 81333
box 0 0 1 1
use contact_32  contact_32_778
timestamp 1624857261
transform 1 0 195432 0 1 81605
box 0 0 1 1
use contact_32  contact_32_777
timestamp 1624857261
transform 1 0 195568 0 1 72901
box 0 0 1 1
use contact_32  contact_32_776
timestamp 1624857261
transform 1 0 195568 0 1 72629
box 0 0 1 1
use contact_32  contact_32_775
timestamp 1624857261
transform 1 0 195432 0 1 115605
box 0 0 1 1
use contact_32  contact_32_774
timestamp 1624857261
transform 1 0 195432 0 1 115333
box 0 0 1 1
use contact_32  contact_32_773
timestamp 1624857261
transform 1 0 195432 0 1 103773
box 0 0 1 1
use contact_32  contact_32_772
timestamp 1624857261
transform 1 0 195432 0 1 103501
box 0 0 1 1
use contact_32  contact_32_771
timestamp 1624857261
transform 1 0 195568 0 1 103909
box 0 0 1 1
use contact_32  contact_32_770
timestamp 1624857261
transform 1 0 195568 0 1 104181
box 0 0 1 1
use contact_32  contact_32_769
timestamp 1624857261
transform 1 0 195432 0 1 66781
box 0 0 1 1
use contact_32  contact_32_768
timestamp 1624857261
transform 1 0 195432 0 1 67053
box 0 0 1 1
use contact_32  contact_32_767
timestamp 1624857261
transform 1 0 195432 0 1 66645
box 0 0 1 1
use contact_32  contact_32_766
timestamp 1624857261
transform 1 0 195432 0 1 66373
box 0 0 1 1
use contact_32  contact_32_765
timestamp 1624857261
transform 1 0 195568 0 1 53317
box 0 0 1 1
use contact_32  contact_32_764
timestamp 1624857261
transform 1 0 195568 0 1 53589
box 0 0 1 1
use contact_32  contact_32_763
timestamp 1624857261
transform 1 0 195432 0 1 53181
box 0 0 1 1
use contact_32  contact_32_762
timestamp 1624857261
transform 1 0 195432 0 1 52909
box 0 0 1 1
use contact_32  contact_32_761
timestamp 1624857261
transform 1 0 195432 0 1 122813
box 0 0 1 1
use contact_32  contact_32_760
timestamp 1624857261
transform 1 0 195432 0 1 123085
box 0 0 1 1
use contact_32  contact_32_759
timestamp 1624857261
transform 1 0 195432 0 1 85277
box 0 0 1 1
use contact_32  contact_32_758
timestamp 1624857261
transform 1 0 195432 0 1 85549
box 0 0 1 1
use contact_32  contact_32_757
timestamp 1624857261
transform 1 0 195568 0 1 85957
box 0 0 1 1
use contact_32  contact_32_756
timestamp 1624857261
transform 1 0 195568 0 1 85685
box 0 0 1 1
use contact_32  contact_32_755
timestamp 1624857261
transform 1 0 195432 0 1 62293
box 0 0 1 1
use contact_32  contact_32_754
timestamp 1624857261
transform 1 0 195432 0 1 62021
box 0 0 1 1
use contact_32  contact_32_753
timestamp 1624857261
transform 1 0 195432 0 1 62429
box 0 0 1 1
use contact_32  contact_32_752
timestamp 1624857261
transform 1 0 195432 0 1 62701
box 0 0 1 1
use contact_32  contact_32_751
timestamp 1624857261
transform 1 0 195568 0 1 39717
box 0 0 1 1
use contact_32  contact_32_750
timestamp 1624857261
transform 1 0 195568 0 1 39445
box 0 0 1 1
use contact_32  contact_32_749
timestamp 1624857261
transform 1 0 195568 0 1 39853
box 0 0 1 1
use contact_32  contact_32_748
timestamp 1624857261
transform 1 0 195568 0 1 40125
box 0 0 1 1
use contact_32  contact_32_747
timestamp 1624857261
transform 1 0 195432 0 1 51957
box 0 0 1 1
use contact_32  contact_32_746
timestamp 1624857261
transform 1 0 195432 0 1 51685
box 0 0 1 1
use contact_32  contact_32_745
timestamp 1624857261
transform 1 0 195432 0 1 52093
box 0 0 1 1
use contact_32  contact_32_744
timestamp 1624857261
transform 1 0 195432 0 1 52365
box 0 0 1 1
use contact_32  contact_32_743
timestamp 1624857261
transform 1 0 195432 0 1 48829
box 0 0 1 1
use contact_32  contact_32_742
timestamp 1624857261
transform 1 0 195432 0 1 48557
box 0 0 1 1
use contact_32  contact_32_741
timestamp 1624857261
transform 1 0 195568 0 1 48965
box 0 0 1 1
use contact_32  contact_32_740
timestamp 1624857261
transform 1 0 195568 0 1 49237
box 0 0 1 1
use contact_32  contact_32_739
timestamp 1624857261
transform 1 0 195432 0 1 37813
box 0 0 1 1
use contact_32  contact_32_738
timestamp 1624857261
transform 1 0 195432 0 1 37541
box 0 0 1 1
use contact_32  contact_32_737
timestamp 1624857261
transform 1 0 195432 0 1 37949
box 0 0 1 1
use contact_32  contact_32_736
timestamp 1624857261
transform 1 0 195432 0 1 38221
box 0 0 1 1
use contact_32  contact_32_735
timestamp 1624857261
transform 1 0 195568 0 1 95885
box 0 0 1 1
use contact_32  contact_32_734
timestamp 1624857261
transform 1 0 195568 0 1 95613
box 0 0 1 1
use contact_32  contact_32_733
timestamp 1624857261
transform 1 0 195432 0 1 65421
box 0 0 1 1
use contact_32  contact_32_732
timestamp 1624857261
transform 1 0 195432 0 1 65149
box 0 0 1 1
use contact_32  contact_32_731
timestamp 1624857261
transform 1 0 195568 0 1 65557
box 0 0 1 1
use contact_32  contact_32_730
timestamp 1624857261
transform 1 0 195568 0 1 65829
box 0 0 1 1
use contact_32  contact_32_729
timestamp 1624857261
transform 1 0 195568 0 1 103365
box 0 0 1 1
use contact_32  contact_32_728
timestamp 1624857261
transform 1 0 195568 0 1 103093
box 0 0 1 1
use contact_32  contact_32_727
timestamp 1624857261
transform 1 0 195432 0 1 124445
box 0 0 1 1
use contact_32  contact_32_726
timestamp 1624857261
transform 1 0 195432 0 1 124717
box 0 0 1 1
use contact_32  contact_32_725
timestamp 1624857261
transform 1 0 195432 0 1 115197
box 0 0 1 1
use contact_32  contact_32_724
timestamp 1624857261
transform 1 0 195432 0 1 114925
box 0 0 1 1
use contact_32  contact_32_723
timestamp 1624857261
transform 1 0 195432 0 1 39037
box 0 0 1 1
use contact_32  contact_32_722
timestamp 1624857261
transform 1 0 195432 0 1 39309
box 0 0 1 1
use contact_32  contact_32_721
timestamp 1624857261
transform 1 0 195432 0 1 29653
box 0 0 1 1
use contact_32  contact_32_720
timestamp 1624857261
transform 1 0 195432 0 1 29925
box 0 0 1 1
use contact_32  contact_32_719
timestamp 1624857261
transform 1 0 195432 0 1 60661
box 0 0 1 1
use contact_32  contact_32_718
timestamp 1624857261
transform 1 0 195432 0 1 60389
box 0 0 1 1
use contact_32  contact_32_717
timestamp 1624857261
transform 1 0 195432 0 1 60797
box 0 0 1 1
use contact_32  contact_32_716
timestamp 1624857261
transform 1 0 195432 0 1 61069
box 0 0 1 1
use contact_32  contact_32_715
timestamp 1624857261
transform 1 0 195568 0 1 123493
box 0 0 1 1
use contact_32  contact_32_714
timestamp 1624857261
transform 1 0 195568 0 1 123221
box 0 0 1 1
use contact_32  contact_32_713
timestamp 1624857261
transform 1 0 195432 0 1 50461
box 0 0 1 1
use contact_32  contact_32_712
timestamp 1624857261
transform 1 0 195432 0 1 50189
box 0 0 1 1
use contact_32  contact_32_711
timestamp 1624857261
transform 1 0 195568 0 1 41349
box 0 0 1 1
use contact_32  contact_32_710
timestamp 1624857261
transform 1 0 195568 0 1 41077
box 0 0 1 1
use contact_32  contact_32_709
timestamp 1624857261
transform 1 0 195432 0 1 101325
box 0 0 1 1
use contact_32  contact_32_708
timestamp 1624857261
transform 1 0 195432 0 1 101053
box 0 0 1 1
use contact_32  contact_32_707
timestamp 1624857261
transform 1 0 195432 0 1 101461
box 0 0 1 1
use contact_32  contact_32_706
timestamp 1624857261
transform 1 0 195432 0 1 101733
box 0 0 1 1
use contact_32  contact_32_705
timestamp 1624857261
transform 1 0 195568 0 1 98605
box 0 0 1 1
use contact_32  contact_32_704
timestamp 1624857261
transform 1 0 195568 0 1 98333
box 0 0 1 1
use contact_32  contact_32_703
timestamp 1624857261
transform 1 0 195432 0 1 68957
box 0 0 1 1
use contact_32  contact_32_702
timestamp 1624857261
transform 1 0 195432 0 1 68685
box 0 0 1 1
use contact_32  contact_32_701
timestamp 1624857261
transform 1 0 195568 0 1 69093
box 0 0 1 1
use contact_32  contact_32_700
timestamp 1624857261
transform 1 0 195568 0 1 69365
box 0 0 1 1
use contact_32  contact_32_699
timestamp 1624857261
transform 1 0 195568 0 1 107717
box 0 0 1 1
use contact_32  contact_32_698
timestamp 1624857261
transform 1 0 195568 0 1 107445
box 0 0 1 1
use contact_32  contact_32_697
timestamp 1624857261
transform 1 0 195568 0 1 37133
box 0 0 1 1
use contact_32  contact_32_696
timestamp 1624857261
transform 1 0 195568 0 1 37405
box 0 0 1 1
use contact_32  contact_32_695
timestamp 1624857261
transform 1 0 195568 0 1 36997
box 0 0 1 1
use contact_32  contact_32_694
timestamp 1624857261
transform 1 0 195568 0 1 36725
box 0 0 1 1
use contact_32  contact_32_693
timestamp 1624857261
transform 1 0 195568 0 1 32781
box 0 0 1 1
use contact_32  contact_32_692
timestamp 1624857261
transform 1 0 195568 0 1 33053
box 0 0 1 1
use contact_32  contact_32_691
timestamp 1624857261
transform 1 0 195432 0 1 35773
box 0 0 1 1
use contact_32  contact_32_690
timestamp 1624857261
transform 1 0 195432 0 1 35501
box 0 0 1 1
use contact_32  contact_32_689
timestamp 1624857261
transform 1 0 195432 0 1 76981
box 0 0 1 1
use contact_32  contact_32_688
timestamp 1624857261
transform 1 0 195432 0 1 77253
box 0 0 1 1
use contact_32  contact_32_687
timestamp 1624857261
transform 1 0 195432 0 1 76845
box 0 0 1 1
use contact_32  contact_32_686
timestamp 1624857261
transform 1 0 195432 0 1 76573
box 0 0 1 1
use contact_32  contact_32_685
timestamp 1624857261
transform 1 0 195432 0 1 52501
box 0 0 1 1
use contact_32  contact_32_684
timestamp 1624857261
transform 1 0 195432 0 1 52773
box 0 0 1 1
use contact_32  contact_32_683
timestamp 1624857261
transform 1 0 195568 0 1 102277
box 0 0 1 1
use contact_32  contact_32_682
timestamp 1624857261
transform 1 0 195568 0 1 102549
box 0 0 1 1
use contact_32  contact_32_681
timestamp 1624857261
transform 1 0 195432 0 1 102141
box 0 0 1 1
use contact_32  contact_32_680
timestamp 1624857261
transform 1 0 195432 0 1 101869
box 0 0 1 1
use contact_32  contact_32_679
timestamp 1624857261
transform 1 0 195432 0 1 82557
box 0 0 1 1
use contact_32  contact_32_678
timestamp 1624857261
transform 1 0 195432 0 1 82829
box 0 0 1 1
use contact_32  contact_32_677
timestamp 1624857261
transform 1 0 195432 0 1 82421
box 0 0 1 1
use contact_32  contact_32_676
timestamp 1624857261
transform 1 0 195432 0 1 82149
box 0 0 1 1
use contact_32  contact_32_675
timestamp 1624857261
transform 1 0 195568 0 1 90445
box 0 0 1 1
use contact_32  contact_32_674
timestamp 1624857261
transform 1 0 195568 0 1 90717
box 0 0 1 1
use contact_32  contact_32_673
timestamp 1624857261
transform 1 0 195568 0 1 90309
box 0 0 1 1
use contact_32  contact_32_672
timestamp 1624857261
transform 1 0 195568 0 1 90037
box 0 0 1 1
use contact_32  contact_32_671
timestamp 1624857261
transform 1 0 195432 0 1 102685
box 0 0 1 1
use contact_32  contact_32_670
timestamp 1624857261
transform 1 0 195432 0 1 102957
box 0 0 1 1
use contact_32  contact_32_669
timestamp 1624857261
transform 1 0 195568 0 1 43661
box 0 0 1 1
use contact_32  contact_32_668
timestamp 1624857261
transform 1 0 195568 0 1 43389
box 0 0 1 1
use contact_32  contact_32_667
timestamp 1624857261
transform 1 0 195568 0 1 80517
box 0 0 1 1
use contact_32  contact_32_666
timestamp 1624857261
transform 1 0 195568 0 1 80789
box 0 0 1 1
use contact_32  contact_32_665
timestamp 1624857261
transform 1 0 195432 0 1 25301
box 0 0 1 1
use contact_32  contact_32_664
timestamp 1624857261
transform 1 0 195432 0 1 25573
box 0 0 1 1
use contact_32  contact_32_663
timestamp 1624857261
transform 1 0 195432 0 1 87181
box 0 0 1 1
use contact_32  contact_32_662
timestamp 1624857261
transform 1 0 195432 0 1 86909
box 0 0 1 1
use contact_32  contact_32_661
timestamp 1624857261
transform 1 0 195568 0 1 90853
box 0 0 1 1
use contact_32  contact_32_660
timestamp 1624857261
transform 1 0 195568 0 1 91125
box 0 0 1 1
use contact_32  contact_32_659
timestamp 1624857261
transform 1 0 195432 0 1 69773
box 0 0 1 1
use contact_32  contact_32_658
timestamp 1624857261
transform 1 0 195432 0 1 69501
box 0 0 1 1
use contact_32  contact_32_657
timestamp 1624857261
transform 1 0 195432 0 1 69909
box 0 0 1 1
use contact_32  contact_32_656
timestamp 1624857261
transform 1 0 195432 0 1 70181
box 0 0 1 1
use contact_32  contact_32_655
timestamp 1624857261
transform 1 0 195432 0 1 78069
box 0 0 1 1
use contact_32  contact_32_654
timestamp 1624857261
transform 1 0 195432 0 1 77797
box 0 0 1 1
use contact_32  contact_32_653
timestamp 1624857261
transform 1 0 195568 0 1 48421
box 0 0 1 1
use contact_32  contact_32_652
timestamp 1624857261
transform 1 0 195568 0 1 48149
box 0 0 1 1
use contact_32  contact_32_651
timestamp 1624857261
transform 1 0 195432 0 1 83645
box 0 0 1 1
use contact_32  contact_32_650
timestamp 1624857261
transform 1 0 195432 0 1 83373
box 0 0 1 1
use contact_32  contact_32_649
timestamp 1624857261
transform 1 0 195432 0 1 77661
box 0 0 1 1
use contact_32  contact_32_648
timestamp 1624857261
transform 1 0 195432 0 1 77389
box 0 0 1 1
use contact_32  contact_32_647
timestamp 1624857261
transform 1 0 195568 0 1 83237
box 0 0 1 1
use contact_32  contact_32_646
timestamp 1624857261
transform 1 0 195568 0 1 82965
box 0 0 1 1
use contact_32  contact_32_645
timestamp 1624857261
transform 1 0 195432 0 1 118869
box 0 0 1 1
use contact_32  contact_32_644
timestamp 1624857261
transform 1 0 195432 0 1 119141
box 0 0 1 1
use contact_32  contact_32_643
timestamp 1624857261
transform 1 0 195432 0 1 72493
box 0 0 1 1
use contact_32  contact_32_642
timestamp 1624857261
transform 1 0 195432 0 1 72221
box 0 0 1 1
use contact_32  contact_32_641
timestamp 1624857261
transform 1 0 195432 0 1 75349
box 0 0 1 1
use contact_32  contact_32_640
timestamp 1624857261
transform 1 0 195432 0 1 75077
box 0 0 1 1
use contact_32  contact_32_639
timestamp 1624857261
transform 1 0 195568 0 1 64197
box 0 0 1 1
use contact_32  contact_32_638
timestamp 1624857261
transform 1 0 195568 0 1 63925
box 0 0 1 1
use contact_32  contact_32_637
timestamp 1624857261
transform 1 0 195568 0 1 64333
box 0 0 1 1
use contact_32  contact_32_636
timestamp 1624857261
transform 1 0 195568 0 1 64605
box 0 0 1 1
use contact_32  contact_32_635
timestamp 1624857261
transform 1 0 195432 0 1 49781
box 0 0 1 1
use contact_32  contact_32_634
timestamp 1624857261
transform 1 0 195432 0 1 50053
box 0 0 1 1
use contact_32  contact_32_633
timestamp 1624857261
transform 1 0 195432 0 1 49645
box 0 0 1 1
use contact_32  contact_32_632
timestamp 1624857261
transform 1 0 195432 0 1 49373
box 0 0 1 1
use contact_32  contact_32_631
timestamp 1624857261
transform 1 0 195568 0 1 114789
box 0 0 1 1
use contact_32  contact_32_630
timestamp 1624857261
transform 1 0 195568 0 1 114517
box 0 0 1 1
use contact_32  contact_32_629
timestamp 1624857261
transform 1 0 195432 0 1 110165
box 0 0 1 1
use contact_32  contact_32_628
timestamp 1624857261
transform 1 0 195432 0 1 110437
box 0 0 1 1
use contact_32  contact_32_627
timestamp 1624857261
transform 1 0 195568 0 1 110029
box 0 0 1 1
use contact_32  contact_32_626
timestamp 1624857261
transform 1 0 195568 0 1 109757
box 0 0 1 1
use contact_32  contact_32_625
timestamp 1624857261
transform 1 0 195432 0 1 105405
box 0 0 1 1
use contact_32  contact_32_624
timestamp 1624857261
transform 1 0 195432 0 1 105677
box 0 0 1 1
use contact_32  contact_32_623
timestamp 1624857261
transform 1 0 195568 0 1 105813
box 0 0 1 1
use contact_32  contact_32_622
timestamp 1624857261
transform 1 0 195568 0 1 106085
box 0 0 1 1
use contact_32  contact_32_621
timestamp 1624857261
transform 1 0 195432 0 1 28701
box 0 0 1 1
use contact_32  contact_32_620
timestamp 1624857261
transform 1 0 195432 0 1 28429
box 0 0 1 1
use contact_32  contact_32_619
timestamp 1624857261
transform 1 0 195568 0 1 113701
box 0 0 1 1
use contact_32  contact_32_618
timestamp 1624857261
transform 1 0 195568 0 1 113973
box 0 0 1 1
use contact_32  contact_32_617
timestamp 1624857261
transform 1 0 195568 0 1 110573
box 0 0 1 1
use contact_32  contact_32_616
timestamp 1624857261
transform 1 0 195568 0 1 110845
box 0 0 1 1
use contact_32  contact_32_615
timestamp 1624857261
transform 1 0 195432 0 1 74941
box 0 0 1 1
use contact_32  contact_32_614
timestamp 1624857261
transform 1 0 195432 0 1 74669
box 0 0 1 1
use contact_32  contact_32_613
timestamp 1624857261
transform 1 0 195432 0 1 74261
box 0 0 1 1
use contact_32  contact_32_612
timestamp 1624857261
transform 1 0 195432 0 1 74533
box 0 0 1 1
use contact_32  contact_32_611
timestamp 1624857261
transform 1 0 195568 0 1 64741
box 0 0 1 1
use contact_32  contact_32_610
timestamp 1624857261
transform 1 0 195568 0 1 65013
box 0 0 1 1
use contact_32  contact_32_609
timestamp 1624857261
transform 1 0 195432 0 1 60253
box 0 0 1 1
use contact_32  contact_32_608
timestamp 1624857261
transform 1 0 195432 0 1 59981
box 0 0 1 1
use contact_32  contact_32_607
timestamp 1624857261
transform 1 0 195568 0 1 68549
box 0 0 1 1
use contact_32  contact_32_606
timestamp 1624857261
transform 1 0 195568 0 1 68277
box 0 0 1 1
use contact_32  contact_32_605
timestamp 1624857261
transform 1 0 195568 0 1 33189
box 0 0 1 1
use contact_32  contact_32_604
timestamp 1624857261
transform 1 0 195568 0 1 33461
box 0 0 1 1
use contact_32  contact_32_603
timestamp 1624857261
transform 1 0 195432 0 1 89085
box 0 0 1 1
use contact_32  contact_32_602
timestamp 1624857261
transform 1 0 195432 0 1 88813
box 0 0 1 1
use contact_32  contact_32_601
timestamp 1624857261
transform 1 0 195432 0 1 66237
box 0 0 1 1
use contact_32  contact_32_600
timestamp 1624857261
transform 1 0 195432 0 1 65965
box 0 0 1 1
use contact_32  contact_32_599
timestamp 1624857261
transform 1 0 195568 0 1 106221
box 0 0 1 1
use contact_32  contact_32_598
timestamp 1624857261
transform 1 0 195568 0 1 106493
box 0 0 1 1
use contact_32  contact_32_597
timestamp 1624857261
transform 1 0 195432 0 1 31421
box 0 0 1 1
use contact_32  contact_32_596
timestamp 1624857261
transform 1 0 195432 0 1 31149
box 0 0 1 1
use contact_32  contact_32_595
timestamp 1624857261
transform 1 0 195568 0 1 109349
box 0 0 1 1
use contact_32  contact_32_594
timestamp 1624857261
transform 1 0 195568 0 1 109621
box 0 0 1 1
use contact_32  contact_32_593
timestamp 1624857261
transform 1 0 195432 0 1 114109
box 0 0 1 1
use contact_32  contact_32_592
timestamp 1624857261
transform 1 0 195432 0 1 114381
box 0 0 1 1
use contact_32  contact_32_591
timestamp 1624857261
transform 1 0 195432 0 1 82013
box 0 0 1 1
use contact_32  contact_32_590
timestamp 1624857261
transform 1 0 195432 0 1 81741
box 0 0 1 1
use contact_32  contact_32_589
timestamp 1624857261
transform 1 0 195568 0 1 26797
box 0 0 1 1
use contact_32  contact_32_588
timestamp 1624857261
transform 1 0 195568 0 1 27069
box 0 0 1 1
use contact_32  contact_32_587
timestamp 1624857261
transform 1 0 196656 0 1 131381
box 0 0 1 1
use contact_32  contact_32_586
timestamp 1624857261
transform 1 0 196656 0 1 134101
box 0 0 1 1
use contact_32  contact_32_585
timestamp 1624857261
transform 1 0 196656 0 1 128389
box 0 0 1 1
use contact_32  contact_32_584
timestamp 1624857261
transform 1 0 196656 0 1 125669
box 0 0 1 1
use contact_32  contact_32_583
timestamp 1624857261
transform 1 0 196656 0 1 83237
box 0 0 1 1
use contact_32  contact_32_582
timestamp 1624857261
transform 1 0 196656 0 1 82965
box 0 0 1 1
use contact_32  contact_32_581
timestamp 1624857261
transform 1 0 196656 0 1 83373
box 0 0 1 1
use contact_32  contact_32_580
timestamp 1624857261
transform 1 0 196656 0 1 83645
box 0 0 1 1
use contact_32  contact_32_579
timestamp 1624857261
transform 1 0 196656 0 1 70181
box 0 0 1 1
use contact_32  contact_32_578
timestamp 1624857261
transform 1 0 196656 0 1 69909
box 0 0 1 1
use contact_32  contact_32_577
timestamp 1624857261
transform 1 0 196656 0 1 70317
box 0 0 1 1
use contact_32  contact_32_576
timestamp 1624857261
transform 1 0 196656 0 1 70589
box 0 0 1 1
use contact_32  contact_32_575
timestamp 1624857261
transform 1 0 196792 0 1 106901
box 0 0 1 1
use contact_32  contact_32_574
timestamp 1624857261
transform 1 0 196792 0 1 106629
box 0 0 1 1
use contact_32  contact_32_573
timestamp 1624857261
transform 1 0 196792 0 1 107037
box 0 0 1 1
use contact_32  contact_32_572
timestamp 1624857261
transform 1 0 196792 0 1 107309
box 0 0 1 1
use contact_32  contact_32_571
timestamp 1624857261
transform 1 0 196656 0 1 73853
box 0 0 1 1
use contact_32  contact_32_570
timestamp 1624857261
transform 1 0 196656 0 1 74125
box 0 0 1 1
use contact_32  contact_32_569
timestamp 1624857261
transform 1 0 196656 0 1 73717
box 0 0 1 1
use contact_32  contact_32_568
timestamp 1624857261
transform 1 0 196656 0 1 73445
box 0 0 1 1
use contact_32  contact_32_567
timestamp 1624857261
transform 1 0 196792 0 1 99421
box 0 0 1 1
use contact_32  contact_32_566
timestamp 1624857261
transform 1 0 196792 0 1 99149
box 0 0 1 1
use contact_32  contact_32_565
timestamp 1624857261
transform 1 0 196656 0 1 99557
box 0 0 1 1
use contact_32  contact_32_564
timestamp 1624857261
transform 1 0 196656 0 1 99829
box 0 0 1 1
use contact_32  contact_32_563
timestamp 1624857261
transform 1 0 196656 0 1 104317
box 0 0 1 1
use contact_32  contact_32_562
timestamp 1624857261
transform 1 0 196656 0 1 104589
box 0 0 1 1
use contact_32  contact_32_561
timestamp 1624857261
transform 1 0 196656 0 1 104181
box 0 0 1 1
use contact_32  contact_32_560
timestamp 1624857261
transform 1 0 196656 0 1 103909
box 0 0 1 1
use contact_32  contact_32_559
timestamp 1624857261
transform 1 0 196792 0 1 107717
box 0 0 1 1
use contact_32  contact_32_558
timestamp 1624857261
transform 1 0 196792 0 1 107445
box 0 0 1 1
use contact_32  contact_32_557
timestamp 1624857261
transform 1 0 196792 0 1 107853
box 0 0 1 1
use contact_32  contact_32_556
timestamp 1624857261
transform 1 0 196792 0 1 108125
box 0 0 1 1
use contact_32  contact_32_555
timestamp 1624857261
transform 1 0 196792 0 1 58757
box 0 0 1 1
use contact_32  contact_32_554
timestamp 1624857261
transform 1 0 196792 0 1 58485
box 0 0 1 1
use contact_32  contact_32_553
timestamp 1624857261
transform 1 0 196792 0 1 58893
box 0 0 1 1
use contact_32  contact_32_552
timestamp 1624857261
transform 1 0 196792 0 1 59165
box 0 0 1 1
use contact_32  contact_32_551
timestamp 1624857261
transform 1 0 196792 0 1 114517
box 0 0 1 1
use contact_32  contact_32_550
timestamp 1624857261
transform 1 0 196792 0 1 114789
box 0 0 1 1
use contact_32  contact_32_549
timestamp 1624857261
transform 1 0 196792 0 1 69773
box 0 0 1 1
use contact_32  contact_32_548
timestamp 1624857261
transform 1 0 196792 0 1 69501
box 0 0 1 1
use contact_32  contact_32_547
timestamp 1624857261
transform 1 0 196792 0 1 121181
box 0 0 1 1
use contact_32  contact_32_546
timestamp 1624857261
transform 1 0 196792 0 1 120909
box 0 0 1 1
use contact_32  contact_32_545
timestamp 1624857261
transform 1 0 196656 0 1 121317
box 0 0 1 1
use contact_32  contact_32_544
timestamp 1624857261
transform 1 0 196656 0 1 121589
box 0 0 1 1
use contact_32  contact_32_543
timestamp 1624857261
transform 1 0 196792 0 1 41349
box 0 0 1 1
use contact_32  contact_32_542
timestamp 1624857261
transform 1 0 196792 0 1 41077
box 0 0 1 1
use contact_32  contact_32_541
timestamp 1624857261
transform 1 0 196792 0 1 41485
box 0 0 1 1
use contact_32  contact_32_540
timestamp 1624857261
transform 1 0 196792 0 1 41757
box 0 0 1 1
use contact_32  contact_32_539
timestamp 1624857261
transform 1 0 196656 0 1 30877
box 0 0 1 1
use contact_32  contact_32_538
timestamp 1624857261
transform 1 0 196656 0 1 31149
box 0 0 1 1
use contact_32  contact_32_537
timestamp 1624857261
transform 1 0 196656 0 1 87725
box 0 0 1 1
use contact_32  contact_32_536
timestamp 1624857261
transform 1 0 196656 0 1 87997
box 0 0 1 1
use contact_32  contact_32_535
timestamp 1624857261
transform 1 0 196656 0 1 87589
box 0 0 1 1
use contact_32  contact_32_534
timestamp 1624857261
transform 1 0 196656 0 1 87317
box 0 0 1 1
use contact_32  contact_32_533
timestamp 1624857261
transform 1 0 196656 0 1 122405
box 0 0 1 1
use contact_32  contact_32_532
timestamp 1624857261
transform 1 0 196656 0 1 122677
box 0 0 1 1
use contact_32  contact_32_531
timestamp 1624857261
transform 1 0 196792 0 1 115333
box 0 0 1 1
use contact_32  contact_32_530
timestamp 1624857261
transform 1 0 196792 0 1 115605
box 0 0 1 1
use contact_32  contact_32_529
timestamp 1624857261
transform 1 0 196656 0 1 115197
box 0 0 1 1
use contact_32  contact_32_528
timestamp 1624857261
transform 1 0 196656 0 1 114925
box 0 0 1 1
use contact_32  contact_32_527
timestamp 1624857261
transform 1 0 196792 0 1 32645
box 0 0 1 1
use contact_32  contact_32_526
timestamp 1624857261
transform 1 0 196792 0 1 32373
box 0 0 1 1
use contact_32  contact_32_525
timestamp 1624857261
transform 1 0 196792 0 1 32781
box 0 0 1 1
use contact_32  contact_32_524
timestamp 1624857261
transform 1 0 196792 0 1 33053
box 0 0 1 1
use contact_32  contact_32_523
timestamp 1624857261
transform 1 0 196656 0 1 31829
box 0 0 1 1
use contact_32  contact_32_522
timestamp 1624857261
transform 1 0 196656 0 1 31557
box 0 0 1 1
use contact_32  contact_32_521
timestamp 1624857261
transform 1 0 196792 0 1 85277
box 0 0 1 1
use contact_32  contact_32_520
timestamp 1624857261
transform 1 0 196792 0 1 85549
box 0 0 1 1
use contact_32  contact_32_519
timestamp 1624857261
transform 1 0 196656 0 1 112885
box 0 0 1 1
use contact_32  contact_32_518
timestamp 1624857261
transform 1 0 196656 0 1 112613
box 0 0 1 1
use contact_32  contact_32_517
timestamp 1624857261
transform 1 0 196656 0 1 113021
box 0 0 1 1
use contact_32  contact_32_516
timestamp 1624857261
transform 1 0 196656 0 1 113293
box 0 0 1 1
use contact_32  contact_32_515
timestamp 1624857261
transform 1 0 196792 0 1 62293
box 0 0 1 1
use contact_32  contact_32_514
timestamp 1624857261
transform 1 0 196792 0 1 62021
box 0 0 1 1
use contact_32  contact_32_513
timestamp 1624857261
transform 1 0 196792 0 1 62429
box 0 0 1 1
use contact_32  contact_32_512
timestamp 1624857261
transform 1 0 196792 0 1 62701
box 0 0 1 1
use contact_32  contact_32_511
timestamp 1624857261
transform 1 0 196792 0 1 84053
box 0 0 1 1
use contact_32  contact_32_510
timestamp 1624857261
transform 1 0 196792 0 1 83781
box 0 0 1 1
use contact_32  contact_32_509
timestamp 1624857261
transform 1 0 196792 0 1 108941
box 0 0 1 1
use contact_32  contact_32_508
timestamp 1624857261
transform 1 0 196792 0 1 108669
box 0 0 1 1
use contact_32  contact_32_507
timestamp 1624857261
transform 1 0 196792 0 1 109077
box 0 0 1 1
use contact_32  contact_32_506
timestamp 1624857261
transform 1 0 196792 0 1 109349
box 0 0 1 1
use contact_32  contact_32_505
timestamp 1624857261
transform 1 0 196792 0 1 104725
box 0 0 1 1
use contact_32  contact_32_504
timestamp 1624857261
transform 1 0 196792 0 1 104997
box 0 0 1 1
use contact_32  contact_32_503
timestamp 1624857261
transform 1 0 196656 0 1 52909
box 0 0 1 1
use contact_32  contact_32_502
timestamp 1624857261
transform 1 0 196656 0 1 53181
box 0 0 1 1
use contact_32  contact_32_501
timestamp 1624857261
transform 1 0 196792 0 1 95069
box 0 0 1 1
use contact_32  contact_32_500
timestamp 1624857261
transform 1 0 196792 0 1 94797
box 0 0 1 1
use contact_32  contact_32_499
timestamp 1624857261
transform 1 0 196656 0 1 95205
box 0 0 1 1
use contact_32  contact_32_498
timestamp 1624857261
transform 1 0 196656 0 1 95477
box 0 0 1 1
use contact_32  contact_32_497
timestamp 1624857261
transform 1 0 196792 0 1 99013
box 0 0 1 1
use contact_32  contact_32_496
timestamp 1624857261
transform 1 0 196792 0 1 98741
box 0 0 1 1
use contact_32  contact_32_495
timestamp 1624857261
transform 1 0 196656 0 1 34685
box 0 0 1 1
use contact_32  contact_32_494
timestamp 1624857261
transform 1 0 196656 0 1 34413
box 0 0 1 1
use contact_32  contact_32_493
timestamp 1624857261
transform 1 0 196792 0 1 34821
box 0 0 1 1
use contact_32  contact_32_492
timestamp 1624857261
transform 1 0 196792 0 1 35093
box 0 0 1 1
use contact_32  contact_32_491
timestamp 1624857261
transform 1 0 196792 0 1 27613
box 0 0 1 1
use contact_32  contact_32_490
timestamp 1624857261
transform 1 0 196792 0 1 27885
box 0 0 1 1
use contact_32  contact_32_489
timestamp 1624857261
transform 1 0 196656 0 1 110845
box 0 0 1 1
use contact_32  contact_32_488
timestamp 1624857261
transform 1 0 196656 0 1 110573
box 0 0 1 1
use contact_32  contact_32_487
timestamp 1624857261
transform 1 0 196792 0 1 110981
box 0 0 1 1
use contact_32  contact_32_486
timestamp 1624857261
transform 1 0 196792 0 1 111253
box 0 0 1 1
use contact_32  contact_32_485
timestamp 1624857261
transform 1 0 196656 0 1 38629
box 0 0 1 1
use contact_32  contact_32_484
timestamp 1624857261
transform 1 0 196656 0 1 38357
box 0 0 1 1
use contact_32  contact_32_483
timestamp 1624857261
transform 1 0 196656 0 1 38765
box 0 0 1 1
use contact_32  contact_32_482
timestamp 1624857261
transform 1 0 196656 0 1 39037
box 0 0 1 1
use contact_32  contact_32_481
timestamp 1624857261
transform 1 0 196792 0 1 124037
box 0 0 1 1
use contact_32  contact_32_480
timestamp 1624857261
transform 1 0 196792 0 1 124309
box 0 0 1 1
use contact_32  contact_32_479
timestamp 1624857261
transform 1 0 196656 0 1 123901
box 0 0 1 1
use contact_32  contact_32_478
timestamp 1624857261
transform 1 0 196656 0 1 123629
box 0 0 1 1
use contact_32  contact_32_477
timestamp 1624857261
transform 1 0 196656 0 1 45293
box 0 0 1 1
use contact_32  contact_32_476
timestamp 1624857261
transform 1 0 196656 0 1 45021
box 0 0 1 1
use contact_32  contact_32_475
timestamp 1624857261
transform 1 0 196656 0 1 45429
box 0 0 1 1
use contact_32  contact_32_474
timestamp 1624857261
transform 1 0 196656 0 1 45701
box 0 0 1 1
use contact_32  contact_32_473
timestamp 1624857261
transform 1 0 196656 0 1 46245
box 0 0 1 1
use contact_32  contact_32_472
timestamp 1624857261
transform 1 0 196656 0 1 46517
box 0 0 1 1
use contact_32  contact_32_471
timestamp 1624857261
transform 1 0 196792 0 1 46109
box 0 0 1 1
use contact_32  contact_32_470
timestamp 1624857261
transform 1 0 196792 0 1 45837
box 0 0 1 1
use contact_32  contact_32_469
timestamp 1624857261
transform 1 0 196792 0 1 28293
box 0 0 1 1
use contact_32  contact_32_468
timestamp 1624857261
transform 1 0 196792 0 1 28021
box 0 0 1 1
use contact_32  contact_32_467
timestamp 1624857261
transform 1 0 196792 0 1 28429
box 0 0 1 1
use contact_32  contact_32_466
timestamp 1624857261
transform 1 0 196792 0 1 28701
box 0 0 1 1
use contact_32  contact_32_465
timestamp 1624857261
transform 1 0 196792 0 1 119957
box 0 0 1 1
use contact_32  contact_32_464
timestamp 1624857261
transform 1 0 196792 0 1 119685
box 0 0 1 1
use contact_32  contact_32_463
timestamp 1624857261
transform 1 0 196792 0 1 120093
box 0 0 1 1
use contact_32  contact_32_462
timestamp 1624857261
transform 1 0 196792 0 1 120365
box 0 0 1 1
use contact_32  contact_32_461
timestamp 1624857261
transform 1 0 196792 0 1 36997
box 0 0 1 1
use contact_32  contact_32_460
timestamp 1624857261
transform 1 0 196792 0 1 36725
box 0 0 1 1
use contact_32  contact_32_459
timestamp 1624857261
transform 1 0 196792 0 1 37133
box 0 0 1 1
use contact_32  contact_32_458
timestamp 1624857261
transform 1 0 196792 0 1 37405
box 0 0 1 1
use contact_32  contact_32_457
timestamp 1624857261
transform 1 0 196792 0 1 112477
box 0 0 1 1
use contact_32  contact_32_456
timestamp 1624857261
transform 1 0 196792 0 1 112205
box 0 0 1 1
use contact_32  contact_32_455
timestamp 1624857261
transform 1 0 196656 0 1 40941
box 0 0 1 1
use contact_32  contact_32_454
timestamp 1624857261
transform 1 0 196656 0 1 40669
box 0 0 1 1
use contact_32  contact_32_453
timestamp 1624857261
transform 1 0 196656 0 1 34277
box 0 0 1 1
use contact_32  contact_32_452
timestamp 1624857261
transform 1 0 196656 0 1 34005
box 0 0 1 1
use contact_32  contact_32_451
timestamp 1624857261
transform 1 0 196656 0 1 80653
box 0 0 1 1
use contact_32  contact_32_450
timestamp 1624857261
transform 1 0 196656 0 1 80925
box 0 0 1 1
use contact_32  contact_32_449
timestamp 1624857261
transform 1 0 196792 0 1 44885
box 0 0 1 1
use contact_32  contact_32_448
timestamp 1624857261
transform 1 0 196792 0 1 44613
box 0 0 1 1
use contact_32  contact_32_447
timestamp 1624857261
transform 1 0 196792 0 1 46925
box 0 0 1 1
use contact_32  contact_32_446
timestamp 1624857261
transform 1 0 196792 0 1 46653
box 0 0 1 1
use contact_32  contact_32_445
timestamp 1624857261
transform 1 0 196656 0 1 91125
box 0 0 1 1
use contact_32  contact_32_444
timestamp 1624857261
transform 1 0 196656 0 1 90853
box 0 0 1 1
use contact_32  contact_32_443
timestamp 1624857261
transform 1 0 196656 0 1 91261
box 0 0 1 1
use contact_32  contact_32_442
timestamp 1624857261
transform 1 0 196656 0 1 91533
box 0 0 1 1
use contact_32  contact_32_441
timestamp 1624857261
transform 1 0 196792 0 1 118733
box 0 0 1 1
use contact_32  contact_32_440
timestamp 1624857261
transform 1 0 196792 0 1 118461
box 0 0 1 1
use contact_32  contact_32_439
timestamp 1624857261
transform 1 0 196656 0 1 86773
box 0 0 1 1
use contact_32  contact_32_438
timestamp 1624857261
transform 1 0 196656 0 1 86501
box 0 0 1 1
use contact_32  contact_32_437
timestamp 1624857261
transform 1 0 196656 0 1 86909
box 0 0 1 1
use contact_32  contact_32_436
timestamp 1624857261
transform 1 0 196656 0 1 87181
box 0 0 1 1
use contact_32  contact_32_435
timestamp 1624857261
transform 1 0 196792 0 1 40261
box 0 0 1 1
use contact_32  contact_32_434
timestamp 1624857261
transform 1 0 196792 0 1 40533
box 0 0 1 1
use contact_32  contact_32_433
timestamp 1624857261
transform 1 0 196792 0 1 71813
box 0 0 1 1
use contact_32  contact_32_432
timestamp 1624857261
transform 1 0 196792 0 1 71541
box 0 0 1 1
use contact_32  contact_32_431
timestamp 1624857261
transform 1 0 196792 0 1 71949
box 0 0 1 1
use contact_32  contact_32_430
timestamp 1624857261
transform 1 0 196792 0 1 72221
box 0 0 1 1
use contact_32  contact_32_429
timestamp 1624857261
transform 1 0 196792 0 1 77389
box 0 0 1 1
use contact_32  contact_32_428
timestamp 1624857261
transform 1 0 196792 0 1 77661
box 0 0 1 1
use contact_32  contact_32_427
timestamp 1624857261
transform 1 0 196656 0 1 100645
box 0 0 1 1
use contact_32  contact_32_426
timestamp 1624857261
transform 1 0 196656 0 1 100373
box 0 0 1 1
use contact_32  contact_32_425
timestamp 1624857261
transform 1 0 196792 0 1 86093
box 0 0 1 1
use contact_32  contact_32_424
timestamp 1624857261
transform 1 0 196792 0 1 86365
box 0 0 1 1
use contact_32  contact_32_423
timestamp 1624857261
transform 1 0 196792 0 1 82829
box 0 0 1 1
use contact_32  contact_32_422
timestamp 1624857261
transform 1 0 196792 0 1 82557
box 0 0 1 1
use contact_32  contact_32_421
timestamp 1624857261
transform 1 0 196792 0 1 115741
box 0 0 1 1
use contact_32  contact_32_420
timestamp 1624857261
transform 1 0 196792 0 1 116013
box 0 0 1 1
use contact_32  contact_32_419
timestamp 1624857261
transform 1 0 196656 0 1 98605
box 0 0 1 1
use contact_32  contact_32_418
timestamp 1624857261
transform 1 0 196656 0 1 98333
box 0 0 1 1
use contact_32  contact_32_417
timestamp 1624857261
transform 1 0 196656 0 1 119277
box 0 0 1 1
use contact_32  contact_32_416
timestamp 1624857261
transform 1 0 196656 0 1 119549
box 0 0 1 1
use contact_32  contact_32_415
timestamp 1624857261
transform 1 0 196792 0 1 50189
box 0 0 1 1
use contact_32  contact_32_414
timestamp 1624857261
transform 1 0 196792 0 1 50461
box 0 0 1 1
use contact_32  contact_32_413
timestamp 1624857261
transform 1 0 196792 0 1 50053
box 0 0 1 1
use contact_32  contact_32_412
timestamp 1624857261
transform 1 0 196792 0 1 49781
box 0 0 1 1
use contact_32  contact_32_411
timestamp 1624857261
transform 1 0 196656 0 1 96293
box 0 0 1 1
use contact_32  contact_32_410
timestamp 1624857261
transform 1 0 196656 0 1 96021
box 0 0 1 1
use contact_32  contact_32_409
timestamp 1624857261
transform 1 0 196656 0 1 96429
box 0 0 1 1
use contact_32  contact_32_408
timestamp 1624857261
transform 1 0 196656 0 1 96701
box 0 0 1 1
use contact_32  contact_32_407
timestamp 1624857261
transform 1 0 196792 0 1 103501
box 0 0 1 1
use contact_32  contact_32_406
timestamp 1624857261
transform 1 0 196792 0 1 103773
box 0 0 1 1
use contact_32  contact_32_405
timestamp 1624857261
transform 1 0 196792 0 1 103365
box 0 0 1 1
use contact_32  contact_32_404
timestamp 1624857261
transform 1 0 196792 0 1 103093
box 0 0 1 1
use contact_32  contact_32_403
timestamp 1624857261
transform 1 0 196656 0 1 101869
box 0 0 1 1
use contact_32  contact_32_402
timestamp 1624857261
transform 1 0 196656 0 1 102141
box 0 0 1 1
use contact_32  contact_32_401
timestamp 1624857261
transform 1 0 196792 0 1 66645
box 0 0 1 1
use contact_32  contact_32_400
timestamp 1624857261
transform 1 0 196792 0 1 66373
box 0 0 1 1
use contact_32  contact_32_399
timestamp 1624857261
transform 1 0 196792 0 1 66781
box 0 0 1 1
use contact_32  contact_32_398
timestamp 1624857261
transform 1 0 196792 0 1 67053
box 0 0 1 1
use contact_32  contact_32_397
timestamp 1624857261
transform 1 0 196792 0 1 74261
box 0 0 1 1
use contact_32  contact_32_396
timestamp 1624857261
transform 1 0 196792 0 1 74533
box 0 0 1 1
use contact_32  contact_32_395
timestamp 1624857261
transform 1 0 196792 0 1 48149
box 0 0 1 1
use contact_32  contact_32_394
timestamp 1624857261
transform 1 0 196792 0 1 48421
box 0 0 1 1
use contact_32  contact_32_393
timestamp 1624857261
transform 1 0 196656 0 1 105133
box 0 0 1 1
use contact_32  contact_32_392
timestamp 1624857261
transform 1 0 196656 0 1 105405
box 0 0 1 1
use contact_32  contact_32_391
timestamp 1624857261
transform 1 0 196656 0 1 64741
box 0 0 1 1
use contact_32  contact_32_390
timestamp 1624857261
transform 1 0 196656 0 1 65013
box 0 0 1 1
use contact_32  contact_32_389
timestamp 1624857261
transform 1 0 196656 0 1 55357
box 0 0 1 1
use contact_32  contact_32_388
timestamp 1624857261
transform 1 0 196656 0 1 55629
box 0 0 1 1
use contact_32  contact_32_387
timestamp 1624857261
transform 1 0 196656 0 1 55221
box 0 0 1 1
use contact_32  contact_32_386
timestamp 1624857261
transform 1 0 196656 0 1 54949
box 0 0 1 1
use contact_32  contact_32_385
timestamp 1624857261
transform 1 0 196792 0 1 70725
box 0 0 1 1
use contact_32  contact_32_384
timestamp 1624857261
transform 1 0 196792 0 1 70997
box 0 0 1 1
use contact_32  contact_32_383
timestamp 1624857261
transform 1 0 196656 0 1 42981
box 0 0 1 1
use contact_32  contact_32_382
timestamp 1624857261
transform 1 0 196656 0 1 42709
box 0 0 1 1
use contact_32  contact_32_381
timestamp 1624857261
transform 1 0 196656 0 1 117237
box 0 0 1 1
use contact_32  contact_32_380
timestamp 1624857261
transform 1 0 196656 0 1 116965
box 0 0 1 1
use contact_32  contact_32_379
timestamp 1624857261
transform 1 0 196656 0 1 58349
box 0 0 1 1
use contact_32  contact_32_378
timestamp 1624857261
transform 1 0 196656 0 1 58077
box 0 0 1 1
use contact_32  contact_32_377
timestamp 1624857261
transform 1 0 196792 0 1 38221
box 0 0 1 1
use contact_32  contact_32_376
timestamp 1624857261
transform 1 0 196792 0 1 37949
box 0 0 1 1
use contact_32  contact_32_375
timestamp 1624857261
transform 1 0 196792 0 1 79701
box 0 0 1 1
use contact_32  contact_32_374
timestamp 1624857261
transform 1 0 196792 0 1 79429
box 0 0 1 1
use contact_32  contact_32_373
timestamp 1624857261
transform 1 0 196792 0 1 79837
box 0 0 1 1
use contact_32  contact_32_372
timestamp 1624857261
transform 1 0 196792 0 1 80109
box 0 0 1 1
use contact_32  contact_32_371
timestamp 1624857261
transform 1 0 196792 0 1 76165
box 0 0 1 1
use contact_32  contact_32_370
timestamp 1624857261
transform 1 0 196792 0 1 75893
box 0 0 1 1
use contact_32  contact_32_369
timestamp 1624857261
transform 1 0 196656 0 1 65965
box 0 0 1 1
use contact_32  contact_32_368
timestamp 1624857261
transform 1 0 196656 0 1 66237
box 0 0 1 1
use contact_32  contact_32_367
timestamp 1624857261
transform 1 0 196656 0 1 65829
box 0 0 1 1
use contact_32  contact_32_366
timestamp 1624857261
transform 1 0 196656 0 1 65557
box 0 0 1 1
use contact_32  contact_32_365
timestamp 1624857261
transform 1 0 196656 0 1 50597
box 0 0 1 1
use contact_32  contact_32_364
timestamp 1624857261
transform 1 0 196656 0 1 50869
box 0 0 1 1
use contact_32  contact_32_363
timestamp 1624857261
transform 1 0 196656 0 1 124853
box 0 0 1 1
use contact_32  contact_32_362
timestamp 1624857261
transform 1 0 196656 0 1 125125
box 0 0 1 1
use contact_32  contact_32_361
timestamp 1624857261
transform 1 0 196656 0 1 124717
box 0 0 1 1
use contact_32  contact_32_360
timestamp 1624857261
transform 1 0 196656 0 1 124445
box 0 0 1 1
use contact_32  contact_32_359
timestamp 1624857261
transform 1 0 196656 0 1 49645
box 0 0 1 1
use contact_32  contact_32_358
timestamp 1624857261
transform 1 0 196656 0 1 49373
box 0 0 1 1
use contact_32  contact_32_357
timestamp 1624857261
transform 1 0 196792 0 1 101461
box 0 0 1 1
use contact_32  contact_32_356
timestamp 1624857261
transform 1 0 196792 0 1 101189
box 0 0 1 1
use contact_32  contact_32_355
timestamp 1624857261
transform 1 0 196792 0 1 63517
box 0 0 1 1
use contact_32  contact_32_354
timestamp 1624857261
transform 1 0 196792 0 1 63245
box 0 0 1 1
use contact_32  contact_32_353
timestamp 1624857261
transform 1 0 196656 0 1 37813
box 0 0 1 1
use contact_32  contact_32_352
timestamp 1624857261
transform 1 0 196656 0 1 37541
box 0 0 1 1
use contact_32  contact_32_351
timestamp 1624857261
transform 1 0 196792 0 1 121997
box 0 0 1 1
use contact_32  contact_32_350
timestamp 1624857261
transform 1 0 196792 0 1 121725
box 0 0 1 1
use contact_32  contact_32_349
timestamp 1624857261
transform 1 0 196656 0 1 82421
box 0 0 1 1
use contact_32  contact_32_348
timestamp 1624857261
transform 1 0 196656 0 1 82149
box 0 0 1 1
use contact_32  contact_32_347
timestamp 1624857261
transform 1 0 196656 0 1 61885
box 0 0 1 1
use contact_32  contact_32_346
timestamp 1624857261
transform 1 0 196656 0 1 61613
box 0 0 1 1
use contact_32  contact_32_345
timestamp 1624857261
transform 1 0 196792 0 1 36317
box 0 0 1 1
use contact_32  contact_32_344
timestamp 1624857261
transform 1 0 196792 0 1 36589
box 0 0 1 1
use contact_32  contact_32_343
timestamp 1624857261
transform 1 0 196792 0 1 90445
box 0 0 1 1
use contact_32  contact_32_342
timestamp 1624857261
transform 1 0 196792 0 1 90717
box 0 0 1 1
use contact_32  contact_32_341
timestamp 1624857261
transform 1 0 196792 0 1 90309
box 0 0 1 1
use contact_32  contact_32_340
timestamp 1624857261
transform 1 0 196792 0 1 90037
box 0 0 1 1
use contact_32  contact_32_339
timestamp 1624857261
transform 1 0 196656 0 1 42301
box 0 0 1 1
use contact_32  contact_32_338
timestamp 1624857261
transform 1 0 196656 0 1 42573
box 0 0 1 1
use contact_32  contact_32_337
timestamp 1624857261
transform 1 0 196656 0 1 42165
box 0 0 1 1
use contact_32  contact_32_336
timestamp 1624857261
transform 1 0 196656 0 1 41893
box 0 0 1 1
use contact_32  contact_32_335
timestamp 1624857261
transform 1 0 196656 0 1 108261
box 0 0 1 1
use contact_32  contact_32_334
timestamp 1624857261
transform 1 0 196656 0 1 108533
box 0 0 1 1
use contact_32  contact_32_333
timestamp 1624857261
transform 1 0 196792 0 1 54541
box 0 0 1 1
use contact_32  contact_32_332
timestamp 1624857261
transform 1 0 196792 0 1 54813
box 0 0 1 1
use contact_32  contact_32_331
timestamp 1624857261
transform 1 0 196792 0 1 54405
box 0 0 1 1
use contact_32  contact_32_330
timestamp 1624857261
transform 1 0 196792 0 1 54133
box 0 0 1 1
use contact_32  contact_32_329
timestamp 1624857261
transform 1 0 196656 0 1 59301
box 0 0 1 1
use contact_32  contact_32_328
timestamp 1624857261
transform 1 0 196656 0 1 59573
box 0 0 1 1
use contact_32  contact_32_327
timestamp 1624857261
transform 1 0 196656 0 1 111661
box 0 0 1 1
use contact_32  contact_32_326
timestamp 1624857261
transform 1 0 196656 0 1 111389
box 0 0 1 1
use contact_32  contact_32_325
timestamp 1624857261
transform 1 0 196656 0 1 111797
box 0 0 1 1
use contact_32  contact_32_324
timestamp 1624857261
transform 1 0 196656 0 1 112069
box 0 0 1 1
use contact_32  contact_32_323
timestamp 1624857261
transform 1 0 196792 0 1 84869
box 0 0 1 1
use contact_32  contact_32_322
timestamp 1624857261
transform 1 0 196792 0 1 84597
box 0 0 1 1
use contact_32  contact_32_321
timestamp 1624857261
transform 1 0 196656 0 1 57533
box 0 0 1 1
use contact_32  contact_32_320
timestamp 1624857261
transform 1 0 196656 0 1 57261
box 0 0 1 1
use contact_32  contact_32_319
timestamp 1624857261
transform 1 0 196792 0 1 57669
box 0 0 1 1
use contact_32  contact_32_318
timestamp 1624857261
transform 1 0 196792 0 1 57941
box 0 0 1 1
use contact_32  contact_32_317
timestamp 1624857261
transform 1 0 196656 0 1 74941
box 0 0 1 1
use contact_32  contact_32_316
timestamp 1624857261
transform 1 0 196656 0 1 74669
box 0 0 1 1
use contact_32  contact_32_315
timestamp 1624857261
transform 1 0 196792 0 1 75077
box 0 0 1 1
use contact_32  contact_32_314
timestamp 1624857261
transform 1 0 196792 0 1 75349
box 0 0 1 1
use contact_32  contact_32_313
timestamp 1624857261
transform 1 0 196792 0 1 123221
box 0 0 1 1
use contact_32  contact_32_312
timestamp 1624857261
transform 1 0 196792 0 1 123493
box 0 0 1 1
use contact_32  contact_32_311
timestamp 1624857261
transform 1 0 196792 0 1 95885
box 0 0 1 1
use contact_32  contact_32_310
timestamp 1624857261
transform 1 0 196792 0 1 95613
box 0 0 1 1
use contact_32  contact_32_309
timestamp 1624857261
transform 1 0 196656 0 1 44477
box 0 0 1 1
use contact_32  contact_32_308
timestamp 1624857261
transform 1 0 196656 0 1 44205
box 0 0 1 1
use contact_32  contact_32_307
timestamp 1624857261
transform 1 0 196792 0 1 100237
box 0 0 1 1
use contact_32  contact_32_306
timestamp 1624857261
transform 1 0 196792 0 1 99965
box 0 0 1 1
use contact_32  contact_32_305
timestamp 1624857261
transform 1 0 196792 0 1 88133
box 0 0 1 1
use contact_32  contact_32_304
timestamp 1624857261
transform 1 0 196792 0 1 88405
box 0 0 1 1
use contact_32  contact_32_303
timestamp 1624857261
transform 1 0 196656 0 1 61477
box 0 0 1 1
use contact_32  contact_32_302
timestamp 1624857261
transform 1 0 196656 0 1 61205
box 0 0 1 1
use contact_32  contact_32_301
timestamp 1624857261
transform 1 0 196792 0 1 97925
box 0 0 1 1
use contact_32  contact_32_300
timestamp 1624857261
transform 1 0 196792 0 1 98197
box 0 0 1 1
use contact_32  contact_32_299
timestamp 1624857261
transform 1 0 196656 0 1 88813
box 0 0 1 1
use contact_32  contact_32_298
timestamp 1624857261
transform 1 0 196656 0 1 88541
box 0 0 1 1
use contact_32  contact_32_297
timestamp 1624857261
transform 1 0 196656 0 1 81333
box 0 0 1 1
use contact_32  contact_32_296
timestamp 1624857261
transform 1 0 196656 0 1 81605
box 0 0 1 1
use contact_32  contact_32_295
timestamp 1624857261
transform 1 0 196656 0 1 29245
box 0 0 1 1
use contact_32  contact_32_294
timestamp 1624857261
transform 1 0 196656 0 1 29517
box 0 0 1 1
use contact_32  contact_32_293
timestamp 1624857261
transform 1 0 196656 0 1 29109
box 0 0 1 1
use contact_32  contact_32_292
timestamp 1624857261
transform 1 0 196656 0 1 28837
box 0 0 1 1
use contact_32  contact_32_291
timestamp 1624857261
transform 1 0 196792 0 1 27205
box 0 0 1 1
use contact_32  contact_32_290
timestamp 1624857261
transform 1 0 196792 0 1 26933
box 0 0 1 1
use contact_32  contact_32_289
timestamp 1624857261
transform 1 0 196656 0 1 67189
box 0 0 1 1
use contact_32  contact_32_288
timestamp 1624857261
transform 1 0 196656 0 1 67461
box 0 0 1 1
use contact_32  contact_32_287
timestamp 1624857261
transform 1 0 196792 0 1 64061
box 0 0 1 1
use contact_32  contact_32_286
timestamp 1624857261
transform 1 0 196792 0 1 64333
box 0 0 1 1
use contact_32  contact_32_285
timestamp 1624857261
transform 1 0 196792 0 1 29653
box 0 0 1 1
use contact_32  contact_32_284
timestamp 1624857261
transform 1 0 196792 0 1 29925
box 0 0 1 1
use contact_32  contact_32_283
timestamp 1624857261
transform 1 0 199104 0 1 29653
box 0 0 1 1
use contact_32  contact_32_282
timestamp 1624857261
transform 1 0 199104 0 1 29925
box 0 0 1 1
use contact_32  contact_32_281
timestamp 1624857261
transform 1 0 196656 0 1 94253
box 0 0 1 1
use contact_32  contact_32_280
timestamp 1624857261
transform 1 0 196656 0 1 93981
box 0 0 1 1
use contact_32  contact_32_279
timestamp 1624857261
transform 1 0 196656 0 1 94389
box 0 0 1 1
use contact_32  contact_32_278
timestamp 1624857261
transform 1 0 196656 0 1 94661
box 0 0 1 1
use contact_32  contact_32_277
timestamp 1624857261
transform 1 0 196792 0 1 56853
box 0 0 1 1
use contact_32  contact_32_276
timestamp 1624857261
transform 1 0 196792 0 1 57125
box 0 0 1 1
use contact_32  contact_32_275
timestamp 1624857261
transform 1 0 196656 0 1 51005
box 0 0 1 1
use contact_32  contact_32_274
timestamp 1624857261
transform 1 0 196656 0 1 51277
box 0 0 1 1
use contact_32  contact_32_273
timestamp 1624857261
transform 1 0 196656 0 1 77797
box 0 0 1 1
use contact_32  contact_32_272
timestamp 1624857261
transform 1 0 196656 0 1 78069
box 0 0 1 1
use contact_32  contact_32_271
timestamp 1624857261
transform 1 0 196656 0 1 51685
box 0 0 1 1
use contact_32  contact_32_270
timestamp 1624857261
transform 1 0 196656 0 1 51413
box 0 0 1 1
use contact_32  contact_32_269
timestamp 1624857261
transform 1 0 196656 0 1 79293
box 0 0 1 1
use contact_32  contact_32_268
timestamp 1624857261
transform 1 0 196656 0 1 79021
box 0 0 1 1
use contact_32  contact_32_267
timestamp 1624857261
transform 1 0 196656 0 1 25573
box 0 0 1 1
use contact_32  contact_32_266
timestamp 1624857261
transform 1 0 196656 0 1 25301
box 0 0 1 1
use contact_32  contact_32_265
timestamp 1624857261
transform 1 0 196656 0 1 25709
box 0 0 1 1
use contact_32  contact_32_264
timestamp 1624857261
transform 1 0 196656 0 1 25981
box 0 0 1 1
use contact_32  contact_32_263
timestamp 1624857261
transform 1 0 196792 0 1 53589
box 0 0 1 1
use contact_32  contact_32_262
timestamp 1624857261
transform 1 0 196792 0 1 53317
box 0 0 1 1
use contact_32  contact_32_261
timestamp 1624857261
transform 1 0 196792 0 1 53725
box 0 0 1 1
use contact_32  contact_32_260
timestamp 1624857261
transform 1 0 196792 0 1 53997
box 0 0 1 1
use contact_32  contact_32_259
timestamp 1624857261
transform 1 0 196656 0 1 118053
box 0 0 1 1
use contact_32  contact_32_258
timestamp 1624857261
transform 1 0 196656 0 1 117781
box 0 0 1 1
use contact_32  contact_32_257
timestamp 1624857261
transform 1 0 196792 0 1 102685
box 0 0 1 1
use contact_32  contact_32_256
timestamp 1624857261
transform 1 0 196792 0 1 102957
box 0 0 1 1
use contact_32  contact_32_255
timestamp 1624857261
transform 1 0 196792 0 1 92757
box 0 0 1 1
use contact_32  contact_32_254
timestamp 1624857261
transform 1 0 196792 0 1 92485
box 0 0 1 1
use contact_32  contact_32_253
timestamp 1624857261
transform 1 0 196656 0 1 71405
box 0 0 1 1
use contact_32  contact_32_252
timestamp 1624857261
transform 1 0 196656 0 1 71133
box 0 0 1 1
use contact_32  contact_32_251
timestamp 1624857261
transform 1 0 196792 0 1 125261
box 0 0 1 1
use contact_32  contact_32_250
timestamp 1624857261
transform 1 0 196792 0 1 125533
box 0 0 1 1
use contact_32  contact_32_249
timestamp 1624857261
transform 1 0 196656 0 1 30061
box 0 0 1 1
use contact_32  contact_32_248
timestamp 1624857261
transform 1 0 196656 0 1 30333
box 0 0 1 1
use contact_32  contact_32_247
timestamp 1624857261
transform 1 0 196792 0 1 26389
box 0 0 1 1
use contact_32  contact_32_246
timestamp 1624857261
transform 1 0 196792 0 1 26117
box 0 0 1 1
use contact_32  contact_32_245
timestamp 1624857261
transform 1 0 196792 0 1 49237
box 0 0 1 1
use contact_32  contact_32_244
timestamp 1624857261
transform 1 0 196792 0 1 48965
box 0 0 1 1
use contact_32  contact_32_243
timestamp 1624857261
transform 1 0 196656 0 1 62837
box 0 0 1 1
use contact_32  contact_32_242
timestamp 1624857261
transform 1 0 196656 0 1 63109
box 0 0 1 1
use contact_32  contact_32_241
timestamp 1624857261
transform 1 0 196656 0 1 33597
box 0 0 1 1
use contact_32  contact_32_240
timestamp 1624857261
transform 1 0 196656 0 1 33869
box 0 0 1 1
use contact_32  contact_32_239
timestamp 1624857261
transform 1 0 196656 0 1 33461
box 0 0 1 1
use contact_32  contact_32_238
timestamp 1624857261
transform 1 0 196656 0 1 33189
box 0 0 1 1
use contact_32  contact_32_237
timestamp 1624857261
transform 1 0 196656 0 1 120501
box 0 0 1 1
use contact_32  contact_32_236
timestamp 1624857261
transform 1 0 196656 0 1 120773
box 0 0 1 1
use contact_32  contact_32_235
timestamp 1624857261
transform 1 0 196656 0 1 75757
box 0 0 1 1
use contact_32  contact_32_234
timestamp 1624857261
transform 1 0 196656 0 1 75485
box 0 0 1 1
use contact_32  contact_32_233
timestamp 1624857261
transform 1 0 196656 0 1 47469
box 0 0 1 1
use contact_32  contact_32_232
timestamp 1624857261
transform 1 0 196656 0 1 47741
box 0 0 1 1
use contact_32  contact_32_231
timestamp 1624857261
transform 1 0 196656 0 1 60797
box 0 0 1 1
use contact_32  contact_32_230
timestamp 1624857261
transform 1 0 196656 0 1 61069
box 0 0 1 1
use contact_32  contact_32_229
timestamp 1624857261
transform 1 0 196792 0 1 68957
box 0 0 1 1
use contact_32  contact_32_228
timestamp 1624857261
transform 1 0 196792 0 1 68685
box 0 0 1 1
use contact_32  contact_32_227
timestamp 1624857261
transform 1 0 196792 0 1 78613
box 0 0 1 1
use contact_32  contact_32_226
timestamp 1624857261
transform 1 0 196792 0 1 78885
box 0 0 1 1
use contact_32  contact_32_225
timestamp 1624857261
transform 1 0 196792 0 1 78477
box 0 0 1 1
use contact_32  contact_32_224
timestamp 1624857261
transform 1 0 196792 0 1 78205
box 0 0 1 1
use contact_32  contact_32_223
timestamp 1624857261
transform 1 0 196792 0 1 67597
box 0 0 1 1
use contact_32  contact_32_222
timestamp 1624857261
transform 1 0 196792 0 1 67869
box 0 0 1 1
use contact_32  contact_32_221
timestamp 1624857261
transform 1 0 196792 0 1 116421
box 0 0 1 1
use contact_32  contact_32_220
timestamp 1624857261
transform 1 0 196792 0 1 116149
box 0 0 1 1
use contact_32  contact_32_219
timestamp 1624857261
transform 1 0 196792 0 1 116557
box 0 0 1 1
use contact_32  contact_32_218
timestamp 1624857261
transform 1 0 196792 0 1 116829
box 0 0 1 1
use contact_32  contact_32_217
timestamp 1624857261
transform 1 0 196792 0 1 81741
box 0 0 1 1
use contact_32  contact_32_216
timestamp 1624857261
transform 1 0 196792 0 1 82013
box 0 0 1 1
use contact_32  contact_32_215
timestamp 1624857261
transform 1 0 196656 0 1 68005
box 0 0 1 1
use contact_32  contact_32_214
timestamp 1624857261
transform 1 0 196656 0 1 68277
box 0 0 1 1
use contact_32  contact_32_213
timestamp 1624857261
transform 1 0 196792 0 1 91669
box 0 0 1 1
use contact_32  contact_32_212
timestamp 1624857261
transform 1 0 196792 0 1 91941
box 0 0 1 1
use contact_32  contact_32_211
timestamp 1624857261
transform 1 0 196656 0 1 92349
box 0 0 1 1
use contact_32  contact_32_210
timestamp 1624857261
transform 1 0 196656 0 1 92077
box 0 0 1 1
use contact_32  contact_32_209
timestamp 1624857261
transform 1 0 196928 0 1 142397
box 0 0 1 1
use contact_32  contact_32_208
timestamp 1624857261
transform 1 0 196928 0 1 142805
box 0 0 1 1
use contact_32  contact_32_207
timestamp 1624857261
transform 1 0 196928 0 1 1773
box 0 0 1 1
use contact_32  contact_32_206
timestamp 1624857261
transform 1 0 196928 0 1 1229
box 0 0 1 1
use contact_32  contact_32_205
timestamp 1624857261
transform 1 0 197880 0 1 128525
box 0 0 1 1
use contact_32  contact_32_204
timestamp 1624857261
transform 1 0 197880 0 1 131245
box 0 0 1 1
use contact_32  contact_32_203
timestamp 1624857261
transform 1 0 197880 0 1 139677
box 0 0 1 1
use contact_32  contact_32_202
timestamp 1624857261
transform 1 0 197880 0 1 137093
box 0 0 1 1
use contact_32  contact_32_201
timestamp 1624857261
transform 1 0 198288 0 1 139813
box 0 0 1 1
use contact_32  contact_32_200
timestamp 1624857261
transform 1 0 198288 0 1 141853
box 0 0 1 1
use contact_32  contact_32_199
timestamp 1624857261
transform 1 0 197880 0 1 134237
box 0 0 1 1
use contact_32  contact_32_198
timestamp 1624857261
transform 1 0 197880 0 1 136821
box 0 0 1 1
use contact_32  contact_32_197
timestamp 1624857261
transform 1 0 203456 0 1 131381
box 0 0 1 1
use contact_32  contact_32_196
timestamp 1624857261
transform 1 0 203456 0 1 132469
box 0 0 1 1
use contact_32  contact_32_195
timestamp 1624857261
transform 1 0 199240 0 1 142261
box 0 0 1 1
use contact_32  contact_32_194
timestamp 1624857261
transform 1 0 199240 0 1 141989
box 0 0 1 1
use contact_32  contact_32_193
timestamp 1624857261
transform 1 0 198832 0 1 142397
box 0 0 1 1
use contact_32  contact_32_192
timestamp 1624857261
transform 1 0 198832 0 1 142805
box 0 0 1 1
use contact_32  contact_32_191
timestamp 1624857261
transform 1 0 198696 0 1 1773
box 0 0 1 1
use contact_32  contact_32_190
timestamp 1624857261
transform 1 0 198696 0 1 1229
box 0 0 1 1
use contact_32  contact_32_189
timestamp 1624857261
transform 1 0 199240 0 1 32237
box 0 0 1 1
use contact_32  contact_32_188
timestamp 1624857261
transform 1 0 199240 0 1 31557
box 0 0 1 1
use contact_32  contact_32_187
timestamp 1624857261
transform 1 0 199104 0 1 32373
box 0 0 1 1
use contact_32  contact_32_186
timestamp 1624857261
transform 1 0 199104 0 1 33053
box 0 0 1 1
use contact_32  contact_32_185
timestamp 1624857261
transform 1 0 199376 0 1 28293
box 0 0 1 1
use contact_32  contact_32_184
timestamp 1624857261
transform 1 0 199376 0 1 27613
box 0 0 1 1
use contact_32  contact_32_183
timestamp 1624857261
transform 1 0 199240 0 1 28429
box 0 0 1 1
use contact_32  contact_32_182
timestamp 1624857261
transform 1 0 199240 0 1 29109
box 0 0 1 1
use contact_32  contact_32_181
timestamp 1624857261
transform 1 0 199104 0 1 33869
box 0 0 1 1
use contact_32  contact_32_180
timestamp 1624857261
transform 1 0 199104 0 1 33189
box 0 0 1 1
use contact_32  contact_32_179
timestamp 1624857261
transform 1 0 199104 0 1 31421
box 0 0 1 1
use contact_32  contact_32_178
timestamp 1624857261
transform 1 0 199104 0 1 30061
box 0 0 1 1
use contact_32  contact_32_177
timestamp 1624857261
transform 1 0 199376 0 1 25301
box 0 0 1 1
use contact_32  contact_32_176
timestamp 1624857261
transform 1 0 199376 0 1 25845
box 0 0 1 1
use contact_32  contact_32_175
timestamp 1624857261
transform 1 0 199376 0 1 25165
box 0 0 1 1
use contact_32  contact_32_174
timestamp 1624857261
transform 1 0 199376 0 1 24893
box 0 0 1 1
use contact_32  contact_32_173
timestamp 1624857261
transform 1 0 199920 0 1 24893
box 0 0 1 1
use contact_32  contact_32_172
timestamp 1624857261
transform 1 0 199920 0 1 25165
box 0 0 1 1
use contact_32  contact_32_171
timestamp 1624857261
transform 1 0 199376 0 1 29925
box 0 0 1 1
use contact_32  contact_32_170
timestamp 1624857261
transform 1 0 199376 0 1 29245
box 0 0 1 1
use contact_32  contact_32_169
timestamp 1624857261
transform 1 0 200192 0 1 25301
box 0 0 1 1
use contact_32  contact_32_168
timestamp 1624857261
transform 1 0 200192 0 1 25981
box 0 0 1 1
use contact_32  contact_32_167
timestamp 1624857261
transform 1 0 200464 0 1 26117
box 0 0 1 1
use contact_32  contact_32_166
timestamp 1624857261
transform 1 0 200464 0 1 27477
box 0 0 1 1
use contact_32  contact_32_165
timestamp 1624857261
transform 1 0 201280 0 1 25981
box 0 0 1 1
use contact_32  contact_32_164
timestamp 1624857261
transform 1 0 201280 0 1 25301
box 0 0 1 1
use contact_32  contact_32_163
timestamp 1624857261
transform 1 0 200192 0 1 1773
box 0 0 1 1
use contact_32  contact_32_162
timestamp 1624857261
transform 1 0 200192 0 1 1229
box 0 0 1 1
use contact_32  contact_32_161
timestamp 1624857261
transform 1 0 200464 0 1 142261
box 0 0 1 1
use contact_32  contact_32_160
timestamp 1624857261
transform 1 0 200464 0 1 141989
box 0 0 1 1
use contact_32  contact_32_159
timestamp 1624857261
transform 1 0 200192 0 1 142397
box 0 0 1 1
use contact_32  contact_32_158
timestamp 1624857261
transform 1 0 200192 0 1 142805
box 0 0 1 1
use contact_32  contact_32_157
timestamp 1624857261
transform 1 0 200464 0 1 33869
box 0 0 1 1
use contact_32  contact_32_156
timestamp 1624857261
transform 1 0 200464 0 1 33189
box 0 0 1 1
use contact_32  contact_32_155
timestamp 1624857261
transform 1 0 200464 0 1 31557
box 0 0 1 1
use contact_32  contact_32_154
timestamp 1624857261
transform 1 0 200464 0 1 32237
box 0 0 1 1
use contact_32  contact_32_153
timestamp 1624857261
transform 1 0 200464 0 1 33053
box 0 0 1 1
use contact_32  contact_32_152
timestamp 1624857261
transform 1 0 200464 0 1 32373
box 0 0 1 1
use contact_32  contact_32_151
timestamp 1624857261
transform 1 0 200600 0 1 29925
box 0 0 1 1
use contact_32  contact_32_150
timestamp 1624857261
transform 1 0 200600 0 1 29245
box 0 0 1 1
use contact_32  contact_32_149
timestamp 1624857261
transform 1 0 201824 0 1 32237
box 0 0 1 1
use contact_32  contact_32_148
timestamp 1624857261
transform 1 0 201824 0 1 31557
box 0 0 1 1
use contact_32  contact_32_147
timestamp 1624857261
transform 1 0 200464 0 1 27613
box 0 0 1 1
use contact_32  contact_32_146
timestamp 1624857261
transform 1 0 200464 0 1 28293
box 0 0 1 1
use contact_32  contact_32_145
timestamp 1624857261
transform 1 0 200464 0 1 28429
box 0 0 1 1
use contact_32  contact_32_144
timestamp 1624857261
transform 1 0 200464 0 1 29109
box 0 0 1 1
use contact_32  contact_32_143
timestamp 1624857261
transform 1 0 204000 0 1 25165
box 0 0 1 1
use contact_32  contact_32_142
timestamp 1624857261
transform 1 0 204000 0 1 24893
box 0 0 1 1
use contact_32  contact_32_141
timestamp 1624857261
transform 1 0 201960 0 1 142397
box 0 0 1 1
use contact_32  contact_32_140
timestamp 1624857261
transform 1 0 201960 0 1 142805
box 0 0 1 1
use contact_32  contact_32_139
timestamp 1624857261
transform 1 0 201960 0 1 1773
box 0 0 1 1
use contact_32  contact_32_138
timestamp 1624857261
transform 1 0 201960 0 1 1229
box 0 0 1 1
use contact_32  contact_32_137
timestamp 1624857261
transform 1 0 203320 0 1 132469
box 0 0 1 1
use contact_32  contact_32_136
timestamp 1624857261
transform 1 0 203320 0 1 129749
box 0 0 1 1
use contact_32  contact_32_135
timestamp 1624857261
transform 1 0 203320 0 1 132605
box 0 0 1 1
use contact_32  contact_32_134
timestamp 1624857261
transform 1 0 203320 0 1 135189
box 0 0 1 1
use contact_32  contact_32_133
timestamp 1624857261
transform 1 0 203456 0 1 129613
box 0 0 1 1
use contact_32  contact_32_132
timestamp 1624857261
transform 1 0 203456 0 1 126893
box 0 0 1 1
use contact_32  contact_32_131
timestamp 1624857261
transform 1 0 203592 0 1 142397
box 0 0 1 1
use contact_32  contact_32_130
timestamp 1624857261
transform 1 0 203592 0 1 142805
box 0 0 1 1
use contact_32  contact_32_129
timestamp 1624857261
transform 1 0 203592 0 1 1773
box 0 0 1 1
use contact_32  contact_32_128
timestamp 1624857261
transform 1 0 203592 0 1 1229
box 0 0 1 1
use contact_32  contact_32_127
timestamp 1624857261
transform 1 0 204136 0 1 19181
box 0 0 1 1
use contact_32  contact_32_126
timestamp 1624857261
transform 1 0 204136 0 1 21901
box 0 0 1 1
use contact_32  contact_32_125
timestamp 1624857261
transform 1 0 204272 0 1 19045
box 0 0 1 1
use contact_32  contact_32_124
timestamp 1624857261
transform 1 0 204272 0 1 16461
box 0 0 1 1
use contact_32  contact_32_123
timestamp 1624857261
transform 1 0 204000 0 1 13605
box 0 0 1 1
use contact_32  contact_32_122
timestamp 1624857261
transform 1 0 204000 0 1 16189
box 0 0 1 1
use contact_32  contact_32_121
timestamp 1624857261
transform 1 0 204136 0 1 22037
box 0 0 1 1
use contact_32  contact_32_120
timestamp 1624857261
transform 1 0 204136 0 1 24757
box 0 0 1 1
use contact_32  contact_32_119
timestamp 1624857261
transform 1 0 205224 0 1 142397
box 0 0 1 1
use contact_32  contact_32_118
timestamp 1624857261
transform 1 0 205224 0 1 142805
box 0 0 1 1
use contact_32  contact_32_117
timestamp 1624857261
transform 1 0 205224 0 1 1773
box 0 0 1 1
use contact_32  contact_32_116
timestamp 1624857261
transform 1 0 205224 0 1 1229
box 0 0 1 1
use contact_32  contact_32_115
timestamp 1624857261
transform 1 0 207128 0 1 1773
box 0 0 1 1
use contact_32  contact_32_114
timestamp 1624857261
transform 1 0 207128 0 1 1229
box 0 0 1 1
use contact_32  contact_32_113
timestamp 1624857261
transform 1 0 206856 0 1 142397
box 0 0 1 1
use contact_32  contact_32_112
timestamp 1624857261
transform 1 0 206856 0 1 142805
box 0 0 1 1
use contact_32  contact_32_111
timestamp 1624857261
transform 1 0 208624 0 1 1773
box 0 0 1 1
use contact_32  contact_32_110
timestamp 1624857261
transform 1 0 208624 0 1 1229
box 0 0 1 1
use contact_32  contact_32_109
timestamp 1624857261
transform 1 0 208624 0 1 142397
box 0 0 1 1
use contact_32  contact_32_108
timestamp 1624857261
transform 1 0 208624 0 1 142805
box 0 0 1 1
use contact_32  contact_32_107
timestamp 1624857261
transform 1 0 210392 0 1 1773
box 0 0 1 1
use contact_32  contact_32_106
timestamp 1624857261
transform 1 0 210392 0 1 1229
box 0 0 1 1
use contact_32  contact_32_105
timestamp 1624857261
transform 1 0 210392 0 1 142397
box 0 0 1 1
use contact_32  contact_32_104
timestamp 1624857261
transform 1 0 210392 0 1 142805
box 0 0 1 1
use contact_32  contact_32_103
timestamp 1624857261
transform 1 0 211888 0 1 1773
box 0 0 1 1
use contact_32  contact_32_102
timestamp 1624857261
transform 1 0 211888 0 1 1229
box 0 0 1 1
use contact_32  contact_32_101
timestamp 1624857261
transform 1 0 212024 0 1 142397
box 0 0 1 1
use contact_32  contact_32_100
timestamp 1624857261
transform 1 0 212024 0 1 142805
box 0 0 1 1
use contact_32  contact_32_99
timestamp 1624857261
transform 1 0 213656 0 1 1773
box 0 0 1 1
use contact_32  contact_32_98
timestamp 1624857261
transform 1 0 213656 0 1 1229
box 0 0 1 1
use contact_32  contact_32_97
timestamp 1624857261
transform 1 0 213656 0 1 142397
box 0 0 1 1
use contact_32  contact_32_96
timestamp 1624857261
transform 1 0 213656 0 1 142805
box 0 0 1 1
use contact_32  contact_32_95
timestamp 1624857261
transform 1 0 215424 0 1 1773
box 0 0 1 1
use contact_32  contact_32_94
timestamp 1624857261
transform 1 0 215424 0 1 1229
box 0 0 1 1
use contact_32  contact_32_93
timestamp 1624857261
transform 1 0 215424 0 1 142397
box 0 0 1 1
use contact_32  contact_32_92
timestamp 1624857261
transform 1 0 215424 0 1 142805
box 0 0 1 1
use contact_32  contact_32_91
timestamp 1624857261
transform 1 0 216784 0 1 116829
box 0 0 1 1
use contact_32  contact_32_90
timestamp 1624857261
transform 1 0 216784 0 1 116421
box 0 0 1 1
use contact_32  contact_32_89
timestamp 1624857261
transform 1 0 216784 0 1 125397
box 0 0 1 1
use contact_32  contact_32_88
timestamp 1624857261
transform 1 0 216784 0 1 124853
box 0 0 1 1
use contact_32  contact_32_87
timestamp 1624857261
transform 1 0 216784 0 1 122677
box 0 0 1 1
use contact_32  contact_32_86
timestamp 1624857261
transform 1 0 216784 0 1 123085
box 0 0 1 1
use contact_32  contact_32_85
timestamp 1624857261
transform 1 0 216784 0 1 135189
box 0 0 1 1
use contact_32  contact_32_84
timestamp 1624857261
transform 1 0 216784 0 1 134917
box 0 0 1 1
use contact_32  contact_32_83
timestamp 1624857261
transform 1 0 217464 0 1 108125
box 0 0 1 1
use contact_32  contact_32_82
timestamp 1624857261
transform 1 0 217464 0 1 69229
box 0 0 1 1
use contact_32  contact_32_81
timestamp 1624857261
transform 1 0 217464 0 1 119821
box 0 0 1 1
use contact_32  contact_32_80
timestamp 1624857261
transform 1 0 217464 0 1 77797
box 0 0 1 1
use contact_32  contact_32_79
timestamp 1624857261
transform 1 0 217464 0 1 101325
box 0 0 1 1
use contact_32  contact_32_78
timestamp 1624857261
transform 1 0 217464 0 1 45973
box 0 0 1 1
use contact_32  contact_32_77
timestamp 1624857261
transform 1 0 217464 0 1 12109
box 0 0 1 1
use contact_32  contact_32_76
timestamp 1624857261
transform 1 0 217464 0 1 129885
box 0 0 1 1
use contact_32  contact_32_75
timestamp 1624857261
transform 1 0 217464 0 1 50733
box 0 0 1 1
use contact_32  contact_32_74
timestamp 1624857261
transform 1 0 217464 0 1 102957
box 0 0 1 1
use contact_32  contact_32_73
timestamp 1624857261
transform 1 0 217464 0 1 126349
box 0 0 1 1
use contact_32  contact_32_72
timestamp 1624857261
transform 1 0 217464 0 1 49101
box 0 0 1 1
use contact_32  contact_32_71
timestamp 1624857261
transform 1 0 217464 0 1 27341
box 0 0 1 1
use contact_32  contact_32_70
timestamp 1624857261
transform 1 0 217464 0 1 10477
box 0 0 1 1
use contact_32  contact_32_69
timestamp 1624857261
transform 1 0 217464 0 1 59301
box 0 0 1 1
use contact_32  contact_32_68
timestamp 1624857261
transform 1 0 217464 0 1 72765
box 0 0 1 1
use contact_32  contact_32_67
timestamp 1624857261
transform 1 0 217464 0 1 5581
box 0 0 1 1
use contact_32  contact_32_66
timestamp 1624857261
transform 1 0 217464 0 1 28973
box 0 0 1 1
use contact_32  contact_32_65
timestamp 1624857261
transform 1 0 217464 0 1 97789
box 0 0 1 1
use contact_32  contact_32_64
timestamp 1624857261
transform 1 0 217464 0 1 131517
box 0 0 1 1
use contact_32  contact_32_63
timestamp 1624857261
transform 1 0 217464 0 1 47469
box 0 0 1 1
use contact_32  contact_32_62
timestamp 1624857261
transform 1 0 217464 0 1 54269
box 0 0 1 1
use contact_32  contact_32_61
timestamp 1624857261
transform 1 0 217464 0 1 94525
box 0 0 1 1
use contact_32  contact_32_60
timestamp 1624857261
transform 1 0 217464 0 1 2045
box 0 0 1 1
use contact_32  contact_32_59
timestamp 1624857261
transform 1 0 217464 0 1 82829
box 0 0 1 1
use contact_32  contact_32_58
timestamp 1624857261
transform 1 0 217464 0 1 81197
box 0 0 1 1
use contact_32  contact_32_57
timestamp 1624857261
transform 1 0 217464 0 1 141717
box 0 0 1 1
use contact_32  contact_32_56
timestamp 1624857261
transform 1 0 217464 0 1 136549
box 0 0 1 1
use contact_32  contact_32_55
timestamp 1624857261
transform 1 0 217464 0 1 109757
box 0 0 1 1
use contact_32  contact_32_54
timestamp 1624857261
transform 1 0 217464 0 1 84325
box 0 0 1 1
use contact_32  contact_32_53
timestamp 1624857261
transform 1 0 217464 0 1 22309
box 0 0 1 1
use contact_32  contact_32_52
timestamp 1624857261
transform 1 0 217464 0 1 86093
box 0 0 1 1
use contact_32  contact_32_51
timestamp 1624857261
transform 1 0 217464 0 1 74533
box 0 0 1 1
use contact_32  contact_32_50
timestamp 1624857261
transform 1 0 217464 0 1 65965
box 0 0 1 1
use contact_32  contact_32_49
timestamp 1624857261
transform 1 0 217464 0 1 106221
box 0 0 1 1
use contact_32  contact_32_48
timestamp 1624857261
transform 1 0 217464 0 1 42573
box 0 0 1 1
use contact_32  contact_32_47
timestamp 1624857261
transform 1 0 217464 0 1 138317
box 0 0 1 1
use contact_32  contact_32_46
timestamp 1624857261
transform 1 0 217464 0 1 17141
box 0 0 1 1
use contact_32  contact_32_45
timestamp 1624857261
transform 1 0 217464 0 1 134781
box 0 0 1 1
use contact_32  contact_32_44
timestamp 1624857261
transform 1 0 217464 0 1 15645
box 0 0 1 1
use contact_32  contact_32_43
timestamp 1624857261
transform 1 0 217464 0 1 55901
box 0 0 1 1
use contact_32  contact_32_42
timestamp 1624857261
transform 1 0 217464 0 1 20541
box 0 0 1 1
use contact_32  contact_32_41
timestamp 1624857261
transform 1 0 217464 0 1 57533
box 0 0 1 1
use contact_32  contact_32_40
timestamp 1624857261
transform 1 0 217464 0 1 64333
box 0 0 1 1
use contact_32  contact_32_39
timestamp 1624857261
transform 1 0 217464 0 1 111389
box 0 0 1 1
use contact_32  contact_32_38
timestamp 1624857261
transform 1 0 217464 0 1 52637
box 0 0 1 1
use contact_32  contact_32_37
timestamp 1624857261
transform 1 0 217464 0 1 139949
box 0 0 1 1
use contact_32  contact_32_36
timestamp 1624857261
transform 1 0 217464 0 1 19045
box 0 0 1 1
use contact_32  contact_32_35
timestamp 1624857261
transform 1 0 217464 0 1 25709
box 0 0 1 1
use contact_32  contact_32_34
timestamp 1624857261
transform 1 0 217464 0 1 96293
box 0 0 1 1
use contact_32  contact_32_33
timestamp 1624857261
transform 1 0 217464 0 1 37541
box 0 0 1 1
use contact_32  contact_32_32
timestamp 1624857261
transform 1 0 217464 0 1 133285
box 0 0 1 1
use contact_32  contact_32_31
timestamp 1624857261
transform 1 0 217464 0 1 118189
box 0 0 1 1
use contact_32  contact_32_30
timestamp 1624857261
transform 1 0 217464 0 1 30605
box 0 0 1 1
use contact_32  contact_32_29
timestamp 1624857261
transform 1 0 217464 0 1 76029
box 0 0 1 1
use contact_32  contact_32_28
timestamp 1624857261
transform 1 0 217464 0 1 62701
box 0 0 1 1
use contact_32  contact_32_27
timestamp 1624857261
transform 1 0 217464 0 1 91261
box 0 0 1 1
use contact_32  contact_32_26
timestamp 1624857261
transform 1 0 217464 0 1 67597
box 0 0 1 1
use contact_32  contact_32_25
timestamp 1624857261
transform 1 0 217464 0 1 121453
box 0 0 1 1
use contact_32  contact_32_24
timestamp 1624857261
transform 1 0 217464 0 1 40805
box 0 0 1 1
use contact_32  contact_32_23
timestamp 1624857261
transform 1 0 217464 0 1 24077
box 0 0 1 1
use contact_32  contact_32_22
timestamp 1624857261
transform 1 0 217464 0 1 92893
box 0 0 1 1
use contact_32  contact_32_21
timestamp 1624857261
transform 1 0 217464 0 1 35773
box 0 0 1 1
use contact_32  contact_32_20
timestamp 1624857261
transform 1 0 217464 0 1 34141
box 0 0 1 1
use contact_32  contact_32_19
timestamp 1624857261
transform 1 0 217464 0 1 44205
box 0 0 1 1
use contact_32  contact_32_18
timestamp 1624857261
transform 1 0 217464 0 1 79293
box 0 0 1 1
use contact_32  contact_32_17
timestamp 1624857261
transform 1 0 217464 0 1 104589
box 0 0 1 1
use contact_32  contact_32_16
timestamp 1624857261
transform 1 0 217464 0 1 14013
box 0 0 1 1
use contact_32  contact_32_15
timestamp 1624857261
transform 1 0 217464 0 1 61069
box 0 0 1 1
use contact_32  contact_32_14
timestamp 1624857261
transform 1 0 217464 0 1 123085
box 0 0 1 1
use contact_32  contact_32_13
timestamp 1624857261
transform 1 0 217464 0 1 3949
box 0 0 1 1
use contact_32  contact_32_12
timestamp 1624857261
transform 1 0 217464 0 1 7213
box 0 0 1 1
use contact_32  contact_32_11
timestamp 1624857261
transform 1 0 217464 0 1 99693
box 0 0 1 1
use contact_32  contact_32_10
timestamp 1624857261
transform 1 0 217464 0 1 71133
box 0 0 1 1
use contact_32  contact_32_9
timestamp 1624857261
transform 1 0 217464 0 1 128253
box 0 0 1 1
use contact_32  contact_32_8
timestamp 1624857261
transform 1 0 217464 0 1 124717
box 0 0 1 1
use contact_32  contact_32_7
timestamp 1624857261
transform 1 0 217464 0 1 112885
box 0 0 1 1
use contact_32  contact_32_6
timestamp 1624857261
transform 1 0 217464 0 1 8845
box 0 0 1 1
use contact_32  contact_32_5
timestamp 1624857261
transform 1 0 217464 0 1 39037
box 0 0 1 1
use contact_32  contact_32_4
timestamp 1624857261
transform 1 0 217464 0 1 87725
box 0 0 1 1
use contact_32  contact_32_3
timestamp 1624857261
transform 1 0 217464 0 1 116285
box 0 0 1 1
use contact_32  contact_32_2
timestamp 1624857261
transform 1 0 217464 0 1 89629
box 0 0 1 1
use contact_32  contact_32_1
timestamp 1624857261
transform 1 0 217464 0 1 32509
box 0 0 1 1
use contact_32  contact_32_0
timestamp 1624857261
transform 1 0 217464 0 1 114789
box 0 0 1 1
use contact_37  contact_37_0
timestamp 1624857261
transform 1 0 1634 0 1 142248
box 0 0 192 192
use contact_37  contact_37_1
timestamp 1624857261
transform 1 0 216840 0 1 142248
box 0 0 192 192
use contact_37  contact_37_2
timestamp 1624857261
transform 1 0 216840 0 1 1752
box 0 0 192 192
use contact_37  contact_37_3
timestamp 1624857261
transform 1 0 1634 0 1 1752
box 0 0 192 192
use contact_31  contact_31_0
timestamp 1624857261
transform 1 0 203395 0 1 141663
box 0 0 1 1
use contact_31  contact_31_1
timestamp 1624857261
transform 1 0 203395 0 1 24492
box 0 0 1 1
use contact_31  contact_31_2
timestamp 1624857261
transform 1 0 15289 0 1 2455
box 0 0 1 1
use contact_31  contact_31_3
timestamp 1624857261
transform 1 0 15289 0 1 34588
box 0 0 1 1
<< labels >>
rlabel metal3 s 0 13192 76 13268 4 csb0
port 54 nsew default input
rlabel metal3 s 0 14960 76 15036 4 web0
port 56 nsew default input
rlabel metal3 s 0 13328 76 13404 4 clk0
port 57 nsew default input
rlabel metal4 s 24616 0 24692 76 4 din0[0]
port 0 nsew default input
rlabel metal4 s 25976 0 26052 76 4 din0[1]
port 1 nsew default input
rlabel metal4 s 27064 0 27140 76 4 din0[2]
port 2 nsew default input
rlabel metal4 s 28288 0 28364 76 4 din0[3]
port 3 nsew default input
rlabel metal4 s 29240 0 29316 76 4 din0[4]
port 4 nsew default input
rlabel metal4 s 30600 0 30676 76 4 din0[5]
port 5 nsew default input
rlabel metal4 s 31688 0 31764 76 4 din0[6]
port 6 nsew default input
rlabel metal4 s 32776 0 32852 76 4 din0[7]
port 7 nsew default input
rlabel metal4 s 34000 0 34076 76 4 din0[8]
port 8 nsew default input
rlabel metal4 s 35088 0 35164 76 4 din0[9]
port 9 nsew default input
rlabel metal4 s 36448 0 36524 76 4 din0[10]
port 10 nsew default input
rlabel metal4 s 37536 0 37612 76 4 din0[11]
port 11 nsew default input
rlabel metal4 s 38624 0 38700 76 4 din0[12]
port 12 nsew default input
rlabel metal4 s 39848 0 39924 76 4 din0[13]
port 13 nsew default input
rlabel metal4 s 40936 0 41012 76 4 din0[14]
port 14 nsew default input
rlabel metal4 s 42296 0 42372 76 4 din0[15]
port 15 nsew default input
rlabel metal4 s 43384 0 43460 76 4 din0[16]
port 16 nsew default input
rlabel metal4 s 44608 0 44684 76 4 din0[17]
port 17 nsew default input
rlabel metal4 s 45832 0 45908 76 4 din0[18]
port 18 nsew default input
rlabel metal4 s 46920 0 46996 76 4 din0[19]
port 19 nsew default input
rlabel metal4 s 48008 0 48084 76 4 din0[20]
port 20 nsew default input
rlabel metal4 s 49096 0 49172 76 4 din0[21]
port 21 nsew default input
rlabel metal4 s 50320 0 50396 76 4 din0[22]
port 22 nsew default input
rlabel metal4 s 51544 0 51620 76 4 din0[23]
port 23 nsew default input
rlabel metal4 s 52768 0 52844 76 4 din0[24]
port 24 nsew default input
rlabel metal4 s 53856 0 53932 76 4 din0[25]
port 25 nsew default input
rlabel metal4 s 54944 0 55020 76 4 din0[26]
port 26 nsew default input
rlabel metal4 s 56168 0 56244 76 4 din0[27]
port 27 nsew default input
rlabel metal4 s 57392 0 57468 76 4 din0[28]
port 28 nsew default input
rlabel metal4 s 58616 0 58692 76 4 din0[29]
port 29 nsew default input
rlabel metal4 s 59840 0 59916 76 4 din0[30]
port 30 nsew default input
rlabel metal4 s 60792 0 60868 76 4 din0[31]
port 31 nsew default input
rlabel metal4 s 28968 0 29044 76 4 dout0[0]
port 63 nsew default output
rlabel metal4 s 34544 0 34620 76 4 dout0[1]
port 64 nsew default output
rlabel metal4 s 39440 0 39516 76 4 dout0[2]
port 65 nsew default output
rlabel metal4 s 44200 0 44276 76 4 dout0[3]
port 66 nsew default output
rlabel metal4 s 49504 0 49580 76 4 dout0[4]
port 67 nsew default output
rlabel metal4 s 54536 0 54612 76 4 dout0[5]
port 68 nsew default output
rlabel metal4 s 59296 0 59372 76 4 dout0[6]
port 69 nsew default output
rlabel metal4 s 64464 0 64540 76 4 dout0[7]
port 70 nsew default output
rlabel metal4 s 69496 0 69572 76 4 dout0[8]
port 71 nsew default output
rlabel metal4 s 74392 0 74468 76 4 dout0[9]
port 72 nsew default output
rlabel metal4 s 79424 0 79500 76 4 dout0[10]
port 73 nsew default output
rlabel metal4 s 84320 0 84396 76 4 dout0[11]
port 74 nsew default output
rlabel metal4 s 89352 0 89428 76 4 dout0[12]
port 75 nsew default output
rlabel metal4 s 94384 0 94460 76 4 dout0[13]
port 76 nsew default output
rlabel metal4 s 99416 0 99492 76 4 dout0[14]
port 77 nsew default output
rlabel metal4 s 104312 0 104388 76 4 dout0[15]
port 78 nsew default output
rlabel metal4 s 109072 0 109148 76 4 dout0[16]
port 79 nsew default output
rlabel metal4 s 114376 0 114452 76 4 dout0[17]
port 80 nsew default output
rlabel metal4 s 119272 0 119348 76 4 dout0[18]
port 81 nsew default output
rlabel metal4 s 124304 0 124380 76 4 dout0[19]
port 82 nsew default output
rlabel metal4 s 129336 0 129412 76 4 dout0[20]
port 83 nsew default output
rlabel metal4 s 134368 0 134444 76 4 dout0[21]
port 84 nsew default output
rlabel metal4 s 139264 0 139340 76 4 dout0[22]
port 85 nsew default output
rlabel metal4 s 144296 0 144372 76 4 dout0[23]
port 86 nsew default output
rlabel metal4 s 149056 0 149132 76 4 dout0[24]
port 87 nsew default output
rlabel metal4 s 154224 0 154300 76 4 dout0[25]
port 88 nsew default output
rlabel metal4 s 159256 0 159332 76 4 dout0[26]
port 89 nsew default output
rlabel metal4 s 164288 0 164364 76 4 dout0[27]
port 90 nsew default output
rlabel metal4 s 169184 0 169260 76 4 dout0[28]
port 91 nsew default output
rlabel metal4 s 174216 0 174292 76 4 dout0[29]
port 92 nsew default output
rlabel metal4 s 179248 0 179324 76 4 dout0[30]
port 93 nsew default output
rlabel metal4 s 184280 0 184356 76 4 dout0[31]
port 94 nsew default output
rlabel metal4 s 16456 0 16532 76 4 addr0[0]
port 32 nsew default input
rlabel metal4 s 17680 0 17756 76 4 addr0[1]
port 33 nsew default input
rlabel metal4 s 18768 0 18844 76 4 addr0[2]
port 34 nsew default input
rlabel metal3 s 0 34816 76 34892 4 addr0[3]
port 35 nsew default input
rlabel metal3 s 0 36448 76 36524 4 addr0[4]
port 36 nsew default input
rlabel metal3 s 0 37808 76 37884 4 addr0[5]
port 37 nsew default input
rlabel metal3 s 0 39440 76 39516 4 addr0[6]
port 38 nsew default input
rlabel metal3 s 0 40528 76 40604 4 addr0[7]
port 39 nsew default input
rlabel metal3 s 0 42160 76 42236 4 addr0[8]
port 40 nsew default input
rlabel metal3 s 0 43248 76 43324 4 addr0[9]
port 41 nsew default input
rlabel metal3 s 0 45152 76 45228 4 addr0[10]
port 42 nsew default input
rlabel metal4 s 19992 0 20068 76 4 wmask0[0]
port 59 nsew default input
rlabel metal4 s 21080 0 21156 76 4 wmask0[1]
port 60 nsew default input
rlabel metal4 s 22304 0 22380 76 4 wmask0[2]
port 61 nsew default input
rlabel metal4 s 23528 0 23604 76 4 wmask0[3]
port 62 nsew default input
rlabel metal3 s 218688 134640 218764 134716 4 csb1
port 55 nsew default input
rlabel metal3 s 218688 134504 218764 134580 4 clk1
port 58 nsew default input
rlabel metal4 s 29512 144024 29588 144100 4 dout1[0]
port 95 nsew default output
rlabel metal4 s 34408 144024 34484 144100 4 dout1[1]
port 96 nsew default output
rlabel metal4 s 39440 144024 39516 144100 4 dout1[2]
port 97 nsew default output
rlabel metal4 s 44472 144024 44548 144100 4 dout1[3]
port 98 nsew default output
rlabel metal4 s 49504 144024 49580 144100 4 dout1[4]
port 99 nsew default output
rlabel metal4 s 54536 144024 54612 144100 4 dout1[5]
port 100 nsew default output
rlabel metal4 s 59432 144024 59508 144100 4 dout1[6]
port 101 nsew default output
rlabel metal4 s 64464 144024 64540 144100 4 dout1[7]
port 102 nsew default output
rlabel metal4 s 69496 144024 69572 144100 4 dout1[8]
port 103 nsew default output
rlabel metal4 s 74528 144024 74604 144100 4 dout1[9]
port 104 nsew default output
rlabel metal4 s 79560 144024 79636 144100 4 dout1[10]
port 105 nsew default output
rlabel metal4 s 84320 144024 84396 144100 4 dout1[11]
port 106 nsew default output
rlabel metal4 s 89352 144024 89428 144100 4 dout1[12]
port 107 nsew default output
rlabel metal4 s 94520 144024 94596 144100 4 dout1[13]
port 108 nsew default output
rlabel metal4 s 99416 144024 99492 144100 4 dout1[14]
port 109 nsew default output
rlabel metal4 s 104312 144024 104388 144100 4 dout1[15]
port 110 nsew default output
rlabel metal4 s 109344 144024 109420 144100 4 dout1[16]
port 111 nsew default output
rlabel metal4 s 114376 144024 114452 144100 4 dout1[17]
port 112 nsew default output
rlabel metal4 s 119272 144024 119348 144100 4 dout1[18]
port 113 nsew default output
rlabel metal4 s 124304 144024 124380 144100 4 dout1[19]
port 114 nsew default output
rlabel metal4 s 129336 144024 129412 144100 4 dout1[20]
port 115 nsew default output
rlabel metal4 s 134368 144024 134444 144100 4 dout1[21]
port 116 nsew default output
rlabel metal4 s 139400 144024 139476 144100 4 dout1[22]
port 117 nsew default output
rlabel metal4 s 144296 144024 144372 144100 4 dout1[23]
port 118 nsew default output
rlabel metal4 s 149328 144024 149404 144100 4 dout1[24]
port 119 nsew default output
rlabel metal4 s 154360 144024 154436 144100 4 dout1[25]
port 120 nsew default output
rlabel metal4 s 159392 144024 159468 144100 4 dout1[26]
port 121 nsew default output
rlabel metal4 s 164424 144024 164500 144100 4 dout1[27]
port 122 nsew default output
rlabel metal4 s 169184 144024 169260 144100 4 dout1[28]
port 123 nsew default output
rlabel metal4 s 174216 144024 174292 144100 4 dout1[29]
port 124 nsew default output
rlabel metal4 s 179384 144024 179460 144100 4 dout1[30]
port 125 nsew default output
rlabel metal4 s 184280 144024 184356 144100 4 dout1[31]
port 126 nsew default output
rlabel metal4 s 201008 144024 201084 144100 4 addr1[0]
port 43 nsew default input
rlabel metal4 s 199920 144024 199996 144100 4 addr1[1]
port 44 nsew default input
rlabel metal4 s 198560 144024 198636 144100 4 addr1[2]
port 45 nsew default input
rlabel metal3 s 218688 24208 218764 24284 4 addr1[3]
port 46 nsew default input
rlabel metal3 s 218688 22576 218764 22652 4 addr1[4]
port 47 nsew default input
rlabel metal3 s 218688 21488 218764 21564 4 addr1[5]
port 48 nsew default input
rlabel metal3 s 218688 19584 218764 19660 4 addr1[6]
port 49 nsew default input
rlabel metal3 s 218688 18496 218764 18572 4 addr1[7]
port 50 nsew default input
rlabel metal3 s 218688 16864 218764 16940 4 addr1[8]
port 51 nsew default input
rlabel metal3 s 218688 15776 218764 15852 4 addr1[9]
port 52 nsew default input
rlabel metal3 s 218688 14144 218764 14220 4 addr1[10]
port 53 nsew default input
rlabel metal3 s 272 272 218492 620 4 vccd1
port 127 nsew power bidirectional abutment
rlabel metal4 s 272 272 620 143828 4 vccd1
port 128 nsew power bidirectional abutment
rlabel metal3 s 272 143480 218492 143828 4 vccd1
port 129 nsew power bidirectional abutment
rlabel metal4 s 218144 272 218492 143828 4 vccd1
port 130 nsew power bidirectional abutment
rlabel metal3 s 952 142800 217812 143148 4 vssd1
port 131 nsew ground bidirectional abutment
rlabel metal4 s 217464 952 217812 143148 4 vssd1
port 132 nsew ground bidirectional abutment
rlabel metal3 s 952 952 217812 1300 4 vssd1
port 133 nsew ground bidirectional abutment
rlabel metal4 s 952 952 1300 143148 4 vssd1
port 134 nsew ground bidirectional abutment
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 218764 144100
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_8kbyte_1rw1r_32x2048_8.gds
string LEFsymmetry X Y R90
string GDS_END 2994894
string GDS_START 134
<< end >>
