magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1319 -1314 1469 1424
<< nwell >>
rect -54 139 204 164
rect -59 -29 209 139
rect -54 -54 204 -29
<< scpmos >>
rect 60 0 90 110
<< pdiff >>
rect 0 72 60 110
rect 0 38 8 72
rect 42 38 60 72
rect 0 0 60 38
rect 90 72 150 110
rect 90 38 108 72
rect 142 38 150 72
rect 90 0 150 38
<< pdiffc >>
rect 8 38 42 72
rect 108 38 142 72
<< poly >>
rect 60 110 90 136
rect 60 -26 90 0
<< locali >>
rect 8 72 42 88
rect 8 22 42 38
rect 108 72 142 88
rect 108 22 142 38
use contact_12  contact_12_0
timestamp 1624857261
transform 1 0 100 0 1 22
box 0 0 1 1
use contact_12  contact_12_1
timestamp 1624857261
transform 1 0 0 0 1 22
box 0 0 1 1
<< labels >>
rlabel poly s 75 55 75 55 4 G
rlabel locali s 25 55 25 55 4 S
rlabel locali s 125 55 125 55 4 D
<< properties >>
string FIXED_BBOX -54 -54 204 -29
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 7704856
string GDS_START 7704064
<< end >>
