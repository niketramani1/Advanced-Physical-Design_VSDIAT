magic
tech sky130A
magscale 1 2
timestamp 1624855602
<< nwell >>
rect -66 377 4098 897
rect 3281 344 3619 377
<< pwell >>
rect 0 -17 4032 17
<< locali >>
rect 303 567 353 599
rect 303 533 608 567
rect 131 259 197 393
rect 163 87 197 259
rect 313 325 466 427
rect 742 431 808 496
rect 742 395 941 431
rect 697 289 839 359
rect 303 255 839 289
rect 875 259 941 395
rect 303 87 337 255
rect 1047 424 1127 430
rect 1047 390 1087 424
rect 1121 390 1127 424
rect 1047 259 1127 390
rect 1174 370 1240 504
rect 163 53 337 87
rect 2137 424 2249 427
rect 2137 390 2143 424
rect 2177 390 2249 424
rect 2137 325 2249 390
rect 3001 390 3007 424
rect 3041 390 3137 424
rect 3001 285 3137 390
rect 3487 103 3567 714
rect 3940 137 4008 751
<< viali >>
rect 1087 390 1121 424
rect 2143 390 2177 424
rect 3007 390 3041 424
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
rect 18 735 197 741
rect 18 701 19 735
rect 53 701 91 735
rect 125 701 163 735
rect 18 641 197 701
rect 233 641 283 741
rect 335 647 423 747
rect 509 735 699 747
rect 509 701 515 735
rect 549 701 587 735
rect 621 701 659 735
rect 693 701 699 735
rect 509 673 699 701
rect 233 497 267 641
rect 389 637 423 647
rect 931 637 981 747
rect 1017 735 1195 751
rect 1051 701 1089 735
rect 1123 701 1161 735
rect 1017 673 1195 701
rect 1231 727 1405 761
rect 1231 637 1265 727
rect 389 603 1265 637
rect 654 533 936 567
rect 654 497 688 533
rect 233 463 688 497
rect 18 113 127 223
rect 18 79 19 113
rect 53 79 91 113
rect 125 79 127 113
rect 18 73 127 79
rect 233 123 267 463
rect 546 325 612 463
rect 870 465 936 533
rect 977 219 1011 603
rect 1301 335 1335 691
rect 1371 405 1405 727
rect 1441 735 1475 741
rect 1441 441 1475 701
rect 1655 685 1721 751
rect 1511 651 1791 685
rect 1511 405 1545 651
rect 1671 603 1721 615
rect 1371 371 1545 405
rect 1581 445 1721 603
rect 1301 301 1539 335
rect 373 87 423 199
rect 655 185 1011 219
rect 655 123 721 185
rect 953 87 1019 151
rect 373 53 1019 87
rect 1055 113 1245 199
rect 1055 79 1061 113
rect 1095 79 1133 113
rect 1167 79 1205 113
rect 1239 79 1245 113
rect 1301 99 1335 301
rect 1473 269 1539 301
rect 1581 199 1630 445
rect 1757 199 1791 651
rect 1374 113 1544 183
rect 1055 73 1245 79
rect 1374 79 1390 113
rect 1424 79 1494 113
rect 1528 79 1544 113
rect 1374 73 1544 79
rect 1580 87 1630 199
rect 1682 123 1791 199
rect 1827 615 1877 751
rect 1985 735 2175 751
rect 1985 701 1991 735
rect 2025 701 2063 735
rect 2097 701 2135 735
rect 2169 701 2175 735
rect 1985 651 2175 701
rect 2265 615 2355 747
rect 1827 581 2355 615
rect 2391 735 2509 747
rect 2391 701 2397 735
rect 2431 701 2469 735
rect 2503 701 2509 735
rect 2391 603 2509 701
rect 1827 199 1861 581
rect 2265 567 2355 581
rect 1902 497 1968 535
rect 2265 533 2389 567
rect 1902 463 2319 497
rect 1902 401 1968 463
rect 1940 219 1995 351
rect 2045 289 2101 389
rect 2285 409 2319 463
rect 2355 445 2389 533
rect 2547 539 2597 751
rect 2687 609 2753 751
rect 2960 735 3144 741
rect 2960 701 2963 735
rect 2997 701 3035 735
rect 3069 701 3107 735
rect 3141 701 3144 735
rect 2687 575 2924 609
rect 2547 505 2714 539
rect 2425 435 2644 469
rect 2425 409 2459 435
rect 2285 375 2459 409
rect 2680 399 2714 505
rect 2495 365 2714 399
rect 2495 289 2529 365
rect 2045 255 2529 289
rect 1827 123 1904 199
rect 1940 185 2429 219
rect 1940 87 1995 185
rect 1580 53 1995 87
rect 2154 113 2361 149
rect 2154 79 2160 113
rect 2194 79 2232 113
rect 2266 79 2304 113
rect 2338 79 2361 113
rect 2154 73 2361 79
rect 2395 87 2429 185
rect 2463 123 2529 255
rect 2565 295 2631 329
rect 2565 87 2599 295
rect 2750 259 2784 575
rect 2635 225 2784 259
rect 2635 123 2685 225
rect 2820 87 2854 511
rect 2890 249 2924 575
rect 2960 535 3144 701
rect 3266 735 3451 741
rect 3266 701 3269 735
rect 3303 701 3341 735
rect 3375 701 3413 735
rect 3447 701 3451 735
rect 3707 735 3897 751
rect 3180 499 3230 635
rect 2960 460 3230 499
rect 3196 401 3230 460
rect 3266 437 3451 701
rect 3196 367 3309 401
rect 3173 249 3239 331
rect 2890 215 3239 249
rect 3275 179 3309 367
rect 2395 53 2854 87
rect 2890 113 3080 179
rect 2890 79 2896 113
rect 2930 79 2968 113
rect 3002 79 3040 113
rect 3074 79 3080 113
rect 3235 103 3309 179
rect 3345 113 3451 261
rect 2890 73 3080 79
rect 3379 79 3417 113
rect 3707 701 3713 735
rect 3747 701 3785 735
rect 3819 701 3857 735
rect 3891 701 3897 735
rect 3605 397 3671 597
rect 3707 435 3897 701
rect 3605 331 3904 397
rect 3605 137 3677 331
rect 3713 113 3903 295
rect 3345 73 3451 79
rect 3713 79 3719 113
rect 3753 79 3791 113
rect 3825 79 3863 113
rect 3897 79 3903 113
rect 3713 73 3903 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
rect 19 701 53 735
rect 91 701 125 735
rect 163 701 197 735
rect 515 701 549 735
rect 587 701 621 735
rect 659 701 693 735
rect 1017 701 1051 735
rect 1089 701 1123 735
rect 1161 701 1195 735
rect 19 79 53 113
rect 91 79 125 113
rect 1441 701 1475 735
rect 1061 79 1095 113
rect 1133 79 1167 113
rect 1205 79 1239 113
rect 1390 79 1424 113
rect 1494 79 1528 113
rect 1991 701 2025 735
rect 2063 701 2097 735
rect 2135 701 2169 735
rect 2397 701 2431 735
rect 2469 701 2503 735
rect 2963 701 2997 735
rect 3035 701 3069 735
rect 3107 701 3141 735
rect 2160 79 2194 113
rect 2232 79 2266 113
rect 2304 79 2338 113
rect 3269 701 3303 735
rect 3341 701 3375 735
rect 3413 701 3447 735
rect 2896 79 2930 113
rect 2968 79 3002 113
rect 3040 79 3074 113
rect 3345 79 3379 113
rect 3417 79 3451 113
rect 3713 701 3747 735
rect 3785 701 3819 735
rect 3857 701 3891 735
rect 3719 79 3753 113
rect 3791 79 3825 113
rect 3863 79 3897 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
<< metal1 >>
rect 0 831 4032 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
rect 0 791 4032 797
rect 0 735 4032 763
rect 0 701 19 735
rect 53 701 91 735
rect 125 701 163 735
rect 197 701 515 735
rect 549 701 587 735
rect 621 701 659 735
rect 693 701 1017 735
rect 1051 701 1089 735
rect 1123 701 1161 735
rect 1195 701 1441 735
rect 1475 701 1991 735
rect 2025 701 2063 735
rect 2097 701 2135 735
rect 2169 701 2397 735
rect 2431 701 2469 735
rect 2503 701 2963 735
rect 2997 701 3035 735
rect 3069 701 3107 735
rect 3141 701 3269 735
rect 3303 701 3341 735
rect 3375 701 3413 735
rect 3447 701 3713 735
rect 3747 701 3785 735
rect 3819 701 3857 735
rect 3891 701 4032 735
rect 0 689 4032 701
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1121 393 2143 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 2131 390 2143 393
rect 2177 421 2189 424
rect 2995 424 3053 430
rect 2995 421 3007 424
rect 2177 393 3007 421
rect 2177 390 2189 393
rect 2131 384 2189 390
rect 2995 390 3007 393
rect 3041 390 3053 424
rect 2995 384 3053 390
rect 0 113 4032 125
rect 0 79 19 113
rect 53 79 91 113
rect 125 79 1061 113
rect 1095 79 1133 113
rect 1167 79 1205 113
rect 1239 79 1390 113
rect 1424 79 1494 113
rect 1528 79 2160 113
rect 2194 79 2232 113
rect 2266 79 2304 113
rect 2338 79 2896 113
rect 2930 79 2968 113
rect 3002 79 3040 113
rect 3074 79 3345 113
rect 3379 79 3417 113
rect 3451 79 3719 113
rect 3753 79 3791 113
rect 3825 79 3863 113
rect 3897 79 4032 113
rect 0 51 4032 79
rect 0 17 4032 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
rect 0 -23 4032 -17
<< labels >>
rlabel locali s 313 325 466 427 6 D
port 2 nsew signal input
rlabel locali s 3940 137 4008 751 6 Q
port 10 nsew signal output
rlabel locali s 3487 103 3567 714 6 Q_N
port 11 nsew signal output
rlabel viali s 2143 390 2177 424 6 RESET_B
port 3 nsew signal input
rlabel viali s 1087 390 1121 424 6 RESET_B
port 3 nsew signal input
rlabel locali s 2137 325 2249 427 6 RESET_B
port 3 nsew signal input
rlabel locali s 1047 259 1127 430 6 RESET_B
port 3 nsew signal input
rlabel viali s 3007 390 3041 424 6 RESET_B
port 3 nsew signal input
rlabel locali s 3001 285 3137 424 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2995 421 3053 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2995 384 3053 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2131 421 2189 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2131 384 2189 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1075 421 1133 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1075 393 3053 421 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1075 384 1133 393 6 RESET_B
port 3 nsew signal input
rlabel locali s 875 259 941 395 6 SCD
port 4 nsew signal input
rlabel locali s 742 431 808 496 6 SCD
port 4 nsew signal input
rlabel locali s 742 395 941 431 6 SCD
port 4 nsew signal input
rlabel locali s 697 289 839 359 6 SCE
port 5 nsew signal input
rlabel locali s 303 567 353 599 6 SCE
port 5 nsew signal input
rlabel locali s 303 533 608 567 6 SCE
port 5 nsew signal input
rlabel locali s 303 255 839 289 6 SCE
port 5 nsew signal input
rlabel locali s 303 87 337 255 6 SCE
port 5 nsew signal input
rlabel locali s 163 87 197 259 6 SCE
port 5 nsew signal input
rlabel locali s 163 53 337 87 6 SCE
port 5 nsew signal input
rlabel locali s 131 259 197 393 6 SCE
port 5 nsew signal input
rlabel locali s 1174 370 1240 504 6 CLK
port 1 nsew clock input
rlabel metal1 s 0 51 4032 125 6 VGND
port 6 nsew ground bidirectional
rlabel pwell s 0 -17 4032 17 8 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 -23 4032 23 8 VNB
port 7 nsew ground bidirectional
rlabel nwell s 3281 344 3619 377 6 VPB
port 8 nsew power bidirectional
rlabel nwell s -66 377 4098 897 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 791 4032 837 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 689 4032 763 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 4032 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 1008942
string GDS_START 974848
<< end >>
