magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1260 -1260 140056 135024
<< dnwell >>
rect 1826 1724 136972 132033
<< nwell >>
rect 1742 131949 137056 132117
rect 1742 1808 1910 131949
rect 136888 1808 137056 131949
rect 1742 1640 137056 1808
<< nsubdiff >>
rect 2137 132050 2187 132074
rect 2137 132016 2145 132050
rect 2179 132016 2187 132050
rect 2137 131992 2187 132016
rect 2473 132050 2523 132074
rect 2473 132016 2481 132050
rect 2515 132016 2523 132050
rect 2473 131992 2523 132016
rect 2809 132050 2859 132074
rect 2809 132016 2817 132050
rect 2851 132016 2859 132050
rect 2809 131992 2859 132016
rect 3145 132050 3195 132074
rect 3145 132016 3153 132050
rect 3187 132016 3195 132050
rect 3145 131992 3195 132016
rect 3481 132050 3531 132074
rect 3481 132016 3489 132050
rect 3523 132016 3531 132050
rect 3481 131992 3531 132016
rect 3817 132050 3867 132074
rect 3817 132016 3825 132050
rect 3859 132016 3867 132050
rect 3817 131992 3867 132016
rect 4153 132050 4203 132074
rect 4153 132016 4161 132050
rect 4195 132016 4203 132050
rect 4153 131992 4203 132016
rect 4489 132050 4539 132074
rect 4489 132016 4497 132050
rect 4531 132016 4539 132050
rect 4489 131992 4539 132016
rect 4825 132050 4875 132074
rect 4825 132016 4833 132050
rect 4867 132016 4875 132050
rect 4825 131992 4875 132016
rect 5161 132050 5211 132074
rect 5161 132016 5169 132050
rect 5203 132016 5211 132050
rect 5161 131992 5211 132016
rect 5497 132050 5547 132074
rect 5497 132016 5505 132050
rect 5539 132016 5547 132050
rect 5497 131992 5547 132016
rect 5833 132050 5883 132074
rect 5833 132016 5841 132050
rect 5875 132016 5883 132050
rect 5833 131992 5883 132016
rect 6169 132050 6219 132074
rect 6169 132016 6177 132050
rect 6211 132016 6219 132050
rect 6169 131992 6219 132016
rect 6505 132050 6555 132074
rect 6505 132016 6513 132050
rect 6547 132016 6555 132050
rect 6505 131992 6555 132016
rect 6841 132050 6891 132074
rect 6841 132016 6849 132050
rect 6883 132016 6891 132050
rect 6841 131992 6891 132016
rect 7177 132050 7227 132074
rect 7177 132016 7185 132050
rect 7219 132016 7227 132050
rect 7177 131992 7227 132016
rect 7513 132050 7563 132074
rect 7513 132016 7521 132050
rect 7555 132016 7563 132050
rect 7513 131992 7563 132016
rect 7849 132050 7899 132074
rect 7849 132016 7857 132050
rect 7891 132016 7899 132050
rect 7849 131992 7899 132016
rect 8185 132050 8235 132074
rect 8185 132016 8193 132050
rect 8227 132016 8235 132050
rect 8185 131992 8235 132016
rect 8521 132050 8571 132074
rect 8521 132016 8529 132050
rect 8563 132016 8571 132050
rect 8521 131992 8571 132016
rect 8857 132050 8907 132074
rect 8857 132016 8865 132050
rect 8899 132016 8907 132050
rect 8857 131992 8907 132016
rect 9193 132050 9243 132074
rect 9193 132016 9201 132050
rect 9235 132016 9243 132050
rect 9193 131992 9243 132016
rect 9529 132050 9579 132074
rect 9529 132016 9537 132050
rect 9571 132016 9579 132050
rect 9529 131992 9579 132016
rect 9865 132050 9915 132074
rect 9865 132016 9873 132050
rect 9907 132016 9915 132050
rect 9865 131992 9915 132016
rect 10201 132050 10251 132074
rect 10201 132016 10209 132050
rect 10243 132016 10251 132050
rect 10201 131992 10251 132016
rect 10537 132050 10587 132074
rect 10537 132016 10545 132050
rect 10579 132016 10587 132050
rect 10537 131992 10587 132016
rect 10873 132050 10923 132074
rect 10873 132016 10881 132050
rect 10915 132016 10923 132050
rect 10873 131992 10923 132016
rect 11209 132050 11259 132074
rect 11209 132016 11217 132050
rect 11251 132016 11259 132050
rect 11209 131992 11259 132016
rect 11545 132050 11595 132074
rect 11545 132016 11553 132050
rect 11587 132016 11595 132050
rect 11545 131992 11595 132016
rect 11881 132050 11931 132074
rect 11881 132016 11889 132050
rect 11923 132016 11931 132050
rect 11881 131992 11931 132016
rect 12217 132050 12267 132074
rect 12217 132016 12225 132050
rect 12259 132016 12267 132050
rect 12217 131992 12267 132016
rect 12553 132050 12603 132074
rect 12553 132016 12561 132050
rect 12595 132016 12603 132050
rect 12553 131992 12603 132016
rect 12889 132050 12939 132074
rect 12889 132016 12897 132050
rect 12931 132016 12939 132050
rect 12889 131992 12939 132016
rect 13225 132050 13275 132074
rect 13225 132016 13233 132050
rect 13267 132016 13275 132050
rect 13225 131992 13275 132016
rect 13561 132050 13611 132074
rect 13561 132016 13569 132050
rect 13603 132016 13611 132050
rect 13561 131992 13611 132016
rect 13897 132050 13947 132074
rect 13897 132016 13905 132050
rect 13939 132016 13947 132050
rect 13897 131992 13947 132016
rect 14233 132050 14283 132074
rect 14233 132016 14241 132050
rect 14275 132016 14283 132050
rect 14233 131992 14283 132016
rect 14569 132050 14619 132074
rect 14569 132016 14577 132050
rect 14611 132016 14619 132050
rect 14569 131992 14619 132016
rect 14905 132050 14955 132074
rect 14905 132016 14913 132050
rect 14947 132016 14955 132050
rect 14905 131992 14955 132016
rect 15241 132050 15291 132074
rect 15241 132016 15249 132050
rect 15283 132016 15291 132050
rect 15241 131992 15291 132016
rect 15577 132050 15627 132074
rect 15577 132016 15585 132050
rect 15619 132016 15627 132050
rect 15577 131992 15627 132016
rect 15913 132050 15963 132074
rect 15913 132016 15921 132050
rect 15955 132016 15963 132050
rect 15913 131992 15963 132016
rect 16249 132050 16299 132074
rect 16249 132016 16257 132050
rect 16291 132016 16299 132050
rect 16249 131992 16299 132016
rect 16585 132050 16635 132074
rect 16585 132016 16593 132050
rect 16627 132016 16635 132050
rect 16585 131992 16635 132016
rect 16921 132050 16971 132074
rect 16921 132016 16929 132050
rect 16963 132016 16971 132050
rect 16921 131992 16971 132016
rect 17257 132050 17307 132074
rect 17257 132016 17265 132050
rect 17299 132016 17307 132050
rect 17257 131992 17307 132016
rect 17593 132050 17643 132074
rect 17593 132016 17601 132050
rect 17635 132016 17643 132050
rect 17593 131992 17643 132016
rect 17929 132050 17979 132074
rect 17929 132016 17937 132050
rect 17971 132016 17979 132050
rect 17929 131992 17979 132016
rect 18265 132050 18315 132074
rect 18265 132016 18273 132050
rect 18307 132016 18315 132050
rect 18265 131992 18315 132016
rect 18601 132050 18651 132074
rect 18601 132016 18609 132050
rect 18643 132016 18651 132050
rect 18601 131992 18651 132016
rect 18937 132050 18987 132074
rect 18937 132016 18945 132050
rect 18979 132016 18987 132050
rect 18937 131992 18987 132016
rect 19273 132050 19323 132074
rect 19273 132016 19281 132050
rect 19315 132016 19323 132050
rect 19273 131992 19323 132016
rect 19609 132050 19659 132074
rect 19609 132016 19617 132050
rect 19651 132016 19659 132050
rect 19609 131992 19659 132016
rect 19945 132050 19995 132074
rect 19945 132016 19953 132050
rect 19987 132016 19995 132050
rect 19945 131992 19995 132016
rect 20281 132050 20331 132074
rect 20281 132016 20289 132050
rect 20323 132016 20331 132050
rect 20281 131992 20331 132016
rect 20617 132050 20667 132074
rect 20617 132016 20625 132050
rect 20659 132016 20667 132050
rect 20617 131992 20667 132016
rect 20953 132050 21003 132074
rect 20953 132016 20961 132050
rect 20995 132016 21003 132050
rect 20953 131992 21003 132016
rect 21289 132050 21339 132074
rect 21289 132016 21297 132050
rect 21331 132016 21339 132050
rect 21289 131992 21339 132016
rect 21625 132050 21675 132074
rect 21625 132016 21633 132050
rect 21667 132016 21675 132050
rect 21625 131992 21675 132016
rect 21961 132050 22011 132074
rect 21961 132016 21969 132050
rect 22003 132016 22011 132050
rect 21961 131992 22011 132016
rect 22297 132050 22347 132074
rect 22297 132016 22305 132050
rect 22339 132016 22347 132050
rect 22297 131992 22347 132016
rect 22633 132050 22683 132074
rect 22633 132016 22641 132050
rect 22675 132016 22683 132050
rect 22633 131992 22683 132016
rect 22969 132050 23019 132074
rect 22969 132016 22977 132050
rect 23011 132016 23019 132050
rect 22969 131992 23019 132016
rect 23305 132050 23355 132074
rect 23305 132016 23313 132050
rect 23347 132016 23355 132050
rect 23305 131992 23355 132016
rect 23641 132050 23691 132074
rect 23641 132016 23649 132050
rect 23683 132016 23691 132050
rect 23641 131992 23691 132016
rect 23977 132050 24027 132074
rect 23977 132016 23985 132050
rect 24019 132016 24027 132050
rect 23977 131992 24027 132016
rect 24313 132050 24363 132074
rect 24313 132016 24321 132050
rect 24355 132016 24363 132050
rect 24313 131992 24363 132016
rect 24649 132050 24699 132074
rect 24649 132016 24657 132050
rect 24691 132016 24699 132050
rect 24649 131992 24699 132016
rect 24985 132050 25035 132074
rect 24985 132016 24993 132050
rect 25027 132016 25035 132050
rect 24985 131992 25035 132016
rect 25321 132050 25371 132074
rect 25321 132016 25329 132050
rect 25363 132016 25371 132050
rect 25321 131992 25371 132016
rect 25657 132050 25707 132074
rect 25657 132016 25665 132050
rect 25699 132016 25707 132050
rect 25657 131992 25707 132016
rect 25993 132050 26043 132074
rect 25993 132016 26001 132050
rect 26035 132016 26043 132050
rect 25993 131992 26043 132016
rect 26329 132050 26379 132074
rect 26329 132016 26337 132050
rect 26371 132016 26379 132050
rect 26329 131992 26379 132016
rect 26665 132050 26715 132074
rect 26665 132016 26673 132050
rect 26707 132016 26715 132050
rect 26665 131992 26715 132016
rect 27001 132050 27051 132074
rect 27001 132016 27009 132050
rect 27043 132016 27051 132050
rect 27001 131992 27051 132016
rect 27337 132050 27387 132074
rect 27337 132016 27345 132050
rect 27379 132016 27387 132050
rect 27337 131992 27387 132016
rect 27673 132050 27723 132074
rect 27673 132016 27681 132050
rect 27715 132016 27723 132050
rect 27673 131992 27723 132016
rect 28009 132050 28059 132074
rect 28009 132016 28017 132050
rect 28051 132016 28059 132050
rect 28009 131992 28059 132016
rect 28345 132050 28395 132074
rect 28345 132016 28353 132050
rect 28387 132016 28395 132050
rect 28345 131992 28395 132016
rect 28681 132050 28731 132074
rect 28681 132016 28689 132050
rect 28723 132016 28731 132050
rect 28681 131992 28731 132016
rect 29017 132050 29067 132074
rect 29017 132016 29025 132050
rect 29059 132016 29067 132050
rect 29017 131992 29067 132016
rect 29353 132050 29403 132074
rect 29353 132016 29361 132050
rect 29395 132016 29403 132050
rect 29353 131992 29403 132016
rect 29689 132050 29739 132074
rect 29689 132016 29697 132050
rect 29731 132016 29739 132050
rect 29689 131992 29739 132016
rect 30025 132050 30075 132074
rect 30025 132016 30033 132050
rect 30067 132016 30075 132050
rect 30025 131992 30075 132016
rect 30361 132050 30411 132074
rect 30361 132016 30369 132050
rect 30403 132016 30411 132050
rect 30361 131992 30411 132016
rect 30697 132050 30747 132074
rect 30697 132016 30705 132050
rect 30739 132016 30747 132050
rect 30697 131992 30747 132016
rect 31033 132050 31083 132074
rect 31033 132016 31041 132050
rect 31075 132016 31083 132050
rect 31033 131992 31083 132016
rect 31369 132050 31419 132074
rect 31369 132016 31377 132050
rect 31411 132016 31419 132050
rect 31369 131992 31419 132016
rect 31705 132050 31755 132074
rect 31705 132016 31713 132050
rect 31747 132016 31755 132050
rect 31705 131992 31755 132016
rect 32041 132050 32091 132074
rect 32041 132016 32049 132050
rect 32083 132016 32091 132050
rect 32041 131992 32091 132016
rect 32377 132050 32427 132074
rect 32377 132016 32385 132050
rect 32419 132016 32427 132050
rect 32377 131992 32427 132016
rect 32713 132050 32763 132074
rect 32713 132016 32721 132050
rect 32755 132016 32763 132050
rect 32713 131992 32763 132016
rect 33049 132050 33099 132074
rect 33049 132016 33057 132050
rect 33091 132016 33099 132050
rect 33049 131992 33099 132016
rect 33385 132050 33435 132074
rect 33385 132016 33393 132050
rect 33427 132016 33435 132050
rect 33385 131992 33435 132016
rect 33721 132050 33771 132074
rect 33721 132016 33729 132050
rect 33763 132016 33771 132050
rect 33721 131992 33771 132016
rect 34057 132050 34107 132074
rect 34057 132016 34065 132050
rect 34099 132016 34107 132050
rect 34057 131992 34107 132016
rect 34393 132050 34443 132074
rect 34393 132016 34401 132050
rect 34435 132016 34443 132050
rect 34393 131992 34443 132016
rect 34729 132050 34779 132074
rect 34729 132016 34737 132050
rect 34771 132016 34779 132050
rect 34729 131992 34779 132016
rect 35065 132050 35115 132074
rect 35065 132016 35073 132050
rect 35107 132016 35115 132050
rect 35065 131992 35115 132016
rect 35401 132050 35451 132074
rect 35401 132016 35409 132050
rect 35443 132016 35451 132050
rect 35401 131992 35451 132016
rect 35737 132050 35787 132074
rect 35737 132016 35745 132050
rect 35779 132016 35787 132050
rect 35737 131992 35787 132016
rect 36073 132050 36123 132074
rect 36073 132016 36081 132050
rect 36115 132016 36123 132050
rect 36073 131992 36123 132016
rect 36409 132050 36459 132074
rect 36409 132016 36417 132050
rect 36451 132016 36459 132050
rect 36409 131992 36459 132016
rect 36745 132050 36795 132074
rect 36745 132016 36753 132050
rect 36787 132016 36795 132050
rect 36745 131992 36795 132016
rect 37081 132050 37131 132074
rect 37081 132016 37089 132050
rect 37123 132016 37131 132050
rect 37081 131992 37131 132016
rect 37417 132050 37467 132074
rect 37417 132016 37425 132050
rect 37459 132016 37467 132050
rect 37417 131992 37467 132016
rect 37753 132050 37803 132074
rect 37753 132016 37761 132050
rect 37795 132016 37803 132050
rect 37753 131992 37803 132016
rect 38089 132050 38139 132074
rect 38089 132016 38097 132050
rect 38131 132016 38139 132050
rect 38089 131992 38139 132016
rect 38425 132050 38475 132074
rect 38425 132016 38433 132050
rect 38467 132016 38475 132050
rect 38425 131992 38475 132016
rect 38761 132050 38811 132074
rect 38761 132016 38769 132050
rect 38803 132016 38811 132050
rect 38761 131992 38811 132016
rect 39097 132050 39147 132074
rect 39097 132016 39105 132050
rect 39139 132016 39147 132050
rect 39097 131992 39147 132016
rect 39433 132050 39483 132074
rect 39433 132016 39441 132050
rect 39475 132016 39483 132050
rect 39433 131992 39483 132016
rect 39769 132050 39819 132074
rect 39769 132016 39777 132050
rect 39811 132016 39819 132050
rect 39769 131992 39819 132016
rect 40105 132050 40155 132074
rect 40105 132016 40113 132050
rect 40147 132016 40155 132050
rect 40105 131992 40155 132016
rect 40441 132050 40491 132074
rect 40441 132016 40449 132050
rect 40483 132016 40491 132050
rect 40441 131992 40491 132016
rect 40777 132050 40827 132074
rect 40777 132016 40785 132050
rect 40819 132016 40827 132050
rect 40777 131992 40827 132016
rect 41113 132050 41163 132074
rect 41113 132016 41121 132050
rect 41155 132016 41163 132050
rect 41113 131992 41163 132016
rect 41449 132050 41499 132074
rect 41449 132016 41457 132050
rect 41491 132016 41499 132050
rect 41449 131992 41499 132016
rect 41785 132050 41835 132074
rect 41785 132016 41793 132050
rect 41827 132016 41835 132050
rect 41785 131992 41835 132016
rect 42121 132050 42171 132074
rect 42121 132016 42129 132050
rect 42163 132016 42171 132050
rect 42121 131992 42171 132016
rect 42457 132050 42507 132074
rect 42457 132016 42465 132050
rect 42499 132016 42507 132050
rect 42457 131992 42507 132016
rect 42793 132050 42843 132074
rect 42793 132016 42801 132050
rect 42835 132016 42843 132050
rect 42793 131992 42843 132016
rect 43129 132050 43179 132074
rect 43129 132016 43137 132050
rect 43171 132016 43179 132050
rect 43129 131992 43179 132016
rect 43465 132050 43515 132074
rect 43465 132016 43473 132050
rect 43507 132016 43515 132050
rect 43465 131992 43515 132016
rect 43801 132050 43851 132074
rect 43801 132016 43809 132050
rect 43843 132016 43851 132050
rect 43801 131992 43851 132016
rect 44137 132050 44187 132074
rect 44137 132016 44145 132050
rect 44179 132016 44187 132050
rect 44137 131992 44187 132016
rect 44473 132050 44523 132074
rect 44473 132016 44481 132050
rect 44515 132016 44523 132050
rect 44473 131992 44523 132016
rect 44809 132050 44859 132074
rect 44809 132016 44817 132050
rect 44851 132016 44859 132050
rect 44809 131992 44859 132016
rect 45145 132050 45195 132074
rect 45145 132016 45153 132050
rect 45187 132016 45195 132050
rect 45145 131992 45195 132016
rect 45481 132050 45531 132074
rect 45481 132016 45489 132050
rect 45523 132016 45531 132050
rect 45481 131992 45531 132016
rect 45817 132050 45867 132074
rect 45817 132016 45825 132050
rect 45859 132016 45867 132050
rect 45817 131992 45867 132016
rect 46153 132050 46203 132074
rect 46153 132016 46161 132050
rect 46195 132016 46203 132050
rect 46153 131992 46203 132016
rect 46489 132050 46539 132074
rect 46489 132016 46497 132050
rect 46531 132016 46539 132050
rect 46489 131992 46539 132016
rect 46825 132050 46875 132074
rect 46825 132016 46833 132050
rect 46867 132016 46875 132050
rect 46825 131992 46875 132016
rect 47161 132050 47211 132074
rect 47161 132016 47169 132050
rect 47203 132016 47211 132050
rect 47161 131992 47211 132016
rect 47497 132050 47547 132074
rect 47497 132016 47505 132050
rect 47539 132016 47547 132050
rect 47497 131992 47547 132016
rect 47833 132050 47883 132074
rect 47833 132016 47841 132050
rect 47875 132016 47883 132050
rect 47833 131992 47883 132016
rect 48169 132050 48219 132074
rect 48169 132016 48177 132050
rect 48211 132016 48219 132050
rect 48169 131992 48219 132016
rect 48505 132050 48555 132074
rect 48505 132016 48513 132050
rect 48547 132016 48555 132050
rect 48505 131992 48555 132016
rect 48841 132050 48891 132074
rect 48841 132016 48849 132050
rect 48883 132016 48891 132050
rect 48841 131992 48891 132016
rect 49177 132050 49227 132074
rect 49177 132016 49185 132050
rect 49219 132016 49227 132050
rect 49177 131992 49227 132016
rect 49513 132050 49563 132074
rect 49513 132016 49521 132050
rect 49555 132016 49563 132050
rect 49513 131992 49563 132016
rect 49849 132050 49899 132074
rect 49849 132016 49857 132050
rect 49891 132016 49899 132050
rect 49849 131992 49899 132016
rect 50185 132050 50235 132074
rect 50185 132016 50193 132050
rect 50227 132016 50235 132050
rect 50185 131992 50235 132016
rect 50521 132050 50571 132074
rect 50521 132016 50529 132050
rect 50563 132016 50571 132050
rect 50521 131992 50571 132016
rect 50857 132050 50907 132074
rect 50857 132016 50865 132050
rect 50899 132016 50907 132050
rect 50857 131992 50907 132016
rect 51193 132050 51243 132074
rect 51193 132016 51201 132050
rect 51235 132016 51243 132050
rect 51193 131992 51243 132016
rect 51529 132050 51579 132074
rect 51529 132016 51537 132050
rect 51571 132016 51579 132050
rect 51529 131992 51579 132016
rect 51865 132050 51915 132074
rect 51865 132016 51873 132050
rect 51907 132016 51915 132050
rect 51865 131992 51915 132016
rect 52201 132050 52251 132074
rect 52201 132016 52209 132050
rect 52243 132016 52251 132050
rect 52201 131992 52251 132016
rect 52537 132050 52587 132074
rect 52537 132016 52545 132050
rect 52579 132016 52587 132050
rect 52537 131992 52587 132016
rect 52873 132050 52923 132074
rect 52873 132016 52881 132050
rect 52915 132016 52923 132050
rect 52873 131992 52923 132016
rect 53209 132050 53259 132074
rect 53209 132016 53217 132050
rect 53251 132016 53259 132050
rect 53209 131992 53259 132016
rect 53545 132050 53595 132074
rect 53545 132016 53553 132050
rect 53587 132016 53595 132050
rect 53545 131992 53595 132016
rect 53881 132050 53931 132074
rect 53881 132016 53889 132050
rect 53923 132016 53931 132050
rect 53881 131992 53931 132016
rect 54217 132050 54267 132074
rect 54217 132016 54225 132050
rect 54259 132016 54267 132050
rect 54217 131992 54267 132016
rect 54553 132050 54603 132074
rect 54553 132016 54561 132050
rect 54595 132016 54603 132050
rect 54553 131992 54603 132016
rect 54889 132050 54939 132074
rect 54889 132016 54897 132050
rect 54931 132016 54939 132050
rect 54889 131992 54939 132016
rect 55225 132050 55275 132074
rect 55225 132016 55233 132050
rect 55267 132016 55275 132050
rect 55225 131992 55275 132016
rect 55561 132050 55611 132074
rect 55561 132016 55569 132050
rect 55603 132016 55611 132050
rect 55561 131992 55611 132016
rect 55897 132050 55947 132074
rect 55897 132016 55905 132050
rect 55939 132016 55947 132050
rect 55897 131992 55947 132016
rect 56233 132050 56283 132074
rect 56233 132016 56241 132050
rect 56275 132016 56283 132050
rect 56233 131992 56283 132016
rect 56569 132050 56619 132074
rect 56569 132016 56577 132050
rect 56611 132016 56619 132050
rect 56569 131992 56619 132016
rect 56905 132050 56955 132074
rect 56905 132016 56913 132050
rect 56947 132016 56955 132050
rect 56905 131992 56955 132016
rect 57241 132050 57291 132074
rect 57241 132016 57249 132050
rect 57283 132016 57291 132050
rect 57241 131992 57291 132016
rect 57577 132050 57627 132074
rect 57577 132016 57585 132050
rect 57619 132016 57627 132050
rect 57577 131992 57627 132016
rect 57913 132050 57963 132074
rect 57913 132016 57921 132050
rect 57955 132016 57963 132050
rect 57913 131992 57963 132016
rect 58249 132050 58299 132074
rect 58249 132016 58257 132050
rect 58291 132016 58299 132050
rect 58249 131992 58299 132016
rect 58585 132050 58635 132074
rect 58585 132016 58593 132050
rect 58627 132016 58635 132050
rect 58585 131992 58635 132016
rect 58921 132050 58971 132074
rect 58921 132016 58929 132050
rect 58963 132016 58971 132050
rect 58921 131992 58971 132016
rect 59257 132050 59307 132074
rect 59257 132016 59265 132050
rect 59299 132016 59307 132050
rect 59257 131992 59307 132016
rect 59593 132050 59643 132074
rect 59593 132016 59601 132050
rect 59635 132016 59643 132050
rect 59593 131992 59643 132016
rect 59929 132050 59979 132074
rect 59929 132016 59937 132050
rect 59971 132016 59979 132050
rect 59929 131992 59979 132016
rect 60265 132050 60315 132074
rect 60265 132016 60273 132050
rect 60307 132016 60315 132050
rect 60265 131992 60315 132016
rect 60601 132050 60651 132074
rect 60601 132016 60609 132050
rect 60643 132016 60651 132050
rect 60601 131992 60651 132016
rect 60937 132050 60987 132074
rect 60937 132016 60945 132050
rect 60979 132016 60987 132050
rect 60937 131992 60987 132016
rect 61273 132050 61323 132074
rect 61273 132016 61281 132050
rect 61315 132016 61323 132050
rect 61273 131992 61323 132016
rect 61609 132050 61659 132074
rect 61609 132016 61617 132050
rect 61651 132016 61659 132050
rect 61609 131992 61659 132016
rect 61945 132050 61995 132074
rect 61945 132016 61953 132050
rect 61987 132016 61995 132050
rect 61945 131992 61995 132016
rect 62281 132050 62331 132074
rect 62281 132016 62289 132050
rect 62323 132016 62331 132050
rect 62281 131992 62331 132016
rect 62617 132050 62667 132074
rect 62617 132016 62625 132050
rect 62659 132016 62667 132050
rect 62617 131992 62667 132016
rect 62953 132050 63003 132074
rect 62953 132016 62961 132050
rect 62995 132016 63003 132050
rect 62953 131992 63003 132016
rect 63289 132050 63339 132074
rect 63289 132016 63297 132050
rect 63331 132016 63339 132050
rect 63289 131992 63339 132016
rect 63625 132050 63675 132074
rect 63625 132016 63633 132050
rect 63667 132016 63675 132050
rect 63625 131992 63675 132016
rect 63961 132050 64011 132074
rect 63961 132016 63969 132050
rect 64003 132016 64011 132050
rect 63961 131992 64011 132016
rect 64297 132050 64347 132074
rect 64297 132016 64305 132050
rect 64339 132016 64347 132050
rect 64297 131992 64347 132016
rect 64633 132050 64683 132074
rect 64633 132016 64641 132050
rect 64675 132016 64683 132050
rect 64633 131992 64683 132016
rect 64969 132050 65019 132074
rect 64969 132016 64977 132050
rect 65011 132016 65019 132050
rect 64969 131992 65019 132016
rect 65305 132050 65355 132074
rect 65305 132016 65313 132050
rect 65347 132016 65355 132050
rect 65305 131992 65355 132016
rect 65641 132050 65691 132074
rect 65641 132016 65649 132050
rect 65683 132016 65691 132050
rect 65641 131992 65691 132016
rect 65977 132050 66027 132074
rect 65977 132016 65985 132050
rect 66019 132016 66027 132050
rect 65977 131992 66027 132016
rect 66313 132050 66363 132074
rect 66313 132016 66321 132050
rect 66355 132016 66363 132050
rect 66313 131992 66363 132016
rect 66649 132050 66699 132074
rect 66649 132016 66657 132050
rect 66691 132016 66699 132050
rect 66649 131992 66699 132016
rect 66985 132050 67035 132074
rect 66985 132016 66993 132050
rect 67027 132016 67035 132050
rect 66985 131992 67035 132016
rect 67321 132050 67371 132074
rect 67321 132016 67329 132050
rect 67363 132016 67371 132050
rect 67321 131992 67371 132016
rect 67657 132050 67707 132074
rect 67657 132016 67665 132050
rect 67699 132016 67707 132050
rect 67657 131992 67707 132016
rect 67993 132050 68043 132074
rect 67993 132016 68001 132050
rect 68035 132016 68043 132050
rect 67993 131992 68043 132016
rect 68329 132050 68379 132074
rect 68329 132016 68337 132050
rect 68371 132016 68379 132050
rect 68329 131992 68379 132016
rect 68665 132050 68715 132074
rect 68665 132016 68673 132050
rect 68707 132016 68715 132050
rect 68665 131992 68715 132016
rect 69001 132050 69051 132074
rect 69001 132016 69009 132050
rect 69043 132016 69051 132050
rect 69001 131992 69051 132016
rect 69337 132050 69387 132074
rect 69337 132016 69345 132050
rect 69379 132016 69387 132050
rect 69337 131992 69387 132016
rect 69673 132050 69723 132074
rect 69673 132016 69681 132050
rect 69715 132016 69723 132050
rect 69673 131992 69723 132016
rect 70009 132050 70059 132074
rect 70009 132016 70017 132050
rect 70051 132016 70059 132050
rect 70009 131992 70059 132016
rect 70345 132050 70395 132074
rect 70345 132016 70353 132050
rect 70387 132016 70395 132050
rect 70345 131992 70395 132016
rect 70681 132050 70731 132074
rect 70681 132016 70689 132050
rect 70723 132016 70731 132050
rect 70681 131992 70731 132016
rect 71017 132050 71067 132074
rect 71017 132016 71025 132050
rect 71059 132016 71067 132050
rect 71017 131992 71067 132016
rect 71353 132050 71403 132074
rect 71353 132016 71361 132050
rect 71395 132016 71403 132050
rect 71353 131992 71403 132016
rect 71689 132050 71739 132074
rect 71689 132016 71697 132050
rect 71731 132016 71739 132050
rect 71689 131992 71739 132016
rect 72025 132050 72075 132074
rect 72025 132016 72033 132050
rect 72067 132016 72075 132050
rect 72025 131992 72075 132016
rect 72361 132050 72411 132074
rect 72361 132016 72369 132050
rect 72403 132016 72411 132050
rect 72361 131992 72411 132016
rect 72697 132050 72747 132074
rect 72697 132016 72705 132050
rect 72739 132016 72747 132050
rect 72697 131992 72747 132016
rect 73033 132050 73083 132074
rect 73033 132016 73041 132050
rect 73075 132016 73083 132050
rect 73033 131992 73083 132016
rect 73369 132050 73419 132074
rect 73369 132016 73377 132050
rect 73411 132016 73419 132050
rect 73369 131992 73419 132016
rect 73705 132050 73755 132074
rect 73705 132016 73713 132050
rect 73747 132016 73755 132050
rect 73705 131992 73755 132016
rect 74041 132050 74091 132074
rect 74041 132016 74049 132050
rect 74083 132016 74091 132050
rect 74041 131992 74091 132016
rect 74377 132050 74427 132074
rect 74377 132016 74385 132050
rect 74419 132016 74427 132050
rect 74377 131992 74427 132016
rect 74713 132050 74763 132074
rect 74713 132016 74721 132050
rect 74755 132016 74763 132050
rect 74713 131992 74763 132016
rect 75049 132050 75099 132074
rect 75049 132016 75057 132050
rect 75091 132016 75099 132050
rect 75049 131992 75099 132016
rect 75385 132050 75435 132074
rect 75385 132016 75393 132050
rect 75427 132016 75435 132050
rect 75385 131992 75435 132016
rect 75721 132050 75771 132074
rect 75721 132016 75729 132050
rect 75763 132016 75771 132050
rect 75721 131992 75771 132016
rect 76057 132050 76107 132074
rect 76057 132016 76065 132050
rect 76099 132016 76107 132050
rect 76057 131992 76107 132016
rect 76393 132050 76443 132074
rect 76393 132016 76401 132050
rect 76435 132016 76443 132050
rect 76393 131992 76443 132016
rect 76729 132050 76779 132074
rect 76729 132016 76737 132050
rect 76771 132016 76779 132050
rect 76729 131992 76779 132016
rect 77065 132050 77115 132074
rect 77065 132016 77073 132050
rect 77107 132016 77115 132050
rect 77065 131992 77115 132016
rect 77401 132050 77451 132074
rect 77401 132016 77409 132050
rect 77443 132016 77451 132050
rect 77401 131992 77451 132016
rect 77737 132050 77787 132074
rect 77737 132016 77745 132050
rect 77779 132016 77787 132050
rect 77737 131992 77787 132016
rect 78073 132050 78123 132074
rect 78073 132016 78081 132050
rect 78115 132016 78123 132050
rect 78073 131992 78123 132016
rect 78409 132050 78459 132074
rect 78409 132016 78417 132050
rect 78451 132016 78459 132050
rect 78409 131992 78459 132016
rect 78745 132050 78795 132074
rect 78745 132016 78753 132050
rect 78787 132016 78795 132050
rect 78745 131992 78795 132016
rect 79081 132050 79131 132074
rect 79081 132016 79089 132050
rect 79123 132016 79131 132050
rect 79081 131992 79131 132016
rect 79417 132050 79467 132074
rect 79417 132016 79425 132050
rect 79459 132016 79467 132050
rect 79417 131992 79467 132016
rect 79753 132050 79803 132074
rect 79753 132016 79761 132050
rect 79795 132016 79803 132050
rect 79753 131992 79803 132016
rect 80089 132050 80139 132074
rect 80089 132016 80097 132050
rect 80131 132016 80139 132050
rect 80089 131992 80139 132016
rect 80425 132050 80475 132074
rect 80425 132016 80433 132050
rect 80467 132016 80475 132050
rect 80425 131992 80475 132016
rect 80761 132050 80811 132074
rect 80761 132016 80769 132050
rect 80803 132016 80811 132050
rect 80761 131992 80811 132016
rect 81097 132050 81147 132074
rect 81097 132016 81105 132050
rect 81139 132016 81147 132050
rect 81097 131992 81147 132016
rect 81433 132050 81483 132074
rect 81433 132016 81441 132050
rect 81475 132016 81483 132050
rect 81433 131992 81483 132016
rect 81769 132050 81819 132074
rect 81769 132016 81777 132050
rect 81811 132016 81819 132050
rect 81769 131992 81819 132016
rect 82105 132050 82155 132074
rect 82105 132016 82113 132050
rect 82147 132016 82155 132050
rect 82105 131992 82155 132016
rect 82441 132050 82491 132074
rect 82441 132016 82449 132050
rect 82483 132016 82491 132050
rect 82441 131992 82491 132016
rect 82777 132050 82827 132074
rect 82777 132016 82785 132050
rect 82819 132016 82827 132050
rect 82777 131992 82827 132016
rect 83113 132050 83163 132074
rect 83113 132016 83121 132050
rect 83155 132016 83163 132050
rect 83113 131992 83163 132016
rect 83449 132050 83499 132074
rect 83449 132016 83457 132050
rect 83491 132016 83499 132050
rect 83449 131992 83499 132016
rect 83785 132050 83835 132074
rect 83785 132016 83793 132050
rect 83827 132016 83835 132050
rect 83785 131992 83835 132016
rect 84121 132050 84171 132074
rect 84121 132016 84129 132050
rect 84163 132016 84171 132050
rect 84121 131992 84171 132016
rect 84457 132050 84507 132074
rect 84457 132016 84465 132050
rect 84499 132016 84507 132050
rect 84457 131992 84507 132016
rect 84793 132050 84843 132074
rect 84793 132016 84801 132050
rect 84835 132016 84843 132050
rect 84793 131992 84843 132016
rect 85129 132050 85179 132074
rect 85129 132016 85137 132050
rect 85171 132016 85179 132050
rect 85129 131992 85179 132016
rect 85465 132050 85515 132074
rect 85465 132016 85473 132050
rect 85507 132016 85515 132050
rect 85465 131992 85515 132016
rect 85801 132050 85851 132074
rect 85801 132016 85809 132050
rect 85843 132016 85851 132050
rect 85801 131992 85851 132016
rect 86137 132050 86187 132074
rect 86137 132016 86145 132050
rect 86179 132016 86187 132050
rect 86137 131992 86187 132016
rect 86473 132050 86523 132074
rect 86473 132016 86481 132050
rect 86515 132016 86523 132050
rect 86473 131992 86523 132016
rect 86809 132050 86859 132074
rect 86809 132016 86817 132050
rect 86851 132016 86859 132050
rect 86809 131992 86859 132016
rect 87145 132050 87195 132074
rect 87145 132016 87153 132050
rect 87187 132016 87195 132050
rect 87145 131992 87195 132016
rect 87481 132050 87531 132074
rect 87481 132016 87489 132050
rect 87523 132016 87531 132050
rect 87481 131992 87531 132016
rect 87817 132050 87867 132074
rect 87817 132016 87825 132050
rect 87859 132016 87867 132050
rect 87817 131992 87867 132016
rect 88153 132050 88203 132074
rect 88153 132016 88161 132050
rect 88195 132016 88203 132050
rect 88153 131992 88203 132016
rect 88489 132050 88539 132074
rect 88489 132016 88497 132050
rect 88531 132016 88539 132050
rect 88489 131992 88539 132016
rect 88825 132050 88875 132074
rect 88825 132016 88833 132050
rect 88867 132016 88875 132050
rect 88825 131992 88875 132016
rect 89161 132050 89211 132074
rect 89161 132016 89169 132050
rect 89203 132016 89211 132050
rect 89161 131992 89211 132016
rect 89497 132050 89547 132074
rect 89497 132016 89505 132050
rect 89539 132016 89547 132050
rect 89497 131992 89547 132016
rect 89833 132050 89883 132074
rect 89833 132016 89841 132050
rect 89875 132016 89883 132050
rect 89833 131992 89883 132016
rect 90169 132050 90219 132074
rect 90169 132016 90177 132050
rect 90211 132016 90219 132050
rect 90169 131992 90219 132016
rect 90505 132050 90555 132074
rect 90505 132016 90513 132050
rect 90547 132016 90555 132050
rect 90505 131992 90555 132016
rect 90841 132050 90891 132074
rect 90841 132016 90849 132050
rect 90883 132016 90891 132050
rect 90841 131992 90891 132016
rect 91177 132050 91227 132074
rect 91177 132016 91185 132050
rect 91219 132016 91227 132050
rect 91177 131992 91227 132016
rect 91513 132050 91563 132074
rect 91513 132016 91521 132050
rect 91555 132016 91563 132050
rect 91513 131992 91563 132016
rect 91849 132050 91899 132074
rect 91849 132016 91857 132050
rect 91891 132016 91899 132050
rect 91849 131992 91899 132016
rect 92185 132050 92235 132074
rect 92185 132016 92193 132050
rect 92227 132016 92235 132050
rect 92185 131992 92235 132016
rect 92521 132050 92571 132074
rect 92521 132016 92529 132050
rect 92563 132016 92571 132050
rect 92521 131992 92571 132016
rect 92857 132050 92907 132074
rect 92857 132016 92865 132050
rect 92899 132016 92907 132050
rect 92857 131992 92907 132016
rect 93193 132050 93243 132074
rect 93193 132016 93201 132050
rect 93235 132016 93243 132050
rect 93193 131992 93243 132016
rect 93529 132050 93579 132074
rect 93529 132016 93537 132050
rect 93571 132016 93579 132050
rect 93529 131992 93579 132016
rect 93865 132050 93915 132074
rect 93865 132016 93873 132050
rect 93907 132016 93915 132050
rect 93865 131992 93915 132016
rect 94201 132050 94251 132074
rect 94201 132016 94209 132050
rect 94243 132016 94251 132050
rect 94201 131992 94251 132016
rect 94537 132050 94587 132074
rect 94537 132016 94545 132050
rect 94579 132016 94587 132050
rect 94537 131992 94587 132016
rect 94873 132050 94923 132074
rect 94873 132016 94881 132050
rect 94915 132016 94923 132050
rect 94873 131992 94923 132016
rect 95209 132050 95259 132074
rect 95209 132016 95217 132050
rect 95251 132016 95259 132050
rect 95209 131992 95259 132016
rect 95545 132050 95595 132074
rect 95545 132016 95553 132050
rect 95587 132016 95595 132050
rect 95545 131992 95595 132016
rect 95881 132050 95931 132074
rect 95881 132016 95889 132050
rect 95923 132016 95931 132050
rect 95881 131992 95931 132016
rect 96217 132050 96267 132074
rect 96217 132016 96225 132050
rect 96259 132016 96267 132050
rect 96217 131992 96267 132016
rect 96553 132050 96603 132074
rect 96553 132016 96561 132050
rect 96595 132016 96603 132050
rect 96553 131992 96603 132016
rect 96889 132050 96939 132074
rect 96889 132016 96897 132050
rect 96931 132016 96939 132050
rect 96889 131992 96939 132016
rect 97225 132050 97275 132074
rect 97225 132016 97233 132050
rect 97267 132016 97275 132050
rect 97225 131992 97275 132016
rect 97561 132050 97611 132074
rect 97561 132016 97569 132050
rect 97603 132016 97611 132050
rect 97561 131992 97611 132016
rect 97897 132050 97947 132074
rect 97897 132016 97905 132050
rect 97939 132016 97947 132050
rect 97897 131992 97947 132016
rect 98233 132050 98283 132074
rect 98233 132016 98241 132050
rect 98275 132016 98283 132050
rect 98233 131992 98283 132016
rect 98569 132050 98619 132074
rect 98569 132016 98577 132050
rect 98611 132016 98619 132050
rect 98569 131992 98619 132016
rect 98905 132050 98955 132074
rect 98905 132016 98913 132050
rect 98947 132016 98955 132050
rect 98905 131992 98955 132016
rect 99241 132050 99291 132074
rect 99241 132016 99249 132050
rect 99283 132016 99291 132050
rect 99241 131992 99291 132016
rect 99577 132050 99627 132074
rect 99577 132016 99585 132050
rect 99619 132016 99627 132050
rect 99577 131992 99627 132016
rect 99913 132050 99963 132074
rect 99913 132016 99921 132050
rect 99955 132016 99963 132050
rect 99913 131992 99963 132016
rect 100249 132050 100299 132074
rect 100249 132016 100257 132050
rect 100291 132016 100299 132050
rect 100249 131992 100299 132016
rect 100585 132050 100635 132074
rect 100585 132016 100593 132050
rect 100627 132016 100635 132050
rect 100585 131992 100635 132016
rect 100921 132050 100971 132074
rect 100921 132016 100929 132050
rect 100963 132016 100971 132050
rect 100921 131992 100971 132016
rect 101257 132050 101307 132074
rect 101257 132016 101265 132050
rect 101299 132016 101307 132050
rect 101257 131992 101307 132016
rect 101593 132050 101643 132074
rect 101593 132016 101601 132050
rect 101635 132016 101643 132050
rect 101593 131992 101643 132016
rect 101929 132050 101979 132074
rect 101929 132016 101937 132050
rect 101971 132016 101979 132050
rect 101929 131992 101979 132016
rect 102265 132050 102315 132074
rect 102265 132016 102273 132050
rect 102307 132016 102315 132050
rect 102265 131992 102315 132016
rect 102601 132050 102651 132074
rect 102601 132016 102609 132050
rect 102643 132016 102651 132050
rect 102601 131992 102651 132016
rect 102937 132050 102987 132074
rect 102937 132016 102945 132050
rect 102979 132016 102987 132050
rect 102937 131992 102987 132016
rect 103273 132050 103323 132074
rect 103273 132016 103281 132050
rect 103315 132016 103323 132050
rect 103273 131992 103323 132016
rect 103609 132050 103659 132074
rect 103609 132016 103617 132050
rect 103651 132016 103659 132050
rect 103609 131992 103659 132016
rect 103945 132050 103995 132074
rect 103945 132016 103953 132050
rect 103987 132016 103995 132050
rect 103945 131992 103995 132016
rect 104281 132050 104331 132074
rect 104281 132016 104289 132050
rect 104323 132016 104331 132050
rect 104281 131992 104331 132016
rect 104617 132050 104667 132074
rect 104617 132016 104625 132050
rect 104659 132016 104667 132050
rect 104617 131992 104667 132016
rect 104953 132050 105003 132074
rect 104953 132016 104961 132050
rect 104995 132016 105003 132050
rect 104953 131992 105003 132016
rect 105289 132050 105339 132074
rect 105289 132016 105297 132050
rect 105331 132016 105339 132050
rect 105289 131992 105339 132016
rect 105625 132050 105675 132074
rect 105625 132016 105633 132050
rect 105667 132016 105675 132050
rect 105625 131992 105675 132016
rect 105961 132050 106011 132074
rect 105961 132016 105969 132050
rect 106003 132016 106011 132050
rect 105961 131992 106011 132016
rect 106297 132050 106347 132074
rect 106297 132016 106305 132050
rect 106339 132016 106347 132050
rect 106297 131992 106347 132016
rect 106633 132050 106683 132074
rect 106633 132016 106641 132050
rect 106675 132016 106683 132050
rect 106633 131992 106683 132016
rect 106969 132050 107019 132074
rect 106969 132016 106977 132050
rect 107011 132016 107019 132050
rect 106969 131992 107019 132016
rect 107305 132050 107355 132074
rect 107305 132016 107313 132050
rect 107347 132016 107355 132050
rect 107305 131992 107355 132016
rect 107641 132050 107691 132074
rect 107641 132016 107649 132050
rect 107683 132016 107691 132050
rect 107641 131992 107691 132016
rect 107977 132050 108027 132074
rect 107977 132016 107985 132050
rect 108019 132016 108027 132050
rect 107977 131992 108027 132016
rect 108313 132050 108363 132074
rect 108313 132016 108321 132050
rect 108355 132016 108363 132050
rect 108313 131992 108363 132016
rect 108649 132050 108699 132074
rect 108649 132016 108657 132050
rect 108691 132016 108699 132050
rect 108649 131992 108699 132016
rect 108985 132050 109035 132074
rect 108985 132016 108993 132050
rect 109027 132016 109035 132050
rect 108985 131992 109035 132016
rect 109321 132050 109371 132074
rect 109321 132016 109329 132050
rect 109363 132016 109371 132050
rect 109321 131992 109371 132016
rect 109657 132050 109707 132074
rect 109657 132016 109665 132050
rect 109699 132016 109707 132050
rect 109657 131992 109707 132016
rect 109993 132050 110043 132074
rect 109993 132016 110001 132050
rect 110035 132016 110043 132050
rect 109993 131992 110043 132016
rect 110329 132050 110379 132074
rect 110329 132016 110337 132050
rect 110371 132016 110379 132050
rect 110329 131992 110379 132016
rect 110665 132050 110715 132074
rect 110665 132016 110673 132050
rect 110707 132016 110715 132050
rect 110665 131992 110715 132016
rect 111001 132050 111051 132074
rect 111001 132016 111009 132050
rect 111043 132016 111051 132050
rect 111001 131992 111051 132016
rect 111337 132050 111387 132074
rect 111337 132016 111345 132050
rect 111379 132016 111387 132050
rect 111337 131992 111387 132016
rect 111673 132050 111723 132074
rect 111673 132016 111681 132050
rect 111715 132016 111723 132050
rect 111673 131992 111723 132016
rect 112009 132050 112059 132074
rect 112009 132016 112017 132050
rect 112051 132016 112059 132050
rect 112009 131992 112059 132016
rect 112345 132050 112395 132074
rect 112345 132016 112353 132050
rect 112387 132016 112395 132050
rect 112345 131992 112395 132016
rect 112681 132050 112731 132074
rect 112681 132016 112689 132050
rect 112723 132016 112731 132050
rect 112681 131992 112731 132016
rect 113017 132050 113067 132074
rect 113017 132016 113025 132050
rect 113059 132016 113067 132050
rect 113017 131992 113067 132016
rect 113353 132050 113403 132074
rect 113353 132016 113361 132050
rect 113395 132016 113403 132050
rect 113353 131992 113403 132016
rect 113689 132050 113739 132074
rect 113689 132016 113697 132050
rect 113731 132016 113739 132050
rect 113689 131992 113739 132016
rect 114025 132050 114075 132074
rect 114025 132016 114033 132050
rect 114067 132016 114075 132050
rect 114025 131992 114075 132016
rect 114361 132050 114411 132074
rect 114361 132016 114369 132050
rect 114403 132016 114411 132050
rect 114361 131992 114411 132016
rect 114697 132050 114747 132074
rect 114697 132016 114705 132050
rect 114739 132016 114747 132050
rect 114697 131992 114747 132016
rect 115033 132050 115083 132074
rect 115033 132016 115041 132050
rect 115075 132016 115083 132050
rect 115033 131992 115083 132016
rect 115369 132050 115419 132074
rect 115369 132016 115377 132050
rect 115411 132016 115419 132050
rect 115369 131992 115419 132016
rect 115705 132050 115755 132074
rect 115705 132016 115713 132050
rect 115747 132016 115755 132050
rect 115705 131992 115755 132016
rect 116041 132050 116091 132074
rect 116041 132016 116049 132050
rect 116083 132016 116091 132050
rect 116041 131992 116091 132016
rect 116377 132050 116427 132074
rect 116377 132016 116385 132050
rect 116419 132016 116427 132050
rect 116377 131992 116427 132016
rect 116713 132050 116763 132074
rect 116713 132016 116721 132050
rect 116755 132016 116763 132050
rect 116713 131992 116763 132016
rect 117049 132050 117099 132074
rect 117049 132016 117057 132050
rect 117091 132016 117099 132050
rect 117049 131992 117099 132016
rect 117385 132050 117435 132074
rect 117385 132016 117393 132050
rect 117427 132016 117435 132050
rect 117385 131992 117435 132016
rect 117721 132050 117771 132074
rect 117721 132016 117729 132050
rect 117763 132016 117771 132050
rect 117721 131992 117771 132016
rect 118057 132050 118107 132074
rect 118057 132016 118065 132050
rect 118099 132016 118107 132050
rect 118057 131992 118107 132016
rect 118393 132050 118443 132074
rect 118393 132016 118401 132050
rect 118435 132016 118443 132050
rect 118393 131992 118443 132016
rect 118729 132050 118779 132074
rect 118729 132016 118737 132050
rect 118771 132016 118779 132050
rect 118729 131992 118779 132016
rect 119065 132050 119115 132074
rect 119065 132016 119073 132050
rect 119107 132016 119115 132050
rect 119065 131992 119115 132016
rect 119401 132050 119451 132074
rect 119401 132016 119409 132050
rect 119443 132016 119451 132050
rect 119401 131992 119451 132016
rect 119737 132050 119787 132074
rect 119737 132016 119745 132050
rect 119779 132016 119787 132050
rect 119737 131992 119787 132016
rect 120073 132050 120123 132074
rect 120073 132016 120081 132050
rect 120115 132016 120123 132050
rect 120073 131992 120123 132016
rect 120409 132050 120459 132074
rect 120409 132016 120417 132050
rect 120451 132016 120459 132050
rect 120409 131992 120459 132016
rect 120745 132050 120795 132074
rect 120745 132016 120753 132050
rect 120787 132016 120795 132050
rect 120745 131992 120795 132016
rect 121081 132050 121131 132074
rect 121081 132016 121089 132050
rect 121123 132016 121131 132050
rect 121081 131992 121131 132016
rect 121417 132050 121467 132074
rect 121417 132016 121425 132050
rect 121459 132016 121467 132050
rect 121417 131992 121467 132016
rect 121753 132050 121803 132074
rect 121753 132016 121761 132050
rect 121795 132016 121803 132050
rect 121753 131992 121803 132016
rect 122089 132050 122139 132074
rect 122089 132016 122097 132050
rect 122131 132016 122139 132050
rect 122089 131992 122139 132016
rect 122425 132050 122475 132074
rect 122425 132016 122433 132050
rect 122467 132016 122475 132050
rect 122425 131992 122475 132016
rect 122761 132050 122811 132074
rect 122761 132016 122769 132050
rect 122803 132016 122811 132050
rect 122761 131992 122811 132016
rect 123097 132050 123147 132074
rect 123097 132016 123105 132050
rect 123139 132016 123147 132050
rect 123097 131992 123147 132016
rect 123433 132050 123483 132074
rect 123433 132016 123441 132050
rect 123475 132016 123483 132050
rect 123433 131992 123483 132016
rect 123769 132050 123819 132074
rect 123769 132016 123777 132050
rect 123811 132016 123819 132050
rect 123769 131992 123819 132016
rect 124105 132050 124155 132074
rect 124105 132016 124113 132050
rect 124147 132016 124155 132050
rect 124105 131992 124155 132016
rect 124441 132050 124491 132074
rect 124441 132016 124449 132050
rect 124483 132016 124491 132050
rect 124441 131992 124491 132016
rect 124777 132050 124827 132074
rect 124777 132016 124785 132050
rect 124819 132016 124827 132050
rect 124777 131992 124827 132016
rect 125113 132050 125163 132074
rect 125113 132016 125121 132050
rect 125155 132016 125163 132050
rect 125113 131992 125163 132016
rect 125449 132050 125499 132074
rect 125449 132016 125457 132050
rect 125491 132016 125499 132050
rect 125449 131992 125499 132016
rect 125785 132050 125835 132074
rect 125785 132016 125793 132050
rect 125827 132016 125835 132050
rect 125785 131992 125835 132016
rect 126121 132050 126171 132074
rect 126121 132016 126129 132050
rect 126163 132016 126171 132050
rect 126121 131992 126171 132016
rect 126457 132050 126507 132074
rect 126457 132016 126465 132050
rect 126499 132016 126507 132050
rect 126457 131992 126507 132016
rect 126793 132050 126843 132074
rect 126793 132016 126801 132050
rect 126835 132016 126843 132050
rect 126793 131992 126843 132016
rect 127129 132050 127179 132074
rect 127129 132016 127137 132050
rect 127171 132016 127179 132050
rect 127129 131992 127179 132016
rect 127465 132050 127515 132074
rect 127465 132016 127473 132050
rect 127507 132016 127515 132050
rect 127465 131992 127515 132016
rect 127801 132050 127851 132074
rect 127801 132016 127809 132050
rect 127843 132016 127851 132050
rect 127801 131992 127851 132016
rect 128137 132050 128187 132074
rect 128137 132016 128145 132050
rect 128179 132016 128187 132050
rect 128137 131992 128187 132016
rect 128473 132050 128523 132074
rect 128473 132016 128481 132050
rect 128515 132016 128523 132050
rect 128473 131992 128523 132016
rect 128809 132050 128859 132074
rect 128809 132016 128817 132050
rect 128851 132016 128859 132050
rect 128809 131992 128859 132016
rect 129145 132050 129195 132074
rect 129145 132016 129153 132050
rect 129187 132016 129195 132050
rect 129145 131992 129195 132016
rect 129481 132050 129531 132074
rect 129481 132016 129489 132050
rect 129523 132016 129531 132050
rect 129481 131992 129531 132016
rect 129817 132050 129867 132074
rect 129817 132016 129825 132050
rect 129859 132016 129867 132050
rect 129817 131992 129867 132016
rect 130153 132050 130203 132074
rect 130153 132016 130161 132050
rect 130195 132016 130203 132050
rect 130153 131992 130203 132016
rect 130489 132050 130539 132074
rect 130489 132016 130497 132050
rect 130531 132016 130539 132050
rect 130489 131992 130539 132016
rect 130825 132050 130875 132074
rect 130825 132016 130833 132050
rect 130867 132016 130875 132050
rect 130825 131992 130875 132016
rect 131161 132050 131211 132074
rect 131161 132016 131169 132050
rect 131203 132016 131211 132050
rect 131161 131992 131211 132016
rect 131497 132050 131547 132074
rect 131497 132016 131505 132050
rect 131539 132016 131547 132050
rect 131497 131992 131547 132016
rect 131833 132050 131883 132074
rect 131833 132016 131841 132050
rect 131875 132016 131883 132050
rect 131833 131992 131883 132016
rect 132169 132050 132219 132074
rect 132169 132016 132177 132050
rect 132211 132016 132219 132050
rect 132169 131992 132219 132016
rect 132505 132050 132555 132074
rect 132505 132016 132513 132050
rect 132547 132016 132555 132050
rect 132505 131992 132555 132016
rect 132841 132050 132891 132074
rect 132841 132016 132849 132050
rect 132883 132016 132891 132050
rect 132841 131992 132891 132016
rect 133177 132050 133227 132074
rect 133177 132016 133185 132050
rect 133219 132016 133227 132050
rect 133177 131992 133227 132016
rect 133513 132050 133563 132074
rect 133513 132016 133521 132050
rect 133555 132016 133563 132050
rect 133513 131992 133563 132016
rect 133849 132050 133899 132074
rect 133849 132016 133857 132050
rect 133891 132016 133899 132050
rect 133849 131992 133899 132016
rect 134185 132050 134235 132074
rect 134185 132016 134193 132050
rect 134227 132016 134235 132050
rect 134185 131992 134235 132016
rect 134521 132050 134571 132074
rect 134521 132016 134529 132050
rect 134563 132016 134571 132050
rect 134521 131992 134571 132016
rect 134857 132050 134907 132074
rect 134857 132016 134865 132050
rect 134899 132016 134907 132050
rect 134857 131992 134907 132016
rect 135193 132050 135243 132074
rect 135193 132016 135201 132050
rect 135235 132016 135243 132050
rect 135193 131992 135243 132016
rect 135529 132050 135579 132074
rect 135529 132016 135537 132050
rect 135571 132016 135579 132050
rect 135529 131992 135579 132016
rect 135865 132050 135915 132074
rect 135865 132016 135873 132050
rect 135907 132016 135915 132050
rect 135865 131992 135915 132016
rect 136201 132050 136251 132074
rect 136201 132016 136209 132050
rect 136243 132016 136251 132050
rect 136201 131992 136251 132016
rect 136537 132050 136587 132074
rect 136537 132016 136545 132050
rect 136579 132016 136587 132050
rect 136537 131992 136587 132016
rect 1801 131437 1851 131461
rect 1801 131403 1809 131437
rect 1843 131403 1851 131437
rect 1801 131379 1851 131403
rect 136947 131437 136997 131461
rect 136947 131403 136955 131437
rect 136989 131403 136997 131437
rect 136947 131379 136997 131403
rect 1801 131101 1851 131125
rect 1801 131067 1809 131101
rect 1843 131067 1851 131101
rect 1801 131043 1851 131067
rect 136947 131101 136997 131125
rect 136947 131067 136955 131101
rect 136989 131067 136997 131101
rect 136947 131043 136997 131067
rect 1801 130765 1851 130789
rect 1801 130731 1809 130765
rect 1843 130731 1851 130765
rect 1801 130707 1851 130731
rect 136947 130765 136997 130789
rect 136947 130731 136955 130765
rect 136989 130731 136997 130765
rect 136947 130707 136997 130731
rect 1801 130429 1851 130453
rect 1801 130395 1809 130429
rect 1843 130395 1851 130429
rect 1801 130371 1851 130395
rect 136947 130429 136997 130453
rect 136947 130395 136955 130429
rect 136989 130395 136997 130429
rect 136947 130371 136997 130395
rect 1801 130093 1851 130117
rect 1801 130059 1809 130093
rect 1843 130059 1851 130093
rect 1801 130035 1851 130059
rect 136947 130093 136997 130117
rect 136947 130059 136955 130093
rect 136989 130059 136997 130093
rect 136947 130035 136997 130059
rect 1801 129757 1851 129781
rect 1801 129723 1809 129757
rect 1843 129723 1851 129757
rect 1801 129699 1851 129723
rect 136947 129757 136997 129781
rect 136947 129723 136955 129757
rect 136989 129723 136997 129757
rect 136947 129699 136997 129723
rect 1801 129421 1851 129445
rect 1801 129387 1809 129421
rect 1843 129387 1851 129421
rect 1801 129363 1851 129387
rect 136947 129421 136997 129445
rect 136947 129387 136955 129421
rect 136989 129387 136997 129421
rect 136947 129363 136997 129387
rect 1801 129085 1851 129109
rect 1801 129051 1809 129085
rect 1843 129051 1851 129085
rect 1801 129027 1851 129051
rect 136947 129085 136997 129109
rect 136947 129051 136955 129085
rect 136989 129051 136997 129085
rect 136947 129027 136997 129051
rect 1801 128749 1851 128773
rect 1801 128715 1809 128749
rect 1843 128715 1851 128749
rect 1801 128691 1851 128715
rect 136947 128749 136997 128773
rect 136947 128715 136955 128749
rect 136989 128715 136997 128749
rect 136947 128691 136997 128715
rect 1801 128413 1851 128437
rect 1801 128379 1809 128413
rect 1843 128379 1851 128413
rect 1801 128355 1851 128379
rect 136947 128413 136997 128437
rect 136947 128379 136955 128413
rect 136989 128379 136997 128413
rect 136947 128355 136997 128379
rect 1801 128077 1851 128101
rect 1801 128043 1809 128077
rect 1843 128043 1851 128077
rect 1801 128019 1851 128043
rect 136947 128077 136997 128101
rect 136947 128043 136955 128077
rect 136989 128043 136997 128077
rect 136947 128019 136997 128043
rect 1801 127741 1851 127765
rect 1801 127707 1809 127741
rect 1843 127707 1851 127741
rect 1801 127683 1851 127707
rect 136947 127741 136997 127765
rect 136947 127707 136955 127741
rect 136989 127707 136997 127741
rect 136947 127683 136997 127707
rect 1801 127405 1851 127429
rect 1801 127371 1809 127405
rect 1843 127371 1851 127405
rect 1801 127347 1851 127371
rect 136947 127405 136997 127429
rect 136947 127371 136955 127405
rect 136989 127371 136997 127405
rect 136947 127347 136997 127371
rect 1801 127069 1851 127093
rect 1801 127035 1809 127069
rect 1843 127035 1851 127069
rect 1801 127011 1851 127035
rect 136947 127069 136997 127093
rect 136947 127035 136955 127069
rect 136989 127035 136997 127069
rect 136947 127011 136997 127035
rect 1801 126733 1851 126757
rect 1801 126699 1809 126733
rect 1843 126699 1851 126733
rect 1801 126675 1851 126699
rect 136947 126733 136997 126757
rect 136947 126699 136955 126733
rect 136989 126699 136997 126733
rect 136947 126675 136997 126699
rect 1801 126397 1851 126421
rect 1801 126363 1809 126397
rect 1843 126363 1851 126397
rect 1801 126339 1851 126363
rect 136947 126397 136997 126421
rect 136947 126363 136955 126397
rect 136989 126363 136997 126397
rect 136947 126339 136997 126363
rect 1801 126061 1851 126085
rect 1801 126027 1809 126061
rect 1843 126027 1851 126061
rect 1801 126003 1851 126027
rect 136947 126061 136997 126085
rect 136947 126027 136955 126061
rect 136989 126027 136997 126061
rect 136947 126003 136997 126027
rect 1801 125725 1851 125749
rect 1801 125691 1809 125725
rect 1843 125691 1851 125725
rect 1801 125667 1851 125691
rect 136947 125725 136997 125749
rect 136947 125691 136955 125725
rect 136989 125691 136997 125725
rect 136947 125667 136997 125691
rect 1801 125389 1851 125413
rect 1801 125355 1809 125389
rect 1843 125355 1851 125389
rect 1801 125331 1851 125355
rect 136947 125389 136997 125413
rect 136947 125355 136955 125389
rect 136989 125355 136997 125389
rect 136947 125331 136997 125355
rect 1801 125053 1851 125077
rect 1801 125019 1809 125053
rect 1843 125019 1851 125053
rect 1801 124995 1851 125019
rect 136947 125053 136997 125077
rect 136947 125019 136955 125053
rect 136989 125019 136997 125053
rect 136947 124995 136997 125019
rect 1801 124717 1851 124741
rect 1801 124683 1809 124717
rect 1843 124683 1851 124717
rect 1801 124659 1851 124683
rect 136947 124717 136997 124741
rect 136947 124683 136955 124717
rect 136989 124683 136997 124717
rect 136947 124659 136997 124683
rect 1801 124381 1851 124405
rect 1801 124347 1809 124381
rect 1843 124347 1851 124381
rect 1801 124323 1851 124347
rect 136947 124381 136997 124405
rect 136947 124347 136955 124381
rect 136989 124347 136997 124381
rect 136947 124323 136997 124347
rect 1801 124045 1851 124069
rect 1801 124011 1809 124045
rect 1843 124011 1851 124045
rect 1801 123987 1851 124011
rect 136947 124045 136997 124069
rect 136947 124011 136955 124045
rect 136989 124011 136997 124045
rect 136947 123987 136997 124011
rect 1801 123709 1851 123733
rect 1801 123675 1809 123709
rect 1843 123675 1851 123709
rect 1801 123651 1851 123675
rect 136947 123709 136997 123733
rect 136947 123675 136955 123709
rect 136989 123675 136997 123709
rect 136947 123651 136997 123675
rect 1801 123373 1851 123397
rect 1801 123339 1809 123373
rect 1843 123339 1851 123373
rect 1801 123315 1851 123339
rect 136947 123373 136997 123397
rect 136947 123339 136955 123373
rect 136989 123339 136997 123373
rect 136947 123315 136997 123339
rect 1801 123037 1851 123061
rect 1801 123003 1809 123037
rect 1843 123003 1851 123037
rect 1801 122979 1851 123003
rect 136947 123037 136997 123061
rect 136947 123003 136955 123037
rect 136989 123003 136997 123037
rect 136947 122979 136997 123003
rect 1801 122701 1851 122725
rect 1801 122667 1809 122701
rect 1843 122667 1851 122701
rect 1801 122643 1851 122667
rect 136947 122701 136997 122725
rect 136947 122667 136955 122701
rect 136989 122667 136997 122701
rect 136947 122643 136997 122667
rect 1801 122365 1851 122389
rect 1801 122331 1809 122365
rect 1843 122331 1851 122365
rect 1801 122307 1851 122331
rect 136947 122365 136997 122389
rect 136947 122331 136955 122365
rect 136989 122331 136997 122365
rect 136947 122307 136997 122331
rect 1801 122029 1851 122053
rect 1801 121995 1809 122029
rect 1843 121995 1851 122029
rect 1801 121971 1851 121995
rect 136947 122029 136997 122053
rect 136947 121995 136955 122029
rect 136989 121995 136997 122029
rect 136947 121971 136997 121995
rect 1801 121693 1851 121717
rect 1801 121659 1809 121693
rect 1843 121659 1851 121693
rect 1801 121635 1851 121659
rect 136947 121693 136997 121717
rect 136947 121659 136955 121693
rect 136989 121659 136997 121693
rect 136947 121635 136997 121659
rect 1801 121357 1851 121381
rect 1801 121323 1809 121357
rect 1843 121323 1851 121357
rect 1801 121299 1851 121323
rect 136947 121357 136997 121381
rect 136947 121323 136955 121357
rect 136989 121323 136997 121357
rect 136947 121299 136997 121323
rect 1801 121021 1851 121045
rect 1801 120987 1809 121021
rect 1843 120987 1851 121021
rect 1801 120963 1851 120987
rect 136947 121021 136997 121045
rect 136947 120987 136955 121021
rect 136989 120987 136997 121021
rect 136947 120963 136997 120987
rect 1801 120685 1851 120709
rect 1801 120651 1809 120685
rect 1843 120651 1851 120685
rect 1801 120627 1851 120651
rect 136947 120685 136997 120709
rect 136947 120651 136955 120685
rect 136989 120651 136997 120685
rect 136947 120627 136997 120651
rect 1801 120349 1851 120373
rect 1801 120315 1809 120349
rect 1843 120315 1851 120349
rect 1801 120291 1851 120315
rect 136947 120349 136997 120373
rect 136947 120315 136955 120349
rect 136989 120315 136997 120349
rect 136947 120291 136997 120315
rect 1801 120013 1851 120037
rect 1801 119979 1809 120013
rect 1843 119979 1851 120013
rect 1801 119955 1851 119979
rect 136947 120013 136997 120037
rect 136947 119979 136955 120013
rect 136989 119979 136997 120013
rect 136947 119955 136997 119979
rect 1801 119677 1851 119701
rect 1801 119643 1809 119677
rect 1843 119643 1851 119677
rect 1801 119619 1851 119643
rect 136947 119677 136997 119701
rect 136947 119643 136955 119677
rect 136989 119643 136997 119677
rect 136947 119619 136997 119643
rect 1801 119341 1851 119365
rect 1801 119307 1809 119341
rect 1843 119307 1851 119341
rect 1801 119283 1851 119307
rect 136947 119341 136997 119365
rect 136947 119307 136955 119341
rect 136989 119307 136997 119341
rect 136947 119283 136997 119307
rect 1801 119005 1851 119029
rect 1801 118971 1809 119005
rect 1843 118971 1851 119005
rect 1801 118947 1851 118971
rect 136947 119005 136997 119029
rect 136947 118971 136955 119005
rect 136989 118971 136997 119005
rect 136947 118947 136997 118971
rect 1801 118669 1851 118693
rect 1801 118635 1809 118669
rect 1843 118635 1851 118669
rect 1801 118611 1851 118635
rect 136947 118669 136997 118693
rect 136947 118635 136955 118669
rect 136989 118635 136997 118669
rect 136947 118611 136997 118635
rect 1801 118333 1851 118357
rect 1801 118299 1809 118333
rect 1843 118299 1851 118333
rect 1801 118275 1851 118299
rect 136947 118333 136997 118357
rect 136947 118299 136955 118333
rect 136989 118299 136997 118333
rect 136947 118275 136997 118299
rect 1801 117997 1851 118021
rect 1801 117963 1809 117997
rect 1843 117963 1851 117997
rect 1801 117939 1851 117963
rect 136947 117997 136997 118021
rect 136947 117963 136955 117997
rect 136989 117963 136997 117997
rect 136947 117939 136997 117963
rect 1801 117661 1851 117685
rect 1801 117627 1809 117661
rect 1843 117627 1851 117661
rect 1801 117603 1851 117627
rect 136947 117661 136997 117685
rect 136947 117627 136955 117661
rect 136989 117627 136997 117661
rect 136947 117603 136997 117627
rect 1801 117325 1851 117349
rect 1801 117291 1809 117325
rect 1843 117291 1851 117325
rect 1801 117267 1851 117291
rect 136947 117325 136997 117349
rect 136947 117291 136955 117325
rect 136989 117291 136997 117325
rect 136947 117267 136997 117291
rect 1801 116989 1851 117013
rect 1801 116955 1809 116989
rect 1843 116955 1851 116989
rect 1801 116931 1851 116955
rect 136947 116989 136997 117013
rect 136947 116955 136955 116989
rect 136989 116955 136997 116989
rect 136947 116931 136997 116955
rect 1801 116653 1851 116677
rect 1801 116619 1809 116653
rect 1843 116619 1851 116653
rect 1801 116595 1851 116619
rect 136947 116653 136997 116677
rect 136947 116619 136955 116653
rect 136989 116619 136997 116653
rect 136947 116595 136997 116619
rect 1801 116317 1851 116341
rect 1801 116283 1809 116317
rect 1843 116283 1851 116317
rect 1801 116259 1851 116283
rect 136947 116317 136997 116341
rect 136947 116283 136955 116317
rect 136989 116283 136997 116317
rect 136947 116259 136997 116283
rect 1801 115981 1851 116005
rect 1801 115947 1809 115981
rect 1843 115947 1851 115981
rect 1801 115923 1851 115947
rect 136947 115981 136997 116005
rect 136947 115947 136955 115981
rect 136989 115947 136997 115981
rect 136947 115923 136997 115947
rect 1801 115645 1851 115669
rect 1801 115611 1809 115645
rect 1843 115611 1851 115645
rect 1801 115587 1851 115611
rect 136947 115645 136997 115669
rect 136947 115611 136955 115645
rect 136989 115611 136997 115645
rect 136947 115587 136997 115611
rect 1801 115309 1851 115333
rect 1801 115275 1809 115309
rect 1843 115275 1851 115309
rect 1801 115251 1851 115275
rect 136947 115309 136997 115333
rect 136947 115275 136955 115309
rect 136989 115275 136997 115309
rect 136947 115251 136997 115275
rect 1801 114973 1851 114997
rect 1801 114939 1809 114973
rect 1843 114939 1851 114973
rect 1801 114915 1851 114939
rect 136947 114973 136997 114997
rect 136947 114939 136955 114973
rect 136989 114939 136997 114973
rect 136947 114915 136997 114939
rect 1801 114637 1851 114661
rect 1801 114603 1809 114637
rect 1843 114603 1851 114637
rect 1801 114579 1851 114603
rect 136947 114637 136997 114661
rect 136947 114603 136955 114637
rect 136989 114603 136997 114637
rect 136947 114579 136997 114603
rect 1801 114301 1851 114325
rect 1801 114267 1809 114301
rect 1843 114267 1851 114301
rect 1801 114243 1851 114267
rect 136947 114301 136997 114325
rect 136947 114267 136955 114301
rect 136989 114267 136997 114301
rect 136947 114243 136997 114267
rect 1801 113965 1851 113989
rect 1801 113931 1809 113965
rect 1843 113931 1851 113965
rect 1801 113907 1851 113931
rect 136947 113965 136997 113989
rect 136947 113931 136955 113965
rect 136989 113931 136997 113965
rect 136947 113907 136997 113931
rect 1801 113629 1851 113653
rect 1801 113595 1809 113629
rect 1843 113595 1851 113629
rect 1801 113571 1851 113595
rect 136947 113629 136997 113653
rect 136947 113595 136955 113629
rect 136989 113595 136997 113629
rect 136947 113571 136997 113595
rect 1801 113293 1851 113317
rect 1801 113259 1809 113293
rect 1843 113259 1851 113293
rect 1801 113235 1851 113259
rect 136947 113293 136997 113317
rect 136947 113259 136955 113293
rect 136989 113259 136997 113293
rect 136947 113235 136997 113259
rect 1801 112957 1851 112981
rect 1801 112923 1809 112957
rect 1843 112923 1851 112957
rect 1801 112899 1851 112923
rect 136947 112957 136997 112981
rect 136947 112923 136955 112957
rect 136989 112923 136997 112957
rect 136947 112899 136997 112923
rect 1801 112621 1851 112645
rect 1801 112587 1809 112621
rect 1843 112587 1851 112621
rect 1801 112563 1851 112587
rect 136947 112621 136997 112645
rect 136947 112587 136955 112621
rect 136989 112587 136997 112621
rect 136947 112563 136997 112587
rect 1801 112285 1851 112309
rect 1801 112251 1809 112285
rect 1843 112251 1851 112285
rect 1801 112227 1851 112251
rect 136947 112285 136997 112309
rect 136947 112251 136955 112285
rect 136989 112251 136997 112285
rect 136947 112227 136997 112251
rect 1801 111949 1851 111973
rect 1801 111915 1809 111949
rect 1843 111915 1851 111949
rect 1801 111891 1851 111915
rect 136947 111949 136997 111973
rect 136947 111915 136955 111949
rect 136989 111915 136997 111949
rect 136947 111891 136997 111915
rect 1801 111613 1851 111637
rect 1801 111579 1809 111613
rect 1843 111579 1851 111613
rect 1801 111555 1851 111579
rect 136947 111613 136997 111637
rect 136947 111579 136955 111613
rect 136989 111579 136997 111613
rect 136947 111555 136997 111579
rect 1801 111277 1851 111301
rect 1801 111243 1809 111277
rect 1843 111243 1851 111277
rect 1801 111219 1851 111243
rect 136947 111277 136997 111301
rect 136947 111243 136955 111277
rect 136989 111243 136997 111277
rect 136947 111219 136997 111243
rect 1801 110941 1851 110965
rect 1801 110907 1809 110941
rect 1843 110907 1851 110941
rect 1801 110883 1851 110907
rect 136947 110941 136997 110965
rect 136947 110907 136955 110941
rect 136989 110907 136997 110941
rect 136947 110883 136997 110907
rect 1801 110605 1851 110629
rect 1801 110571 1809 110605
rect 1843 110571 1851 110605
rect 1801 110547 1851 110571
rect 136947 110605 136997 110629
rect 136947 110571 136955 110605
rect 136989 110571 136997 110605
rect 136947 110547 136997 110571
rect 1801 110269 1851 110293
rect 1801 110235 1809 110269
rect 1843 110235 1851 110269
rect 1801 110211 1851 110235
rect 136947 110269 136997 110293
rect 136947 110235 136955 110269
rect 136989 110235 136997 110269
rect 136947 110211 136997 110235
rect 1801 109933 1851 109957
rect 1801 109899 1809 109933
rect 1843 109899 1851 109933
rect 1801 109875 1851 109899
rect 136947 109933 136997 109957
rect 136947 109899 136955 109933
rect 136989 109899 136997 109933
rect 136947 109875 136997 109899
rect 1801 109597 1851 109621
rect 1801 109563 1809 109597
rect 1843 109563 1851 109597
rect 1801 109539 1851 109563
rect 136947 109597 136997 109621
rect 136947 109563 136955 109597
rect 136989 109563 136997 109597
rect 136947 109539 136997 109563
rect 1801 109261 1851 109285
rect 1801 109227 1809 109261
rect 1843 109227 1851 109261
rect 1801 109203 1851 109227
rect 136947 109261 136997 109285
rect 136947 109227 136955 109261
rect 136989 109227 136997 109261
rect 136947 109203 136997 109227
rect 1801 108925 1851 108949
rect 1801 108891 1809 108925
rect 1843 108891 1851 108925
rect 1801 108867 1851 108891
rect 136947 108925 136997 108949
rect 136947 108891 136955 108925
rect 136989 108891 136997 108925
rect 136947 108867 136997 108891
rect 1801 108589 1851 108613
rect 1801 108555 1809 108589
rect 1843 108555 1851 108589
rect 1801 108531 1851 108555
rect 136947 108589 136997 108613
rect 136947 108555 136955 108589
rect 136989 108555 136997 108589
rect 136947 108531 136997 108555
rect 1801 108253 1851 108277
rect 1801 108219 1809 108253
rect 1843 108219 1851 108253
rect 1801 108195 1851 108219
rect 136947 108253 136997 108277
rect 136947 108219 136955 108253
rect 136989 108219 136997 108253
rect 136947 108195 136997 108219
rect 1801 107917 1851 107941
rect 1801 107883 1809 107917
rect 1843 107883 1851 107917
rect 1801 107859 1851 107883
rect 136947 107917 136997 107941
rect 136947 107883 136955 107917
rect 136989 107883 136997 107917
rect 136947 107859 136997 107883
rect 1801 107581 1851 107605
rect 1801 107547 1809 107581
rect 1843 107547 1851 107581
rect 1801 107523 1851 107547
rect 136947 107581 136997 107605
rect 136947 107547 136955 107581
rect 136989 107547 136997 107581
rect 136947 107523 136997 107547
rect 1801 107245 1851 107269
rect 1801 107211 1809 107245
rect 1843 107211 1851 107245
rect 1801 107187 1851 107211
rect 136947 107245 136997 107269
rect 136947 107211 136955 107245
rect 136989 107211 136997 107245
rect 136947 107187 136997 107211
rect 1801 106909 1851 106933
rect 1801 106875 1809 106909
rect 1843 106875 1851 106909
rect 1801 106851 1851 106875
rect 136947 106909 136997 106933
rect 136947 106875 136955 106909
rect 136989 106875 136997 106909
rect 136947 106851 136997 106875
rect 1801 106573 1851 106597
rect 1801 106539 1809 106573
rect 1843 106539 1851 106573
rect 1801 106515 1851 106539
rect 136947 106573 136997 106597
rect 136947 106539 136955 106573
rect 136989 106539 136997 106573
rect 136947 106515 136997 106539
rect 1801 106237 1851 106261
rect 1801 106203 1809 106237
rect 1843 106203 1851 106237
rect 1801 106179 1851 106203
rect 136947 106237 136997 106261
rect 136947 106203 136955 106237
rect 136989 106203 136997 106237
rect 136947 106179 136997 106203
rect 1801 105901 1851 105925
rect 1801 105867 1809 105901
rect 1843 105867 1851 105901
rect 1801 105843 1851 105867
rect 136947 105901 136997 105925
rect 136947 105867 136955 105901
rect 136989 105867 136997 105901
rect 136947 105843 136997 105867
rect 1801 105565 1851 105589
rect 1801 105531 1809 105565
rect 1843 105531 1851 105565
rect 1801 105507 1851 105531
rect 136947 105565 136997 105589
rect 136947 105531 136955 105565
rect 136989 105531 136997 105565
rect 136947 105507 136997 105531
rect 1801 105229 1851 105253
rect 1801 105195 1809 105229
rect 1843 105195 1851 105229
rect 1801 105171 1851 105195
rect 136947 105229 136997 105253
rect 136947 105195 136955 105229
rect 136989 105195 136997 105229
rect 136947 105171 136997 105195
rect 1801 104893 1851 104917
rect 1801 104859 1809 104893
rect 1843 104859 1851 104893
rect 1801 104835 1851 104859
rect 136947 104893 136997 104917
rect 136947 104859 136955 104893
rect 136989 104859 136997 104893
rect 136947 104835 136997 104859
rect 1801 104557 1851 104581
rect 1801 104523 1809 104557
rect 1843 104523 1851 104557
rect 1801 104499 1851 104523
rect 136947 104557 136997 104581
rect 136947 104523 136955 104557
rect 136989 104523 136997 104557
rect 136947 104499 136997 104523
rect 1801 104221 1851 104245
rect 1801 104187 1809 104221
rect 1843 104187 1851 104221
rect 1801 104163 1851 104187
rect 136947 104221 136997 104245
rect 136947 104187 136955 104221
rect 136989 104187 136997 104221
rect 136947 104163 136997 104187
rect 1801 103885 1851 103909
rect 1801 103851 1809 103885
rect 1843 103851 1851 103885
rect 1801 103827 1851 103851
rect 136947 103885 136997 103909
rect 136947 103851 136955 103885
rect 136989 103851 136997 103885
rect 136947 103827 136997 103851
rect 1801 103549 1851 103573
rect 1801 103515 1809 103549
rect 1843 103515 1851 103549
rect 1801 103491 1851 103515
rect 136947 103549 136997 103573
rect 136947 103515 136955 103549
rect 136989 103515 136997 103549
rect 136947 103491 136997 103515
rect 1801 103213 1851 103237
rect 1801 103179 1809 103213
rect 1843 103179 1851 103213
rect 1801 103155 1851 103179
rect 136947 103213 136997 103237
rect 136947 103179 136955 103213
rect 136989 103179 136997 103213
rect 136947 103155 136997 103179
rect 1801 102877 1851 102901
rect 1801 102843 1809 102877
rect 1843 102843 1851 102877
rect 1801 102819 1851 102843
rect 136947 102877 136997 102901
rect 136947 102843 136955 102877
rect 136989 102843 136997 102877
rect 136947 102819 136997 102843
rect 1801 102541 1851 102565
rect 1801 102507 1809 102541
rect 1843 102507 1851 102541
rect 1801 102483 1851 102507
rect 136947 102541 136997 102565
rect 136947 102507 136955 102541
rect 136989 102507 136997 102541
rect 136947 102483 136997 102507
rect 1801 102205 1851 102229
rect 1801 102171 1809 102205
rect 1843 102171 1851 102205
rect 1801 102147 1851 102171
rect 136947 102205 136997 102229
rect 136947 102171 136955 102205
rect 136989 102171 136997 102205
rect 136947 102147 136997 102171
rect 1801 101869 1851 101893
rect 1801 101835 1809 101869
rect 1843 101835 1851 101869
rect 1801 101811 1851 101835
rect 136947 101869 136997 101893
rect 136947 101835 136955 101869
rect 136989 101835 136997 101869
rect 136947 101811 136997 101835
rect 1801 101533 1851 101557
rect 1801 101499 1809 101533
rect 1843 101499 1851 101533
rect 1801 101475 1851 101499
rect 136947 101533 136997 101557
rect 136947 101499 136955 101533
rect 136989 101499 136997 101533
rect 136947 101475 136997 101499
rect 1801 101197 1851 101221
rect 1801 101163 1809 101197
rect 1843 101163 1851 101197
rect 1801 101139 1851 101163
rect 136947 101197 136997 101221
rect 136947 101163 136955 101197
rect 136989 101163 136997 101197
rect 136947 101139 136997 101163
rect 1801 100861 1851 100885
rect 1801 100827 1809 100861
rect 1843 100827 1851 100861
rect 1801 100803 1851 100827
rect 136947 100861 136997 100885
rect 136947 100827 136955 100861
rect 136989 100827 136997 100861
rect 136947 100803 136997 100827
rect 1801 100525 1851 100549
rect 1801 100491 1809 100525
rect 1843 100491 1851 100525
rect 1801 100467 1851 100491
rect 136947 100525 136997 100549
rect 136947 100491 136955 100525
rect 136989 100491 136997 100525
rect 136947 100467 136997 100491
rect 1801 100189 1851 100213
rect 1801 100155 1809 100189
rect 1843 100155 1851 100189
rect 1801 100131 1851 100155
rect 136947 100189 136997 100213
rect 136947 100155 136955 100189
rect 136989 100155 136997 100189
rect 136947 100131 136997 100155
rect 1801 99853 1851 99877
rect 1801 99819 1809 99853
rect 1843 99819 1851 99853
rect 1801 99795 1851 99819
rect 136947 99853 136997 99877
rect 136947 99819 136955 99853
rect 136989 99819 136997 99853
rect 136947 99795 136997 99819
rect 1801 99517 1851 99541
rect 1801 99483 1809 99517
rect 1843 99483 1851 99517
rect 1801 99459 1851 99483
rect 136947 99517 136997 99541
rect 136947 99483 136955 99517
rect 136989 99483 136997 99517
rect 136947 99459 136997 99483
rect 1801 99181 1851 99205
rect 1801 99147 1809 99181
rect 1843 99147 1851 99181
rect 1801 99123 1851 99147
rect 136947 99181 136997 99205
rect 136947 99147 136955 99181
rect 136989 99147 136997 99181
rect 136947 99123 136997 99147
rect 1801 98845 1851 98869
rect 1801 98811 1809 98845
rect 1843 98811 1851 98845
rect 1801 98787 1851 98811
rect 136947 98845 136997 98869
rect 136947 98811 136955 98845
rect 136989 98811 136997 98845
rect 136947 98787 136997 98811
rect 1801 98509 1851 98533
rect 1801 98475 1809 98509
rect 1843 98475 1851 98509
rect 1801 98451 1851 98475
rect 136947 98509 136997 98533
rect 136947 98475 136955 98509
rect 136989 98475 136997 98509
rect 136947 98451 136997 98475
rect 1801 98173 1851 98197
rect 1801 98139 1809 98173
rect 1843 98139 1851 98173
rect 1801 98115 1851 98139
rect 136947 98173 136997 98197
rect 136947 98139 136955 98173
rect 136989 98139 136997 98173
rect 136947 98115 136997 98139
rect 1801 97837 1851 97861
rect 1801 97803 1809 97837
rect 1843 97803 1851 97837
rect 1801 97779 1851 97803
rect 136947 97837 136997 97861
rect 136947 97803 136955 97837
rect 136989 97803 136997 97837
rect 136947 97779 136997 97803
rect 1801 97501 1851 97525
rect 1801 97467 1809 97501
rect 1843 97467 1851 97501
rect 1801 97443 1851 97467
rect 136947 97501 136997 97525
rect 136947 97467 136955 97501
rect 136989 97467 136997 97501
rect 136947 97443 136997 97467
rect 1801 97165 1851 97189
rect 1801 97131 1809 97165
rect 1843 97131 1851 97165
rect 1801 97107 1851 97131
rect 136947 97165 136997 97189
rect 136947 97131 136955 97165
rect 136989 97131 136997 97165
rect 136947 97107 136997 97131
rect 1801 96829 1851 96853
rect 1801 96795 1809 96829
rect 1843 96795 1851 96829
rect 1801 96771 1851 96795
rect 136947 96829 136997 96853
rect 136947 96795 136955 96829
rect 136989 96795 136997 96829
rect 136947 96771 136997 96795
rect 1801 96493 1851 96517
rect 1801 96459 1809 96493
rect 1843 96459 1851 96493
rect 1801 96435 1851 96459
rect 136947 96493 136997 96517
rect 136947 96459 136955 96493
rect 136989 96459 136997 96493
rect 136947 96435 136997 96459
rect 1801 96157 1851 96181
rect 1801 96123 1809 96157
rect 1843 96123 1851 96157
rect 1801 96099 1851 96123
rect 136947 96157 136997 96181
rect 136947 96123 136955 96157
rect 136989 96123 136997 96157
rect 136947 96099 136997 96123
rect 1801 95821 1851 95845
rect 1801 95787 1809 95821
rect 1843 95787 1851 95821
rect 1801 95763 1851 95787
rect 136947 95821 136997 95845
rect 136947 95787 136955 95821
rect 136989 95787 136997 95821
rect 136947 95763 136997 95787
rect 1801 95485 1851 95509
rect 1801 95451 1809 95485
rect 1843 95451 1851 95485
rect 1801 95427 1851 95451
rect 136947 95485 136997 95509
rect 136947 95451 136955 95485
rect 136989 95451 136997 95485
rect 136947 95427 136997 95451
rect 1801 95149 1851 95173
rect 1801 95115 1809 95149
rect 1843 95115 1851 95149
rect 1801 95091 1851 95115
rect 136947 95149 136997 95173
rect 136947 95115 136955 95149
rect 136989 95115 136997 95149
rect 136947 95091 136997 95115
rect 1801 94813 1851 94837
rect 1801 94779 1809 94813
rect 1843 94779 1851 94813
rect 1801 94755 1851 94779
rect 136947 94813 136997 94837
rect 136947 94779 136955 94813
rect 136989 94779 136997 94813
rect 136947 94755 136997 94779
rect 1801 94477 1851 94501
rect 1801 94443 1809 94477
rect 1843 94443 1851 94477
rect 1801 94419 1851 94443
rect 136947 94477 136997 94501
rect 136947 94443 136955 94477
rect 136989 94443 136997 94477
rect 136947 94419 136997 94443
rect 1801 94141 1851 94165
rect 1801 94107 1809 94141
rect 1843 94107 1851 94141
rect 1801 94083 1851 94107
rect 136947 94141 136997 94165
rect 136947 94107 136955 94141
rect 136989 94107 136997 94141
rect 136947 94083 136997 94107
rect 1801 93805 1851 93829
rect 1801 93771 1809 93805
rect 1843 93771 1851 93805
rect 1801 93747 1851 93771
rect 136947 93805 136997 93829
rect 136947 93771 136955 93805
rect 136989 93771 136997 93805
rect 136947 93747 136997 93771
rect 1801 93469 1851 93493
rect 1801 93435 1809 93469
rect 1843 93435 1851 93469
rect 1801 93411 1851 93435
rect 136947 93469 136997 93493
rect 136947 93435 136955 93469
rect 136989 93435 136997 93469
rect 136947 93411 136997 93435
rect 1801 93133 1851 93157
rect 1801 93099 1809 93133
rect 1843 93099 1851 93133
rect 1801 93075 1851 93099
rect 136947 93133 136997 93157
rect 136947 93099 136955 93133
rect 136989 93099 136997 93133
rect 136947 93075 136997 93099
rect 1801 92797 1851 92821
rect 1801 92763 1809 92797
rect 1843 92763 1851 92797
rect 1801 92739 1851 92763
rect 136947 92797 136997 92821
rect 136947 92763 136955 92797
rect 136989 92763 136997 92797
rect 136947 92739 136997 92763
rect 1801 92461 1851 92485
rect 1801 92427 1809 92461
rect 1843 92427 1851 92461
rect 1801 92403 1851 92427
rect 136947 92461 136997 92485
rect 136947 92427 136955 92461
rect 136989 92427 136997 92461
rect 136947 92403 136997 92427
rect 1801 92125 1851 92149
rect 1801 92091 1809 92125
rect 1843 92091 1851 92125
rect 1801 92067 1851 92091
rect 136947 92125 136997 92149
rect 136947 92091 136955 92125
rect 136989 92091 136997 92125
rect 136947 92067 136997 92091
rect 1801 91789 1851 91813
rect 1801 91755 1809 91789
rect 1843 91755 1851 91789
rect 1801 91731 1851 91755
rect 136947 91789 136997 91813
rect 136947 91755 136955 91789
rect 136989 91755 136997 91789
rect 136947 91731 136997 91755
rect 1801 91453 1851 91477
rect 1801 91419 1809 91453
rect 1843 91419 1851 91453
rect 1801 91395 1851 91419
rect 136947 91453 136997 91477
rect 136947 91419 136955 91453
rect 136989 91419 136997 91453
rect 136947 91395 136997 91419
rect 1801 91117 1851 91141
rect 1801 91083 1809 91117
rect 1843 91083 1851 91117
rect 1801 91059 1851 91083
rect 136947 91117 136997 91141
rect 136947 91083 136955 91117
rect 136989 91083 136997 91117
rect 136947 91059 136997 91083
rect 1801 90781 1851 90805
rect 1801 90747 1809 90781
rect 1843 90747 1851 90781
rect 1801 90723 1851 90747
rect 136947 90781 136997 90805
rect 136947 90747 136955 90781
rect 136989 90747 136997 90781
rect 136947 90723 136997 90747
rect 1801 90445 1851 90469
rect 1801 90411 1809 90445
rect 1843 90411 1851 90445
rect 1801 90387 1851 90411
rect 136947 90445 136997 90469
rect 136947 90411 136955 90445
rect 136989 90411 136997 90445
rect 136947 90387 136997 90411
rect 1801 90109 1851 90133
rect 1801 90075 1809 90109
rect 1843 90075 1851 90109
rect 1801 90051 1851 90075
rect 136947 90109 136997 90133
rect 136947 90075 136955 90109
rect 136989 90075 136997 90109
rect 136947 90051 136997 90075
rect 1801 89773 1851 89797
rect 1801 89739 1809 89773
rect 1843 89739 1851 89773
rect 1801 89715 1851 89739
rect 136947 89773 136997 89797
rect 136947 89739 136955 89773
rect 136989 89739 136997 89773
rect 136947 89715 136997 89739
rect 1801 89437 1851 89461
rect 1801 89403 1809 89437
rect 1843 89403 1851 89437
rect 1801 89379 1851 89403
rect 136947 89437 136997 89461
rect 136947 89403 136955 89437
rect 136989 89403 136997 89437
rect 136947 89379 136997 89403
rect 1801 89101 1851 89125
rect 1801 89067 1809 89101
rect 1843 89067 1851 89101
rect 1801 89043 1851 89067
rect 136947 89101 136997 89125
rect 136947 89067 136955 89101
rect 136989 89067 136997 89101
rect 136947 89043 136997 89067
rect 1801 88765 1851 88789
rect 1801 88731 1809 88765
rect 1843 88731 1851 88765
rect 1801 88707 1851 88731
rect 136947 88765 136997 88789
rect 136947 88731 136955 88765
rect 136989 88731 136997 88765
rect 136947 88707 136997 88731
rect 1801 88429 1851 88453
rect 1801 88395 1809 88429
rect 1843 88395 1851 88429
rect 1801 88371 1851 88395
rect 136947 88429 136997 88453
rect 136947 88395 136955 88429
rect 136989 88395 136997 88429
rect 136947 88371 136997 88395
rect 1801 88093 1851 88117
rect 1801 88059 1809 88093
rect 1843 88059 1851 88093
rect 1801 88035 1851 88059
rect 136947 88093 136997 88117
rect 136947 88059 136955 88093
rect 136989 88059 136997 88093
rect 136947 88035 136997 88059
rect 1801 87757 1851 87781
rect 1801 87723 1809 87757
rect 1843 87723 1851 87757
rect 1801 87699 1851 87723
rect 136947 87757 136997 87781
rect 136947 87723 136955 87757
rect 136989 87723 136997 87757
rect 136947 87699 136997 87723
rect 1801 87421 1851 87445
rect 1801 87387 1809 87421
rect 1843 87387 1851 87421
rect 1801 87363 1851 87387
rect 136947 87421 136997 87445
rect 136947 87387 136955 87421
rect 136989 87387 136997 87421
rect 136947 87363 136997 87387
rect 1801 87085 1851 87109
rect 1801 87051 1809 87085
rect 1843 87051 1851 87085
rect 1801 87027 1851 87051
rect 136947 87085 136997 87109
rect 136947 87051 136955 87085
rect 136989 87051 136997 87085
rect 136947 87027 136997 87051
rect 1801 86749 1851 86773
rect 1801 86715 1809 86749
rect 1843 86715 1851 86749
rect 1801 86691 1851 86715
rect 136947 86749 136997 86773
rect 136947 86715 136955 86749
rect 136989 86715 136997 86749
rect 136947 86691 136997 86715
rect 1801 86413 1851 86437
rect 1801 86379 1809 86413
rect 1843 86379 1851 86413
rect 1801 86355 1851 86379
rect 136947 86413 136997 86437
rect 136947 86379 136955 86413
rect 136989 86379 136997 86413
rect 136947 86355 136997 86379
rect 1801 86077 1851 86101
rect 1801 86043 1809 86077
rect 1843 86043 1851 86077
rect 1801 86019 1851 86043
rect 136947 86077 136997 86101
rect 136947 86043 136955 86077
rect 136989 86043 136997 86077
rect 136947 86019 136997 86043
rect 1801 85741 1851 85765
rect 1801 85707 1809 85741
rect 1843 85707 1851 85741
rect 1801 85683 1851 85707
rect 136947 85741 136997 85765
rect 136947 85707 136955 85741
rect 136989 85707 136997 85741
rect 136947 85683 136997 85707
rect 1801 85405 1851 85429
rect 1801 85371 1809 85405
rect 1843 85371 1851 85405
rect 1801 85347 1851 85371
rect 136947 85405 136997 85429
rect 136947 85371 136955 85405
rect 136989 85371 136997 85405
rect 136947 85347 136997 85371
rect 1801 85069 1851 85093
rect 1801 85035 1809 85069
rect 1843 85035 1851 85069
rect 1801 85011 1851 85035
rect 136947 85069 136997 85093
rect 136947 85035 136955 85069
rect 136989 85035 136997 85069
rect 136947 85011 136997 85035
rect 1801 84733 1851 84757
rect 1801 84699 1809 84733
rect 1843 84699 1851 84733
rect 1801 84675 1851 84699
rect 136947 84733 136997 84757
rect 136947 84699 136955 84733
rect 136989 84699 136997 84733
rect 136947 84675 136997 84699
rect 1801 84397 1851 84421
rect 1801 84363 1809 84397
rect 1843 84363 1851 84397
rect 1801 84339 1851 84363
rect 136947 84397 136997 84421
rect 136947 84363 136955 84397
rect 136989 84363 136997 84397
rect 136947 84339 136997 84363
rect 1801 84061 1851 84085
rect 1801 84027 1809 84061
rect 1843 84027 1851 84061
rect 1801 84003 1851 84027
rect 136947 84061 136997 84085
rect 136947 84027 136955 84061
rect 136989 84027 136997 84061
rect 136947 84003 136997 84027
rect 1801 83725 1851 83749
rect 1801 83691 1809 83725
rect 1843 83691 1851 83725
rect 1801 83667 1851 83691
rect 136947 83725 136997 83749
rect 136947 83691 136955 83725
rect 136989 83691 136997 83725
rect 136947 83667 136997 83691
rect 1801 83389 1851 83413
rect 1801 83355 1809 83389
rect 1843 83355 1851 83389
rect 1801 83331 1851 83355
rect 136947 83389 136997 83413
rect 136947 83355 136955 83389
rect 136989 83355 136997 83389
rect 136947 83331 136997 83355
rect 1801 83053 1851 83077
rect 1801 83019 1809 83053
rect 1843 83019 1851 83053
rect 1801 82995 1851 83019
rect 136947 83053 136997 83077
rect 136947 83019 136955 83053
rect 136989 83019 136997 83053
rect 136947 82995 136997 83019
rect 1801 82717 1851 82741
rect 1801 82683 1809 82717
rect 1843 82683 1851 82717
rect 1801 82659 1851 82683
rect 136947 82717 136997 82741
rect 136947 82683 136955 82717
rect 136989 82683 136997 82717
rect 136947 82659 136997 82683
rect 1801 82381 1851 82405
rect 1801 82347 1809 82381
rect 1843 82347 1851 82381
rect 1801 82323 1851 82347
rect 136947 82381 136997 82405
rect 136947 82347 136955 82381
rect 136989 82347 136997 82381
rect 136947 82323 136997 82347
rect 1801 82045 1851 82069
rect 1801 82011 1809 82045
rect 1843 82011 1851 82045
rect 1801 81987 1851 82011
rect 136947 82045 136997 82069
rect 136947 82011 136955 82045
rect 136989 82011 136997 82045
rect 136947 81987 136997 82011
rect 1801 81709 1851 81733
rect 1801 81675 1809 81709
rect 1843 81675 1851 81709
rect 1801 81651 1851 81675
rect 136947 81709 136997 81733
rect 136947 81675 136955 81709
rect 136989 81675 136997 81709
rect 136947 81651 136997 81675
rect 1801 81373 1851 81397
rect 1801 81339 1809 81373
rect 1843 81339 1851 81373
rect 1801 81315 1851 81339
rect 136947 81373 136997 81397
rect 136947 81339 136955 81373
rect 136989 81339 136997 81373
rect 136947 81315 136997 81339
rect 1801 81037 1851 81061
rect 1801 81003 1809 81037
rect 1843 81003 1851 81037
rect 1801 80979 1851 81003
rect 136947 81037 136997 81061
rect 136947 81003 136955 81037
rect 136989 81003 136997 81037
rect 136947 80979 136997 81003
rect 1801 80701 1851 80725
rect 1801 80667 1809 80701
rect 1843 80667 1851 80701
rect 1801 80643 1851 80667
rect 136947 80701 136997 80725
rect 136947 80667 136955 80701
rect 136989 80667 136997 80701
rect 136947 80643 136997 80667
rect 1801 80365 1851 80389
rect 1801 80331 1809 80365
rect 1843 80331 1851 80365
rect 1801 80307 1851 80331
rect 136947 80365 136997 80389
rect 136947 80331 136955 80365
rect 136989 80331 136997 80365
rect 136947 80307 136997 80331
rect 1801 80029 1851 80053
rect 1801 79995 1809 80029
rect 1843 79995 1851 80029
rect 1801 79971 1851 79995
rect 136947 80029 136997 80053
rect 136947 79995 136955 80029
rect 136989 79995 136997 80029
rect 136947 79971 136997 79995
rect 1801 79693 1851 79717
rect 1801 79659 1809 79693
rect 1843 79659 1851 79693
rect 1801 79635 1851 79659
rect 136947 79693 136997 79717
rect 136947 79659 136955 79693
rect 136989 79659 136997 79693
rect 136947 79635 136997 79659
rect 1801 79357 1851 79381
rect 1801 79323 1809 79357
rect 1843 79323 1851 79357
rect 1801 79299 1851 79323
rect 136947 79357 136997 79381
rect 136947 79323 136955 79357
rect 136989 79323 136997 79357
rect 136947 79299 136997 79323
rect 1801 79021 1851 79045
rect 1801 78987 1809 79021
rect 1843 78987 1851 79021
rect 1801 78963 1851 78987
rect 136947 79021 136997 79045
rect 136947 78987 136955 79021
rect 136989 78987 136997 79021
rect 136947 78963 136997 78987
rect 1801 78685 1851 78709
rect 1801 78651 1809 78685
rect 1843 78651 1851 78685
rect 1801 78627 1851 78651
rect 136947 78685 136997 78709
rect 136947 78651 136955 78685
rect 136989 78651 136997 78685
rect 136947 78627 136997 78651
rect 1801 78349 1851 78373
rect 1801 78315 1809 78349
rect 1843 78315 1851 78349
rect 1801 78291 1851 78315
rect 136947 78349 136997 78373
rect 136947 78315 136955 78349
rect 136989 78315 136997 78349
rect 136947 78291 136997 78315
rect 1801 78013 1851 78037
rect 1801 77979 1809 78013
rect 1843 77979 1851 78013
rect 1801 77955 1851 77979
rect 136947 78013 136997 78037
rect 136947 77979 136955 78013
rect 136989 77979 136997 78013
rect 136947 77955 136997 77979
rect 1801 77677 1851 77701
rect 1801 77643 1809 77677
rect 1843 77643 1851 77677
rect 1801 77619 1851 77643
rect 136947 77677 136997 77701
rect 136947 77643 136955 77677
rect 136989 77643 136997 77677
rect 136947 77619 136997 77643
rect 1801 77341 1851 77365
rect 1801 77307 1809 77341
rect 1843 77307 1851 77341
rect 1801 77283 1851 77307
rect 136947 77341 136997 77365
rect 136947 77307 136955 77341
rect 136989 77307 136997 77341
rect 136947 77283 136997 77307
rect 1801 77005 1851 77029
rect 1801 76971 1809 77005
rect 1843 76971 1851 77005
rect 1801 76947 1851 76971
rect 136947 77005 136997 77029
rect 136947 76971 136955 77005
rect 136989 76971 136997 77005
rect 136947 76947 136997 76971
rect 1801 76669 1851 76693
rect 1801 76635 1809 76669
rect 1843 76635 1851 76669
rect 1801 76611 1851 76635
rect 136947 76669 136997 76693
rect 136947 76635 136955 76669
rect 136989 76635 136997 76669
rect 136947 76611 136997 76635
rect 1801 76333 1851 76357
rect 1801 76299 1809 76333
rect 1843 76299 1851 76333
rect 1801 76275 1851 76299
rect 136947 76333 136997 76357
rect 136947 76299 136955 76333
rect 136989 76299 136997 76333
rect 136947 76275 136997 76299
rect 1801 75997 1851 76021
rect 1801 75963 1809 75997
rect 1843 75963 1851 75997
rect 1801 75939 1851 75963
rect 136947 75997 136997 76021
rect 136947 75963 136955 75997
rect 136989 75963 136997 75997
rect 136947 75939 136997 75963
rect 1801 75661 1851 75685
rect 1801 75627 1809 75661
rect 1843 75627 1851 75661
rect 1801 75603 1851 75627
rect 136947 75661 136997 75685
rect 136947 75627 136955 75661
rect 136989 75627 136997 75661
rect 136947 75603 136997 75627
rect 1801 75325 1851 75349
rect 1801 75291 1809 75325
rect 1843 75291 1851 75325
rect 1801 75267 1851 75291
rect 136947 75325 136997 75349
rect 136947 75291 136955 75325
rect 136989 75291 136997 75325
rect 136947 75267 136997 75291
rect 1801 74989 1851 75013
rect 1801 74955 1809 74989
rect 1843 74955 1851 74989
rect 1801 74931 1851 74955
rect 136947 74989 136997 75013
rect 136947 74955 136955 74989
rect 136989 74955 136997 74989
rect 136947 74931 136997 74955
rect 1801 74653 1851 74677
rect 1801 74619 1809 74653
rect 1843 74619 1851 74653
rect 1801 74595 1851 74619
rect 136947 74653 136997 74677
rect 136947 74619 136955 74653
rect 136989 74619 136997 74653
rect 136947 74595 136997 74619
rect 1801 74317 1851 74341
rect 1801 74283 1809 74317
rect 1843 74283 1851 74317
rect 1801 74259 1851 74283
rect 136947 74317 136997 74341
rect 136947 74283 136955 74317
rect 136989 74283 136997 74317
rect 136947 74259 136997 74283
rect 1801 73981 1851 74005
rect 1801 73947 1809 73981
rect 1843 73947 1851 73981
rect 1801 73923 1851 73947
rect 136947 73981 136997 74005
rect 136947 73947 136955 73981
rect 136989 73947 136997 73981
rect 136947 73923 136997 73947
rect 1801 73645 1851 73669
rect 1801 73611 1809 73645
rect 1843 73611 1851 73645
rect 1801 73587 1851 73611
rect 136947 73645 136997 73669
rect 136947 73611 136955 73645
rect 136989 73611 136997 73645
rect 136947 73587 136997 73611
rect 1801 73309 1851 73333
rect 1801 73275 1809 73309
rect 1843 73275 1851 73309
rect 1801 73251 1851 73275
rect 136947 73309 136997 73333
rect 136947 73275 136955 73309
rect 136989 73275 136997 73309
rect 136947 73251 136997 73275
rect 1801 72973 1851 72997
rect 1801 72939 1809 72973
rect 1843 72939 1851 72973
rect 1801 72915 1851 72939
rect 136947 72973 136997 72997
rect 136947 72939 136955 72973
rect 136989 72939 136997 72973
rect 136947 72915 136997 72939
rect 1801 72637 1851 72661
rect 1801 72603 1809 72637
rect 1843 72603 1851 72637
rect 1801 72579 1851 72603
rect 136947 72637 136997 72661
rect 136947 72603 136955 72637
rect 136989 72603 136997 72637
rect 136947 72579 136997 72603
rect 1801 72301 1851 72325
rect 1801 72267 1809 72301
rect 1843 72267 1851 72301
rect 1801 72243 1851 72267
rect 136947 72301 136997 72325
rect 136947 72267 136955 72301
rect 136989 72267 136997 72301
rect 136947 72243 136997 72267
rect 1801 71965 1851 71989
rect 1801 71931 1809 71965
rect 1843 71931 1851 71965
rect 1801 71907 1851 71931
rect 136947 71965 136997 71989
rect 136947 71931 136955 71965
rect 136989 71931 136997 71965
rect 136947 71907 136997 71931
rect 1801 71629 1851 71653
rect 1801 71595 1809 71629
rect 1843 71595 1851 71629
rect 1801 71571 1851 71595
rect 136947 71629 136997 71653
rect 136947 71595 136955 71629
rect 136989 71595 136997 71629
rect 136947 71571 136997 71595
rect 1801 71293 1851 71317
rect 1801 71259 1809 71293
rect 1843 71259 1851 71293
rect 1801 71235 1851 71259
rect 136947 71293 136997 71317
rect 136947 71259 136955 71293
rect 136989 71259 136997 71293
rect 136947 71235 136997 71259
rect 1801 70957 1851 70981
rect 1801 70923 1809 70957
rect 1843 70923 1851 70957
rect 1801 70899 1851 70923
rect 136947 70957 136997 70981
rect 136947 70923 136955 70957
rect 136989 70923 136997 70957
rect 136947 70899 136997 70923
rect 1801 70621 1851 70645
rect 1801 70587 1809 70621
rect 1843 70587 1851 70621
rect 1801 70563 1851 70587
rect 136947 70621 136997 70645
rect 136947 70587 136955 70621
rect 136989 70587 136997 70621
rect 136947 70563 136997 70587
rect 1801 70285 1851 70309
rect 1801 70251 1809 70285
rect 1843 70251 1851 70285
rect 1801 70227 1851 70251
rect 136947 70285 136997 70309
rect 136947 70251 136955 70285
rect 136989 70251 136997 70285
rect 136947 70227 136997 70251
rect 1801 69949 1851 69973
rect 1801 69915 1809 69949
rect 1843 69915 1851 69949
rect 1801 69891 1851 69915
rect 136947 69949 136997 69973
rect 136947 69915 136955 69949
rect 136989 69915 136997 69949
rect 136947 69891 136997 69915
rect 1801 69613 1851 69637
rect 1801 69579 1809 69613
rect 1843 69579 1851 69613
rect 1801 69555 1851 69579
rect 136947 69613 136997 69637
rect 136947 69579 136955 69613
rect 136989 69579 136997 69613
rect 136947 69555 136997 69579
rect 1801 69277 1851 69301
rect 1801 69243 1809 69277
rect 1843 69243 1851 69277
rect 1801 69219 1851 69243
rect 136947 69277 136997 69301
rect 136947 69243 136955 69277
rect 136989 69243 136997 69277
rect 136947 69219 136997 69243
rect 1801 68941 1851 68965
rect 1801 68907 1809 68941
rect 1843 68907 1851 68941
rect 1801 68883 1851 68907
rect 136947 68941 136997 68965
rect 136947 68907 136955 68941
rect 136989 68907 136997 68941
rect 136947 68883 136997 68907
rect 1801 68605 1851 68629
rect 1801 68571 1809 68605
rect 1843 68571 1851 68605
rect 1801 68547 1851 68571
rect 136947 68605 136997 68629
rect 136947 68571 136955 68605
rect 136989 68571 136997 68605
rect 136947 68547 136997 68571
rect 1801 68269 1851 68293
rect 1801 68235 1809 68269
rect 1843 68235 1851 68269
rect 1801 68211 1851 68235
rect 136947 68269 136997 68293
rect 136947 68235 136955 68269
rect 136989 68235 136997 68269
rect 136947 68211 136997 68235
rect 1801 67933 1851 67957
rect 1801 67899 1809 67933
rect 1843 67899 1851 67933
rect 1801 67875 1851 67899
rect 136947 67933 136997 67957
rect 136947 67899 136955 67933
rect 136989 67899 136997 67933
rect 136947 67875 136997 67899
rect 1801 67597 1851 67621
rect 1801 67563 1809 67597
rect 1843 67563 1851 67597
rect 1801 67539 1851 67563
rect 136947 67597 136997 67621
rect 136947 67563 136955 67597
rect 136989 67563 136997 67597
rect 136947 67539 136997 67563
rect 1801 67261 1851 67285
rect 1801 67227 1809 67261
rect 1843 67227 1851 67261
rect 1801 67203 1851 67227
rect 136947 67261 136997 67285
rect 136947 67227 136955 67261
rect 136989 67227 136997 67261
rect 136947 67203 136997 67227
rect 1801 66925 1851 66949
rect 1801 66891 1809 66925
rect 1843 66891 1851 66925
rect 1801 66867 1851 66891
rect 136947 66925 136997 66949
rect 136947 66891 136955 66925
rect 136989 66891 136997 66925
rect 136947 66867 136997 66891
rect 1801 66589 1851 66613
rect 1801 66555 1809 66589
rect 1843 66555 1851 66589
rect 1801 66531 1851 66555
rect 136947 66589 136997 66613
rect 136947 66555 136955 66589
rect 136989 66555 136997 66589
rect 136947 66531 136997 66555
rect 1801 66253 1851 66277
rect 1801 66219 1809 66253
rect 1843 66219 1851 66253
rect 1801 66195 1851 66219
rect 136947 66253 136997 66277
rect 136947 66219 136955 66253
rect 136989 66219 136997 66253
rect 136947 66195 136997 66219
rect 1801 65917 1851 65941
rect 1801 65883 1809 65917
rect 1843 65883 1851 65917
rect 1801 65859 1851 65883
rect 136947 65917 136997 65941
rect 136947 65883 136955 65917
rect 136989 65883 136997 65917
rect 136947 65859 136997 65883
rect 1801 65581 1851 65605
rect 1801 65547 1809 65581
rect 1843 65547 1851 65581
rect 1801 65523 1851 65547
rect 136947 65581 136997 65605
rect 136947 65547 136955 65581
rect 136989 65547 136997 65581
rect 136947 65523 136997 65547
rect 1801 65245 1851 65269
rect 1801 65211 1809 65245
rect 1843 65211 1851 65245
rect 1801 65187 1851 65211
rect 136947 65245 136997 65269
rect 136947 65211 136955 65245
rect 136989 65211 136997 65245
rect 136947 65187 136997 65211
rect 1801 64909 1851 64933
rect 1801 64875 1809 64909
rect 1843 64875 1851 64909
rect 1801 64851 1851 64875
rect 136947 64909 136997 64933
rect 136947 64875 136955 64909
rect 136989 64875 136997 64909
rect 136947 64851 136997 64875
rect 1801 64573 1851 64597
rect 1801 64539 1809 64573
rect 1843 64539 1851 64573
rect 1801 64515 1851 64539
rect 136947 64573 136997 64597
rect 136947 64539 136955 64573
rect 136989 64539 136997 64573
rect 136947 64515 136997 64539
rect 1801 64237 1851 64261
rect 1801 64203 1809 64237
rect 1843 64203 1851 64237
rect 1801 64179 1851 64203
rect 136947 64237 136997 64261
rect 136947 64203 136955 64237
rect 136989 64203 136997 64237
rect 136947 64179 136997 64203
rect 1801 63901 1851 63925
rect 1801 63867 1809 63901
rect 1843 63867 1851 63901
rect 1801 63843 1851 63867
rect 136947 63901 136997 63925
rect 136947 63867 136955 63901
rect 136989 63867 136997 63901
rect 136947 63843 136997 63867
rect 1801 63565 1851 63589
rect 1801 63531 1809 63565
rect 1843 63531 1851 63565
rect 1801 63507 1851 63531
rect 136947 63565 136997 63589
rect 136947 63531 136955 63565
rect 136989 63531 136997 63565
rect 136947 63507 136997 63531
rect 1801 63229 1851 63253
rect 1801 63195 1809 63229
rect 1843 63195 1851 63229
rect 1801 63171 1851 63195
rect 136947 63229 136997 63253
rect 136947 63195 136955 63229
rect 136989 63195 136997 63229
rect 136947 63171 136997 63195
rect 1801 62893 1851 62917
rect 1801 62859 1809 62893
rect 1843 62859 1851 62893
rect 1801 62835 1851 62859
rect 136947 62893 136997 62917
rect 136947 62859 136955 62893
rect 136989 62859 136997 62893
rect 136947 62835 136997 62859
rect 1801 62557 1851 62581
rect 1801 62523 1809 62557
rect 1843 62523 1851 62557
rect 1801 62499 1851 62523
rect 136947 62557 136997 62581
rect 136947 62523 136955 62557
rect 136989 62523 136997 62557
rect 136947 62499 136997 62523
rect 1801 62221 1851 62245
rect 1801 62187 1809 62221
rect 1843 62187 1851 62221
rect 1801 62163 1851 62187
rect 136947 62221 136997 62245
rect 136947 62187 136955 62221
rect 136989 62187 136997 62221
rect 136947 62163 136997 62187
rect 1801 61885 1851 61909
rect 1801 61851 1809 61885
rect 1843 61851 1851 61885
rect 1801 61827 1851 61851
rect 136947 61885 136997 61909
rect 136947 61851 136955 61885
rect 136989 61851 136997 61885
rect 136947 61827 136997 61851
rect 1801 61549 1851 61573
rect 1801 61515 1809 61549
rect 1843 61515 1851 61549
rect 1801 61491 1851 61515
rect 136947 61549 136997 61573
rect 136947 61515 136955 61549
rect 136989 61515 136997 61549
rect 136947 61491 136997 61515
rect 1801 61213 1851 61237
rect 1801 61179 1809 61213
rect 1843 61179 1851 61213
rect 1801 61155 1851 61179
rect 136947 61213 136997 61237
rect 136947 61179 136955 61213
rect 136989 61179 136997 61213
rect 136947 61155 136997 61179
rect 1801 60877 1851 60901
rect 1801 60843 1809 60877
rect 1843 60843 1851 60877
rect 1801 60819 1851 60843
rect 136947 60877 136997 60901
rect 136947 60843 136955 60877
rect 136989 60843 136997 60877
rect 136947 60819 136997 60843
rect 1801 60541 1851 60565
rect 1801 60507 1809 60541
rect 1843 60507 1851 60541
rect 1801 60483 1851 60507
rect 136947 60541 136997 60565
rect 136947 60507 136955 60541
rect 136989 60507 136997 60541
rect 136947 60483 136997 60507
rect 1801 60205 1851 60229
rect 1801 60171 1809 60205
rect 1843 60171 1851 60205
rect 1801 60147 1851 60171
rect 136947 60205 136997 60229
rect 136947 60171 136955 60205
rect 136989 60171 136997 60205
rect 136947 60147 136997 60171
rect 1801 59869 1851 59893
rect 1801 59835 1809 59869
rect 1843 59835 1851 59869
rect 1801 59811 1851 59835
rect 136947 59869 136997 59893
rect 136947 59835 136955 59869
rect 136989 59835 136997 59869
rect 136947 59811 136997 59835
rect 1801 59533 1851 59557
rect 1801 59499 1809 59533
rect 1843 59499 1851 59533
rect 1801 59475 1851 59499
rect 136947 59533 136997 59557
rect 136947 59499 136955 59533
rect 136989 59499 136997 59533
rect 136947 59475 136997 59499
rect 1801 59197 1851 59221
rect 1801 59163 1809 59197
rect 1843 59163 1851 59197
rect 1801 59139 1851 59163
rect 136947 59197 136997 59221
rect 136947 59163 136955 59197
rect 136989 59163 136997 59197
rect 136947 59139 136997 59163
rect 1801 58861 1851 58885
rect 1801 58827 1809 58861
rect 1843 58827 1851 58861
rect 1801 58803 1851 58827
rect 136947 58861 136997 58885
rect 136947 58827 136955 58861
rect 136989 58827 136997 58861
rect 136947 58803 136997 58827
rect 1801 58525 1851 58549
rect 1801 58491 1809 58525
rect 1843 58491 1851 58525
rect 1801 58467 1851 58491
rect 136947 58525 136997 58549
rect 136947 58491 136955 58525
rect 136989 58491 136997 58525
rect 136947 58467 136997 58491
rect 1801 58189 1851 58213
rect 1801 58155 1809 58189
rect 1843 58155 1851 58189
rect 1801 58131 1851 58155
rect 136947 58189 136997 58213
rect 136947 58155 136955 58189
rect 136989 58155 136997 58189
rect 136947 58131 136997 58155
rect 1801 57853 1851 57877
rect 1801 57819 1809 57853
rect 1843 57819 1851 57853
rect 1801 57795 1851 57819
rect 136947 57853 136997 57877
rect 136947 57819 136955 57853
rect 136989 57819 136997 57853
rect 136947 57795 136997 57819
rect 1801 57517 1851 57541
rect 1801 57483 1809 57517
rect 1843 57483 1851 57517
rect 1801 57459 1851 57483
rect 136947 57517 136997 57541
rect 136947 57483 136955 57517
rect 136989 57483 136997 57517
rect 136947 57459 136997 57483
rect 1801 57181 1851 57205
rect 1801 57147 1809 57181
rect 1843 57147 1851 57181
rect 1801 57123 1851 57147
rect 136947 57181 136997 57205
rect 136947 57147 136955 57181
rect 136989 57147 136997 57181
rect 136947 57123 136997 57147
rect 1801 56845 1851 56869
rect 1801 56811 1809 56845
rect 1843 56811 1851 56845
rect 1801 56787 1851 56811
rect 136947 56845 136997 56869
rect 136947 56811 136955 56845
rect 136989 56811 136997 56845
rect 136947 56787 136997 56811
rect 1801 56509 1851 56533
rect 1801 56475 1809 56509
rect 1843 56475 1851 56509
rect 1801 56451 1851 56475
rect 136947 56509 136997 56533
rect 136947 56475 136955 56509
rect 136989 56475 136997 56509
rect 136947 56451 136997 56475
rect 1801 56173 1851 56197
rect 1801 56139 1809 56173
rect 1843 56139 1851 56173
rect 1801 56115 1851 56139
rect 136947 56173 136997 56197
rect 136947 56139 136955 56173
rect 136989 56139 136997 56173
rect 136947 56115 136997 56139
rect 1801 55837 1851 55861
rect 1801 55803 1809 55837
rect 1843 55803 1851 55837
rect 1801 55779 1851 55803
rect 136947 55837 136997 55861
rect 136947 55803 136955 55837
rect 136989 55803 136997 55837
rect 136947 55779 136997 55803
rect 1801 55501 1851 55525
rect 1801 55467 1809 55501
rect 1843 55467 1851 55501
rect 1801 55443 1851 55467
rect 136947 55501 136997 55525
rect 136947 55467 136955 55501
rect 136989 55467 136997 55501
rect 136947 55443 136997 55467
rect 1801 55165 1851 55189
rect 1801 55131 1809 55165
rect 1843 55131 1851 55165
rect 1801 55107 1851 55131
rect 136947 55165 136997 55189
rect 136947 55131 136955 55165
rect 136989 55131 136997 55165
rect 136947 55107 136997 55131
rect 1801 54829 1851 54853
rect 1801 54795 1809 54829
rect 1843 54795 1851 54829
rect 1801 54771 1851 54795
rect 136947 54829 136997 54853
rect 136947 54795 136955 54829
rect 136989 54795 136997 54829
rect 136947 54771 136997 54795
rect 1801 54493 1851 54517
rect 1801 54459 1809 54493
rect 1843 54459 1851 54493
rect 1801 54435 1851 54459
rect 136947 54493 136997 54517
rect 136947 54459 136955 54493
rect 136989 54459 136997 54493
rect 136947 54435 136997 54459
rect 1801 54157 1851 54181
rect 1801 54123 1809 54157
rect 1843 54123 1851 54157
rect 1801 54099 1851 54123
rect 136947 54157 136997 54181
rect 136947 54123 136955 54157
rect 136989 54123 136997 54157
rect 136947 54099 136997 54123
rect 1801 53821 1851 53845
rect 1801 53787 1809 53821
rect 1843 53787 1851 53821
rect 1801 53763 1851 53787
rect 136947 53821 136997 53845
rect 136947 53787 136955 53821
rect 136989 53787 136997 53821
rect 136947 53763 136997 53787
rect 1801 53485 1851 53509
rect 1801 53451 1809 53485
rect 1843 53451 1851 53485
rect 1801 53427 1851 53451
rect 136947 53485 136997 53509
rect 136947 53451 136955 53485
rect 136989 53451 136997 53485
rect 136947 53427 136997 53451
rect 1801 53149 1851 53173
rect 1801 53115 1809 53149
rect 1843 53115 1851 53149
rect 1801 53091 1851 53115
rect 136947 53149 136997 53173
rect 136947 53115 136955 53149
rect 136989 53115 136997 53149
rect 136947 53091 136997 53115
rect 1801 52813 1851 52837
rect 1801 52779 1809 52813
rect 1843 52779 1851 52813
rect 1801 52755 1851 52779
rect 136947 52813 136997 52837
rect 136947 52779 136955 52813
rect 136989 52779 136997 52813
rect 136947 52755 136997 52779
rect 1801 52477 1851 52501
rect 1801 52443 1809 52477
rect 1843 52443 1851 52477
rect 1801 52419 1851 52443
rect 136947 52477 136997 52501
rect 136947 52443 136955 52477
rect 136989 52443 136997 52477
rect 136947 52419 136997 52443
rect 1801 52141 1851 52165
rect 1801 52107 1809 52141
rect 1843 52107 1851 52141
rect 1801 52083 1851 52107
rect 136947 52141 136997 52165
rect 136947 52107 136955 52141
rect 136989 52107 136997 52141
rect 136947 52083 136997 52107
rect 1801 51805 1851 51829
rect 1801 51771 1809 51805
rect 1843 51771 1851 51805
rect 1801 51747 1851 51771
rect 136947 51805 136997 51829
rect 136947 51771 136955 51805
rect 136989 51771 136997 51805
rect 136947 51747 136997 51771
rect 1801 51469 1851 51493
rect 1801 51435 1809 51469
rect 1843 51435 1851 51469
rect 1801 51411 1851 51435
rect 136947 51469 136997 51493
rect 136947 51435 136955 51469
rect 136989 51435 136997 51469
rect 136947 51411 136997 51435
rect 1801 51133 1851 51157
rect 1801 51099 1809 51133
rect 1843 51099 1851 51133
rect 1801 51075 1851 51099
rect 136947 51133 136997 51157
rect 136947 51099 136955 51133
rect 136989 51099 136997 51133
rect 136947 51075 136997 51099
rect 1801 50797 1851 50821
rect 1801 50763 1809 50797
rect 1843 50763 1851 50797
rect 1801 50739 1851 50763
rect 136947 50797 136997 50821
rect 136947 50763 136955 50797
rect 136989 50763 136997 50797
rect 136947 50739 136997 50763
rect 1801 50461 1851 50485
rect 1801 50427 1809 50461
rect 1843 50427 1851 50461
rect 1801 50403 1851 50427
rect 136947 50461 136997 50485
rect 136947 50427 136955 50461
rect 136989 50427 136997 50461
rect 136947 50403 136997 50427
rect 1801 50125 1851 50149
rect 1801 50091 1809 50125
rect 1843 50091 1851 50125
rect 1801 50067 1851 50091
rect 136947 50125 136997 50149
rect 136947 50091 136955 50125
rect 136989 50091 136997 50125
rect 136947 50067 136997 50091
rect 1801 49789 1851 49813
rect 1801 49755 1809 49789
rect 1843 49755 1851 49789
rect 1801 49731 1851 49755
rect 136947 49789 136997 49813
rect 136947 49755 136955 49789
rect 136989 49755 136997 49789
rect 136947 49731 136997 49755
rect 1801 49453 1851 49477
rect 1801 49419 1809 49453
rect 1843 49419 1851 49453
rect 1801 49395 1851 49419
rect 136947 49453 136997 49477
rect 136947 49419 136955 49453
rect 136989 49419 136997 49453
rect 136947 49395 136997 49419
rect 1801 49117 1851 49141
rect 1801 49083 1809 49117
rect 1843 49083 1851 49117
rect 1801 49059 1851 49083
rect 136947 49117 136997 49141
rect 136947 49083 136955 49117
rect 136989 49083 136997 49117
rect 136947 49059 136997 49083
rect 1801 48781 1851 48805
rect 1801 48747 1809 48781
rect 1843 48747 1851 48781
rect 1801 48723 1851 48747
rect 136947 48781 136997 48805
rect 136947 48747 136955 48781
rect 136989 48747 136997 48781
rect 136947 48723 136997 48747
rect 1801 48445 1851 48469
rect 1801 48411 1809 48445
rect 1843 48411 1851 48445
rect 1801 48387 1851 48411
rect 136947 48445 136997 48469
rect 136947 48411 136955 48445
rect 136989 48411 136997 48445
rect 136947 48387 136997 48411
rect 1801 48109 1851 48133
rect 1801 48075 1809 48109
rect 1843 48075 1851 48109
rect 1801 48051 1851 48075
rect 136947 48109 136997 48133
rect 136947 48075 136955 48109
rect 136989 48075 136997 48109
rect 136947 48051 136997 48075
rect 1801 47773 1851 47797
rect 1801 47739 1809 47773
rect 1843 47739 1851 47773
rect 1801 47715 1851 47739
rect 136947 47773 136997 47797
rect 136947 47739 136955 47773
rect 136989 47739 136997 47773
rect 136947 47715 136997 47739
rect 1801 47437 1851 47461
rect 1801 47403 1809 47437
rect 1843 47403 1851 47437
rect 1801 47379 1851 47403
rect 136947 47437 136997 47461
rect 136947 47403 136955 47437
rect 136989 47403 136997 47437
rect 136947 47379 136997 47403
rect 1801 47101 1851 47125
rect 1801 47067 1809 47101
rect 1843 47067 1851 47101
rect 1801 47043 1851 47067
rect 136947 47101 136997 47125
rect 136947 47067 136955 47101
rect 136989 47067 136997 47101
rect 136947 47043 136997 47067
rect 1801 46765 1851 46789
rect 1801 46731 1809 46765
rect 1843 46731 1851 46765
rect 1801 46707 1851 46731
rect 136947 46765 136997 46789
rect 136947 46731 136955 46765
rect 136989 46731 136997 46765
rect 136947 46707 136997 46731
rect 1801 46429 1851 46453
rect 1801 46395 1809 46429
rect 1843 46395 1851 46429
rect 1801 46371 1851 46395
rect 136947 46429 136997 46453
rect 136947 46395 136955 46429
rect 136989 46395 136997 46429
rect 136947 46371 136997 46395
rect 1801 46093 1851 46117
rect 1801 46059 1809 46093
rect 1843 46059 1851 46093
rect 1801 46035 1851 46059
rect 136947 46093 136997 46117
rect 136947 46059 136955 46093
rect 136989 46059 136997 46093
rect 136947 46035 136997 46059
rect 1801 45757 1851 45781
rect 1801 45723 1809 45757
rect 1843 45723 1851 45757
rect 1801 45699 1851 45723
rect 136947 45757 136997 45781
rect 136947 45723 136955 45757
rect 136989 45723 136997 45757
rect 136947 45699 136997 45723
rect 1801 45421 1851 45445
rect 1801 45387 1809 45421
rect 1843 45387 1851 45421
rect 1801 45363 1851 45387
rect 136947 45421 136997 45445
rect 136947 45387 136955 45421
rect 136989 45387 136997 45421
rect 136947 45363 136997 45387
rect 1801 45085 1851 45109
rect 1801 45051 1809 45085
rect 1843 45051 1851 45085
rect 1801 45027 1851 45051
rect 136947 45085 136997 45109
rect 136947 45051 136955 45085
rect 136989 45051 136997 45085
rect 136947 45027 136997 45051
rect 1801 44749 1851 44773
rect 1801 44715 1809 44749
rect 1843 44715 1851 44749
rect 1801 44691 1851 44715
rect 136947 44749 136997 44773
rect 136947 44715 136955 44749
rect 136989 44715 136997 44749
rect 136947 44691 136997 44715
rect 1801 44413 1851 44437
rect 1801 44379 1809 44413
rect 1843 44379 1851 44413
rect 1801 44355 1851 44379
rect 136947 44413 136997 44437
rect 136947 44379 136955 44413
rect 136989 44379 136997 44413
rect 136947 44355 136997 44379
rect 1801 44077 1851 44101
rect 1801 44043 1809 44077
rect 1843 44043 1851 44077
rect 1801 44019 1851 44043
rect 136947 44077 136997 44101
rect 136947 44043 136955 44077
rect 136989 44043 136997 44077
rect 136947 44019 136997 44043
rect 1801 43741 1851 43765
rect 1801 43707 1809 43741
rect 1843 43707 1851 43741
rect 1801 43683 1851 43707
rect 136947 43741 136997 43765
rect 136947 43707 136955 43741
rect 136989 43707 136997 43741
rect 136947 43683 136997 43707
rect 1801 43405 1851 43429
rect 1801 43371 1809 43405
rect 1843 43371 1851 43405
rect 1801 43347 1851 43371
rect 136947 43405 136997 43429
rect 136947 43371 136955 43405
rect 136989 43371 136997 43405
rect 136947 43347 136997 43371
rect 1801 43069 1851 43093
rect 1801 43035 1809 43069
rect 1843 43035 1851 43069
rect 1801 43011 1851 43035
rect 136947 43069 136997 43093
rect 136947 43035 136955 43069
rect 136989 43035 136997 43069
rect 136947 43011 136997 43035
rect 1801 42733 1851 42757
rect 1801 42699 1809 42733
rect 1843 42699 1851 42733
rect 1801 42675 1851 42699
rect 136947 42733 136997 42757
rect 136947 42699 136955 42733
rect 136989 42699 136997 42733
rect 136947 42675 136997 42699
rect 1801 42397 1851 42421
rect 1801 42363 1809 42397
rect 1843 42363 1851 42397
rect 1801 42339 1851 42363
rect 136947 42397 136997 42421
rect 136947 42363 136955 42397
rect 136989 42363 136997 42397
rect 136947 42339 136997 42363
rect 1801 42061 1851 42085
rect 1801 42027 1809 42061
rect 1843 42027 1851 42061
rect 1801 42003 1851 42027
rect 136947 42061 136997 42085
rect 136947 42027 136955 42061
rect 136989 42027 136997 42061
rect 136947 42003 136997 42027
rect 1801 41725 1851 41749
rect 1801 41691 1809 41725
rect 1843 41691 1851 41725
rect 1801 41667 1851 41691
rect 136947 41725 136997 41749
rect 136947 41691 136955 41725
rect 136989 41691 136997 41725
rect 136947 41667 136997 41691
rect 1801 41389 1851 41413
rect 1801 41355 1809 41389
rect 1843 41355 1851 41389
rect 1801 41331 1851 41355
rect 136947 41389 136997 41413
rect 136947 41355 136955 41389
rect 136989 41355 136997 41389
rect 136947 41331 136997 41355
rect 1801 41053 1851 41077
rect 1801 41019 1809 41053
rect 1843 41019 1851 41053
rect 1801 40995 1851 41019
rect 136947 41053 136997 41077
rect 136947 41019 136955 41053
rect 136989 41019 136997 41053
rect 136947 40995 136997 41019
rect 1801 40717 1851 40741
rect 1801 40683 1809 40717
rect 1843 40683 1851 40717
rect 1801 40659 1851 40683
rect 136947 40717 136997 40741
rect 136947 40683 136955 40717
rect 136989 40683 136997 40717
rect 136947 40659 136997 40683
rect 1801 40381 1851 40405
rect 1801 40347 1809 40381
rect 1843 40347 1851 40381
rect 1801 40323 1851 40347
rect 136947 40381 136997 40405
rect 136947 40347 136955 40381
rect 136989 40347 136997 40381
rect 136947 40323 136997 40347
rect 1801 40045 1851 40069
rect 1801 40011 1809 40045
rect 1843 40011 1851 40045
rect 1801 39987 1851 40011
rect 136947 40045 136997 40069
rect 136947 40011 136955 40045
rect 136989 40011 136997 40045
rect 136947 39987 136997 40011
rect 1801 39709 1851 39733
rect 1801 39675 1809 39709
rect 1843 39675 1851 39709
rect 1801 39651 1851 39675
rect 136947 39709 136997 39733
rect 136947 39675 136955 39709
rect 136989 39675 136997 39709
rect 136947 39651 136997 39675
rect 1801 39373 1851 39397
rect 1801 39339 1809 39373
rect 1843 39339 1851 39373
rect 1801 39315 1851 39339
rect 136947 39373 136997 39397
rect 136947 39339 136955 39373
rect 136989 39339 136997 39373
rect 136947 39315 136997 39339
rect 1801 39037 1851 39061
rect 1801 39003 1809 39037
rect 1843 39003 1851 39037
rect 1801 38979 1851 39003
rect 136947 39037 136997 39061
rect 136947 39003 136955 39037
rect 136989 39003 136997 39037
rect 136947 38979 136997 39003
rect 1801 38701 1851 38725
rect 1801 38667 1809 38701
rect 1843 38667 1851 38701
rect 1801 38643 1851 38667
rect 136947 38701 136997 38725
rect 136947 38667 136955 38701
rect 136989 38667 136997 38701
rect 136947 38643 136997 38667
rect 1801 38365 1851 38389
rect 1801 38331 1809 38365
rect 1843 38331 1851 38365
rect 1801 38307 1851 38331
rect 136947 38365 136997 38389
rect 136947 38331 136955 38365
rect 136989 38331 136997 38365
rect 136947 38307 136997 38331
rect 1801 38029 1851 38053
rect 1801 37995 1809 38029
rect 1843 37995 1851 38029
rect 1801 37971 1851 37995
rect 136947 38029 136997 38053
rect 136947 37995 136955 38029
rect 136989 37995 136997 38029
rect 136947 37971 136997 37995
rect 1801 37693 1851 37717
rect 1801 37659 1809 37693
rect 1843 37659 1851 37693
rect 1801 37635 1851 37659
rect 136947 37693 136997 37717
rect 136947 37659 136955 37693
rect 136989 37659 136997 37693
rect 136947 37635 136997 37659
rect 1801 37357 1851 37381
rect 1801 37323 1809 37357
rect 1843 37323 1851 37357
rect 1801 37299 1851 37323
rect 136947 37357 136997 37381
rect 136947 37323 136955 37357
rect 136989 37323 136997 37357
rect 136947 37299 136997 37323
rect 1801 37021 1851 37045
rect 1801 36987 1809 37021
rect 1843 36987 1851 37021
rect 1801 36963 1851 36987
rect 136947 37021 136997 37045
rect 136947 36987 136955 37021
rect 136989 36987 136997 37021
rect 136947 36963 136997 36987
rect 1801 36685 1851 36709
rect 1801 36651 1809 36685
rect 1843 36651 1851 36685
rect 1801 36627 1851 36651
rect 136947 36685 136997 36709
rect 136947 36651 136955 36685
rect 136989 36651 136997 36685
rect 136947 36627 136997 36651
rect 1801 36349 1851 36373
rect 1801 36315 1809 36349
rect 1843 36315 1851 36349
rect 1801 36291 1851 36315
rect 136947 36349 136997 36373
rect 136947 36315 136955 36349
rect 136989 36315 136997 36349
rect 136947 36291 136997 36315
rect 1801 36013 1851 36037
rect 1801 35979 1809 36013
rect 1843 35979 1851 36013
rect 1801 35955 1851 35979
rect 136947 36013 136997 36037
rect 136947 35979 136955 36013
rect 136989 35979 136997 36013
rect 136947 35955 136997 35979
rect 1801 35677 1851 35701
rect 1801 35643 1809 35677
rect 1843 35643 1851 35677
rect 1801 35619 1851 35643
rect 136947 35677 136997 35701
rect 136947 35643 136955 35677
rect 136989 35643 136997 35677
rect 136947 35619 136997 35643
rect 1801 35341 1851 35365
rect 1801 35307 1809 35341
rect 1843 35307 1851 35341
rect 1801 35283 1851 35307
rect 136947 35341 136997 35365
rect 136947 35307 136955 35341
rect 136989 35307 136997 35341
rect 136947 35283 136997 35307
rect 1801 35005 1851 35029
rect 1801 34971 1809 35005
rect 1843 34971 1851 35005
rect 1801 34947 1851 34971
rect 136947 35005 136997 35029
rect 136947 34971 136955 35005
rect 136989 34971 136997 35005
rect 136947 34947 136997 34971
rect 1801 34669 1851 34693
rect 1801 34635 1809 34669
rect 1843 34635 1851 34669
rect 1801 34611 1851 34635
rect 136947 34669 136997 34693
rect 136947 34635 136955 34669
rect 136989 34635 136997 34669
rect 136947 34611 136997 34635
rect 1801 34333 1851 34357
rect 1801 34299 1809 34333
rect 1843 34299 1851 34333
rect 1801 34275 1851 34299
rect 136947 34333 136997 34357
rect 136947 34299 136955 34333
rect 136989 34299 136997 34333
rect 136947 34275 136997 34299
rect 1801 33997 1851 34021
rect 1801 33963 1809 33997
rect 1843 33963 1851 33997
rect 1801 33939 1851 33963
rect 136947 33997 136997 34021
rect 136947 33963 136955 33997
rect 136989 33963 136997 33997
rect 136947 33939 136997 33963
rect 1801 33661 1851 33685
rect 1801 33627 1809 33661
rect 1843 33627 1851 33661
rect 1801 33603 1851 33627
rect 136947 33661 136997 33685
rect 136947 33627 136955 33661
rect 136989 33627 136997 33661
rect 136947 33603 136997 33627
rect 1801 33325 1851 33349
rect 1801 33291 1809 33325
rect 1843 33291 1851 33325
rect 1801 33267 1851 33291
rect 136947 33325 136997 33349
rect 136947 33291 136955 33325
rect 136989 33291 136997 33325
rect 136947 33267 136997 33291
rect 1801 32989 1851 33013
rect 1801 32955 1809 32989
rect 1843 32955 1851 32989
rect 1801 32931 1851 32955
rect 136947 32989 136997 33013
rect 136947 32955 136955 32989
rect 136989 32955 136997 32989
rect 136947 32931 136997 32955
rect 1801 32653 1851 32677
rect 1801 32619 1809 32653
rect 1843 32619 1851 32653
rect 1801 32595 1851 32619
rect 136947 32653 136997 32677
rect 136947 32619 136955 32653
rect 136989 32619 136997 32653
rect 136947 32595 136997 32619
rect 1801 32317 1851 32341
rect 1801 32283 1809 32317
rect 1843 32283 1851 32317
rect 1801 32259 1851 32283
rect 136947 32317 136997 32341
rect 136947 32283 136955 32317
rect 136989 32283 136997 32317
rect 136947 32259 136997 32283
rect 1801 31981 1851 32005
rect 1801 31947 1809 31981
rect 1843 31947 1851 31981
rect 1801 31923 1851 31947
rect 136947 31981 136997 32005
rect 136947 31947 136955 31981
rect 136989 31947 136997 31981
rect 136947 31923 136997 31947
rect 1801 31645 1851 31669
rect 1801 31611 1809 31645
rect 1843 31611 1851 31645
rect 1801 31587 1851 31611
rect 136947 31645 136997 31669
rect 136947 31611 136955 31645
rect 136989 31611 136997 31645
rect 136947 31587 136997 31611
rect 1801 31309 1851 31333
rect 1801 31275 1809 31309
rect 1843 31275 1851 31309
rect 1801 31251 1851 31275
rect 136947 31309 136997 31333
rect 136947 31275 136955 31309
rect 136989 31275 136997 31309
rect 136947 31251 136997 31275
rect 1801 30973 1851 30997
rect 1801 30939 1809 30973
rect 1843 30939 1851 30973
rect 1801 30915 1851 30939
rect 136947 30973 136997 30997
rect 136947 30939 136955 30973
rect 136989 30939 136997 30973
rect 136947 30915 136997 30939
rect 1801 30637 1851 30661
rect 1801 30603 1809 30637
rect 1843 30603 1851 30637
rect 1801 30579 1851 30603
rect 136947 30637 136997 30661
rect 136947 30603 136955 30637
rect 136989 30603 136997 30637
rect 136947 30579 136997 30603
rect 1801 30301 1851 30325
rect 1801 30267 1809 30301
rect 1843 30267 1851 30301
rect 1801 30243 1851 30267
rect 136947 30301 136997 30325
rect 136947 30267 136955 30301
rect 136989 30267 136997 30301
rect 136947 30243 136997 30267
rect 1801 29965 1851 29989
rect 1801 29931 1809 29965
rect 1843 29931 1851 29965
rect 1801 29907 1851 29931
rect 136947 29965 136997 29989
rect 136947 29931 136955 29965
rect 136989 29931 136997 29965
rect 136947 29907 136997 29931
rect 1801 29629 1851 29653
rect 1801 29595 1809 29629
rect 1843 29595 1851 29629
rect 1801 29571 1851 29595
rect 136947 29629 136997 29653
rect 136947 29595 136955 29629
rect 136989 29595 136997 29629
rect 136947 29571 136997 29595
rect 1801 29293 1851 29317
rect 1801 29259 1809 29293
rect 1843 29259 1851 29293
rect 1801 29235 1851 29259
rect 136947 29293 136997 29317
rect 136947 29259 136955 29293
rect 136989 29259 136997 29293
rect 136947 29235 136997 29259
rect 1801 28957 1851 28981
rect 1801 28923 1809 28957
rect 1843 28923 1851 28957
rect 1801 28899 1851 28923
rect 136947 28957 136997 28981
rect 136947 28923 136955 28957
rect 136989 28923 136997 28957
rect 136947 28899 136997 28923
rect 1801 28621 1851 28645
rect 1801 28587 1809 28621
rect 1843 28587 1851 28621
rect 1801 28563 1851 28587
rect 136947 28621 136997 28645
rect 136947 28587 136955 28621
rect 136989 28587 136997 28621
rect 136947 28563 136997 28587
rect 1801 28285 1851 28309
rect 1801 28251 1809 28285
rect 1843 28251 1851 28285
rect 1801 28227 1851 28251
rect 136947 28285 136997 28309
rect 136947 28251 136955 28285
rect 136989 28251 136997 28285
rect 136947 28227 136997 28251
rect 1801 27949 1851 27973
rect 1801 27915 1809 27949
rect 1843 27915 1851 27949
rect 1801 27891 1851 27915
rect 136947 27949 136997 27973
rect 136947 27915 136955 27949
rect 136989 27915 136997 27949
rect 136947 27891 136997 27915
rect 1801 27613 1851 27637
rect 1801 27579 1809 27613
rect 1843 27579 1851 27613
rect 1801 27555 1851 27579
rect 136947 27613 136997 27637
rect 136947 27579 136955 27613
rect 136989 27579 136997 27613
rect 136947 27555 136997 27579
rect 1801 27277 1851 27301
rect 1801 27243 1809 27277
rect 1843 27243 1851 27277
rect 1801 27219 1851 27243
rect 136947 27277 136997 27301
rect 136947 27243 136955 27277
rect 136989 27243 136997 27277
rect 136947 27219 136997 27243
rect 1801 26941 1851 26965
rect 1801 26907 1809 26941
rect 1843 26907 1851 26941
rect 1801 26883 1851 26907
rect 136947 26941 136997 26965
rect 136947 26907 136955 26941
rect 136989 26907 136997 26941
rect 136947 26883 136997 26907
rect 1801 26605 1851 26629
rect 1801 26571 1809 26605
rect 1843 26571 1851 26605
rect 1801 26547 1851 26571
rect 136947 26605 136997 26629
rect 136947 26571 136955 26605
rect 136989 26571 136997 26605
rect 136947 26547 136997 26571
rect 1801 26269 1851 26293
rect 1801 26235 1809 26269
rect 1843 26235 1851 26269
rect 1801 26211 1851 26235
rect 136947 26269 136997 26293
rect 136947 26235 136955 26269
rect 136989 26235 136997 26269
rect 136947 26211 136997 26235
rect 1801 25933 1851 25957
rect 1801 25899 1809 25933
rect 1843 25899 1851 25933
rect 1801 25875 1851 25899
rect 136947 25933 136997 25957
rect 136947 25899 136955 25933
rect 136989 25899 136997 25933
rect 136947 25875 136997 25899
rect 1801 25597 1851 25621
rect 1801 25563 1809 25597
rect 1843 25563 1851 25597
rect 1801 25539 1851 25563
rect 136947 25597 136997 25621
rect 136947 25563 136955 25597
rect 136989 25563 136997 25597
rect 136947 25539 136997 25563
rect 1801 25261 1851 25285
rect 1801 25227 1809 25261
rect 1843 25227 1851 25261
rect 1801 25203 1851 25227
rect 136947 25261 136997 25285
rect 136947 25227 136955 25261
rect 136989 25227 136997 25261
rect 136947 25203 136997 25227
rect 1801 24925 1851 24949
rect 1801 24891 1809 24925
rect 1843 24891 1851 24925
rect 1801 24867 1851 24891
rect 136947 24925 136997 24949
rect 136947 24891 136955 24925
rect 136989 24891 136997 24925
rect 136947 24867 136997 24891
rect 1801 24589 1851 24613
rect 1801 24555 1809 24589
rect 1843 24555 1851 24589
rect 1801 24531 1851 24555
rect 136947 24589 136997 24613
rect 136947 24555 136955 24589
rect 136989 24555 136997 24589
rect 136947 24531 136997 24555
rect 1801 24253 1851 24277
rect 1801 24219 1809 24253
rect 1843 24219 1851 24253
rect 1801 24195 1851 24219
rect 136947 24253 136997 24277
rect 136947 24219 136955 24253
rect 136989 24219 136997 24253
rect 136947 24195 136997 24219
rect 1801 23917 1851 23941
rect 1801 23883 1809 23917
rect 1843 23883 1851 23917
rect 1801 23859 1851 23883
rect 136947 23917 136997 23941
rect 136947 23883 136955 23917
rect 136989 23883 136997 23917
rect 136947 23859 136997 23883
rect 1801 23581 1851 23605
rect 1801 23547 1809 23581
rect 1843 23547 1851 23581
rect 1801 23523 1851 23547
rect 136947 23581 136997 23605
rect 136947 23547 136955 23581
rect 136989 23547 136997 23581
rect 136947 23523 136997 23547
rect 1801 23245 1851 23269
rect 1801 23211 1809 23245
rect 1843 23211 1851 23245
rect 1801 23187 1851 23211
rect 136947 23245 136997 23269
rect 136947 23211 136955 23245
rect 136989 23211 136997 23245
rect 136947 23187 136997 23211
rect 1801 22909 1851 22933
rect 1801 22875 1809 22909
rect 1843 22875 1851 22909
rect 1801 22851 1851 22875
rect 136947 22909 136997 22933
rect 136947 22875 136955 22909
rect 136989 22875 136997 22909
rect 136947 22851 136997 22875
rect 1801 22573 1851 22597
rect 1801 22539 1809 22573
rect 1843 22539 1851 22573
rect 1801 22515 1851 22539
rect 136947 22573 136997 22597
rect 136947 22539 136955 22573
rect 136989 22539 136997 22573
rect 136947 22515 136997 22539
rect 1801 22237 1851 22261
rect 1801 22203 1809 22237
rect 1843 22203 1851 22237
rect 1801 22179 1851 22203
rect 136947 22237 136997 22261
rect 136947 22203 136955 22237
rect 136989 22203 136997 22237
rect 136947 22179 136997 22203
rect 1801 21901 1851 21925
rect 1801 21867 1809 21901
rect 1843 21867 1851 21901
rect 1801 21843 1851 21867
rect 136947 21901 136997 21925
rect 136947 21867 136955 21901
rect 136989 21867 136997 21901
rect 136947 21843 136997 21867
rect 1801 21565 1851 21589
rect 1801 21531 1809 21565
rect 1843 21531 1851 21565
rect 1801 21507 1851 21531
rect 136947 21565 136997 21589
rect 136947 21531 136955 21565
rect 136989 21531 136997 21565
rect 136947 21507 136997 21531
rect 1801 21229 1851 21253
rect 1801 21195 1809 21229
rect 1843 21195 1851 21229
rect 1801 21171 1851 21195
rect 136947 21229 136997 21253
rect 136947 21195 136955 21229
rect 136989 21195 136997 21229
rect 136947 21171 136997 21195
rect 1801 20893 1851 20917
rect 1801 20859 1809 20893
rect 1843 20859 1851 20893
rect 1801 20835 1851 20859
rect 136947 20893 136997 20917
rect 136947 20859 136955 20893
rect 136989 20859 136997 20893
rect 136947 20835 136997 20859
rect 1801 20557 1851 20581
rect 1801 20523 1809 20557
rect 1843 20523 1851 20557
rect 1801 20499 1851 20523
rect 136947 20557 136997 20581
rect 136947 20523 136955 20557
rect 136989 20523 136997 20557
rect 136947 20499 136997 20523
rect 1801 20221 1851 20245
rect 1801 20187 1809 20221
rect 1843 20187 1851 20221
rect 1801 20163 1851 20187
rect 136947 20221 136997 20245
rect 136947 20187 136955 20221
rect 136989 20187 136997 20221
rect 136947 20163 136997 20187
rect 1801 19885 1851 19909
rect 1801 19851 1809 19885
rect 1843 19851 1851 19885
rect 1801 19827 1851 19851
rect 136947 19885 136997 19909
rect 136947 19851 136955 19885
rect 136989 19851 136997 19885
rect 136947 19827 136997 19851
rect 1801 19549 1851 19573
rect 1801 19515 1809 19549
rect 1843 19515 1851 19549
rect 1801 19491 1851 19515
rect 136947 19549 136997 19573
rect 136947 19515 136955 19549
rect 136989 19515 136997 19549
rect 136947 19491 136997 19515
rect 1801 19213 1851 19237
rect 1801 19179 1809 19213
rect 1843 19179 1851 19213
rect 1801 19155 1851 19179
rect 136947 19213 136997 19237
rect 136947 19179 136955 19213
rect 136989 19179 136997 19213
rect 136947 19155 136997 19179
rect 1801 18877 1851 18901
rect 1801 18843 1809 18877
rect 1843 18843 1851 18877
rect 1801 18819 1851 18843
rect 136947 18877 136997 18901
rect 136947 18843 136955 18877
rect 136989 18843 136997 18877
rect 136947 18819 136997 18843
rect 1801 18541 1851 18565
rect 1801 18507 1809 18541
rect 1843 18507 1851 18541
rect 1801 18483 1851 18507
rect 136947 18541 136997 18565
rect 136947 18507 136955 18541
rect 136989 18507 136997 18541
rect 136947 18483 136997 18507
rect 1801 18205 1851 18229
rect 1801 18171 1809 18205
rect 1843 18171 1851 18205
rect 1801 18147 1851 18171
rect 136947 18205 136997 18229
rect 136947 18171 136955 18205
rect 136989 18171 136997 18205
rect 136947 18147 136997 18171
rect 1801 17869 1851 17893
rect 1801 17835 1809 17869
rect 1843 17835 1851 17869
rect 1801 17811 1851 17835
rect 136947 17869 136997 17893
rect 136947 17835 136955 17869
rect 136989 17835 136997 17869
rect 136947 17811 136997 17835
rect 1801 17533 1851 17557
rect 1801 17499 1809 17533
rect 1843 17499 1851 17533
rect 1801 17475 1851 17499
rect 136947 17533 136997 17557
rect 136947 17499 136955 17533
rect 136989 17499 136997 17533
rect 136947 17475 136997 17499
rect 1801 17197 1851 17221
rect 1801 17163 1809 17197
rect 1843 17163 1851 17197
rect 1801 17139 1851 17163
rect 136947 17197 136997 17221
rect 136947 17163 136955 17197
rect 136989 17163 136997 17197
rect 136947 17139 136997 17163
rect 1801 16861 1851 16885
rect 1801 16827 1809 16861
rect 1843 16827 1851 16861
rect 1801 16803 1851 16827
rect 136947 16861 136997 16885
rect 136947 16827 136955 16861
rect 136989 16827 136997 16861
rect 136947 16803 136997 16827
rect 1801 16525 1851 16549
rect 1801 16491 1809 16525
rect 1843 16491 1851 16525
rect 1801 16467 1851 16491
rect 136947 16525 136997 16549
rect 136947 16491 136955 16525
rect 136989 16491 136997 16525
rect 136947 16467 136997 16491
rect 1801 16189 1851 16213
rect 1801 16155 1809 16189
rect 1843 16155 1851 16189
rect 1801 16131 1851 16155
rect 136947 16189 136997 16213
rect 136947 16155 136955 16189
rect 136989 16155 136997 16189
rect 136947 16131 136997 16155
rect 1801 15853 1851 15877
rect 1801 15819 1809 15853
rect 1843 15819 1851 15853
rect 1801 15795 1851 15819
rect 136947 15853 136997 15877
rect 136947 15819 136955 15853
rect 136989 15819 136997 15853
rect 136947 15795 136997 15819
rect 1801 15517 1851 15541
rect 1801 15483 1809 15517
rect 1843 15483 1851 15517
rect 1801 15459 1851 15483
rect 136947 15517 136997 15541
rect 136947 15483 136955 15517
rect 136989 15483 136997 15517
rect 136947 15459 136997 15483
rect 1801 15181 1851 15205
rect 1801 15147 1809 15181
rect 1843 15147 1851 15181
rect 1801 15123 1851 15147
rect 136947 15181 136997 15205
rect 136947 15147 136955 15181
rect 136989 15147 136997 15181
rect 136947 15123 136997 15147
rect 1801 14845 1851 14869
rect 1801 14811 1809 14845
rect 1843 14811 1851 14845
rect 1801 14787 1851 14811
rect 136947 14845 136997 14869
rect 136947 14811 136955 14845
rect 136989 14811 136997 14845
rect 136947 14787 136997 14811
rect 1801 14509 1851 14533
rect 1801 14475 1809 14509
rect 1843 14475 1851 14509
rect 1801 14451 1851 14475
rect 136947 14509 136997 14533
rect 136947 14475 136955 14509
rect 136989 14475 136997 14509
rect 136947 14451 136997 14475
rect 1801 14173 1851 14197
rect 1801 14139 1809 14173
rect 1843 14139 1851 14173
rect 1801 14115 1851 14139
rect 136947 14173 136997 14197
rect 136947 14139 136955 14173
rect 136989 14139 136997 14173
rect 136947 14115 136997 14139
rect 1801 13837 1851 13861
rect 1801 13803 1809 13837
rect 1843 13803 1851 13837
rect 1801 13779 1851 13803
rect 136947 13837 136997 13861
rect 136947 13803 136955 13837
rect 136989 13803 136997 13837
rect 136947 13779 136997 13803
rect 1801 13501 1851 13525
rect 1801 13467 1809 13501
rect 1843 13467 1851 13501
rect 1801 13443 1851 13467
rect 136947 13501 136997 13525
rect 136947 13467 136955 13501
rect 136989 13467 136997 13501
rect 136947 13443 136997 13467
rect 1801 13165 1851 13189
rect 1801 13131 1809 13165
rect 1843 13131 1851 13165
rect 1801 13107 1851 13131
rect 136947 13165 136997 13189
rect 136947 13131 136955 13165
rect 136989 13131 136997 13165
rect 136947 13107 136997 13131
rect 1801 12829 1851 12853
rect 1801 12795 1809 12829
rect 1843 12795 1851 12829
rect 1801 12771 1851 12795
rect 136947 12829 136997 12853
rect 136947 12795 136955 12829
rect 136989 12795 136997 12829
rect 136947 12771 136997 12795
rect 1801 12493 1851 12517
rect 1801 12459 1809 12493
rect 1843 12459 1851 12493
rect 1801 12435 1851 12459
rect 136947 12493 136997 12517
rect 136947 12459 136955 12493
rect 136989 12459 136997 12493
rect 136947 12435 136997 12459
rect 1801 12157 1851 12181
rect 1801 12123 1809 12157
rect 1843 12123 1851 12157
rect 1801 12099 1851 12123
rect 136947 12157 136997 12181
rect 136947 12123 136955 12157
rect 136989 12123 136997 12157
rect 136947 12099 136997 12123
rect 1801 11821 1851 11845
rect 1801 11787 1809 11821
rect 1843 11787 1851 11821
rect 1801 11763 1851 11787
rect 136947 11821 136997 11845
rect 136947 11787 136955 11821
rect 136989 11787 136997 11821
rect 136947 11763 136997 11787
rect 1801 11485 1851 11509
rect 1801 11451 1809 11485
rect 1843 11451 1851 11485
rect 1801 11427 1851 11451
rect 136947 11485 136997 11509
rect 136947 11451 136955 11485
rect 136989 11451 136997 11485
rect 136947 11427 136997 11451
rect 1801 11149 1851 11173
rect 1801 11115 1809 11149
rect 1843 11115 1851 11149
rect 1801 11091 1851 11115
rect 136947 11149 136997 11173
rect 136947 11115 136955 11149
rect 136989 11115 136997 11149
rect 136947 11091 136997 11115
rect 1801 10813 1851 10837
rect 1801 10779 1809 10813
rect 1843 10779 1851 10813
rect 1801 10755 1851 10779
rect 136947 10813 136997 10837
rect 136947 10779 136955 10813
rect 136989 10779 136997 10813
rect 136947 10755 136997 10779
rect 1801 10477 1851 10501
rect 1801 10443 1809 10477
rect 1843 10443 1851 10477
rect 1801 10419 1851 10443
rect 136947 10477 136997 10501
rect 136947 10443 136955 10477
rect 136989 10443 136997 10477
rect 136947 10419 136997 10443
rect 1801 10141 1851 10165
rect 1801 10107 1809 10141
rect 1843 10107 1851 10141
rect 1801 10083 1851 10107
rect 136947 10141 136997 10165
rect 136947 10107 136955 10141
rect 136989 10107 136997 10141
rect 136947 10083 136997 10107
rect 1801 9805 1851 9829
rect 1801 9771 1809 9805
rect 1843 9771 1851 9805
rect 1801 9747 1851 9771
rect 136947 9805 136997 9829
rect 136947 9771 136955 9805
rect 136989 9771 136997 9805
rect 136947 9747 136997 9771
rect 1801 9469 1851 9493
rect 1801 9435 1809 9469
rect 1843 9435 1851 9469
rect 1801 9411 1851 9435
rect 136947 9469 136997 9493
rect 136947 9435 136955 9469
rect 136989 9435 136997 9469
rect 136947 9411 136997 9435
rect 1801 9133 1851 9157
rect 1801 9099 1809 9133
rect 1843 9099 1851 9133
rect 1801 9075 1851 9099
rect 136947 9133 136997 9157
rect 136947 9099 136955 9133
rect 136989 9099 136997 9133
rect 136947 9075 136997 9099
rect 1801 8797 1851 8821
rect 1801 8763 1809 8797
rect 1843 8763 1851 8797
rect 1801 8739 1851 8763
rect 136947 8797 136997 8821
rect 136947 8763 136955 8797
rect 136989 8763 136997 8797
rect 136947 8739 136997 8763
rect 1801 8461 1851 8485
rect 1801 8427 1809 8461
rect 1843 8427 1851 8461
rect 1801 8403 1851 8427
rect 136947 8461 136997 8485
rect 136947 8427 136955 8461
rect 136989 8427 136997 8461
rect 136947 8403 136997 8427
rect 1801 8125 1851 8149
rect 1801 8091 1809 8125
rect 1843 8091 1851 8125
rect 1801 8067 1851 8091
rect 136947 8125 136997 8149
rect 136947 8091 136955 8125
rect 136989 8091 136997 8125
rect 136947 8067 136997 8091
rect 1801 7789 1851 7813
rect 1801 7755 1809 7789
rect 1843 7755 1851 7789
rect 1801 7731 1851 7755
rect 136947 7789 136997 7813
rect 136947 7755 136955 7789
rect 136989 7755 136997 7789
rect 136947 7731 136997 7755
rect 1801 7453 1851 7477
rect 1801 7419 1809 7453
rect 1843 7419 1851 7453
rect 1801 7395 1851 7419
rect 136947 7453 136997 7477
rect 136947 7419 136955 7453
rect 136989 7419 136997 7453
rect 136947 7395 136997 7419
rect 1801 7117 1851 7141
rect 1801 7083 1809 7117
rect 1843 7083 1851 7117
rect 1801 7059 1851 7083
rect 136947 7117 136997 7141
rect 136947 7083 136955 7117
rect 136989 7083 136997 7117
rect 136947 7059 136997 7083
rect 1801 6781 1851 6805
rect 1801 6747 1809 6781
rect 1843 6747 1851 6781
rect 1801 6723 1851 6747
rect 136947 6781 136997 6805
rect 136947 6747 136955 6781
rect 136989 6747 136997 6781
rect 136947 6723 136997 6747
rect 1801 6445 1851 6469
rect 1801 6411 1809 6445
rect 1843 6411 1851 6445
rect 1801 6387 1851 6411
rect 136947 6445 136997 6469
rect 136947 6411 136955 6445
rect 136989 6411 136997 6445
rect 136947 6387 136997 6411
rect 1801 6109 1851 6133
rect 1801 6075 1809 6109
rect 1843 6075 1851 6109
rect 1801 6051 1851 6075
rect 136947 6109 136997 6133
rect 136947 6075 136955 6109
rect 136989 6075 136997 6109
rect 136947 6051 136997 6075
rect 1801 5773 1851 5797
rect 1801 5739 1809 5773
rect 1843 5739 1851 5773
rect 1801 5715 1851 5739
rect 136947 5773 136997 5797
rect 136947 5739 136955 5773
rect 136989 5739 136997 5773
rect 136947 5715 136997 5739
rect 1801 5437 1851 5461
rect 1801 5403 1809 5437
rect 1843 5403 1851 5437
rect 1801 5379 1851 5403
rect 136947 5437 136997 5461
rect 136947 5403 136955 5437
rect 136989 5403 136997 5437
rect 136947 5379 136997 5403
rect 1801 5101 1851 5125
rect 1801 5067 1809 5101
rect 1843 5067 1851 5101
rect 1801 5043 1851 5067
rect 136947 5101 136997 5125
rect 136947 5067 136955 5101
rect 136989 5067 136997 5101
rect 136947 5043 136997 5067
rect 1801 4765 1851 4789
rect 1801 4731 1809 4765
rect 1843 4731 1851 4765
rect 1801 4707 1851 4731
rect 136947 4765 136997 4789
rect 136947 4731 136955 4765
rect 136989 4731 136997 4765
rect 136947 4707 136997 4731
rect 1801 4429 1851 4453
rect 1801 4395 1809 4429
rect 1843 4395 1851 4429
rect 1801 4371 1851 4395
rect 136947 4429 136997 4453
rect 136947 4395 136955 4429
rect 136989 4395 136997 4429
rect 136947 4371 136997 4395
rect 1801 4093 1851 4117
rect 1801 4059 1809 4093
rect 1843 4059 1851 4093
rect 1801 4035 1851 4059
rect 136947 4093 136997 4117
rect 136947 4059 136955 4093
rect 136989 4059 136997 4093
rect 136947 4035 136997 4059
rect 1801 3757 1851 3781
rect 1801 3723 1809 3757
rect 1843 3723 1851 3757
rect 1801 3699 1851 3723
rect 136947 3757 136997 3781
rect 136947 3723 136955 3757
rect 136989 3723 136997 3757
rect 136947 3699 136997 3723
rect 1801 3421 1851 3445
rect 1801 3387 1809 3421
rect 1843 3387 1851 3421
rect 1801 3363 1851 3387
rect 136947 3421 136997 3445
rect 136947 3387 136955 3421
rect 136989 3387 136997 3421
rect 136947 3363 136997 3387
rect 1801 3085 1851 3109
rect 1801 3051 1809 3085
rect 1843 3051 1851 3085
rect 1801 3027 1851 3051
rect 136947 3085 136997 3109
rect 136947 3051 136955 3085
rect 136989 3051 136997 3085
rect 136947 3027 136997 3051
rect 1801 2749 1851 2773
rect 1801 2715 1809 2749
rect 1843 2715 1851 2749
rect 1801 2691 1851 2715
rect 136947 2749 136997 2773
rect 136947 2715 136955 2749
rect 136989 2715 136997 2749
rect 136947 2691 136997 2715
rect 1801 2413 1851 2437
rect 1801 2379 1809 2413
rect 1843 2379 1851 2413
rect 1801 2355 1851 2379
rect 136947 2413 136997 2437
rect 136947 2379 136955 2413
rect 136989 2379 136997 2413
rect 136947 2355 136997 2379
rect 1801 2077 1851 2101
rect 1801 2043 1809 2077
rect 1843 2043 1851 2077
rect 1801 2019 1851 2043
rect 136947 2077 136997 2101
rect 136947 2043 136955 2077
rect 136989 2043 136997 2077
rect 136947 2019 136997 2043
rect 2137 1741 2187 1765
rect 2137 1707 2145 1741
rect 2179 1707 2187 1741
rect 2137 1683 2187 1707
rect 2473 1741 2523 1765
rect 2473 1707 2481 1741
rect 2515 1707 2523 1741
rect 2473 1683 2523 1707
rect 2809 1741 2859 1765
rect 2809 1707 2817 1741
rect 2851 1707 2859 1741
rect 2809 1683 2859 1707
rect 3145 1741 3195 1765
rect 3145 1707 3153 1741
rect 3187 1707 3195 1741
rect 3145 1683 3195 1707
rect 3481 1741 3531 1765
rect 3481 1707 3489 1741
rect 3523 1707 3531 1741
rect 3481 1683 3531 1707
rect 3817 1741 3867 1765
rect 3817 1707 3825 1741
rect 3859 1707 3867 1741
rect 3817 1683 3867 1707
rect 4153 1741 4203 1765
rect 4153 1707 4161 1741
rect 4195 1707 4203 1741
rect 4153 1683 4203 1707
rect 4489 1741 4539 1765
rect 4489 1707 4497 1741
rect 4531 1707 4539 1741
rect 4489 1683 4539 1707
rect 4825 1741 4875 1765
rect 4825 1707 4833 1741
rect 4867 1707 4875 1741
rect 4825 1683 4875 1707
rect 5161 1741 5211 1765
rect 5161 1707 5169 1741
rect 5203 1707 5211 1741
rect 5161 1683 5211 1707
rect 5497 1741 5547 1765
rect 5497 1707 5505 1741
rect 5539 1707 5547 1741
rect 5497 1683 5547 1707
rect 5833 1741 5883 1765
rect 5833 1707 5841 1741
rect 5875 1707 5883 1741
rect 5833 1683 5883 1707
rect 6169 1741 6219 1765
rect 6169 1707 6177 1741
rect 6211 1707 6219 1741
rect 6169 1683 6219 1707
rect 6505 1741 6555 1765
rect 6505 1707 6513 1741
rect 6547 1707 6555 1741
rect 6505 1683 6555 1707
rect 6841 1741 6891 1765
rect 6841 1707 6849 1741
rect 6883 1707 6891 1741
rect 6841 1683 6891 1707
rect 7177 1741 7227 1765
rect 7177 1707 7185 1741
rect 7219 1707 7227 1741
rect 7177 1683 7227 1707
rect 7513 1741 7563 1765
rect 7513 1707 7521 1741
rect 7555 1707 7563 1741
rect 7513 1683 7563 1707
rect 7849 1741 7899 1765
rect 7849 1707 7857 1741
rect 7891 1707 7899 1741
rect 7849 1683 7899 1707
rect 8185 1741 8235 1765
rect 8185 1707 8193 1741
rect 8227 1707 8235 1741
rect 8185 1683 8235 1707
rect 8521 1741 8571 1765
rect 8521 1707 8529 1741
rect 8563 1707 8571 1741
rect 8521 1683 8571 1707
rect 8857 1741 8907 1765
rect 8857 1707 8865 1741
rect 8899 1707 8907 1741
rect 8857 1683 8907 1707
rect 9193 1741 9243 1765
rect 9193 1707 9201 1741
rect 9235 1707 9243 1741
rect 9193 1683 9243 1707
rect 9529 1741 9579 1765
rect 9529 1707 9537 1741
rect 9571 1707 9579 1741
rect 9529 1683 9579 1707
rect 9865 1741 9915 1765
rect 9865 1707 9873 1741
rect 9907 1707 9915 1741
rect 9865 1683 9915 1707
rect 10201 1741 10251 1765
rect 10201 1707 10209 1741
rect 10243 1707 10251 1741
rect 10201 1683 10251 1707
rect 10537 1741 10587 1765
rect 10537 1707 10545 1741
rect 10579 1707 10587 1741
rect 10537 1683 10587 1707
rect 10873 1741 10923 1765
rect 10873 1707 10881 1741
rect 10915 1707 10923 1741
rect 10873 1683 10923 1707
rect 11209 1741 11259 1765
rect 11209 1707 11217 1741
rect 11251 1707 11259 1741
rect 11209 1683 11259 1707
rect 11545 1741 11595 1765
rect 11545 1707 11553 1741
rect 11587 1707 11595 1741
rect 11545 1683 11595 1707
rect 11881 1741 11931 1765
rect 11881 1707 11889 1741
rect 11923 1707 11931 1741
rect 11881 1683 11931 1707
rect 12217 1741 12267 1765
rect 12217 1707 12225 1741
rect 12259 1707 12267 1741
rect 12217 1683 12267 1707
rect 12553 1741 12603 1765
rect 12553 1707 12561 1741
rect 12595 1707 12603 1741
rect 12553 1683 12603 1707
rect 12889 1741 12939 1765
rect 12889 1707 12897 1741
rect 12931 1707 12939 1741
rect 12889 1683 12939 1707
rect 13225 1741 13275 1765
rect 13225 1707 13233 1741
rect 13267 1707 13275 1741
rect 13225 1683 13275 1707
rect 13561 1741 13611 1765
rect 13561 1707 13569 1741
rect 13603 1707 13611 1741
rect 13561 1683 13611 1707
rect 13897 1741 13947 1765
rect 13897 1707 13905 1741
rect 13939 1707 13947 1741
rect 13897 1683 13947 1707
rect 14233 1741 14283 1765
rect 14233 1707 14241 1741
rect 14275 1707 14283 1741
rect 14233 1683 14283 1707
rect 14569 1741 14619 1765
rect 14569 1707 14577 1741
rect 14611 1707 14619 1741
rect 14569 1683 14619 1707
rect 14905 1741 14955 1765
rect 14905 1707 14913 1741
rect 14947 1707 14955 1741
rect 14905 1683 14955 1707
rect 15241 1741 15291 1765
rect 15241 1707 15249 1741
rect 15283 1707 15291 1741
rect 15241 1683 15291 1707
rect 15577 1741 15627 1765
rect 15577 1707 15585 1741
rect 15619 1707 15627 1741
rect 15577 1683 15627 1707
rect 15913 1741 15963 1765
rect 15913 1707 15921 1741
rect 15955 1707 15963 1741
rect 15913 1683 15963 1707
rect 16249 1741 16299 1765
rect 16249 1707 16257 1741
rect 16291 1707 16299 1741
rect 16249 1683 16299 1707
rect 16585 1741 16635 1765
rect 16585 1707 16593 1741
rect 16627 1707 16635 1741
rect 16585 1683 16635 1707
rect 16921 1741 16971 1765
rect 16921 1707 16929 1741
rect 16963 1707 16971 1741
rect 16921 1683 16971 1707
rect 17257 1741 17307 1765
rect 17257 1707 17265 1741
rect 17299 1707 17307 1741
rect 17257 1683 17307 1707
rect 17593 1741 17643 1765
rect 17593 1707 17601 1741
rect 17635 1707 17643 1741
rect 17593 1683 17643 1707
rect 17929 1741 17979 1765
rect 17929 1707 17937 1741
rect 17971 1707 17979 1741
rect 17929 1683 17979 1707
rect 18265 1741 18315 1765
rect 18265 1707 18273 1741
rect 18307 1707 18315 1741
rect 18265 1683 18315 1707
rect 18601 1741 18651 1765
rect 18601 1707 18609 1741
rect 18643 1707 18651 1741
rect 18601 1683 18651 1707
rect 18937 1741 18987 1765
rect 18937 1707 18945 1741
rect 18979 1707 18987 1741
rect 18937 1683 18987 1707
rect 19273 1741 19323 1765
rect 19273 1707 19281 1741
rect 19315 1707 19323 1741
rect 19273 1683 19323 1707
rect 19609 1741 19659 1765
rect 19609 1707 19617 1741
rect 19651 1707 19659 1741
rect 19609 1683 19659 1707
rect 19945 1741 19995 1765
rect 19945 1707 19953 1741
rect 19987 1707 19995 1741
rect 19945 1683 19995 1707
rect 20281 1741 20331 1765
rect 20281 1707 20289 1741
rect 20323 1707 20331 1741
rect 20281 1683 20331 1707
rect 20617 1741 20667 1765
rect 20617 1707 20625 1741
rect 20659 1707 20667 1741
rect 20617 1683 20667 1707
rect 20953 1741 21003 1765
rect 20953 1707 20961 1741
rect 20995 1707 21003 1741
rect 20953 1683 21003 1707
rect 21289 1741 21339 1765
rect 21289 1707 21297 1741
rect 21331 1707 21339 1741
rect 21289 1683 21339 1707
rect 21625 1741 21675 1765
rect 21625 1707 21633 1741
rect 21667 1707 21675 1741
rect 21625 1683 21675 1707
rect 21961 1741 22011 1765
rect 21961 1707 21969 1741
rect 22003 1707 22011 1741
rect 21961 1683 22011 1707
rect 22297 1741 22347 1765
rect 22297 1707 22305 1741
rect 22339 1707 22347 1741
rect 22297 1683 22347 1707
rect 22633 1741 22683 1765
rect 22633 1707 22641 1741
rect 22675 1707 22683 1741
rect 22633 1683 22683 1707
rect 22969 1741 23019 1765
rect 22969 1707 22977 1741
rect 23011 1707 23019 1741
rect 22969 1683 23019 1707
rect 23305 1741 23355 1765
rect 23305 1707 23313 1741
rect 23347 1707 23355 1741
rect 23305 1683 23355 1707
rect 23641 1741 23691 1765
rect 23641 1707 23649 1741
rect 23683 1707 23691 1741
rect 23641 1683 23691 1707
rect 23977 1741 24027 1765
rect 23977 1707 23985 1741
rect 24019 1707 24027 1741
rect 23977 1683 24027 1707
rect 24313 1741 24363 1765
rect 24313 1707 24321 1741
rect 24355 1707 24363 1741
rect 24313 1683 24363 1707
rect 24649 1741 24699 1765
rect 24649 1707 24657 1741
rect 24691 1707 24699 1741
rect 24649 1683 24699 1707
rect 24985 1741 25035 1765
rect 24985 1707 24993 1741
rect 25027 1707 25035 1741
rect 24985 1683 25035 1707
rect 25321 1741 25371 1765
rect 25321 1707 25329 1741
rect 25363 1707 25371 1741
rect 25321 1683 25371 1707
rect 25657 1741 25707 1765
rect 25657 1707 25665 1741
rect 25699 1707 25707 1741
rect 25657 1683 25707 1707
rect 25993 1741 26043 1765
rect 25993 1707 26001 1741
rect 26035 1707 26043 1741
rect 25993 1683 26043 1707
rect 26329 1741 26379 1765
rect 26329 1707 26337 1741
rect 26371 1707 26379 1741
rect 26329 1683 26379 1707
rect 26665 1741 26715 1765
rect 26665 1707 26673 1741
rect 26707 1707 26715 1741
rect 26665 1683 26715 1707
rect 27001 1741 27051 1765
rect 27001 1707 27009 1741
rect 27043 1707 27051 1741
rect 27001 1683 27051 1707
rect 27337 1741 27387 1765
rect 27337 1707 27345 1741
rect 27379 1707 27387 1741
rect 27337 1683 27387 1707
rect 27673 1741 27723 1765
rect 27673 1707 27681 1741
rect 27715 1707 27723 1741
rect 27673 1683 27723 1707
rect 28009 1741 28059 1765
rect 28009 1707 28017 1741
rect 28051 1707 28059 1741
rect 28009 1683 28059 1707
rect 28345 1741 28395 1765
rect 28345 1707 28353 1741
rect 28387 1707 28395 1741
rect 28345 1683 28395 1707
rect 28681 1741 28731 1765
rect 28681 1707 28689 1741
rect 28723 1707 28731 1741
rect 28681 1683 28731 1707
rect 29017 1741 29067 1765
rect 29017 1707 29025 1741
rect 29059 1707 29067 1741
rect 29017 1683 29067 1707
rect 29353 1741 29403 1765
rect 29353 1707 29361 1741
rect 29395 1707 29403 1741
rect 29353 1683 29403 1707
rect 29689 1741 29739 1765
rect 29689 1707 29697 1741
rect 29731 1707 29739 1741
rect 29689 1683 29739 1707
rect 30025 1741 30075 1765
rect 30025 1707 30033 1741
rect 30067 1707 30075 1741
rect 30025 1683 30075 1707
rect 30361 1741 30411 1765
rect 30361 1707 30369 1741
rect 30403 1707 30411 1741
rect 30361 1683 30411 1707
rect 30697 1741 30747 1765
rect 30697 1707 30705 1741
rect 30739 1707 30747 1741
rect 30697 1683 30747 1707
rect 31033 1741 31083 1765
rect 31033 1707 31041 1741
rect 31075 1707 31083 1741
rect 31033 1683 31083 1707
rect 31369 1741 31419 1765
rect 31369 1707 31377 1741
rect 31411 1707 31419 1741
rect 31369 1683 31419 1707
rect 31705 1741 31755 1765
rect 31705 1707 31713 1741
rect 31747 1707 31755 1741
rect 31705 1683 31755 1707
rect 32041 1741 32091 1765
rect 32041 1707 32049 1741
rect 32083 1707 32091 1741
rect 32041 1683 32091 1707
rect 32377 1741 32427 1765
rect 32377 1707 32385 1741
rect 32419 1707 32427 1741
rect 32377 1683 32427 1707
rect 32713 1741 32763 1765
rect 32713 1707 32721 1741
rect 32755 1707 32763 1741
rect 32713 1683 32763 1707
rect 33049 1741 33099 1765
rect 33049 1707 33057 1741
rect 33091 1707 33099 1741
rect 33049 1683 33099 1707
rect 33385 1741 33435 1765
rect 33385 1707 33393 1741
rect 33427 1707 33435 1741
rect 33385 1683 33435 1707
rect 33721 1741 33771 1765
rect 33721 1707 33729 1741
rect 33763 1707 33771 1741
rect 33721 1683 33771 1707
rect 34057 1741 34107 1765
rect 34057 1707 34065 1741
rect 34099 1707 34107 1741
rect 34057 1683 34107 1707
rect 34393 1741 34443 1765
rect 34393 1707 34401 1741
rect 34435 1707 34443 1741
rect 34393 1683 34443 1707
rect 34729 1741 34779 1765
rect 34729 1707 34737 1741
rect 34771 1707 34779 1741
rect 34729 1683 34779 1707
rect 35065 1741 35115 1765
rect 35065 1707 35073 1741
rect 35107 1707 35115 1741
rect 35065 1683 35115 1707
rect 35401 1741 35451 1765
rect 35401 1707 35409 1741
rect 35443 1707 35451 1741
rect 35401 1683 35451 1707
rect 35737 1741 35787 1765
rect 35737 1707 35745 1741
rect 35779 1707 35787 1741
rect 35737 1683 35787 1707
rect 36073 1741 36123 1765
rect 36073 1707 36081 1741
rect 36115 1707 36123 1741
rect 36073 1683 36123 1707
rect 36409 1741 36459 1765
rect 36409 1707 36417 1741
rect 36451 1707 36459 1741
rect 36409 1683 36459 1707
rect 36745 1741 36795 1765
rect 36745 1707 36753 1741
rect 36787 1707 36795 1741
rect 36745 1683 36795 1707
rect 37081 1741 37131 1765
rect 37081 1707 37089 1741
rect 37123 1707 37131 1741
rect 37081 1683 37131 1707
rect 37417 1741 37467 1765
rect 37417 1707 37425 1741
rect 37459 1707 37467 1741
rect 37417 1683 37467 1707
rect 37753 1741 37803 1765
rect 37753 1707 37761 1741
rect 37795 1707 37803 1741
rect 37753 1683 37803 1707
rect 38089 1741 38139 1765
rect 38089 1707 38097 1741
rect 38131 1707 38139 1741
rect 38089 1683 38139 1707
rect 38425 1741 38475 1765
rect 38425 1707 38433 1741
rect 38467 1707 38475 1741
rect 38425 1683 38475 1707
rect 38761 1741 38811 1765
rect 38761 1707 38769 1741
rect 38803 1707 38811 1741
rect 38761 1683 38811 1707
rect 39097 1741 39147 1765
rect 39097 1707 39105 1741
rect 39139 1707 39147 1741
rect 39097 1683 39147 1707
rect 39433 1741 39483 1765
rect 39433 1707 39441 1741
rect 39475 1707 39483 1741
rect 39433 1683 39483 1707
rect 39769 1741 39819 1765
rect 39769 1707 39777 1741
rect 39811 1707 39819 1741
rect 39769 1683 39819 1707
rect 40105 1741 40155 1765
rect 40105 1707 40113 1741
rect 40147 1707 40155 1741
rect 40105 1683 40155 1707
rect 40441 1741 40491 1765
rect 40441 1707 40449 1741
rect 40483 1707 40491 1741
rect 40441 1683 40491 1707
rect 40777 1741 40827 1765
rect 40777 1707 40785 1741
rect 40819 1707 40827 1741
rect 40777 1683 40827 1707
rect 41113 1741 41163 1765
rect 41113 1707 41121 1741
rect 41155 1707 41163 1741
rect 41113 1683 41163 1707
rect 41449 1741 41499 1765
rect 41449 1707 41457 1741
rect 41491 1707 41499 1741
rect 41449 1683 41499 1707
rect 41785 1741 41835 1765
rect 41785 1707 41793 1741
rect 41827 1707 41835 1741
rect 41785 1683 41835 1707
rect 42121 1741 42171 1765
rect 42121 1707 42129 1741
rect 42163 1707 42171 1741
rect 42121 1683 42171 1707
rect 42457 1741 42507 1765
rect 42457 1707 42465 1741
rect 42499 1707 42507 1741
rect 42457 1683 42507 1707
rect 42793 1741 42843 1765
rect 42793 1707 42801 1741
rect 42835 1707 42843 1741
rect 42793 1683 42843 1707
rect 43129 1741 43179 1765
rect 43129 1707 43137 1741
rect 43171 1707 43179 1741
rect 43129 1683 43179 1707
rect 43465 1741 43515 1765
rect 43465 1707 43473 1741
rect 43507 1707 43515 1741
rect 43465 1683 43515 1707
rect 43801 1741 43851 1765
rect 43801 1707 43809 1741
rect 43843 1707 43851 1741
rect 43801 1683 43851 1707
rect 44137 1741 44187 1765
rect 44137 1707 44145 1741
rect 44179 1707 44187 1741
rect 44137 1683 44187 1707
rect 44473 1741 44523 1765
rect 44473 1707 44481 1741
rect 44515 1707 44523 1741
rect 44473 1683 44523 1707
rect 44809 1741 44859 1765
rect 44809 1707 44817 1741
rect 44851 1707 44859 1741
rect 44809 1683 44859 1707
rect 45145 1741 45195 1765
rect 45145 1707 45153 1741
rect 45187 1707 45195 1741
rect 45145 1683 45195 1707
rect 45481 1741 45531 1765
rect 45481 1707 45489 1741
rect 45523 1707 45531 1741
rect 45481 1683 45531 1707
rect 45817 1741 45867 1765
rect 45817 1707 45825 1741
rect 45859 1707 45867 1741
rect 45817 1683 45867 1707
rect 46153 1741 46203 1765
rect 46153 1707 46161 1741
rect 46195 1707 46203 1741
rect 46153 1683 46203 1707
rect 46489 1741 46539 1765
rect 46489 1707 46497 1741
rect 46531 1707 46539 1741
rect 46489 1683 46539 1707
rect 46825 1741 46875 1765
rect 46825 1707 46833 1741
rect 46867 1707 46875 1741
rect 46825 1683 46875 1707
rect 47161 1741 47211 1765
rect 47161 1707 47169 1741
rect 47203 1707 47211 1741
rect 47161 1683 47211 1707
rect 47497 1741 47547 1765
rect 47497 1707 47505 1741
rect 47539 1707 47547 1741
rect 47497 1683 47547 1707
rect 47833 1741 47883 1765
rect 47833 1707 47841 1741
rect 47875 1707 47883 1741
rect 47833 1683 47883 1707
rect 48169 1741 48219 1765
rect 48169 1707 48177 1741
rect 48211 1707 48219 1741
rect 48169 1683 48219 1707
rect 48505 1741 48555 1765
rect 48505 1707 48513 1741
rect 48547 1707 48555 1741
rect 48505 1683 48555 1707
rect 48841 1741 48891 1765
rect 48841 1707 48849 1741
rect 48883 1707 48891 1741
rect 48841 1683 48891 1707
rect 49177 1741 49227 1765
rect 49177 1707 49185 1741
rect 49219 1707 49227 1741
rect 49177 1683 49227 1707
rect 49513 1741 49563 1765
rect 49513 1707 49521 1741
rect 49555 1707 49563 1741
rect 49513 1683 49563 1707
rect 49849 1741 49899 1765
rect 49849 1707 49857 1741
rect 49891 1707 49899 1741
rect 49849 1683 49899 1707
rect 50185 1741 50235 1765
rect 50185 1707 50193 1741
rect 50227 1707 50235 1741
rect 50185 1683 50235 1707
rect 50521 1741 50571 1765
rect 50521 1707 50529 1741
rect 50563 1707 50571 1741
rect 50521 1683 50571 1707
rect 50857 1741 50907 1765
rect 50857 1707 50865 1741
rect 50899 1707 50907 1741
rect 50857 1683 50907 1707
rect 51193 1741 51243 1765
rect 51193 1707 51201 1741
rect 51235 1707 51243 1741
rect 51193 1683 51243 1707
rect 51529 1741 51579 1765
rect 51529 1707 51537 1741
rect 51571 1707 51579 1741
rect 51529 1683 51579 1707
rect 51865 1741 51915 1765
rect 51865 1707 51873 1741
rect 51907 1707 51915 1741
rect 51865 1683 51915 1707
rect 52201 1741 52251 1765
rect 52201 1707 52209 1741
rect 52243 1707 52251 1741
rect 52201 1683 52251 1707
rect 52537 1741 52587 1765
rect 52537 1707 52545 1741
rect 52579 1707 52587 1741
rect 52537 1683 52587 1707
rect 52873 1741 52923 1765
rect 52873 1707 52881 1741
rect 52915 1707 52923 1741
rect 52873 1683 52923 1707
rect 53209 1741 53259 1765
rect 53209 1707 53217 1741
rect 53251 1707 53259 1741
rect 53209 1683 53259 1707
rect 53545 1741 53595 1765
rect 53545 1707 53553 1741
rect 53587 1707 53595 1741
rect 53545 1683 53595 1707
rect 53881 1741 53931 1765
rect 53881 1707 53889 1741
rect 53923 1707 53931 1741
rect 53881 1683 53931 1707
rect 54217 1741 54267 1765
rect 54217 1707 54225 1741
rect 54259 1707 54267 1741
rect 54217 1683 54267 1707
rect 54553 1741 54603 1765
rect 54553 1707 54561 1741
rect 54595 1707 54603 1741
rect 54553 1683 54603 1707
rect 54889 1741 54939 1765
rect 54889 1707 54897 1741
rect 54931 1707 54939 1741
rect 54889 1683 54939 1707
rect 55225 1741 55275 1765
rect 55225 1707 55233 1741
rect 55267 1707 55275 1741
rect 55225 1683 55275 1707
rect 55561 1741 55611 1765
rect 55561 1707 55569 1741
rect 55603 1707 55611 1741
rect 55561 1683 55611 1707
rect 55897 1741 55947 1765
rect 55897 1707 55905 1741
rect 55939 1707 55947 1741
rect 55897 1683 55947 1707
rect 56233 1741 56283 1765
rect 56233 1707 56241 1741
rect 56275 1707 56283 1741
rect 56233 1683 56283 1707
rect 56569 1741 56619 1765
rect 56569 1707 56577 1741
rect 56611 1707 56619 1741
rect 56569 1683 56619 1707
rect 56905 1741 56955 1765
rect 56905 1707 56913 1741
rect 56947 1707 56955 1741
rect 56905 1683 56955 1707
rect 57241 1741 57291 1765
rect 57241 1707 57249 1741
rect 57283 1707 57291 1741
rect 57241 1683 57291 1707
rect 57577 1741 57627 1765
rect 57577 1707 57585 1741
rect 57619 1707 57627 1741
rect 57577 1683 57627 1707
rect 57913 1741 57963 1765
rect 57913 1707 57921 1741
rect 57955 1707 57963 1741
rect 57913 1683 57963 1707
rect 58249 1741 58299 1765
rect 58249 1707 58257 1741
rect 58291 1707 58299 1741
rect 58249 1683 58299 1707
rect 58585 1741 58635 1765
rect 58585 1707 58593 1741
rect 58627 1707 58635 1741
rect 58585 1683 58635 1707
rect 58921 1741 58971 1765
rect 58921 1707 58929 1741
rect 58963 1707 58971 1741
rect 58921 1683 58971 1707
rect 59257 1741 59307 1765
rect 59257 1707 59265 1741
rect 59299 1707 59307 1741
rect 59257 1683 59307 1707
rect 59593 1741 59643 1765
rect 59593 1707 59601 1741
rect 59635 1707 59643 1741
rect 59593 1683 59643 1707
rect 59929 1741 59979 1765
rect 59929 1707 59937 1741
rect 59971 1707 59979 1741
rect 59929 1683 59979 1707
rect 60265 1741 60315 1765
rect 60265 1707 60273 1741
rect 60307 1707 60315 1741
rect 60265 1683 60315 1707
rect 60601 1741 60651 1765
rect 60601 1707 60609 1741
rect 60643 1707 60651 1741
rect 60601 1683 60651 1707
rect 60937 1741 60987 1765
rect 60937 1707 60945 1741
rect 60979 1707 60987 1741
rect 60937 1683 60987 1707
rect 61273 1741 61323 1765
rect 61273 1707 61281 1741
rect 61315 1707 61323 1741
rect 61273 1683 61323 1707
rect 61609 1741 61659 1765
rect 61609 1707 61617 1741
rect 61651 1707 61659 1741
rect 61609 1683 61659 1707
rect 61945 1741 61995 1765
rect 61945 1707 61953 1741
rect 61987 1707 61995 1741
rect 61945 1683 61995 1707
rect 62281 1741 62331 1765
rect 62281 1707 62289 1741
rect 62323 1707 62331 1741
rect 62281 1683 62331 1707
rect 62617 1741 62667 1765
rect 62617 1707 62625 1741
rect 62659 1707 62667 1741
rect 62617 1683 62667 1707
rect 62953 1741 63003 1765
rect 62953 1707 62961 1741
rect 62995 1707 63003 1741
rect 62953 1683 63003 1707
rect 63289 1741 63339 1765
rect 63289 1707 63297 1741
rect 63331 1707 63339 1741
rect 63289 1683 63339 1707
rect 63625 1741 63675 1765
rect 63625 1707 63633 1741
rect 63667 1707 63675 1741
rect 63625 1683 63675 1707
rect 63961 1741 64011 1765
rect 63961 1707 63969 1741
rect 64003 1707 64011 1741
rect 63961 1683 64011 1707
rect 64297 1741 64347 1765
rect 64297 1707 64305 1741
rect 64339 1707 64347 1741
rect 64297 1683 64347 1707
rect 64633 1741 64683 1765
rect 64633 1707 64641 1741
rect 64675 1707 64683 1741
rect 64633 1683 64683 1707
rect 64969 1741 65019 1765
rect 64969 1707 64977 1741
rect 65011 1707 65019 1741
rect 64969 1683 65019 1707
rect 65305 1741 65355 1765
rect 65305 1707 65313 1741
rect 65347 1707 65355 1741
rect 65305 1683 65355 1707
rect 65641 1741 65691 1765
rect 65641 1707 65649 1741
rect 65683 1707 65691 1741
rect 65641 1683 65691 1707
rect 65977 1741 66027 1765
rect 65977 1707 65985 1741
rect 66019 1707 66027 1741
rect 65977 1683 66027 1707
rect 66313 1741 66363 1765
rect 66313 1707 66321 1741
rect 66355 1707 66363 1741
rect 66313 1683 66363 1707
rect 66649 1741 66699 1765
rect 66649 1707 66657 1741
rect 66691 1707 66699 1741
rect 66649 1683 66699 1707
rect 66985 1741 67035 1765
rect 66985 1707 66993 1741
rect 67027 1707 67035 1741
rect 66985 1683 67035 1707
rect 67321 1741 67371 1765
rect 67321 1707 67329 1741
rect 67363 1707 67371 1741
rect 67321 1683 67371 1707
rect 67657 1741 67707 1765
rect 67657 1707 67665 1741
rect 67699 1707 67707 1741
rect 67657 1683 67707 1707
rect 67993 1741 68043 1765
rect 67993 1707 68001 1741
rect 68035 1707 68043 1741
rect 67993 1683 68043 1707
rect 68329 1741 68379 1765
rect 68329 1707 68337 1741
rect 68371 1707 68379 1741
rect 68329 1683 68379 1707
rect 68665 1741 68715 1765
rect 68665 1707 68673 1741
rect 68707 1707 68715 1741
rect 68665 1683 68715 1707
rect 69001 1741 69051 1765
rect 69001 1707 69009 1741
rect 69043 1707 69051 1741
rect 69001 1683 69051 1707
rect 69337 1741 69387 1765
rect 69337 1707 69345 1741
rect 69379 1707 69387 1741
rect 69337 1683 69387 1707
rect 69673 1741 69723 1765
rect 69673 1707 69681 1741
rect 69715 1707 69723 1741
rect 69673 1683 69723 1707
rect 70009 1741 70059 1765
rect 70009 1707 70017 1741
rect 70051 1707 70059 1741
rect 70009 1683 70059 1707
rect 70345 1741 70395 1765
rect 70345 1707 70353 1741
rect 70387 1707 70395 1741
rect 70345 1683 70395 1707
rect 70681 1741 70731 1765
rect 70681 1707 70689 1741
rect 70723 1707 70731 1741
rect 70681 1683 70731 1707
rect 71017 1741 71067 1765
rect 71017 1707 71025 1741
rect 71059 1707 71067 1741
rect 71017 1683 71067 1707
rect 71353 1741 71403 1765
rect 71353 1707 71361 1741
rect 71395 1707 71403 1741
rect 71353 1683 71403 1707
rect 71689 1741 71739 1765
rect 71689 1707 71697 1741
rect 71731 1707 71739 1741
rect 71689 1683 71739 1707
rect 72025 1741 72075 1765
rect 72025 1707 72033 1741
rect 72067 1707 72075 1741
rect 72025 1683 72075 1707
rect 72361 1741 72411 1765
rect 72361 1707 72369 1741
rect 72403 1707 72411 1741
rect 72361 1683 72411 1707
rect 72697 1741 72747 1765
rect 72697 1707 72705 1741
rect 72739 1707 72747 1741
rect 72697 1683 72747 1707
rect 73033 1741 73083 1765
rect 73033 1707 73041 1741
rect 73075 1707 73083 1741
rect 73033 1683 73083 1707
rect 73369 1741 73419 1765
rect 73369 1707 73377 1741
rect 73411 1707 73419 1741
rect 73369 1683 73419 1707
rect 73705 1741 73755 1765
rect 73705 1707 73713 1741
rect 73747 1707 73755 1741
rect 73705 1683 73755 1707
rect 74041 1741 74091 1765
rect 74041 1707 74049 1741
rect 74083 1707 74091 1741
rect 74041 1683 74091 1707
rect 74377 1741 74427 1765
rect 74377 1707 74385 1741
rect 74419 1707 74427 1741
rect 74377 1683 74427 1707
rect 74713 1741 74763 1765
rect 74713 1707 74721 1741
rect 74755 1707 74763 1741
rect 74713 1683 74763 1707
rect 75049 1741 75099 1765
rect 75049 1707 75057 1741
rect 75091 1707 75099 1741
rect 75049 1683 75099 1707
rect 75385 1741 75435 1765
rect 75385 1707 75393 1741
rect 75427 1707 75435 1741
rect 75385 1683 75435 1707
rect 75721 1741 75771 1765
rect 75721 1707 75729 1741
rect 75763 1707 75771 1741
rect 75721 1683 75771 1707
rect 76057 1741 76107 1765
rect 76057 1707 76065 1741
rect 76099 1707 76107 1741
rect 76057 1683 76107 1707
rect 76393 1741 76443 1765
rect 76393 1707 76401 1741
rect 76435 1707 76443 1741
rect 76393 1683 76443 1707
rect 76729 1741 76779 1765
rect 76729 1707 76737 1741
rect 76771 1707 76779 1741
rect 76729 1683 76779 1707
rect 77065 1741 77115 1765
rect 77065 1707 77073 1741
rect 77107 1707 77115 1741
rect 77065 1683 77115 1707
rect 77401 1741 77451 1765
rect 77401 1707 77409 1741
rect 77443 1707 77451 1741
rect 77401 1683 77451 1707
rect 77737 1741 77787 1765
rect 77737 1707 77745 1741
rect 77779 1707 77787 1741
rect 77737 1683 77787 1707
rect 78073 1741 78123 1765
rect 78073 1707 78081 1741
rect 78115 1707 78123 1741
rect 78073 1683 78123 1707
rect 78409 1741 78459 1765
rect 78409 1707 78417 1741
rect 78451 1707 78459 1741
rect 78409 1683 78459 1707
rect 78745 1741 78795 1765
rect 78745 1707 78753 1741
rect 78787 1707 78795 1741
rect 78745 1683 78795 1707
rect 79081 1741 79131 1765
rect 79081 1707 79089 1741
rect 79123 1707 79131 1741
rect 79081 1683 79131 1707
rect 79417 1741 79467 1765
rect 79417 1707 79425 1741
rect 79459 1707 79467 1741
rect 79417 1683 79467 1707
rect 79753 1741 79803 1765
rect 79753 1707 79761 1741
rect 79795 1707 79803 1741
rect 79753 1683 79803 1707
rect 80089 1741 80139 1765
rect 80089 1707 80097 1741
rect 80131 1707 80139 1741
rect 80089 1683 80139 1707
rect 80425 1741 80475 1765
rect 80425 1707 80433 1741
rect 80467 1707 80475 1741
rect 80425 1683 80475 1707
rect 80761 1741 80811 1765
rect 80761 1707 80769 1741
rect 80803 1707 80811 1741
rect 80761 1683 80811 1707
rect 81097 1741 81147 1765
rect 81097 1707 81105 1741
rect 81139 1707 81147 1741
rect 81097 1683 81147 1707
rect 81433 1741 81483 1765
rect 81433 1707 81441 1741
rect 81475 1707 81483 1741
rect 81433 1683 81483 1707
rect 81769 1741 81819 1765
rect 81769 1707 81777 1741
rect 81811 1707 81819 1741
rect 81769 1683 81819 1707
rect 82105 1741 82155 1765
rect 82105 1707 82113 1741
rect 82147 1707 82155 1741
rect 82105 1683 82155 1707
rect 82441 1741 82491 1765
rect 82441 1707 82449 1741
rect 82483 1707 82491 1741
rect 82441 1683 82491 1707
rect 82777 1741 82827 1765
rect 82777 1707 82785 1741
rect 82819 1707 82827 1741
rect 82777 1683 82827 1707
rect 83113 1741 83163 1765
rect 83113 1707 83121 1741
rect 83155 1707 83163 1741
rect 83113 1683 83163 1707
rect 83449 1741 83499 1765
rect 83449 1707 83457 1741
rect 83491 1707 83499 1741
rect 83449 1683 83499 1707
rect 83785 1741 83835 1765
rect 83785 1707 83793 1741
rect 83827 1707 83835 1741
rect 83785 1683 83835 1707
rect 84121 1741 84171 1765
rect 84121 1707 84129 1741
rect 84163 1707 84171 1741
rect 84121 1683 84171 1707
rect 84457 1741 84507 1765
rect 84457 1707 84465 1741
rect 84499 1707 84507 1741
rect 84457 1683 84507 1707
rect 84793 1741 84843 1765
rect 84793 1707 84801 1741
rect 84835 1707 84843 1741
rect 84793 1683 84843 1707
rect 85129 1741 85179 1765
rect 85129 1707 85137 1741
rect 85171 1707 85179 1741
rect 85129 1683 85179 1707
rect 85465 1741 85515 1765
rect 85465 1707 85473 1741
rect 85507 1707 85515 1741
rect 85465 1683 85515 1707
rect 85801 1741 85851 1765
rect 85801 1707 85809 1741
rect 85843 1707 85851 1741
rect 85801 1683 85851 1707
rect 86137 1741 86187 1765
rect 86137 1707 86145 1741
rect 86179 1707 86187 1741
rect 86137 1683 86187 1707
rect 86473 1741 86523 1765
rect 86473 1707 86481 1741
rect 86515 1707 86523 1741
rect 86473 1683 86523 1707
rect 86809 1741 86859 1765
rect 86809 1707 86817 1741
rect 86851 1707 86859 1741
rect 86809 1683 86859 1707
rect 87145 1741 87195 1765
rect 87145 1707 87153 1741
rect 87187 1707 87195 1741
rect 87145 1683 87195 1707
rect 87481 1741 87531 1765
rect 87481 1707 87489 1741
rect 87523 1707 87531 1741
rect 87481 1683 87531 1707
rect 87817 1741 87867 1765
rect 87817 1707 87825 1741
rect 87859 1707 87867 1741
rect 87817 1683 87867 1707
rect 88153 1741 88203 1765
rect 88153 1707 88161 1741
rect 88195 1707 88203 1741
rect 88153 1683 88203 1707
rect 88489 1741 88539 1765
rect 88489 1707 88497 1741
rect 88531 1707 88539 1741
rect 88489 1683 88539 1707
rect 88825 1741 88875 1765
rect 88825 1707 88833 1741
rect 88867 1707 88875 1741
rect 88825 1683 88875 1707
rect 89161 1741 89211 1765
rect 89161 1707 89169 1741
rect 89203 1707 89211 1741
rect 89161 1683 89211 1707
rect 89497 1741 89547 1765
rect 89497 1707 89505 1741
rect 89539 1707 89547 1741
rect 89497 1683 89547 1707
rect 89833 1741 89883 1765
rect 89833 1707 89841 1741
rect 89875 1707 89883 1741
rect 89833 1683 89883 1707
rect 90169 1741 90219 1765
rect 90169 1707 90177 1741
rect 90211 1707 90219 1741
rect 90169 1683 90219 1707
rect 90505 1741 90555 1765
rect 90505 1707 90513 1741
rect 90547 1707 90555 1741
rect 90505 1683 90555 1707
rect 90841 1741 90891 1765
rect 90841 1707 90849 1741
rect 90883 1707 90891 1741
rect 90841 1683 90891 1707
rect 91177 1741 91227 1765
rect 91177 1707 91185 1741
rect 91219 1707 91227 1741
rect 91177 1683 91227 1707
rect 91513 1741 91563 1765
rect 91513 1707 91521 1741
rect 91555 1707 91563 1741
rect 91513 1683 91563 1707
rect 91849 1741 91899 1765
rect 91849 1707 91857 1741
rect 91891 1707 91899 1741
rect 91849 1683 91899 1707
rect 92185 1741 92235 1765
rect 92185 1707 92193 1741
rect 92227 1707 92235 1741
rect 92185 1683 92235 1707
rect 92521 1741 92571 1765
rect 92521 1707 92529 1741
rect 92563 1707 92571 1741
rect 92521 1683 92571 1707
rect 92857 1741 92907 1765
rect 92857 1707 92865 1741
rect 92899 1707 92907 1741
rect 92857 1683 92907 1707
rect 93193 1741 93243 1765
rect 93193 1707 93201 1741
rect 93235 1707 93243 1741
rect 93193 1683 93243 1707
rect 93529 1741 93579 1765
rect 93529 1707 93537 1741
rect 93571 1707 93579 1741
rect 93529 1683 93579 1707
rect 93865 1741 93915 1765
rect 93865 1707 93873 1741
rect 93907 1707 93915 1741
rect 93865 1683 93915 1707
rect 94201 1741 94251 1765
rect 94201 1707 94209 1741
rect 94243 1707 94251 1741
rect 94201 1683 94251 1707
rect 94537 1741 94587 1765
rect 94537 1707 94545 1741
rect 94579 1707 94587 1741
rect 94537 1683 94587 1707
rect 94873 1741 94923 1765
rect 94873 1707 94881 1741
rect 94915 1707 94923 1741
rect 94873 1683 94923 1707
rect 95209 1741 95259 1765
rect 95209 1707 95217 1741
rect 95251 1707 95259 1741
rect 95209 1683 95259 1707
rect 95545 1741 95595 1765
rect 95545 1707 95553 1741
rect 95587 1707 95595 1741
rect 95545 1683 95595 1707
rect 95881 1741 95931 1765
rect 95881 1707 95889 1741
rect 95923 1707 95931 1741
rect 95881 1683 95931 1707
rect 96217 1741 96267 1765
rect 96217 1707 96225 1741
rect 96259 1707 96267 1741
rect 96217 1683 96267 1707
rect 96553 1741 96603 1765
rect 96553 1707 96561 1741
rect 96595 1707 96603 1741
rect 96553 1683 96603 1707
rect 96889 1741 96939 1765
rect 96889 1707 96897 1741
rect 96931 1707 96939 1741
rect 96889 1683 96939 1707
rect 97225 1741 97275 1765
rect 97225 1707 97233 1741
rect 97267 1707 97275 1741
rect 97225 1683 97275 1707
rect 97561 1741 97611 1765
rect 97561 1707 97569 1741
rect 97603 1707 97611 1741
rect 97561 1683 97611 1707
rect 97897 1741 97947 1765
rect 97897 1707 97905 1741
rect 97939 1707 97947 1741
rect 97897 1683 97947 1707
rect 98233 1741 98283 1765
rect 98233 1707 98241 1741
rect 98275 1707 98283 1741
rect 98233 1683 98283 1707
rect 98569 1741 98619 1765
rect 98569 1707 98577 1741
rect 98611 1707 98619 1741
rect 98569 1683 98619 1707
rect 98905 1741 98955 1765
rect 98905 1707 98913 1741
rect 98947 1707 98955 1741
rect 98905 1683 98955 1707
rect 99241 1741 99291 1765
rect 99241 1707 99249 1741
rect 99283 1707 99291 1741
rect 99241 1683 99291 1707
rect 99577 1741 99627 1765
rect 99577 1707 99585 1741
rect 99619 1707 99627 1741
rect 99577 1683 99627 1707
rect 99913 1741 99963 1765
rect 99913 1707 99921 1741
rect 99955 1707 99963 1741
rect 99913 1683 99963 1707
rect 100249 1741 100299 1765
rect 100249 1707 100257 1741
rect 100291 1707 100299 1741
rect 100249 1683 100299 1707
rect 100585 1741 100635 1765
rect 100585 1707 100593 1741
rect 100627 1707 100635 1741
rect 100585 1683 100635 1707
rect 100921 1741 100971 1765
rect 100921 1707 100929 1741
rect 100963 1707 100971 1741
rect 100921 1683 100971 1707
rect 101257 1741 101307 1765
rect 101257 1707 101265 1741
rect 101299 1707 101307 1741
rect 101257 1683 101307 1707
rect 101593 1741 101643 1765
rect 101593 1707 101601 1741
rect 101635 1707 101643 1741
rect 101593 1683 101643 1707
rect 101929 1741 101979 1765
rect 101929 1707 101937 1741
rect 101971 1707 101979 1741
rect 101929 1683 101979 1707
rect 102265 1741 102315 1765
rect 102265 1707 102273 1741
rect 102307 1707 102315 1741
rect 102265 1683 102315 1707
rect 102601 1741 102651 1765
rect 102601 1707 102609 1741
rect 102643 1707 102651 1741
rect 102601 1683 102651 1707
rect 102937 1741 102987 1765
rect 102937 1707 102945 1741
rect 102979 1707 102987 1741
rect 102937 1683 102987 1707
rect 103273 1741 103323 1765
rect 103273 1707 103281 1741
rect 103315 1707 103323 1741
rect 103273 1683 103323 1707
rect 103609 1741 103659 1765
rect 103609 1707 103617 1741
rect 103651 1707 103659 1741
rect 103609 1683 103659 1707
rect 103945 1741 103995 1765
rect 103945 1707 103953 1741
rect 103987 1707 103995 1741
rect 103945 1683 103995 1707
rect 104281 1741 104331 1765
rect 104281 1707 104289 1741
rect 104323 1707 104331 1741
rect 104281 1683 104331 1707
rect 104617 1741 104667 1765
rect 104617 1707 104625 1741
rect 104659 1707 104667 1741
rect 104617 1683 104667 1707
rect 104953 1741 105003 1765
rect 104953 1707 104961 1741
rect 104995 1707 105003 1741
rect 104953 1683 105003 1707
rect 105289 1741 105339 1765
rect 105289 1707 105297 1741
rect 105331 1707 105339 1741
rect 105289 1683 105339 1707
rect 105625 1741 105675 1765
rect 105625 1707 105633 1741
rect 105667 1707 105675 1741
rect 105625 1683 105675 1707
rect 105961 1741 106011 1765
rect 105961 1707 105969 1741
rect 106003 1707 106011 1741
rect 105961 1683 106011 1707
rect 106297 1741 106347 1765
rect 106297 1707 106305 1741
rect 106339 1707 106347 1741
rect 106297 1683 106347 1707
rect 106633 1741 106683 1765
rect 106633 1707 106641 1741
rect 106675 1707 106683 1741
rect 106633 1683 106683 1707
rect 106969 1741 107019 1765
rect 106969 1707 106977 1741
rect 107011 1707 107019 1741
rect 106969 1683 107019 1707
rect 107305 1741 107355 1765
rect 107305 1707 107313 1741
rect 107347 1707 107355 1741
rect 107305 1683 107355 1707
rect 107641 1741 107691 1765
rect 107641 1707 107649 1741
rect 107683 1707 107691 1741
rect 107641 1683 107691 1707
rect 107977 1741 108027 1765
rect 107977 1707 107985 1741
rect 108019 1707 108027 1741
rect 107977 1683 108027 1707
rect 108313 1741 108363 1765
rect 108313 1707 108321 1741
rect 108355 1707 108363 1741
rect 108313 1683 108363 1707
rect 108649 1741 108699 1765
rect 108649 1707 108657 1741
rect 108691 1707 108699 1741
rect 108649 1683 108699 1707
rect 108985 1741 109035 1765
rect 108985 1707 108993 1741
rect 109027 1707 109035 1741
rect 108985 1683 109035 1707
rect 109321 1741 109371 1765
rect 109321 1707 109329 1741
rect 109363 1707 109371 1741
rect 109321 1683 109371 1707
rect 109657 1741 109707 1765
rect 109657 1707 109665 1741
rect 109699 1707 109707 1741
rect 109657 1683 109707 1707
rect 109993 1741 110043 1765
rect 109993 1707 110001 1741
rect 110035 1707 110043 1741
rect 109993 1683 110043 1707
rect 110329 1741 110379 1765
rect 110329 1707 110337 1741
rect 110371 1707 110379 1741
rect 110329 1683 110379 1707
rect 110665 1741 110715 1765
rect 110665 1707 110673 1741
rect 110707 1707 110715 1741
rect 110665 1683 110715 1707
rect 111001 1741 111051 1765
rect 111001 1707 111009 1741
rect 111043 1707 111051 1741
rect 111001 1683 111051 1707
rect 111337 1741 111387 1765
rect 111337 1707 111345 1741
rect 111379 1707 111387 1741
rect 111337 1683 111387 1707
rect 111673 1741 111723 1765
rect 111673 1707 111681 1741
rect 111715 1707 111723 1741
rect 111673 1683 111723 1707
rect 112009 1741 112059 1765
rect 112009 1707 112017 1741
rect 112051 1707 112059 1741
rect 112009 1683 112059 1707
rect 112345 1741 112395 1765
rect 112345 1707 112353 1741
rect 112387 1707 112395 1741
rect 112345 1683 112395 1707
rect 112681 1741 112731 1765
rect 112681 1707 112689 1741
rect 112723 1707 112731 1741
rect 112681 1683 112731 1707
rect 113017 1741 113067 1765
rect 113017 1707 113025 1741
rect 113059 1707 113067 1741
rect 113017 1683 113067 1707
rect 113353 1741 113403 1765
rect 113353 1707 113361 1741
rect 113395 1707 113403 1741
rect 113353 1683 113403 1707
rect 113689 1741 113739 1765
rect 113689 1707 113697 1741
rect 113731 1707 113739 1741
rect 113689 1683 113739 1707
rect 114025 1741 114075 1765
rect 114025 1707 114033 1741
rect 114067 1707 114075 1741
rect 114025 1683 114075 1707
rect 114361 1741 114411 1765
rect 114361 1707 114369 1741
rect 114403 1707 114411 1741
rect 114361 1683 114411 1707
rect 114697 1741 114747 1765
rect 114697 1707 114705 1741
rect 114739 1707 114747 1741
rect 114697 1683 114747 1707
rect 115033 1741 115083 1765
rect 115033 1707 115041 1741
rect 115075 1707 115083 1741
rect 115033 1683 115083 1707
rect 115369 1741 115419 1765
rect 115369 1707 115377 1741
rect 115411 1707 115419 1741
rect 115369 1683 115419 1707
rect 115705 1741 115755 1765
rect 115705 1707 115713 1741
rect 115747 1707 115755 1741
rect 115705 1683 115755 1707
rect 116041 1741 116091 1765
rect 116041 1707 116049 1741
rect 116083 1707 116091 1741
rect 116041 1683 116091 1707
rect 116377 1741 116427 1765
rect 116377 1707 116385 1741
rect 116419 1707 116427 1741
rect 116377 1683 116427 1707
rect 116713 1741 116763 1765
rect 116713 1707 116721 1741
rect 116755 1707 116763 1741
rect 116713 1683 116763 1707
rect 117049 1741 117099 1765
rect 117049 1707 117057 1741
rect 117091 1707 117099 1741
rect 117049 1683 117099 1707
rect 117385 1741 117435 1765
rect 117385 1707 117393 1741
rect 117427 1707 117435 1741
rect 117385 1683 117435 1707
rect 117721 1741 117771 1765
rect 117721 1707 117729 1741
rect 117763 1707 117771 1741
rect 117721 1683 117771 1707
rect 118057 1741 118107 1765
rect 118057 1707 118065 1741
rect 118099 1707 118107 1741
rect 118057 1683 118107 1707
rect 118393 1741 118443 1765
rect 118393 1707 118401 1741
rect 118435 1707 118443 1741
rect 118393 1683 118443 1707
rect 118729 1741 118779 1765
rect 118729 1707 118737 1741
rect 118771 1707 118779 1741
rect 118729 1683 118779 1707
rect 119065 1741 119115 1765
rect 119065 1707 119073 1741
rect 119107 1707 119115 1741
rect 119065 1683 119115 1707
rect 119401 1741 119451 1765
rect 119401 1707 119409 1741
rect 119443 1707 119451 1741
rect 119401 1683 119451 1707
rect 119737 1741 119787 1765
rect 119737 1707 119745 1741
rect 119779 1707 119787 1741
rect 119737 1683 119787 1707
rect 120073 1741 120123 1765
rect 120073 1707 120081 1741
rect 120115 1707 120123 1741
rect 120073 1683 120123 1707
rect 120409 1741 120459 1765
rect 120409 1707 120417 1741
rect 120451 1707 120459 1741
rect 120409 1683 120459 1707
rect 120745 1741 120795 1765
rect 120745 1707 120753 1741
rect 120787 1707 120795 1741
rect 120745 1683 120795 1707
rect 121081 1741 121131 1765
rect 121081 1707 121089 1741
rect 121123 1707 121131 1741
rect 121081 1683 121131 1707
rect 121417 1741 121467 1765
rect 121417 1707 121425 1741
rect 121459 1707 121467 1741
rect 121417 1683 121467 1707
rect 121753 1741 121803 1765
rect 121753 1707 121761 1741
rect 121795 1707 121803 1741
rect 121753 1683 121803 1707
rect 122089 1741 122139 1765
rect 122089 1707 122097 1741
rect 122131 1707 122139 1741
rect 122089 1683 122139 1707
rect 122425 1741 122475 1765
rect 122425 1707 122433 1741
rect 122467 1707 122475 1741
rect 122425 1683 122475 1707
rect 122761 1741 122811 1765
rect 122761 1707 122769 1741
rect 122803 1707 122811 1741
rect 122761 1683 122811 1707
rect 123097 1741 123147 1765
rect 123097 1707 123105 1741
rect 123139 1707 123147 1741
rect 123097 1683 123147 1707
rect 123433 1741 123483 1765
rect 123433 1707 123441 1741
rect 123475 1707 123483 1741
rect 123433 1683 123483 1707
rect 123769 1741 123819 1765
rect 123769 1707 123777 1741
rect 123811 1707 123819 1741
rect 123769 1683 123819 1707
rect 124105 1741 124155 1765
rect 124105 1707 124113 1741
rect 124147 1707 124155 1741
rect 124105 1683 124155 1707
rect 124441 1741 124491 1765
rect 124441 1707 124449 1741
rect 124483 1707 124491 1741
rect 124441 1683 124491 1707
rect 124777 1741 124827 1765
rect 124777 1707 124785 1741
rect 124819 1707 124827 1741
rect 124777 1683 124827 1707
rect 125113 1741 125163 1765
rect 125113 1707 125121 1741
rect 125155 1707 125163 1741
rect 125113 1683 125163 1707
rect 125449 1741 125499 1765
rect 125449 1707 125457 1741
rect 125491 1707 125499 1741
rect 125449 1683 125499 1707
rect 125785 1741 125835 1765
rect 125785 1707 125793 1741
rect 125827 1707 125835 1741
rect 125785 1683 125835 1707
rect 126121 1741 126171 1765
rect 126121 1707 126129 1741
rect 126163 1707 126171 1741
rect 126121 1683 126171 1707
rect 126457 1741 126507 1765
rect 126457 1707 126465 1741
rect 126499 1707 126507 1741
rect 126457 1683 126507 1707
rect 126793 1741 126843 1765
rect 126793 1707 126801 1741
rect 126835 1707 126843 1741
rect 126793 1683 126843 1707
rect 127129 1741 127179 1765
rect 127129 1707 127137 1741
rect 127171 1707 127179 1741
rect 127129 1683 127179 1707
rect 127465 1741 127515 1765
rect 127465 1707 127473 1741
rect 127507 1707 127515 1741
rect 127465 1683 127515 1707
rect 127801 1741 127851 1765
rect 127801 1707 127809 1741
rect 127843 1707 127851 1741
rect 127801 1683 127851 1707
rect 128137 1741 128187 1765
rect 128137 1707 128145 1741
rect 128179 1707 128187 1741
rect 128137 1683 128187 1707
rect 128473 1741 128523 1765
rect 128473 1707 128481 1741
rect 128515 1707 128523 1741
rect 128473 1683 128523 1707
rect 128809 1741 128859 1765
rect 128809 1707 128817 1741
rect 128851 1707 128859 1741
rect 128809 1683 128859 1707
rect 129145 1741 129195 1765
rect 129145 1707 129153 1741
rect 129187 1707 129195 1741
rect 129145 1683 129195 1707
rect 129481 1741 129531 1765
rect 129481 1707 129489 1741
rect 129523 1707 129531 1741
rect 129481 1683 129531 1707
rect 129817 1741 129867 1765
rect 129817 1707 129825 1741
rect 129859 1707 129867 1741
rect 129817 1683 129867 1707
rect 130153 1741 130203 1765
rect 130153 1707 130161 1741
rect 130195 1707 130203 1741
rect 130153 1683 130203 1707
rect 130489 1741 130539 1765
rect 130489 1707 130497 1741
rect 130531 1707 130539 1741
rect 130489 1683 130539 1707
rect 130825 1741 130875 1765
rect 130825 1707 130833 1741
rect 130867 1707 130875 1741
rect 130825 1683 130875 1707
rect 131161 1741 131211 1765
rect 131161 1707 131169 1741
rect 131203 1707 131211 1741
rect 131161 1683 131211 1707
rect 131497 1741 131547 1765
rect 131497 1707 131505 1741
rect 131539 1707 131547 1741
rect 131497 1683 131547 1707
rect 131833 1741 131883 1765
rect 131833 1707 131841 1741
rect 131875 1707 131883 1741
rect 131833 1683 131883 1707
rect 132169 1741 132219 1765
rect 132169 1707 132177 1741
rect 132211 1707 132219 1741
rect 132169 1683 132219 1707
rect 132505 1741 132555 1765
rect 132505 1707 132513 1741
rect 132547 1707 132555 1741
rect 132505 1683 132555 1707
rect 132841 1741 132891 1765
rect 132841 1707 132849 1741
rect 132883 1707 132891 1741
rect 132841 1683 132891 1707
rect 133177 1741 133227 1765
rect 133177 1707 133185 1741
rect 133219 1707 133227 1741
rect 133177 1683 133227 1707
rect 133513 1741 133563 1765
rect 133513 1707 133521 1741
rect 133555 1707 133563 1741
rect 133513 1683 133563 1707
rect 133849 1741 133899 1765
rect 133849 1707 133857 1741
rect 133891 1707 133899 1741
rect 133849 1683 133899 1707
rect 134185 1741 134235 1765
rect 134185 1707 134193 1741
rect 134227 1707 134235 1741
rect 134185 1683 134235 1707
rect 134521 1741 134571 1765
rect 134521 1707 134529 1741
rect 134563 1707 134571 1741
rect 134521 1683 134571 1707
rect 134857 1741 134907 1765
rect 134857 1707 134865 1741
rect 134899 1707 134907 1741
rect 134857 1683 134907 1707
rect 135193 1741 135243 1765
rect 135193 1707 135201 1741
rect 135235 1707 135243 1741
rect 135193 1683 135243 1707
rect 135529 1741 135579 1765
rect 135529 1707 135537 1741
rect 135571 1707 135579 1741
rect 135529 1683 135579 1707
rect 135865 1741 135915 1765
rect 135865 1707 135873 1741
rect 135907 1707 135915 1741
rect 135865 1683 135915 1707
rect 136201 1741 136251 1765
rect 136201 1707 136209 1741
rect 136243 1707 136251 1741
rect 136201 1683 136251 1707
rect 136537 1741 136587 1765
rect 136537 1707 136545 1741
rect 136579 1707 136587 1741
rect 136537 1683 136587 1707
<< nsubdiffcont >>
rect 2145 132016 2179 132050
rect 2481 132016 2515 132050
rect 2817 132016 2851 132050
rect 3153 132016 3187 132050
rect 3489 132016 3523 132050
rect 3825 132016 3859 132050
rect 4161 132016 4195 132050
rect 4497 132016 4531 132050
rect 4833 132016 4867 132050
rect 5169 132016 5203 132050
rect 5505 132016 5539 132050
rect 5841 132016 5875 132050
rect 6177 132016 6211 132050
rect 6513 132016 6547 132050
rect 6849 132016 6883 132050
rect 7185 132016 7219 132050
rect 7521 132016 7555 132050
rect 7857 132016 7891 132050
rect 8193 132016 8227 132050
rect 8529 132016 8563 132050
rect 8865 132016 8899 132050
rect 9201 132016 9235 132050
rect 9537 132016 9571 132050
rect 9873 132016 9907 132050
rect 10209 132016 10243 132050
rect 10545 132016 10579 132050
rect 10881 132016 10915 132050
rect 11217 132016 11251 132050
rect 11553 132016 11587 132050
rect 11889 132016 11923 132050
rect 12225 132016 12259 132050
rect 12561 132016 12595 132050
rect 12897 132016 12931 132050
rect 13233 132016 13267 132050
rect 13569 132016 13603 132050
rect 13905 132016 13939 132050
rect 14241 132016 14275 132050
rect 14577 132016 14611 132050
rect 14913 132016 14947 132050
rect 15249 132016 15283 132050
rect 15585 132016 15619 132050
rect 15921 132016 15955 132050
rect 16257 132016 16291 132050
rect 16593 132016 16627 132050
rect 16929 132016 16963 132050
rect 17265 132016 17299 132050
rect 17601 132016 17635 132050
rect 17937 132016 17971 132050
rect 18273 132016 18307 132050
rect 18609 132016 18643 132050
rect 18945 132016 18979 132050
rect 19281 132016 19315 132050
rect 19617 132016 19651 132050
rect 19953 132016 19987 132050
rect 20289 132016 20323 132050
rect 20625 132016 20659 132050
rect 20961 132016 20995 132050
rect 21297 132016 21331 132050
rect 21633 132016 21667 132050
rect 21969 132016 22003 132050
rect 22305 132016 22339 132050
rect 22641 132016 22675 132050
rect 22977 132016 23011 132050
rect 23313 132016 23347 132050
rect 23649 132016 23683 132050
rect 23985 132016 24019 132050
rect 24321 132016 24355 132050
rect 24657 132016 24691 132050
rect 24993 132016 25027 132050
rect 25329 132016 25363 132050
rect 25665 132016 25699 132050
rect 26001 132016 26035 132050
rect 26337 132016 26371 132050
rect 26673 132016 26707 132050
rect 27009 132016 27043 132050
rect 27345 132016 27379 132050
rect 27681 132016 27715 132050
rect 28017 132016 28051 132050
rect 28353 132016 28387 132050
rect 28689 132016 28723 132050
rect 29025 132016 29059 132050
rect 29361 132016 29395 132050
rect 29697 132016 29731 132050
rect 30033 132016 30067 132050
rect 30369 132016 30403 132050
rect 30705 132016 30739 132050
rect 31041 132016 31075 132050
rect 31377 132016 31411 132050
rect 31713 132016 31747 132050
rect 32049 132016 32083 132050
rect 32385 132016 32419 132050
rect 32721 132016 32755 132050
rect 33057 132016 33091 132050
rect 33393 132016 33427 132050
rect 33729 132016 33763 132050
rect 34065 132016 34099 132050
rect 34401 132016 34435 132050
rect 34737 132016 34771 132050
rect 35073 132016 35107 132050
rect 35409 132016 35443 132050
rect 35745 132016 35779 132050
rect 36081 132016 36115 132050
rect 36417 132016 36451 132050
rect 36753 132016 36787 132050
rect 37089 132016 37123 132050
rect 37425 132016 37459 132050
rect 37761 132016 37795 132050
rect 38097 132016 38131 132050
rect 38433 132016 38467 132050
rect 38769 132016 38803 132050
rect 39105 132016 39139 132050
rect 39441 132016 39475 132050
rect 39777 132016 39811 132050
rect 40113 132016 40147 132050
rect 40449 132016 40483 132050
rect 40785 132016 40819 132050
rect 41121 132016 41155 132050
rect 41457 132016 41491 132050
rect 41793 132016 41827 132050
rect 42129 132016 42163 132050
rect 42465 132016 42499 132050
rect 42801 132016 42835 132050
rect 43137 132016 43171 132050
rect 43473 132016 43507 132050
rect 43809 132016 43843 132050
rect 44145 132016 44179 132050
rect 44481 132016 44515 132050
rect 44817 132016 44851 132050
rect 45153 132016 45187 132050
rect 45489 132016 45523 132050
rect 45825 132016 45859 132050
rect 46161 132016 46195 132050
rect 46497 132016 46531 132050
rect 46833 132016 46867 132050
rect 47169 132016 47203 132050
rect 47505 132016 47539 132050
rect 47841 132016 47875 132050
rect 48177 132016 48211 132050
rect 48513 132016 48547 132050
rect 48849 132016 48883 132050
rect 49185 132016 49219 132050
rect 49521 132016 49555 132050
rect 49857 132016 49891 132050
rect 50193 132016 50227 132050
rect 50529 132016 50563 132050
rect 50865 132016 50899 132050
rect 51201 132016 51235 132050
rect 51537 132016 51571 132050
rect 51873 132016 51907 132050
rect 52209 132016 52243 132050
rect 52545 132016 52579 132050
rect 52881 132016 52915 132050
rect 53217 132016 53251 132050
rect 53553 132016 53587 132050
rect 53889 132016 53923 132050
rect 54225 132016 54259 132050
rect 54561 132016 54595 132050
rect 54897 132016 54931 132050
rect 55233 132016 55267 132050
rect 55569 132016 55603 132050
rect 55905 132016 55939 132050
rect 56241 132016 56275 132050
rect 56577 132016 56611 132050
rect 56913 132016 56947 132050
rect 57249 132016 57283 132050
rect 57585 132016 57619 132050
rect 57921 132016 57955 132050
rect 58257 132016 58291 132050
rect 58593 132016 58627 132050
rect 58929 132016 58963 132050
rect 59265 132016 59299 132050
rect 59601 132016 59635 132050
rect 59937 132016 59971 132050
rect 60273 132016 60307 132050
rect 60609 132016 60643 132050
rect 60945 132016 60979 132050
rect 61281 132016 61315 132050
rect 61617 132016 61651 132050
rect 61953 132016 61987 132050
rect 62289 132016 62323 132050
rect 62625 132016 62659 132050
rect 62961 132016 62995 132050
rect 63297 132016 63331 132050
rect 63633 132016 63667 132050
rect 63969 132016 64003 132050
rect 64305 132016 64339 132050
rect 64641 132016 64675 132050
rect 64977 132016 65011 132050
rect 65313 132016 65347 132050
rect 65649 132016 65683 132050
rect 65985 132016 66019 132050
rect 66321 132016 66355 132050
rect 66657 132016 66691 132050
rect 66993 132016 67027 132050
rect 67329 132016 67363 132050
rect 67665 132016 67699 132050
rect 68001 132016 68035 132050
rect 68337 132016 68371 132050
rect 68673 132016 68707 132050
rect 69009 132016 69043 132050
rect 69345 132016 69379 132050
rect 69681 132016 69715 132050
rect 70017 132016 70051 132050
rect 70353 132016 70387 132050
rect 70689 132016 70723 132050
rect 71025 132016 71059 132050
rect 71361 132016 71395 132050
rect 71697 132016 71731 132050
rect 72033 132016 72067 132050
rect 72369 132016 72403 132050
rect 72705 132016 72739 132050
rect 73041 132016 73075 132050
rect 73377 132016 73411 132050
rect 73713 132016 73747 132050
rect 74049 132016 74083 132050
rect 74385 132016 74419 132050
rect 74721 132016 74755 132050
rect 75057 132016 75091 132050
rect 75393 132016 75427 132050
rect 75729 132016 75763 132050
rect 76065 132016 76099 132050
rect 76401 132016 76435 132050
rect 76737 132016 76771 132050
rect 77073 132016 77107 132050
rect 77409 132016 77443 132050
rect 77745 132016 77779 132050
rect 78081 132016 78115 132050
rect 78417 132016 78451 132050
rect 78753 132016 78787 132050
rect 79089 132016 79123 132050
rect 79425 132016 79459 132050
rect 79761 132016 79795 132050
rect 80097 132016 80131 132050
rect 80433 132016 80467 132050
rect 80769 132016 80803 132050
rect 81105 132016 81139 132050
rect 81441 132016 81475 132050
rect 81777 132016 81811 132050
rect 82113 132016 82147 132050
rect 82449 132016 82483 132050
rect 82785 132016 82819 132050
rect 83121 132016 83155 132050
rect 83457 132016 83491 132050
rect 83793 132016 83827 132050
rect 84129 132016 84163 132050
rect 84465 132016 84499 132050
rect 84801 132016 84835 132050
rect 85137 132016 85171 132050
rect 85473 132016 85507 132050
rect 85809 132016 85843 132050
rect 86145 132016 86179 132050
rect 86481 132016 86515 132050
rect 86817 132016 86851 132050
rect 87153 132016 87187 132050
rect 87489 132016 87523 132050
rect 87825 132016 87859 132050
rect 88161 132016 88195 132050
rect 88497 132016 88531 132050
rect 88833 132016 88867 132050
rect 89169 132016 89203 132050
rect 89505 132016 89539 132050
rect 89841 132016 89875 132050
rect 90177 132016 90211 132050
rect 90513 132016 90547 132050
rect 90849 132016 90883 132050
rect 91185 132016 91219 132050
rect 91521 132016 91555 132050
rect 91857 132016 91891 132050
rect 92193 132016 92227 132050
rect 92529 132016 92563 132050
rect 92865 132016 92899 132050
rect 93201 132016 93235 132050
rect 93537 132016 93571 132050
rect 93873 132016 93907 132050
rect 94209 132016 94243 132050
rect 94545 132016 94579 132050
rect 94881 132016 94915 132050
rect 95217 132016 95251 132050
rect 95553 132016 95587 132050
rect 95889 132016 95923 132050
rect 96225 132016 96259 132050
rect 96561 132016 96595 132050
rect 96897 132016 96931 132050
rect 97233 132016 97267 132050
rect 97569 132016 97603 132050
rect 97905 132016 97939 132050
rect 98241 132016 98275 132050
rect 98577 132016 98611 132050
rect 98913 132016 98947 132050
rect 99249 132016 99283 132050
rect 99585 132016 99619 132050
rect 99921 132016 99955 132050
rect 100257 132016 100291 132050
rect 100593 132016 100627 132050
rect 100929 132016 100963 132050
rect 101265 132016 101299 132050
rect 101601 132016 101635 132050
rect 101937 132016 101971 132050
rect 102273 132016 102307 132050
rect 102609 132016 102643 132050
rect 102945 132016 102979 132050
rect 103281 132016 103315 132050
rect 103617 132016 103651 132050
rect 103953 132016 103987 132050
rect 104289 132016 104323 132050
rect 104625 132016 104659 132050
rect 104961 132016 104995 132050
rect 105297 132016 105331 132050
rect 105633 132016 105667 132050
rect 105969 132016 106003 132050
rect 106305 132016 106339 132050
rect 106641 132016 106675 132050
rect 106977 132016 107011 132050
rect 107313 132016 107347 132050
rect 107649 132016 107683 132050
rect 107985 132016 108019 132050
rect 108321 132016 108355 132050
rect 108657 132016 108691 132050
rect 108993 132016 109027 132050
rect 109329 132016 109363 132050
rect 109665 132016 109699 132050
rect 110001 132016 110035 132050
rect 110337 132016 110371 132050
rect 110673 132016 110707 132050
rect 111009 132016 111043 132050
rect 111345 132016 111379 132050
rect 111681 132016 111715 132050
rect 112017 132016 112051 132050
rect 112353 132016 112387 132050
rect 112689 132016 112723 132050
rect 113025 132016 113059 132050
rect 113361 132016 113395 132050
rect 113697 132016 113731 132050
rect 114033 132016 114067 132050
rect 114369 132016 114403 132050
rect 114705 132016 114739 132050
rect 115041 132016 115075 132050
rect 115377 132016 115411 132050
rect 115713 132016 115747 132050
rect 116049 132016 116083 132050
rect 116385 132016 116419 132050
rect 116721 132016 116755 132050
rect 117057 132016 117091 132050
rect 117393 132016 117427 132050
rect 117729 132016 117763 132050
rect 118065 132016 118099 132050
rect 118401 132016 118435 132050
rect 118737 132016 118771 132050
rect 119073 132016 119107 132050
rect 119409 132016 119443 132050
rect 119745 132016 119779 132050
rect 120081 132016 120115 132050
rect 120417 132016 120451 132050
rect 120753 132016 120787 132050
rect 121089 132016 121123 132050
rect 121425 132016 121459 132050
rect 121761 132016 121795 132050
rect 122097 132016 122131 132050
rect 122433 132016 122467 132050
rect 122769 132016 122803 132050
rect 123105 132016 123139 132050
rect 123441 132016 123475 132050
rect 123777 132016 123811 132050
rect 124113 132016 124147 132050
rect 124449 132016 124483 132050
rect 124785 132016 124819 132050
rect 125121 132016 125155 132050
rect 125457 132016 125491 132050
rect 125793 132016 125827 132050
rect 126129 132016 126163 132050
rect 126465 132016 126499 132050
rect 126801 132016 126835 132050
rect 127137 132016 127171 132050
rect 127473 132016 127507 132050
rect 127809 132016 127843 132050
rect 128145 132016 128179 132050
rect 128481 132016 128515 132050
rect 128817 132016 128851 132050
rect 129153 132016 129187 132050
rect 129489 132016 129523 132050
rect 129825 132016 129859 132050
rect 130161 132016 130195 132050
rect 130497 132016 130531 132050
rect 130833 132016 130867 132050
rect 131169 132016 131203 132050
rect 131505 132016 131539 132050
rect 131841 132016 131875 132050
rect 132177 132016 132211 132050
rect 132513 132016 132547 132050
rect 132849 132016 132883 132050
rect 133185 132016 133219 132050
rect 133521 132016 133555 132050
rect 133857 132016 133891 132050
rect 134193 132016 134227 132050
rect 134529 132016 134563 132050
rect 134865 132016 134899 132050
rect 135201 132016 135235 132050
rect 135537 132016 135571 132050
rect 135873 132016 135907 132050
rect 136209 132016 136243 132050
rect 136545 132016 136579 132050
rect 1809 131403 1843 131437
rect 136955 131403 136989 131437
rect 1809 131067 1843 131101
rect 136955 131067 136989 131101
rect 1809 130731 1843 130765
rect 136955 130731 136989 130765
rect 1809 130395 1843 130429
rect 136955 130395 136989 130429
rect 1809 130059 1843 130093
rect 136955 130059 136989 130093
rect 1809 129723 1843 129757
rect 136955 129723 136989 129757
rect 1809 129387 1843 129421
rect 136955 129387 136989 129421
rect 1809 129051 1843 129085
rect 136955 129051 136989 129085
rect 1809 128715 1843 128749
rect 136955 128715 136989 128749
rect 1809 128379 1843 128413
rect 136955 128379 136989 128413
rect 1809 128043 1843 128077
rect 136955 128043 136989 128077
rect 1809 127707 1843 127741
rect 136955 127707 136989 127741
rect 1809 127371 1843 127405
rect 136955 127371 136989 127405
rect 1809 127035 1843 127069
rect 136955 127035 136989 127069
rect 1809 126699 1843 126733
rect 136955 126699 136989 126733
rect 1809 126363 1843 126397
rect 136955 126363 136989 126397
rect 1809 126027 1843 126061
rect 136955 126027 136989 126061
rect 1809 125691 1843 125725
rect 136955 125691 136989 125725
rect 1809 125355 1843 125389
rect 136955 125355 136989 125389
rect 1809 125019 1843 125053
rect 136955 125019 136989 125053
rect 1809 124683 1843 124717
rect 136955 124683 136989 124717
rect 1809 124347 1843 124381
rect 136955 124347 136989 124381
rect 1809 124011 1843 124045
rect 136955 124011 136989 124045
rect 1809 123675 1843 123709
rect 136955 123675 136989 123709
rect 1809 123339 1843 123373
rect 136955 123339 136989 123373
rect 1809 123003 1843 123037
rect 136955 123003 136989 123037
rect 1809 122667 1843 122701
rect 136955 122667 136989 122701
rect 1809 122331 1843 122365
rect 136955 122331 136989 122365
rect 1809 121995 1843 122029
rect 136955 121995 136989 122029
rect 1809 121659 1843 121693
rect 136955 121659 136989 121693
rect 1809 121323 1843 121357
rect 136955 121323 136989 121357
rect 1809 120987 1843 121021
rect 136955 120987 136989 121021
rect 1809 120651 1843 120685
rect 136955 120651 136989 120685
rect 1809 120315 1843 120349
rect 136955 120315 136989 120349
rect 1809 119979 1843 120013
rect 136955 119979 136989 120013
rect 1809 119643 1843 119677
rect 136955 119643 136989 119677
rect 1809 119307 1843 119341
rect 136955 119307 136989 119341
rect 1809 118971 1843 119005
rect 136955 118971 136989 119005
rect 1809 118635 1843 118669
rect 136955 118635 136989 118669
rect 1809 118299 1843 118333
rect 136955 118299 136989 118333
rect 1809 117963 1843 117997
rect 136955 117963 136989 117997
rect 1809 117627 1843 117661
rect 136955 117627 136989 117661
rect 1809 117291 1843 117325
rect 136955 117291 136989 117325
rect 1809 116955 1843 116989
rect 136955 116955 136989 116989
rect 1809 116619 1843 116653
rect 136955 116619 136989 116653
rect 1809 116283 1843 116317
rect 136955 116283 136989 116317
rect 1809 115947 1843 115981
rect 136955 115947 136989 115981
rect 1809 115611 1843 115645
rect 136955 115611 136989 115645
rect 1809 115275 1843 115309
rect 136955 115275 136989 115309
rect 1809 114939 1843 114973
rect 136955 114939 136989 114973
rect 1809 114603 1843 114637
rect 136955 114603 136989 114637
rect 1809 114267 1843 114301
rect 136955 114267 136989 114301
rect 1809 113931 1843 113965
rect 136955 113931 136989 113965
rect 1809 113595 1843 113629
rect 136955 113595 136989 113629
rect 1809 113259 1843 113293
rect 136955 113259 136989 113293
rect 1809 112923 1843 112957
rect 136955 112923 136989 112957
rect 1809 112587 1843 112621
rect 136955 112587 136989 112621
rect 1809 112251 1843 112285
rect 136955 112251 136989 112285
rect 1809 111915 1843 111949
rect 136955 111915 136989 111949
rect 1809 111579 1843 111613
rect 136955 111579 136989 111613
rect 1809 111243 1843 111277
rect 136955 111243 136989 111277
rect 1809 110907 1843 110941
rect 136955 110907 136989 110941
rect 1809 110571 1843 110605
rect 136955 110571 136989 110605
rect 1809 110235 1843 110269
rect 136955 110235 136989 110269
rect 1809 109899 1843 109933
rect 136955 109899 136989 109933
rect 1809 109563 1843 109597
rect 136955 109563 136989 109597
rect 1809 109227 1843 109261
rect 136955 109227 136989 109261
rect 1809 108891 1843 108925
rect 136955 108891 136989 108925
rect 1809 108555 1843 108589
rect 136955 108555 136989 108589
rect 1809 108219 1843 108253
rect 136955 108219 136989 108253
rect 1809 107883 1843 107917
rect 136955 107883 136989 107917
rect 1809 107547 1843 107581
rect 136955 107547 136989 107581
rect 1809 107211 1843 107245
rect 136955 107211 136989 107245
rect 1809 106875 1843 106909
rect 136955 106875 136989 106909
rect 1809 106539 1843 106573
rect 136955 106539 136989 106573
rect 1809 106203 1843 106237
rect 136955 106203 136989 106237
rect 1809 105867 1843 105901
rect 136955 105867 136989 105901
rect 1809 105531 1843 105565
rect 136955 105531 136989 105565
rect 1809 105195 1843 105229
rect 136955 105195 136989 105229
rect 1809 104859 1843 104893
rect 136955 104859 136989 104893
rect 1809 104523 1843 104557
rect 136955 104523 136989 104557
rect 1809 104187 1843 104221
rect 136955 104187 136989 104221
rect 1809 103851 1843 103885
rect 136955 103851 136989 103885
rect 1809 103515 1843 103549
rect 136955 103515 136989 103549
rect 1809 103179 1843 103213
rect 136955 103179 136989 103213
rect 1809 102843 1843 102877
rect 136955 102843 136989 102877
rect 1809 102507 1843 102541
rect 136955 102507 136989 102541
rect 1809 102171 1843 102205
rect 136955 102171 136989 102205
rect 1809 101835 1843 101869
rect 136955 101835 136989 101869
rect 1809 101499 1843 101533
rect 136955 101499 136989 101533
rect 1809 101163 1843 101197
rect 136955 101163 136989 101197
rect 1809 100827 1843 100861
rect 136955 100827 136989 100861
rect 1809 100491 1843 100525
rect 136955 100491 136989 100525
rect 1809 100155 1843 100189
rect 136955 100155 136989 100189
rect 1809 99819 1843 99853
rect 136955 99819 136989 99853
rect 1809 99483 1843 99517
rect 136955 99483 136989 99517
rect 1809 99147 1843 99181
rect 136955 99147 136989 99181
rect 1809 98811 1843 98845
rect 136955 98811 136989 98845
rect 1809 98475 1843 98509
rect 136955 98475 136989 98509
rect 1809 98139 1843 98173
rect 136955 98139 136989 98173
rect 1809 97803 1843 97837
rect 136955 97803 136989 97837
rect 1809 97467 1843 97501
rect 136955 97467 136989 97501
rect 1809 97131 1843 97165
rect 136955 97131 136989 97165
rect 1809 96795 1843 96829
rect 136955 96795 136989 96829
rect 1809 96459 1843 96493
rect 136955 96459 136989 96493
rect 1809 96123 1843 96157
rect 136955 96123 136989 96157
rect 1809 95787 1843 95821
rect 136955 95787 136989 95821
rect 1809 95451 1843 95485
rect 136955 95451 136989 95485
rect 1809 95115 1843 95149
rect 136955 95115 136989 95149
rect 1809 94779 1843 94813
rect 136955 94779 136989 94813
rect 1809 94443 1843 94477
rect 136955 94443 136989 94477
rect 1809 94107 1843 94141
rect 136955 94107 136989 94141
rect 1809 93771 1843 93805
rect 136955 93771 136989 93805
rect 1809 93435 1843 93469
rect 136955 93435 136989 93469
rect 1809 93099 1843 93133
rect 136955 93099 136989 93133
rect 1809 92763 1843 92797
rect 136955 92763 136989 92797
rect 1809 92427 1843 92461
rect 136955 92427 136989 92461
rect 1809 92091 1843 92125
rect 136955 92091 136989 92125
rect 1809 91755 1843 91789
rect 136955 91755 136989 91789
rect 1809 91419 1843 91453
rect 136955 91419 136989 91453
rect 1809 91083 1843 91117
rect 136955 91083 136989 91117
rect 1809 90747 1843 90781
rect 136955 90747 136989 90781
rect 1809 90411 1843 90445
rect 136955 90411 136989 90445
rect 1809 90075 1843 90109
rect 136955 90075 136989 90109
rect 1809 89739 1843 89773
rect 136955 89739 136989 89773
rect 1809 89403 1843 89437
rect 136955 89403 136989 89437
rect 1809 89067 1843 89101
rect 136955 89067 136989 89101
rect 1809 88731 1843 88765
rect 136955 88731 136989 88765
rect 1809 88395 1843 88429
rect 136955 88395 136989 88429
rect 1809 88059 1843 88093
rect 136955 88059 136989 88093
rect 1809 87723 1843 87757
rect 136955 87723 136989 87757
rect 1809 87387 1843 87421
rect 136955 87387 136989 87421
rect 1809 87051 1843 87085
rect 136955 87051 136989 87085
rect 1809 86715 1843 86749
rect 136955 86715 136989 86749
rect 1809 86379 1843 86413
rect 136955 86379 136989 86413
rect 1809 86043 1843 86077
rect 136955 86043 136989 86077
rect 1809 85707 1843 85741
rect 136955 85707 136989 85741
rect 1809 85371 1843 85405
rect 136955 85371 136989 85405
rect 1809 85035 1843 85069
rect 136955 85035 136989 85069
rect 1809 84699 1843 84733
rect 136955 84699 136989 84733
rect 1809 84363 1843 84397
rect 136955 84363 136989 84397
rect 1809 84027 1843 84061
rect 136955 84027 136989 84061
rect 1809 83691 1843 83725
rect 136955 83691 136989 83725
rect 1809 83355 1843 83389
rect 136955 83355 136989 83389
rect 1809 83019 1843 83053
rect 136955 83019 136989 83053
rect 1809 82683 1843 82717
rect 136955 82683 136989 82717
rect 1809 82347 1843 82381
rect 136955 82347 136989 82381
rect 1809 82011 1843 82045
rect 136955 82011 136989 82045
rect 1809 81675 1843 81709
rect 136955 81675 136989 81709
rect 1809 81339 1843 81373
rect 136955 81339 136989 81373
rect 1809 81003 1843 81037
rect 136955 81003 136989 81037
rect 1809 80667 1843 80701
rect 136955 80667 136989 80701
rect 1809 80331 1843 80365
rect 136955 80331 136989 80365
rect 1809 79995 1843 80029
rect 136955 79995 136989 80029
rect 1809 79659 1843 79693
rect 136955 79659 136989 79693
rect 1809 79323 1843 79357
rect 136955 79323 136989 79357
rect 1809 78987 1843 79021
rect 136955 78987 136989 79021
rect 1809 78651 1843 78685
rect 136955 78651 136989 78685
rect 1809 78315 1843 78349
rect 136955 78315 136989 78349
rect 1809 77979 1843 78013
rect 136955 77979 136989 78013
rect 1809 77643 1843 77677
rect 136955 77643 136989 77677
rect 1809 77307 1843 77341
rect 136955 77307 136989 77341
rect 1809 76971 1843 77005
rect 136955 76971 136989 77005
rect 1809 76635 1843 76669
rect 136955 76635 136989 76669
rect 1809 76299 1843 76333
rect 136955 76299 136989 76333
rect 1809 75963 1843 75997
rect 136955 75963 136989 75997
rect 1809 75627 1843 75661
rect 136955 75627 136989 75661
rect 1809 75291 1843 75325
rect 136955 75291 136989 75325
rect 1809 74955 1843 74989
rect 136955 74955 136989 74989
rect 1809 74619 1843 74653
rect 136955 74619 136989 74653
rect 1809 74283 1843 74317
rect 136955 74283 136989 74317
rect 1809 73947 1843 73981
rect 136955 73947 136989 73981
rect 1809 73611 1843 73645
rect 136955 73611 136989 73645
rect 1809 73275 1843 73309
rect 136955 73275 136989 73309
rect 1809 72939 1843 72973
rect 136955 72939 136989 72973
rect 1809 72603 1843 72637
rect 136955 72603 136989 72637
rect 1809 72267 1843 72301
rect 136955 72267 136989 72301
rect 1809 71931 1843 71965
rect 136955 71931 136989 71965
rect 1809 71595 1843 71629
rect 136955 71595 136989 71629
rect 1809 71259 1843 71293
rect 136955 71259 136989 71293
rect 1809 70923 1843 70957
rect 136955 70923 136989 70957
rect 1809 70587 1843 70621
rect 136955 70587 136989 70621
rect 1809 70251 1843 70285
rect 136955 70251 136989 70285
rect 1809 69915 1843 69949
rect 136955 69915 136989 69949
rect 1809 69579 1843 69613
rect 136955 69579 136989 69613
rect 1809 69243 1843 69277
rect 136955 69243 136989 69277
rect 1809 68907 1843 68941
rect 136955 68907 136989 68941
rect 1809 68571 1843 68605
rect 136955 68571 136989 68605
rect 1809 68235 1843 68269
rect 136955 68235 136989 68269
rect 1809 67899 1843 67933
rect 136955 67899 136989 67933
rect 1809 67563 1843 67597
rect 136955 67563 136989 67597
rect 1809 67227 1843 67261
rect 136955 67227 136989 67261
rect 1809 66891 1843 66925
rect 136955 66891 136989 66925
rect 1809 66555 1843 66589
rect 136955 66555 136989 66589
rect 1809 66219 1843 66253
rect 136955 66219 136989 66253
rect 1809 65883 1843 65917
rect 136955 65883 136989 65917
rect 1809 65547 1843 65581
rect 136955 65547 136989 65581
rect 1809 65211 1843 65245
rect 136955 65211 136989 65245
rect 1809 64875 1843 64909
rect 136955 64875 136989 64909
rect 1809 64539 1843 64573
rect 136955 64539 136989 64573
rect 1809 64203 1843 64237
rect 136955 64203 136989 64237
rect 1809 63867 1843 63901
rect 136955 63867 136989 63901
rect 1809 63531 1843 63565
rect 136955 63531 136989 63565
rect 1809 63195 1843 63229
rect 136955 63195 136989 63229
rect 1809 62859 1843 62893
rect 136955 62859 136989 62893
rect 1809 62523 1843 62557
rect 136955 62523 136989 62557
rect 1809 62187 1843 62221
rect 136955 62187 136989 62221
rect 1809 61851 1843 61885
rect 136955 61851 136989 61885
rect 1809 61515 1843 61549
rect 136955 61515 136989 61549
rect 1809 61179 1843 61213
rect 136955 61179 136989 61213
rect 1809 60843 1843 60877
rect 136955 60843 136989 60877
rect 1809 60507 1843 60541
rect 136955 60507 136989 60541
rect 1809 60171 1843 60205
rect 136955 60171 136989 60205
rect 1809 59835 1843 59869
rect 136955 59835 136989 59869
rect 1809 59499 1843 59533
rect 136955 59499 136989 59533
rect 1809 59163 1843 59197
rect 136955 59163 136989 59197
rect 1809 58827 1843 58861
rect 136955 58827 136989 58861
rect 1809 58491 1843 58525
rect 136955 58491 136989 58525
rect 1809 58155 1843 58189
rect 136955 58155 136989 58189
rect 1809 57819 1843 57853
rect 136955 57819 136989 57853
rect 1809 57483 1843 57517
rect 136955 57483 136989 57517
rect 1809 57147 1843 57181
rect 136955 57147 136989 57181
rect 1809 56811 1843 56845
rect 136955 56811 136989 56845
rect 1809 56475 1843 56509
rect 136955 56475 136989 56509
rect 1809 56139 1843 56173
rect 136955 56139 136989 56173
rect 1809 55803 1843 55837
rect 136955 55803 136989 55837
rect 1809 55467 1843 55501
rect 136955 55467 136989 55501
rect 1809 55131 1843 55165
rect 136955 55131 136989 55165
rect 1809 54795 1843 54829
rect 136955 54795 136989 54829
rect 1809 54459 1843 54493
rect 136955 54459 136989 54493
rect 1809 54123 1843 54157
rect 136955 54123 136989 54157
rect 1809 53787 1843 53821
rect 136955 53787 136989 53821
rect 1809 53451 1843 53485
rect 136955 53451 136989 53485
rect 1809 53115 1843 53149
rect 136955 53115 136989 53149
rect 1809 52779 1843 52813
rect 136955 52779 136989 52813
rect 1809 52443 1843 52477
rect 136955 52443 136989 52477
rect 1809 52107 1843 52141
rect 136955 52107 136989 52141
rect 1809 51771 1843 51805
rect 136955 51771 136989 51805
rect 1809 51435 1843 51469
rect 136955 51435 136989 51469
rect 1809 51099 1843 51133
rect 136955 51099 136989 51133
rect 1809 50763 1843 50797
rect 136955 50763 136989 50797
rect 1809 50427 1843 50461
rect 136955 50427 136989 50461
rect 1809 50091 1843 50125
rect 136955 50091 136989 50125
rect 1809 49755 1843 49789
rect 136955 49755 136989 49789
rect 1809 49419 1843 49453
rect 136955 49419 136989 49453
rect 1809 49083 1843 49117
rect 136955 49083 136989 49117
rect 1809 48747 1843 48781
rect 136955 48747 136989 48781
rect 1809 48411 1843 48445
rect 136955 48411 136989 48445
rect 1809 48075 1843 48109
rect 136955 48075 136989 48109
rect 1809 47739 1843 47773
rect 136955 47739 136989 47773
rect 1809 47403 1843 47437
rect 136955 47403 136989 47437
rect 1809 47067 1843 47101
rect 136955 47067 136989 47101
rect 1809 46731 1843 46765
rect 136955 46731 136989 46765
rect 1809 46395 1843 46429
rect 136955 46395 136989 46429
rect 1809 46059 1843 46093
rect 136955 46059 136989 46093
rect 1809 45723 1843 45757
rect 136955 45723 136989 45757
rect 1809 45387 1843 45421
rect 136955 45387 136989 45421
rect 1809 45051 1843 45085
rect 136955 45051 136989 45085
rect 1809 44715 1843 44749
rect 136955 44715 136989 44749
rect 1809 44379 1843 44413
rect 136955 44379 136989 44413
rect 1809 44043 1843 44077
rect 136955 44043 136989 44077
rect 1809 43707 1843 43741
rect 136955 43707 136989 43741
rect 1809 43371 1843 43405
rect 136955 43371 136989 43405
rect 1809 43035 1843 43069
rect 136955 43035 136989 43069
rect 1809 42699 1843 42733
rect 136955 42699 136989 42733
rect 1809 42363 1843 42397
rect 136955 42363 136989 42397
rect 1809 42027 1843 42061
rect 136955 42027 136989 42061
rect 1809 41691 1843 41725
rect 136955 41691 136989 41725
rect 1809 41355 1843 41389
rect 136955 41355 136989 41389
rect 1809 41019 1843 41053
rect 136955 41019 136989 41053
rect 1809 40683 1843 40717
rect 136955 40683 136989 40717
rect 1809 40347 1843 40381
rect 136955 40347 136989 40381
rect 1809 40011 1843 40045
rect 136955 40011 136989 40045
rect 1809 39675 1843 39709
rect 136955 39675 136989 39709
rect 1809 39339 1843 39373
rect 136955 39339 136989 39373
rect 1809 39003 1843 39037
rect 136955 39003 136989 39037
rect 1809 38667 1843 38701
rect 136955 38667 136989 38701
rect 1809 38331 1843 38365
rect 136955 38331 136989 38365
rect 1809 37995 1843 38029
rect 136955 37995 136989 38029
rect 1809 37659 1843 37693
rect 136955 37659 136989 37693
rect 1809 37323 1843 37357
rect 136955 37323 136989 37357
rect 1809 36987 1843 37021
rect 136955 36987 136989 37021
rect 1809 36651 1843 36685
rect 136955 36651 136989 36685
rect 1809 36315 1843 36349
rect 136955 36315 136989 36349
rect 1809 35979 1843 36013
rect 136955 35979 136989 36013
rect 1809 35643 1843 35677
rect 136955 35643 136989 35677
rect 1809 35307 1843 35341
rect 136955 35307 136989 35341
rect 1809 34971 1843 35005
rect 136955 34971 136989 35005
rect 1809 34635 1843 34669
rect 136955 34635 136989 34669
rect 1809 34299 1843 34333
rect 136955 34299 136989 34333
rect 1809 33963 1843 33997
rect 136955 33963 136989 33997
rect 1809 33627 1843 33661
rect 136955 33627 136989 33661
rect 1809 33291 1843 33325
rect 136955 33291 136989 33325
rect 1809 32955 1843 32989
rect 136955 32955 136989 32989
rect 1809 32619 1843 32653
rect 136955 32619 136989 32653
rect 1809 32283 1843 32317
rect 136955 32283 136989 32317
rect 1809 31947 1843 31981
rect 136955 31947 136989 31981
rect 1809 31611 1843 31645
rect 136955 31611 136989 31645
rect 1809 31275 1843 31309
rect 136955 31275 136989 31309
rect 1809 30939 1843 30973
rect 136955 30939 136989 30973
rect 1809 30603 1843 30637
rect 136955 30603 136989 30637
rect 1809 30267 1843 30301
rect 136955 30267 136989 30301
rect 1809 29931 1843 29965
rect 136955 29931 136989 29965
rect 1809 29595 1843 29629
rect 136955 29595 136989 29629
rect 1809 29259 1843 29293
rect 136955 29259 136989 29293
rect 1809 28923 1843 28957
rect 136955 28923 136989 28957
rect 1809 28587 1843 28621
rect 136955 28587 136989 28621
rect 1809 28251 1843 28285
rect 136955 28251 136989 28285
rect 1809 27915 1843 27949
rect 136955 27915 136989 27949
rect 1809 27579 1843 27613
rect 136955 27579 136989 27613
rect 1809 27243 1843 27277
rect 136955 27243 136989 27277
rect 1809 26907 1843 26941
rect 136955 26907 136989 26941
rect 1809 26571 1843 26605
rect 136955 26571 136989 26605
rect 1809 26235 1843 26269
rect 136955 26235 136989 26269
rect 1809 25899 1843 25933
rect 136955 25899 136989 25933
rect 1809 25563 1843 25597
rect 136955 25563 136989 25597
rect 1809 25227 1843 25261
rect 136955 25227 136989 25261
rect 1809 24891 1843 24925
rect 136955 24891 136989 24925
rect 1809 24555 1843 24589
rect 136955 24555 136989 24589
rect 1809 24219 1843 24253
rect 136955 24219 136989 24253
rect 1809 23883 1843 23917
rect 136955 23883 136989 23917
rect 1809 23547 1843 23581
rect 136955 23547 136989 23581
rect 1809 23211 1843 23245
rect 136955 23211 136989 23245
rect 1809 22875 1843 22909
rect 136955 22875 136989 22909
rect 1809 22539 1843 22573
rect 136955 22539 136989 22573
rect 1809 22203 1843 22237
rect 136955 22203 136989 22237
rect 1809 21867 1843 21901
rect 136955 21867 136989 21901
rect 1809 21531 1843 21565
rect 136955 21531 136989 21565
rect 1809 21195 1843 21229
rect 136955 21195 136989 21229
rect 1809 20859 1843 20893
rect 136955 20859 136989 20893
rect 1809 20523 1843 20557
rect 136955 20523 136989 20557
rect 1809 20187 1843 20221
rect 136955 20187 136989 20221
rect 1809 19851 1843 19885
rect 136955 19851 136989 19885
rect 1809 19515 1843 19549
rect 136955 19515 136989 19549
rect 1809 19179 1843 19213
rect 136955 19179 136989 19213
rect 1809 18843 1843 18877
rect 136955 18843 136989 18877
rect 1809 18507 1843 18541
rect 136955 18507 136989 18541
rect 1809 18171 1843 18205
rect 136955 18171 136989 18205
rect 1809 17835 1843 17869
rect 136955 17835 136989 17869
rect 1809 17499 1843 17533
rect 136955 17499 136989 17533
rect 1809 17163 1843 17197
rect 136955 17163 136989 17197
rect 1809 16827 1843 16861
rect 136955 16827 136989 16861
rect 1809 16491 1843 16525
rect 136955 16491 136989 16525
rect 1809 16155 1843 16189
rect 136955 16155 136989 16189
rect 1809 15819 1843 15853
rect 136955 15819 136989 15853
rect 1809 15483 1843 15517
rect 136955 15483 136989 15517
rect 1809 15147 1843 15181
rect 136955 15147 136989 15181
rect 1809 14811 1843 14845
rect 136955 14811 136989 14845
rect 1809 14475 1843 14509
rect 136955 14475 136989 14509
rect 1809 14139 1843 14173
rect 136955 14139 136989 14173
rect 1809 13803 1843 13837
rect 136955 13803 136989 13837
rect 1809 13467 1843 13501
rect 136955 13467 136989 13501
rect 1809 13131 1843 13165
rect 136955 13131 136989 13165
rect 1809 12795 1843 12829
rect 136955 12795 136989 12829
rect 1809 12459 1843 12493
rect 136955 12459 136989 12493
rect 1809 12123 1843 12157
rect 136955 12123 136989 12157
rect 1809 11787 1843 11821
rect 136955 11787 136989 11821
rect 1809 11451 1843 11485
rect 136955 11451 136989 11485
rect 1809 11115 1843 11149
rect 136955 11115 136989 11149
rect 1809 10779 1843 10813
rect 136955 10779 136989 10813
rect 1809 10443 1843 10477
rect 136955 10443 136989 10477
rect 1809 10107 1843 10141
rect 136955 10107 136989 10141
rect 1809 9771 1843 9805
rect 136955 9771 136989 9805
rect 1809 9435 1843 9469
rect 136955 9435 136989 9469
rect 1809 9099 1843 9133
rect 136955 9099 136989 9133
rect 1809 8763 1843 8797
rect 136955 8763 136989 8797
rect 1809 8427 1843 8461
rect 136955 8427 136989 8461
rect 1809 8091 1843 8125
rect 136955 8091 136989 8125
rect 1809 7755 1843 7789
rect 136955 7755 136989 7789
rect 1809 7419 1843 7453
rect 136955 7419 136989 7453
rect 1809 7083 1843 7117
rect 136955 7083 136989 7117
rect 1809 6747 1843 6781
rect 136955 6747 136989 6781
rect 1809 6411 1843 6445
rect 136955 6411 136989 6445
rect 1809 6075 1843 6109
rect 136955 6075 136989 6109
rect 1809 5739 1843 5773
rect 136955 5739 136989 5773
rect 1809 5403 1843 5437
rect 136955 5403 136989 5437
rect 1809 5067 1843 5101
rect 136955 5067 136989 5101
rect 1809 4731 1843 4765
rect 136955 4731 136989 4765
rect 1809 4395 1843 4429
rect 136955 4395 136989 4429
rect 1809 4059 1843 4093
rect 136955 4059 136989 4093
rect 1809 3723 1843 3757
rect 136955 3723 136989 3757
rect 1809 3387 1843 3421
rect 136955 3387 136989 3421
rect 1809 3051 1843 3085
rect 136955 3051 136989 3085
rect 1809 2715 1843 2749
rect 136955 2715 136989 2749
rect 1809 2379 1843 2413
rect 136955 2379 136989 2413
rect 1809 2043 1843 2077
rect 136955 2043 136989 2077
rect 2145 1707 2179 1741
rect 2481 1707 2515 1741
rect 2817 1707 2851 1741
rect 3153 1707 3187 1741
rect 3489 1707 3523 1741
rect 3825 1707 3859 1741
rect 4161 1707 4195 1741
rect 4497 1707 4531 1741
rect 4833 1707 4867 1741
rect 5169 1707 5203 1741
rect 5505 1707 5539 1741
rect 5841 1707 5875 1741
rect 6177 1707 6211 1741
rect 6513 1707 6547 1741
rect 6849 1707 6883 1741
rect 7185 1707 7219 1741
rect 7521 1707 7555 1741
rect 7857 1707 7891 1741
rect 8193 1707 8227 1741
rect 8529 1707 8563 1741
rect 8865 1707 8899 1741
rect 9201 1707 9235 1741
rect 9537 1707 9571 1741
rect 9873 1707 9907 1741
rect 10209 1707 10243 1741
rect 10545 1707 10579 1741
rect 10881 1707 10915 1741
rect 11217 1707 11251 1741
rect 11553 1707 11587 1741
rect 11889 1707 11923 1741
rect 12225 1707 12259 1741
rect 12561 1707 12595 1741
rect 12897 1707 12931 1741
rect 13233 1707 13267 1741
rect 13569 1707 13603 1741
rect 13905 1707 13939 1741
rect 14241 1707 14275 1741
rect 14577 1707 14611 1741
rect 14913 1707 14947 1741
rect 15249 1707 15283 1741
rect 15585 1707 15619 1741
rect 15921 1707 15955 1741
rect 16257 1707 16291 1741
rect 16593 1707 16627 1741
rect 16929 1707 16963 1741
rect 17265 1707 17299 1741
rect 17601 1707 17635 1741
rect 17937 1707 17971 1741
rect 18273 1707 18307 1741
rect 18609 1707 18643 1741
rect 18945 1707 18979 1741
rect 19281 1707 19315 1741
rect 19617 1707 19651 1741
rect 19953 1707 19987 1741
rect 20289 1707 20323 1741
rect 20625 1707 20659 1741
rect 20961 1707 20995 1741
rect 21297 1707 21331 1741
rect 21633 1707 21667 1741
rect 21969 1707 22003 1741
rect 22305 1707 22339 1741
rect 22641 1707 22675 1741
rect 22977 1707 23011 1741
rect 23313 1707 23347 1741
rect 23649 1707 23683 1741
rect 23985 1707 24019 1741
rect 24321 1707 24355 1741
rect 24657 1707 24691 1741
rect 24993 1707 25027 1741
rect 25329 1707 25363 1741
rect 25665 1707 25699 1741
rect 26001 1707 26035 1741
rect 26337 1707 26371 1741
rect 26673 1707 26707 1741
rect 27009 1707 27043 1741
rect 27345 1707 27379 1741
rect 27681 1707 27715 1741
rect 28017 1707 28051 1741
rect 28353 1707 28387 1741
rect 28689 1707 28723 1741
rect 29025 1707 29059 1741
rect 29361 1707 29395 1741
rect 29697 1707 29731 1741
rect 30033 1707 30067 1741
rect 30369 1707 30403 1741
rect 30705 1707 30739 1741
rect 31041 1707 31075 1741
rect 31377 1707 31411 1741
rect 31713 1707 31747 1741
rect 32049 1707 32083 1741
rect 32385 1707 32419 1741
rect 32721 1707 32755 1741
rect 33057 1707 33091 1741
rect 33393 1707 33427 1741
rect 33729 1707 33763 1741
rect 34065 1707 34099 1741
rect 34401 1707 34435 1741
rect 34737 1707 34771 1741
rect 35073 1707 35107 1741
rect 35409 1707 35443 1741
rect 35745 1707 35779 1741
rect 36081 1707 36115 1741
rect 36417 1707 36451 1741
rect 36753 1707 36787 1741
rect 37089 1707 37123 1741
rect 37425 1707 37459 1741
rect 37761 1707 37795 1741
rect 38097 1707 38131 1741
rect 38433 1707 38467 1741
rect 38769 1707 38803 1741
rect 39105 1707 39139 1741
rect 39441 1707 39475 1741
rect 39777 1707 39811 1741
rect 40113 1707 40147 1741
rect 40449 1707 40483 1741
rect 40785 1707 40819 1741
rect 41121 1707 41155 1741
rect 41457 1707 41491 1741
rect 41793 1707 41827 1741
rect 42129 1707 42163 1741
rect 42465 1707 42499 1741
rect 42801 1707 42835 1741
rect 43137 1707 43171 1741
rect 43473 1707 43507 1741
rect 43809 1707 43843 1741
rect 44145 1707 44179 1741
rect 44481 1707 44515 1741
rect 44817 1707 44851 1741
rect 45153 1707 45187 1741
rect 45489 1707 45523 1741
rect 45825 1707 45859 1741
rect 46161 1707 46195 1741
rect 46497 1707 46531 1741
rect 46833 1707 46867 1741
rect 47169 1707 47203 1741
rect 47505 1707 47539 1741
rect 47841 1707 47875 1741
rect 48177 1707 48211 1741
rect 48513 1707 48547 1741
rect 48849 1707 48883 1741
rect 49185 1707 49219 1741
rect 49521 1707 49555 1741
rect 49857 1707 49891 1741
rect 50193 1707 50227 1741
rect 50529 1707 50563 1741
rect 50865 1707 50899 1741
rect 51201 1707 51235 1741
rect 51537 1707 51571 1741
rect 51873 1707 51907 1741
rect 52209 1707 52243 1741
rect 52545 1707 52579 1741
rect 52881 1707 52915 1741
rect 53217 1707 53251 1741
rect 53553 1707 53587 1741
rect 53889 1707 53923 1741
rect 54225 1707 54259 1741
rect 54561 1707 54595 1741
rect 54897 1707 54931 1741
rect 55233 1707 55267 1741
rect 55569 1707 55603 1741
rect 55905 1707 55939 1741
rect 56241 1707 56275 1741
rect 56577 1707 56611 1741
rect 56913 1707 56947 1741
rect 57249 1707 57283 1741
rect 57585 1707 57619 1741
rect 57921 1707 57955 1741
rect 58257 1707 58291 1741
rect 58593 1707 58627 1741
rect 58929 1707 58963 1741
rect 59265 1707 59299 1741
rect 59601 1707 59635 1741
rect 59937 1707 59971 1741
rect 60273 1707 60307 1741
rect 60609 1707 60643 1741
rect 60945 1707 60979 1741
rect 61281 1707 61315 1741
rect 61617 1707 61651 1741
rect 61953 1707 61987 1741
rect 62289 1707 62323 1741
rect 62625 1707 62659 1741
rect 62961 1707 62995 1741
rect 63297 1707 63331 1741
rect 63633 1707 63667 1741
rect 63969 1707 64003 1741
rect 64305 1707 64339 1741
rect 64641 1707 64675 1741
rect 64977 1707 65011 1741
rect 65313 1707 65347 1741
rect 65649 1707 65683 1741
rect 65985 1707 66019 1741
rect 66321 1707 66355 1741
rect 66657 1707 66691 1741
rect 66993 1707 67027 1741
rect 67329 1707 67363 1741
rect 67665 1707 67699 1741
rect 68001 1707 68035 1741
rect 68337 1707 68371 1741
rect 68673 1707 68707 1741
rect 69009 1707 69043 1741
rect 69345 1707 69379 1741
rect 69681 1707 69715 1741
rect 70017 1707 70051 1741
rect 70353 1707 70387 1741
rect 70689 1707 70723 1741
rect 71025 1707 71059 1741
rect 71361 1707 71395 1741
rect 71697 1707 71731 1741
rect 72033 1707 72067 1741
rect 72369 1707 72403 1741
rect 72705 1707 72739 1741
rect 73041 1707 73075 1741
rect 73377 1707 73411 1741
rect 73713 1707 73747 1741
rect 74049 1707 74083 1741
rect 74385 1707 74419 1741
rect 74721 1707 74755 1741
rect 75057 1707 75091 1741
rect 75393 1707 75427 1741
rect 75729 1707 75763 1741
rect 76065 1707 76099 1741
rect 76401 1707 76435 1741
rect 76737 1707 76771 1741
rect 77073 1707 77107 1741
rect 77409 1707 77443 1741
rect 77745 1707 77779 1741
rect 78081 1707 78115 1741
rect 78417 1707 78451 1741
rect 78753 1707 78787 1741
rect 79089 1707 79123 1741
rect 79425 1707 79459 1741
rect 79761 1707 79795 1741
rect 80097 1707 80131 1741
rect 80433 1707 80467 1741
rect 80769 1707 80803 1741
rect 81105 1707 81139 1741
rect 81441 1707 81475 1741
rect 81777 1707 81811 1741
rect 82113 1707 82147 1741
rect 82449 1707 82483 1741
rect 82785 1707 82819 1741
rect 83121 1707 83155 1741
rect 83457 1707 83491 1741
rect 83793 1707 83827 1741
rect 84129 1707 84163 1741
rect 84465 1707 84499 1741
rect 84801 1707 84835 1741
rect 85137 1707 85171 1741
rect 85473 1707 85507 1741
rect 85809 1707 85843 1741
rect 86145 1707 86179 1741
rect 86481 1707 86515 1741
rect 86817 1707 86851 1741
rect 87153 1707 87187 1741
rect 87489 1707 87523 1741
rect 87825 1707 87859 1741
rect 88161 1707 88195 1741
rect 88497 1707 88531 1741
rect 88833 1707 88867 1741
rect 89169 1707 89203 1741
rect 89505 1707 89539 1741
rect 89841 1707 89875 1741
rect 90177 1707 90211 1741
rect 90513 1707 90547 1741
rect 90849 1707 90883 1741
rect 91185 1707 91219 1741
rect 91521 1707 91555 1741
rect 91857 1707 91891 1741
rect 92193 1707 92227 1741
rect 92529 1707 92563 1741
rect 92865 1707 92899 1741
rect 93201 1707 93235 1741
rect 93537 1707 93571 1741
rect 93873 1707 93907 1741
rect 94209 1707 94243 1741
rect 94545 1707 94579 1741
rect 94881 1707 94915 1741
rect 95217 1707 95251 1741
rect 95553 1707 95587 1741
rect 95889 1707 95923 1741
rect 96225 1707 96259 1741
rect 96561 1707 96595 1741
rect 96897 1707 96931 1741
rect 97233 1707 97267 1741
rect 97569 1707 97603 1741
rect 97905 1707 97939 1741
rect 98241 1707 98275 1741
rect 98577 1707 98611 1741
rect 98913 1707 98947 1741
rect 99249 1707 99283 1741
rect 99585 1707 99619 1741
rect 99921 1707 99955 1741
rect 100257 1707 100291 1741
rect 100593 1707 100627 1741
rect 100929 1707 100963 1741
rect 101265 1707 101299 1741
rect 101601 1707 101635 1741
rect 101937 1707 101971 1741
rect 102273 1707 102307 1741
rect 102609 1707 102643 1741
rect 102945 1707 102979 1741
rect 103281 1707 103315 1741
rect 103617 1707 103651 1741
rect 103953 1707 103987 1741
rect 104289 1707 104323 1741
rect 104625 1707 104659 1741
rect 104961 1707 104995 1741
rect 105297 1707 105331 1741
rect 105633 1707 105667 1741
rect 105969 1707 106003 1741
rect 106305 1707 106339 1741
rect 106641 1707 106675 1741
rect 106977 1707 107011 1741
rect 107313 1707 107347 1741
rect 107649 1707 107683 1741
rect 107985 1707 108019 1741
rect 108321 1707 108355 1741
rect 108657 1707 108691 1741
rect 108993 1707 109027 1741
rect 109329 1707 109363 1741
rect 109665 1707 109699 1741
rect 110001 1707 110035 1741
rect 110337 1707 110371 1741
rect 110673 1707 110707 1741
rect 111009 1707 111043 1741
rect 111345 1707 111379 1741
rect 111681 1707 111715 1741
rect 112017 1707 112051 1741
rect 112353 1707 112387 1741
rect 112689 1707 112723 1741
rect 113025 1707 113059 1741
rect 113361 1707 113395 1741
rect 113697 1707 113731 1741
rect 114033 1707 114067 1741
rect 114369 1707 114403 1741
rect 114705 1707 114739 1741
rect 115041 1707 115075 1741
rect 115377 1707 115411 1741
rect 115713 1707 115747 1741
rect 116049 1707 116083 1741
rect 116385 1707 116419 1741
rect 116721 1707 116755 1741
rect 117057 1707 117091 1741
rect 117393 1707 117427 1741
rect 117729 1707 117763 1741
rect 118065 1707 118099 1741
rect 118401 1707 118435 1741
rect 118737 1707 118771 1741
rect 119073 1707 119107 1741
rect 119409 1707 119443 1741
rect 119745 1707 119779 1741
rect 120081 1707 120115 1741
rect 120417 1707 120451 1741
rect 120753 1707 120787 1741
rect 121089 1707 121123 1741
rect 121425 1707 121459 1741
rect 121761 1707 121795 1741
rect 122097 1707 122131 1741
rect 122433 1707 122467 1741
rect 122769 1707 122803 1741
rect 123105 1707 123139 1741
rect 123441 1707 123475 1741
rect 123777 1707 123811 1741
rect 124113 1707 124147 1741
rect 124449 1707 124483 1741
rect 124785 1707 124819 1741
rect 125121 1707 125155 1741
rect 125457 1707 125491 1741
rect 125793 1707 125827 1741
rect 126129 1707 126163 1741
rect 126465 1707 126499 1741
rect 126801 1707 126835 1741
rect 127137 1707 127171 1741
rect 127473 1707 127507 1741
rect 127809 1707 127843 1741
rect 128145 1707 128179 1741
rect 128481 1707 128515 1741
rect 128817 1707 128851 1741
rect 129153 1707 129187 1741
rect 129489 1707 129523 1741
rect 129825 1707 129859 1741
rect 130161 1707 130195 1741
rect 130497 1707 130531 1741
rect 130833 1707 130867 1741
rect 131169 1707 131203 1741
rect 131505 1707 131539 1741
rect 131841 1707 131875 1741
rect 132177 1707 132211 1741
rect 132513 1707 132547 1741
rect 132849 1707 132883 1741
rect 133185 1707 133219 1741
rect 133521 1707 133555 1741
rect 133857 1707 133891 1741
rect 134193 1707 134227 1741
rect 134529 1707 134563 1741
rect 134865 1707 134899 1741
rect 135201 1707 135235 1741
rect 135537 1707 135571 1741
rect 135873 1707 135907 1741
rect 136209 1707 136243 1741
rect 136545 1707 136579 1741
<< locali >>
rect 2145 132050 2179 132066
rect 2145 132000 2179 132016
rect 2481 132050 2515 132066
rect 2481 132000 2515 132016
rect 2817 132050 2851 132066
rect 2817 132000 2851 132016
rect 3153 132050 3187 132066
rect 3153 132000 3187 132016
rect 3489 132050 3523 132066
rect 3489 132000 3523 132016
rect 3825 132050 3859 132066
rect 3825 132000 3859 132016
rect 4161 132050 4195 132066
rect 4161 132000 4195 132016
rect 4497 132050 4531 132066
rect 4497 132000 4531 132016
rect 4833 132050 4867 132066
rect 4833 132000 4867 132016
rect 5169 132050 5203 132066
rect 5169 132000 5203 132016
rect 5505 132050 5539 132066
rect 5505 132000 5539 132016
rect 5841 132050 5875 132066
rect 5841 132000 5875 132016
rect 6177 132050 6211 132066
rect 6177 132000 6211 132016
rect 6513 132050 6547 132066
rect 6513 132000 6547 132016
rect 6849 132050 6883 132066
rect 6849 132000 6883 132016
rect 7185 132050 7219 132066
rect 7185 132000 7219 132016
rect 7521 132050 7555 132066
rect 7521 132000 7555 132016
rect 7857 132050 7891 132066
rect 7857 132000 7891 132016
rect 8193 132050 8227 132066
rect 8193 132000 8227 132016
rect 8529 132050 8563 132066
rect 8529 132000 8563 132016
rect 8865 132050 8899 132066
rect 8865 132000 8899 132016
rect 9201 132050 9235 132066
rect 9201 132000 9235 132016
rect 9537 132050 9571 132066
rect 9537 132000 9571 132016
rect 9873 132050 9907 132066
rect 9873 132000 9907 132016
rect 10209 132050 10243 132066
rect 10209 132000 10243 132016
rect 10545 132050 10579 132066
rect 10545 132000 10579 132016
rect 10881 132050 10915 132066
rect 10881 132000 10915 132016
rect 11217 132050 11251 132066
rect 11217 132000 11251 132016
rect 11553 132050 11587 132066
rect 11553 132000 11587 132016
rect 11889 132050 11923 132066
rect 11889 132000 11923 132016
rect 12225 132050 12259 132066
rect 12225 132000 12259 132016
rect 12561 132050 12595 132066
rect 12561 132000 12595 132016
rect 12897 132050 12931 132066
rect 12897 132000 12931 132016
rect 13233 132050 13267 132066
rect 13233 132000 13267 132016
rect 13569 132050 13603 132066
rect 13569 132000 13603 132016
rect 13905 132050 13939 132066
rect 13905 132000 13939 132016
rect 14241 132050 14275 132066
rect 14241 132000 14275 132016
rect 14577 132050 14611 132066
rect 14577 132000 14611 132016
rect 14913 132050 14947 132066
rect 14913 132000 14947 132016
rect 15249 132050 15283 132066
rect 15249 132000 15283 132016
rect 15585 132050 15619 132066
rect 15585 132000 15619 132016
rect 15921 132050 15955 132066
rect 15921 132000 15955 132016
rect 16257 132050 16291 132066
rect 16257 132000 16291 132016
rect 16593 132050 16627 132066
rect 16593 132000 16627 132016
rect 16929 132050 16963 132066
rect 16929 132000 16963 132016
rect 17265 132050 17299 132066
rect 17265 132000 17299 132016
rect 17601 132050 17635 132066
rect 17601 132000 17635 132016
rect 17937 132050 17971 132066
rect 17937 132000 17971 132016
rect 18273 132050 18307 132066
rect 18273 132000 18307 132016
rect 18609 132050 18643 132066
rect 18609 132000 18643 132016
rect 18945 132050 18979 132066
rect 18945 132000 18979 132016
rect 19281 132050 19315 132066
rect 19281 132000 19315 132016
rect 19617 132050 19651 132066
rect 19617 132000 19651 132016
rect 19953 132050 19987 132066
rect 19953 132000 19987 132016
rect 20289 132050 20323 132066
rect 20289 132000 20323 132016
rect 20625 132050 20659 132066
rect 20625 132000 20659 132016
rect 20961 132050 20995 132066
rect 20961 132000 20995 132016
rect 21297 132050 21331 132066
rect 21297 132000 21331 132016
rect 21633 132050 21667 132066
rect 21633 132000 21667 132016
rect 21969 132050 22003 132066
rect 21969 132000 22003 132016
rect 22305 132050 22339 132066
rect 22305 132000 22339 132016
rect 22641 132050 22675 132066
rect 22641 132000 22675 132016
rect 22977 132050 23011 132066
rect 22977 132000 23011 132016
rect 23313 132050 23347 132066
rect 23313 132000 23347 132016
rect 23649 132050 23683 132066
rect 23649 132000 23683 132016
rect 23985 132050 24019 132066
rect 23985 132000 24019 132016
rect 24321 132050 24355 132066
rect 24321 132000 24355 132016
rect 24657 132050 24691 132066
rect 24657 132000 24691 132016
rect 24993 132050 25027 132066
rect 24993 132000 25027 132016
rect 25329 132050 25363 132066
rect 25329 132000 25363 132016
rect 25665 132050 25699 132066
rect 25665 132000 25699 132016
rect 26001 132050 26035 132066
rect 26001 132000 26035 132016
rect 26337 132050 26371 132066
rect 26337 132000 26371 132016
rect 26673 132050 26707 132066
rect 26673 132000 26707 132016
rect 27009 132050 27043 132066
rect 27009 132000 27043 132016
rect 27345 132050 27379 132066
rect 27345 132000 27379 132016
rect 27681 132050 27715 132066
rect 27681 132000 27715 132016
rect 28017 132050 28051 132066
rect 28017 132000 28051 132016
rect 28353 132050 28387 132066
rect 28353 132000 28387 132016
rect 28689 132050 28723 132066
rect 28689 132000 28723 132016
rect 29025 132050 29059 132066
rect 29025 132000 29059 132016
rect 29361 132050 29395 132066
rect 29361 132000 29395 132016
rect 29697 132050 29731 132066
rect 29697 132000 29731 132016
rect 30033 132050 30067 132066
rect 30033 132000 30067 132016
rect 30369 132050 30403 132066
rect 30369 132000 30403 132016
rect 30705 132050 30739 132066
rect 30705 132000 30739 132016
rect 31041 132050 31075 132066
rect 31041 132000 31075 132016
rect 31377 132050 31411 132066
rect 31377 132000 31411 132016
rect 31713 132050 31747 132066
rect 31713 132000 31747 132016
rect 32049 132050 32083 132066
rect 32049 132000 32083 132016
rect 32385 132050 32419 132066
rect 32385 132000 32419 132016
rect 32721 132050 32755 132066
rect 32721 132000 32755 132016
rect 33057 132050 33091 132066
rect 33057 132000 33091 132016
rect 33393 132050 33427 132066
rect 33393 132000 33427 132016
rect 33729 132050 33763 132066
rect 33729 132000 33763 132016
rect 34065 132050 34099 132066
rect 34065 132000 34099 132016
rect 34401 132050 34435 132066
rect 34401 132000 34435 132016
rect 34737 132050 34771 132066
rect 34737 132000 34771 132016
rect 35073 132050 35107 132066
rect 35073 132000 35107 132016
rect 35409 132050 35443 132066
rect 35409 132000 35443 132016
rect 35745 132050 35779 132066
rect 35745 132000 35779 132016
rect 36081 132050 36115 132066
rect 36081 132000 36115 132016
rect 36417 132050 36451 132066
rect 36417 132000 36451 132016
rect 36753 132050 36787 132066
rect 36753 132000 36787 132016
rect 37089 132050 37123 132066
rect 37089 132000 37123 132016
rect 37425 132050 37459 132066
rect 37425 132000 37459 132016
rect 37761 132050 37795 132066
rect 37761 132000 37795 132016
rect 38097 132050 38131 132066
rect 38097 132000 38131 132016
rect 38433 132050 38467 132066
rect 38433 132000 38467 132016
rect 38769 132050 38803 132066
rect 38769 132000 38803 132016
rect 39105 132050 39139 132066
rect 39105 132000 39139 132016
rect 39441 132050 39475 132066
rect 39441 132000 39475 132016
rect 39777 132050 39811 132066
rect 39777 132000 39811 132016
rect 40113 132050 40147 132066
rect 40113 132000 40147 132016
rect 40449 132050 40483 132066
rect 40449 132000 40483 132016
rect 40785 132050 40819 132066
rect 40785 132000 40819 132016
rect 41121 132050 41155 132066
rect 41121 132000 41155 132016
rect 41457 132050 41491 132066
rect 41457 132000 41491 132016
rect 41793 132050 41827 132066
rect 41793 132000 41827 132016
rect 42129 132050 42163 132066
rect 42129 132000 42163 132016
rect 42465 132050 42499 132066
rect 42465 132000 42499 132016
rect 42801 132050 42835 132066
rect 42801 132000 42835 132016
rect 43137 132050 43171 132066
rect 43137 132000 43171 132016
rect 43473 132050 43507 132066
rect 43473 132000 43507 132016
rect 43809 132050 43843 132066
rect 43809 132000 43843 132016
rect 44145 132050 44179 132066
rect 44145 132000 44179 132016
rect 44481 132050 44515 132066
rect 44481 132000 44515 132016
rect 44817 132050 44851 132066
rect 44817 132000 44851 132016
rect 45153 132050 45187 132066
rect 45153 132000 45187 132016
rect 45489 132050 45523 132066
rect 45489 132000 45523 132016
rect 45825 132050 45859 132066
rect 45825 132000 45859 132016
rect 46161 132050 46195 132066
rect 46161 132000 46195 132016
rect 46497 132050 46531 132066
rect 46497 132000 46531 132016
rect 46833 132050 46867 132066
rect 46833 132000 46867 132016
rect 47169 132050 47203 132066
rect 47169 132000 47203 132016
rect 47505 132050 47539 132066
rect 47505 132000 47539 132016
rect 47841 132050 47875 132066
rect 47841 132000 47875 132016
rect 48177 132050 48211 132066
rect 48177 132000 48211 132016
rect 48513 132050 48547 132066
rect 48513 132000 48547 132016
rect 48849 132050 48883 132066
rect 48849 132000 48883 132016
rect 49185 132050 49219 132066
rect 49185 132000 49219 132016
rect 49521 132050 49555 132066
rect 49521 132000 49555 132016
rect 49857 132050 49891 132066
rect 49857 132000 49891 132016
rect 50193 132050 50227 132066
rect 50193 132000 50227 132016
rect 50529 132050 50563 132066
rect 50529 132000 50563 132016
rect 50865 132050 50899 132066
rect 50865 132000 50899 132016
rect 51201 132050 51235 132066
rect 51201 132000 51235 132016
rect 51537 132050 51571 132066
rect 51537 132000 51571 132016
rect 51873 132050 51907 132066
rect 51873 132000 51907 132016
rect 52209 132050 52243 132066
rect 52209 132000 52243 132016
rect 52545 132050 52579 132066
rect 52545 132000 52579 132016
rect 52881 132050 52915 132066
rect 52881 132000 52915 132016
rect 53217 132050 53251 132066
rect 53217 132000 53251 132016
rect 53553 132050 53587 132066
rect 53553 132000 53587 132016
rect 53889 132050 53923 132066
rect 53889 132000 53923 132016
rect 54225 132050 54259 132066
rect 54225 132000 54259 132016
rect 54561 132050 54595 132066
rect 54561 132000 54595 132016
rect 54897 132050 54931 132066
rect 54897 132000 54931 132016
rect 55233 132050 55267 132066
rect 55233 132000 55267 132016
rect 55569 132050 55603 132066
rect 55569 132000 55603 132016
rect 55905 132050 55939 132066
rect 55905 132000 55939 132016
rect 56241 132050 56275 132066
rect 56241 132000 56275 132016
rect 56577 132050 56611 132066
rect 56577 132000 56611 132016
rect 56913 132050 56947 132066
rect 56913 132000 56947 132016
rect 57249 132050 57283 132066
rect 57249 132000 57283 132016
rect 57585 132050 57619 132066
rect 57585 132000 57619 132016
rect 57921 132050 57955 132066
rect 57921 132000 57955 132016
rect 58257 132050 58291 132066
rect 58257 132000 58291 132016
rect 58593 132050 58627 132066
rect 58593 132000 58627 132016
rect 58929 132050 58963 132066
rect 58929 132000 58963 132016
rect 59265 132050 59299 132066
rect 59265 132000 59299 132016
rect 59601 132050 59635 132066
rect 59601 132000 59635 132016
rect 59937 132050 59971 132066
rect 59937 132000 59971 132016
rect 60273 132050 60307 132066
rect 60273 132000 60307 132016
rect 60609 132050 60643 132066
rect 60609 132000 60643 132016
rect 60945 132050 60979 132066
rect 60945 132000 60979 132016
rect 61281 132050 61315 132066
rect 61281 132000 61315 132016
rect 61617 132050 61651 132066
rect 61617 132000 61651 132016
rect 61953 132050 61987 132066
rect 61953 132000 61987 132016
rect 62289 132050 62323 132066
rect 62289 132000 62323 132016
rect 62625 132050 62659 132066
rect 62625 132000 62659 132016
rect 62961 132050 62995 132066
rect 62961 132000 62995 132016
rect 63297 132050 63331 132066
rect 63297 132000 63331 132016
rect 63633 132050 63667 132066
rect 63633 132000 63667 132016
rect 63969 132050 64003 132066
rect 63969 132000 64003 132016
rect 64305 132050 64339 132066
rect 64305 132000 64339 132016
rect 64641 132050 64675 132066
rect 64641 132000 64675 132016
rect 64977 132050 65011 132066
rect 64977 132000 65011 132016
rect 65313 132050 65347 132066
rect 65313 132000 65347 132016
rect 65649 132050 65683 132066
rect 65649 132000 65683 132016
rect 65985 132050 66019 132066
rect 65985 132000 66019 132016
rect 66321 132050 66355 132066
rect 66321 132000 66355 132016
rect 66657 132050 66691 132066
rect 66657 132000 66691 132016
rect 66993 132050 67027 132066
rect 66993 132000 67027 132016
rect 67329 132050 67363 132066
rect 67329 132000 67363 132016
rect 67665 132050 67699 132066
rect 67665 132000 67699 132016
rect 68001 132050 68035 132066
rect 68001 132000 68035 132016
rect 68337 132050 68371 132066
rect 68337 132000 68371 132016
rect 68673 132050 68707 132066
rect 68673 132000 68707 132016
rect 69009 132050 69043 132066
rect 69009 132000 69043 132016
rect 69345 132050 69379 132066
rect 69345 132000 69379 132016
rect 69681 132050 69715 132066
rect 69681 132000 69715 132016
rect 70017 132050 70051 132066
rect 70017 132000 70051 132016
rect 70353 132050 70387 132066
rect 70353 132000 70387 132016
rect 70689 132050 70723 132066
rect 70689 132000 70723 132016
rect 71025 132050 71059 132066
rect 71025 132000 71059 132016
rect 71361 132050 71395 132066
rect 71361 132000 71395 132016
rect 71697 132050 71731 132066
rect 71697 132000 71731 132016
rect 72033 132050 72067 132066
rect 72033 132000 72067 132016
rect 72369 132050 72403 132066
rect 72369 132000 72403 132016
rect 72705 132050 72739 132066
rect 72705 132000 72739 132016
rect 73041 132050 73075 132066
rect 73041 132000 73075 132016
rect 73377 132050 73411 132066
rect 73377 132000 73411 132016
rect 73713 132050 73747 132066
rect 73713 132000 73747 132016
rect 74049 132050 74083 132066
rect 74049 132000 74083 132016
rect 74385 132050 74419 132066
rect 74385 132000 74419 132016
rect 74721 132050 74755 132066
rect 74721 132000 74755 132016
rect 75057 132050 75091 132066
rect 75057 132000 75091 132016
rect 75393 132050 75427 132066
rect 75393 132000 75427 132016
rect 75729 132050 75763 132066
rect 75729 132000 75763 132016
rect 76065 132050 76099 132066
rect 76065 132000 76099 132016
rect 76401 132050 76435 132066
rect 76401 132000 76435 132016
rect 76737 132050 76771 132066
rect 76737 132000 76771 132016
rect 77073 132050 77107 132066
rect 77073 132000 77107 132016
rect 77409 132050 77443 132066
rect 77409 132000 77443 132016
rect 77745 132050 77779 132066
rect 77745 132000 77779 132016
rect 78081 132050 78115 132066
rect 78081 132000 78115 132016
rect 78417 132050 78451 132066
rect 78417 132000 78451 132016
rect 78753 132050 78787 132066
rect 78753 132000 78787 132016
rect 79089 132050 79123 132066
rect 79089 132000 79123 132016
rect 79425 132050 79459 132066
rect 79425 132000 79459 132016
rect 79761 132050 79795 132066
rect 79761 132000 79795 132016
rect 80097 132050 80131 132066
rect 80097 132000 80131 132016
rect 80433 132050 80467 132066
rect 80433 132000 80467 132016
rect 80769 132050 80803 132066
rect 80769 132000 80803 132016
rect 81105 132050 81139 132066
rect 81105 132000 81139 132016
rect 81441 132050 81475 132066
rect 81441 132000 81475 132016
rect 81777 132050 81811 132066
rect 81777 132000 81811 132016
rect 82113 132050 82147 132066
rect 82113 132000 82147 132016
rect 82449 132050 82483 132066
rect 82449 132000 82483 132016
rect 82785 132050 82819 132066
rect 82785 132000 82819 132016
rect 83121 132050 83155 132066
rect 83121 132000 83155 132016
rect 83457 132050 83491 132066
rect 83457 132000 83491 132016
rect 83793 132050 83827 132066
rect 83793 132000 83827 132016
rect 84129 132050 84163 132066
rect 84129 132000 84163 132016
rect 84465 132050 84499 132066
rect 84465 132000 84499 132016
rect 84801 132050 84835 132066
rect 84801 132000 84835 132016
rect 85137 132050 85171 132066
rect 85137 132000 85171 132016
rect 85473 132050 85507 132066
rect 85473 132000 85507 132016
rect 85809 132050 85843 132066
rect 85809 132000 85843 132016
rect 86145 132050 86179 132066
rect 86145 132000 86179 132016
rect 86481 132050 86515 132066
rect 86481 132000 86515 132016
rect 86817 132050 86851 132066
rect 86817 132000 86851 132016
rect 87153 132050 87187 132066
rect 87153 132000 87187 132016
rect 87489 132050 87523 132066
rect 87489 132000 87523 132016
rect 87825 132050 87859 132066
rect 87825 132000 87859 132016
rect 88161 132050 88195 132066
rect 88161 132000 88195 132016
rect 88497 132050 88531 132066
rect 88497 132000 88531 132016
rect 88833 132050 88867 132066
rect 88833 132000 88867 132016
rect 89169 132050 89203 132066
rect 89169 132000 89203 132016
rect 89505 132050 89539 132066
rect 89505 132000 89539 132016
rect 89841 132050 89875 132066
rect 89841 132000 89875 132016
rect 90177 132050 90211 132066
rect 90177 132000 90211 132016
rect 90513 132050 90547 132066
rect 90513 132000 90547 132016
rect 90849 132050 90883 132066
rect 90849 132000 90883 132016
rect 91185 132050 91219 132066
rect 91185 132000 91219 132016
rect 91521 132050 91555 132066
rect 91521 132000 91555 132016
rect 91857 132050 91891 132066
rect 91857 132000 91891 132016
rect 92193 132050 92227 132066
rect 92193 132000 92227 132016
rect 92529 132050 92563 132066
rect 92529 132000 92563 132016
rect 92865 132050 92899 132066
rect 92865 132000 92899 132016
rect 93201 132050 93235 132066
rect 93201 132000 93235 132016
rect 93537 132050 93571 132066
rect 93537 132000 93571 132016
rect 93873 132050 93907 132066
rect 93873 132000 93907 132016
rect 94209 132050 94243 132066
rect 94209 132000 94243 132016
rect 94545 132050 94579 132066
rect 94545 132000 94579 132016
rect 94881 132050 94915 132066
rect 94881 132000 94915 132016
rect 95217 132050 95251 132066
rect 95217 132000 95251 132016
rect 95553 132050 95587 132066
rect 95553 132000 95587 132016
rect 95889 132050 95923 132066
rect 95889 132000 95923 132016
rect 96225 132050 96259 132066
rect 96225 132000 96259 132016
rect 96561 132050 96595 132066
rect 96561 132000 96595 132016
rect 96897 132050 96931 132066
rect 96897 132000 96931 132016
rect 97233 132050 97267 132066
rect 97233 132000 97267 132016
rect 97569 132050 97603 132066
rect 97569 132000 97603 132016
rect 97905 132050 97939 132066
rect 97905 132000 97939 132016
rect 98241 132050 98275 132066
rect 98241 132000 98275 132016
rect 98577 132050 98611 132066
rect 98577 132000 98611 132016
rect 98913 132050 98947 132066
rect 98913 132000 98947 132016
rect 99249 132050 99283 132066
rect 99249 132000 99283 132016
rect 99585 132050 99619 132066
rect 99585 132000 99619 132016
rect 99921 132050 99955 132066
rect 99921 132000 99955 132016
rect 100257 132050 100291 132066
rect 100257 132000 100291 132016
rect 100593 132050 100627 132066
rect 100593 132000 100627 132016
rect 100929 132050 100963 132066
rect 100929 132000 100963 132016
rect 101265 132050 101299 132066
rect 101265 132000 101299 132016
rect 101601 132050 101635 132066
rect 101601 132000 101635 132016
rect 101937 132050 101971 132066
rect 101937 132000 101971 132016
rect 102273 132050 102307 132066
rect 102273 132000 102307 132016
rect 102609 132050 102643 132066
rect 102609 132000 102643 132016
rect 102945 132050 102979 132066
rect 102945 132000 102979 132016
rect 103281 132050 103315 132066
rect 103281 132000 103315 132016
rect 103617 132050 103651 132066
rect 103617 132000 103651 132016
rect 103953 132050 103987 132066
rect 103953 132000 103987 132016
rect 104289 132050 104323 132066
rect 104289 132000 104323 132016
rect 104625 132050 104659 132066
rect 104625 132000 104659 132016
rect 104961 132050 104995 132066
rect 104961 132000 104995 132016
rect 105297 132050 105331 132066
rect 105297 132000 105331 132016
rect 105633 132050 105667 132066
rect 105633 132000 105667 132016
rect 105969 132050 106003 132066
rect 105969 132000 106003 132016
rect 106305 132050 106339 132066
rect 106305 132000 106339 132016
rect 106641 132050 106675 132066
rect 106641 132000 106675 132016
rect 106977 132050 107011 132066
rect 106977 132000 107011 132016
rect 107313 132050 107347 132066
rect 107313 132000 107347 132016
rect 107649 132050 107683 132066
rect 107649 132000 107683 132016
rect 107985 132050 108019 132066
rect 107985 132000 108019 132016
rect 108321 132050 108355 132066
rect 108321 132000 108355 132016
rect 108657 132050 108691 132066
rect 108657 132000 108691 132016
rect 108993 132050 109027 132066
rect 108993 132000 109027 132016
rect 109329 132050 109363 132066
rect 109329 132000 109363 132016
rect 109665 132050 109699 132066
rect 109665 132000 109699 132016
rect 110001 132050 110035 132066
rect 110001 132000 110035 132016
rect 110337 132050 110371 132066
rect 110337 132000 110371 132016
rect 110673 132050 110707 132066
rect 110673 132000 110707 132016
rect 111009 132050 111043 132066
rect 111009 132000 111043 132016
rect 111345 132050 111379 132066
rect 111345 132000 111379 132016
rect 111681 132050 111715 132066
rect 111681 132000 111715 132016
rect 112017 132050 112051 132066
rect 112017 132000 112051 132016
rect 112353 132050 112387 132066
rect 112353 132000 112387 132016
rect 112689 132050 112723 132066
rect 112689 132000 112723 132016
rect 113025 132050 113059 132066
rect 113025 132000 113059 132016
rect 113361 132050 113395 132066
rect 113361 132000 113395 132016
rect 113697 132050 113731 132066
rect 113697 132000 113731 132016
rect 114033 132050 114067 132066
rect 114033 132000 114067 132016
rect 114369 132050 114403 132066
rect 114369 132000 114403 132016
rect 114705 132050 114739 132066
rect 114705 132000 114739 132016
rect 115041 132050 115075 132066
rect 115041 132000 115075 132016
rect 115377 132050 115411 132066
rect 115377 132000 115411 132016
rect 115713 132050 115747 132066
rect 115713 132000 115747 132016
rect 116049 132050 116083 132066
rect 116049 132000 116083 132016
rect 116385 132050 116419 132066
rect 116385 132000 116419 132016
rect 116721 132050 116755 132066
rect 116721 132000 116755 132016
rect 117057 132050 117091 132066
rect 117057 132000 117091 132016
rect 117393 132050 117427 132066
rect 117393 132000 117427 132016
rect 117729 132050 117763 132066
rect 117729 132000 117763 132016
rect 118065 132050 118099 132066
rect 118065 132000 118099 132016
rect 118401 132050 118435 132066
rect 118401 132000 118435 132016
rect 118737 132050 118771 132066
rect 118737 132000 118771 132016
rect 119073 132050 119107 132066
rect 119073 132000 119107 132016
rect 119409 132050 119443 132066
rect 119409 132000 119443 132016
rect 119745 132050 119779 132066
rect 119745 132000 119779 132016
rect 120081 132050 120115 132066
rect 120081 132000 120115 132016
rect 120417 132050 120451 132066
rect 120417 132000 120451 132016
rect 120753 132050 120787 132066
rect 120753 132000 120787 132016
rect 121089 132050 121123 132066
rect 121089 132000 121123 132016
rect 121425 132050 121459 132066
rect 121425 132000 121459 132016
rect 121761 132050 121795 132066
rect 121761 132000 121795 132016
rect 122097 132050 122131 132066
rect 122097 132000 122131 132016
rect 122433 132050 122467 132066
rect 122433 132000 122467 132016
rect 122769 132050 122803 132066
rect 122769 132000 122803 132016
rect 123105 132050 123139 132066
rect 123105 132000 123139 132016
rect 123441 132050 123475 132066
rect 123441 132000 123475 132016
rect 123777 132050 123811 132066
rect 123777 132000 123811 132016
rect 124113 132050 124147 132066
rect 124113 132000 124147 132016
rect 124449 132050 124483 132066
rect 124449 132000 124483 132016
rect 124785 132050 124819 132066
rect 124785 132000 124819 132016
rect 125121 132050 125155 132066
rect 125121 132000 125155 132016
rect 125457 132050 125491 132066
rect 125457 132000 125491 132016
rect 125793 132050 125827 132066
rect 125793 132000 125827 132016
rect 126129 132050 126163 132066
rect 126129 132000 126163 132016
rect 126465 132050 126499 132066
rect 126465 132000 126499 132016
rect 126801 132050 126835 132066
rect 126801 132000 126835 132016
rect 127137 132050 127171 132066
rect 127137 132000 127171 132016
rect 127473 132050 127507 132066
rect 127473 132000 127507 132016
rect 127809 132050 127843 132066
rect 127809 132000 127843 132016
rect 128145 132050 128179 132066
rect 128145 132000 128179 132016
rect 128481 132050 128515 132066
rect 128481 132000 128515 132016
rect 128817 132050 128851 132066
rect 128817 132000 128851 132016
rect 129153 132050 129187 132066
rect 129153 132000 129187 132016
rect 129489 132050 129523 132066
rect 129489 132000 129523 132016
rect 129825 132050 129859 132066
rect 129825 132000 129859 132016
rect 130161 132050 130195 132066
rect 130161 132000 130195 132016
rect 130497 132050 130531 132066
rect 130497 132000 130531 132016
rect 130833 132050 130867 132066
rect 130833 132000 130867 132016
rect 131169 132050 131203 132066
rect 131169 132000 131203 132016
rect 131505 132050 131539 132066
rect 131505 132000 131539 132016
rect 131841 132050 131875 132066
rect 131841 132000 131875 132016
rect 132177 132050 132211 132066
rect 132177 132000 132211 132016
rect 132513 132050 132547 132066
rect 132513 132000 132547 132016
rect 132849 132050 132883 132066
rect 132849 132000 132883 132016
rect 133185 132050 133219 132066
rect 133185 132000 133219 132016
rect 133521 132050 133555 132066
rect 133521 132000 133555 132016
rect 133857 132050 133891 132066
rect 133857 132000 133891 132016
rect 134193 132050 134227 132066
rect 134193 132000 134227 132016
rect 134529 132050 134563 132066
rect 134529 132000 134563 132016
rect 134865 132050 134899 132066
rect 134865 132000 134899 132016
rect 135201 132050 135235 132066
rect 135201 132000 135235 132016
rect 135537 132050 135571 132066
rect 135537 132000 135571 132016
rect 135873 132050 135907 132066
rect 135873 132000 135907 132016
rect 136209 132050 136243 132066
rect 136209 132000 136243 132016
rect 136545 132050 136579 132066
rect 136545 132000 136579 132016
rect 1809 131437 1843 131453
rect 1809 131387 1843 131403
rect 136955 131437 136989 131453
rect 136955 131387 136989 131403
rect 1809 131101 1843 131117
rect 1809 131051 1843 131067
rect 136955 131101 136989 131117
rect 136955 131051 136989 131067
rect 1809 130765 1843 130781
rect 1809 130715 1843 130731
rect 136955 130765 136989 130781
rect 136955 130715 136989 130731
rect 1809 130429 1843 130445
rect 1809 130379 1843 130395
rect 136955 130429 136989 130445
rect 136955 130379 136989 130395
rect 1809 130093 1843 130109
rect 1809 130043 1843 130059
rect 136955 130093 136989 130109
rect 136955 130043 136989 130059
rect 1809 129757 1843 129773
rect 1809 129707 1843 129723
rect 136955 129757 136989 129773
rect 136955 129707 136989 129723
rect 1809 129421 1843 129437
rect 1809 129371 1843 129387
rect 136955 129421 136989 129437
rect 136955 129371 136989 129387
rect 1809 129085 1843 129101
rect 1809 129035 1843 129051
rect 136955 129085 136989 129101
rect 136955 129035 136989 129051
rect 1809 128749 1843 128765
rect 1809 128699 1843 128715
rect 136955 128749 136989 128765
rect 136955 128699 136989 128715
rect 1809 128413 1843 128429
rect 1809 128363 1843 128379
rect 136955 128413 136989 128429
rect 136955 128363 136989 128379
rect 1809 128077 1843 128093
rect 1809 128027 1843 128043
rect 136955 128077 136989 128093
rect 136955 128027 136989 128043
rect 1809 127741 1843 127757
rect 1809 127691 1843 127707
rect 136955 127741 136989 127757
rect 136955 127691 136989 127707
rect 1809 127405 1843 127421
rect 1809 127355 1843 127371
rect 136955 127405 136989 127421
rect 136955 127355 136989 127371
rect 1809 127069 1843 127085
rect 1809 127019 1843 127035
rect 136955 127069 136989 127085
rect 136955 127019 136989 127035
rect 1809 126733 1843 126749
rect 1809 126683 1843 126699
rect 136955 126733 136989 126749
rect 136955 126683 136989 126699
rect 1809 126397 1843 126413
rect 1809 126347 1843 126363
rect 136955 126397 136989 126413
rect 136955 126347 136989 126363
rect 1809 126061 1843 126077
rect 1809 126011 1843 126027
rect 136955 126061 136989 126077
rect 136955 126011 136989 126027
rect 1809 125725 1843 125741
rect 1809 125675 1843 125691
rect 136955 125725 136989 125741
rect 136955 125675 136989 125691
rect 1809 125389 1843 125405
rect 1809 125339 1843 125355
rect 136955 125389 136989 125405
rect 136955 125339 136989 125355
rect 1809 125053 1843 125069
rect 1809 125003 1843 125019
rect 136955 125053 136989 125069
rect 136955 125003 136989 125019
rect 1809 124717 1843 124733
rect 1809 124667 1843 124683
rect 136955 124717 136989 124733
rect 136955 124667 136989 124683
rect 1809 124381 1843 124397
rect 1809 124331 1843 124347
rect 136955 124381 136989 124397
rect 136955 124331 136989 124347
rect 1809 124045 1843 124061
rect 1809 123995 1843 124011
rect 136955 124045 136989 124061
rect 136955 123995 136989 124011
rect 1809 123709 1843 123725
rect 1809 123659 1843 123675
rect 136955 123709 136989 123725
rect 136955 123659 136989 123675
rect 1809 123373 1843 123389
rect 1809 123323 1843 123339
rect 136955 123373 136989 123389
rect 136955 123323 136989 123339
rect 1809 123037 1843 123053
rect 1809 122987 1843 123003
rect 136955 123037 136989 123053
rect 136955 122987 136989 123003
rect 1809 122701 1843 122717
rect 1809 122651 1843 122667
rect 136955 122701 136989 122717
rect 136955 122651 136989 122667
rect 1809 122365 1843 122381
rect 1809 122315 1843 122331
rect 136955 122365 136989 122381
rect 136955 122315 136989 122331
rect 1809 122029 1843 122045
rect 1809 121979 1843 121995
rect 136955 122029 136989 122045
rect 136955 121979 136989 121995
rect 1809 121693 1843 121709
rect 1809 121643 1843 121659
rect 136955 121693 136989 121709
rect 136955 121643 136989 121659
rect 1809 121357 1843 121373
rect 1809 121307 1843 121323
rect 136955 121357 136989 121373
rect 136955 121307 136989 121323
rect 1809 121021 1843 121037
rect 1809 120971 1843 120987
rect 136955 121021 136989 121037
rect 136955 120971 136989 120987
rect 1809 120685 1843 120701
rect 1809 120635 1843 120651
rect 136955 120685 136989 120701
rect 136955 120635 136989 120651
rect 1809 120349 1843 120365
rect 1809 120299 1843 120315
rect 136955 120349 136989 120365
rect 136955 120299 136989 120315
rect 1809 120013 1843 120029
rect 1809 119963 1843 119979
rect 136955 120013 136989 120029
rect 136955 119963 136989 119979
rect 1809 119677 1843 119693
rect 1809 119627 1843 119643
rect 136955 119677 136989 119693
rect 136955 119627 136989 119643
rect 1809 119341 1843 119357
rect 1809 119291 1843 119307
rect 136955 119341 136989 119357
rect 136955 119291 136989 119307
rect 1809 119005 1843 119021
rect 1809 118955 1843 118971
rect 136955 119005 136989 119021
rect 136955 118955 136989 118971
rect 1809 118669 1843 118685
rect 1809 118619 1843 118635
rect 136955 118669 136989 118685
rect 136955 118619 136989 118635
rect 1809 118333 1843 118349
rect 1809 118283 1843 118299
rect 136955 118333 136989 118349
rect 136955 118283 136989 118299
rect 1809 117997 1843 118013
rect 1809 117947 1843 117963
rect 136955 117997 136989 118013
rect 136955 117947 136989 117963
rect 1809 117661 1843 117677
rect 1809 117611 1843 117627
rect 136955 117661 136989 117677
rect 136955 117611 136989 117627
rect 1809 117325 1843 117341
rect 1809 117275 1843 117291
rect 136955 117325 136989 117341
rect 136955 117275 136989 117291
rect 1809 116989 1843 117005
rect 1809 116939 1843 116955
rect 136955 116989 136989 117005
rect 136955 116939 136989 116955
rect 1809 116653 1843 116669
rect 1809 116603 1843 116619
rect 136955 116653 136989 116669
rect 136955 116603 136989 116619
rect 1809 116317 1843 116333
rect 1809 116267 1843 116283
rect 136955 116317 136989 116333
rect 136955 116267 136989 116283
rect 1809 115981 1843 115997
rect 1809 115931 1843 115947
rect 136955 115981 136989 115997
rect 136955 115931 136989 115947
rect 1809 115645 1843 115661
rect 1809 115595 1843 115611
rect 136955 115645 136989 115661
rect 136955 115595 136989 115611
rect 1809 115309 1843 115325
rect 1809 115259 1843 115275
rect 136955 115309 136989 115325
rect 136955 115259 136989 115275
rect 1809 114973 1843 114989
rect 1809 114923 1843 114939
rect 136955 114973 136989 114989
rect 136955 114923 136989 114939
rect 1809 114637 1843 114653
rect 1809 114587 1843 114603
rect 136955 114637 136989 114653
rect 136955 114587 136989 114603
rect 1809 114301 1843 114317
rect 1809 114251 1843 114267
rect 136955 114301 136989 114317
rect 136955 114251 136989 114267
rect 1809 113965 1843 113981
rect 1809 113915 1843 113931
rect 136955 113965 136989 113981
rect 136955 113915 136989 113931
rect 1809 113629 1843 113645
rect 1809 113579 1843 113595
rect 136955 113629 136989 113645
rect 136955 113579 136989 113595
rect 1809 113293 1843 113309
rect 1809 113243 1843 113259
rect 136955 113293 136989 113309
rect 136955 113243 136989 113259
rect 1809 112957 1843 112973
rect 1809 112907 1843 112923
rect 136955 112957 136989 112973
rect 136955 112907 136989 112923
rect 1809 112621 1843 112637
rect 1809 112571 1843 112587
rect 136955 112621 136989 112637
rect 136955 112571 136989 112587
rect 1809 112285 1843 112301
rect 1809 112235 1843 112251
rect 136955 112285 136989 112301
rect 136955 112235 136989 112251
rect 1809 111949 1843 111965
rect 1809 111899 1843 111915
rect 136955 111949 136989 111965
rect 136955 111899 136989 111915
rect 1809 111613 1843 111629
rect 1809 111563 1843 111579
rect 136955 111613 136989 111629
rect 136955 111563 136989 111579
rect 1809 111277 1843 111293
rect 1809 111227 1843 111243
rect 136955 111277 136989 111293
rect 136955 111227 136989 111243
rect 1809 110941 1843 110957
rect 1809 110891 1843 110907
rect 136955 110941 136989 110957
rect 136955 110891 136989 110907
rect 1809 110605 1843 110621
rect 1809 110555 1843 110571
rect 136955 110605 136989 110621
rect 136955 110555 136989 110571
rect 1809 110269 1843 110285
rect 1809 110219 1843 110235
rect 136955 110269 136989 110285
rect 136955 110219 136989 110235
rect 1809 109933 1843 109949
rect 1809 109883 1843 109899
rect 136955 109933 136989 109949
rect 136955 109883 136989 109899
rect 1809 109597 1843 109613
rect 1809 109547 1843 109563
rect 136955 109597 136989 109613
rect 136955 109547 136989 109563
rect 1809 109261 1843 109277
rect 1809 109211 1843 109227
rect 136955 109261 136989 109277
rect 136955 109211 136989 109227
rect 1809 108925 1843 108941
rect 1809 108875 1843 108891
rect 136955 108925 136989 108941
rect 136955 108875 136989 108891
rect 1809 108589 1843 108605
rect 1809 108539 1843 108555
rect 136955 108589 136989 108605
rect 136955 108539 136989 108555
rect 1809 108253 1843 108269
rect 1809 108203 1843 108219
rect 136955 108253 136989 108269
rect 136955 108203 136989 108219
rect 1809 107917 1843 107933
rect 1809 107867 1843 107883
rect 136955 107917 136989 107933
rect 136955 107867 136989 107883
rect 1809 107581 1843 107597
rect 1809 107531 1843 107547
rect 136955 107581 136989 107597
rect 136955 107531 136989 107547
rect 1809 107245 1843 107261
rect 1809 107195 1843 107211
rect 136955 107245 136989 107261
rect 136955 107195 136989 107211
rect 1809 106909 1843 106925
rect 1809 106859 1843 106875
rect 136955 106909 136989 106925
rect 136955 106859 136989 106875
rect 1809 106573 1843 106589
rect 1809 106523 1843 106539
rect 136955 106573 136989 106589
rect 136955 106523 136989 106539
rect 1809 106237 1843 106253
rect 1809 106187 1843 106203
rect 136955 106237 136989 106253
rect 136955 106187 136989 106203
rect 1809 105901 1843 105917
rect 1809 105851 1843 105867
rect 136955 105901 136989 105917
rect 136955 105851 136989 105867
rect 1809 105565 1843 105581
rect 1809 105515 1843 105531
rect 136955 105565 136989 105581
rect 136955 105515 136989 105531
rect 1809 105229 1843 105245
rect 1809 105179 1843 105195
rect 136955 105229 136989 105245
rect 136955 105179 136989 105195
rect 1809 104893 1843 104909
rect 1809 104843 1843 104859
rect 136955 104893 136989 104909
rect 136955 104843 136989 104859
rect 1809 104557 1843 104573
rect 1809 104507 1843 104523
rect 136955 104557 136989 104573
rect 136955 104507 136989 104523
rect 1809 104221 1843 104237
rect 1809 104171 1843 104187
rect 136955 104221 136989 104237
rect 136955 104171 136989 104187
rect 1809 103885 1843 103901
rect 1809 103835 1843 103851
rect 136955 103885 136989 103901
rect 136955 103835 136989 103851
rect 1809 103549 1843 103565
rect 1809 103499 1843 103515
rect 136955 103549 136989 103565
rect 136955 103499 136989 103515
rect 1809 103213 1843 103229
rect 1809 103163 1843 103179
rect 136955 103213 136989 103229
rect 136955 103163 136989 103179
rect 1809 102877 1843 102893
rect 1809 102827 1843 102843
rect 136955 102877 136989 102893
rect 136955 102827 136989 102843
rect 1809 102541 1843 102557
rect 1809 102491 1843 102507
rect 136955 102541 136989 102557
rect 136955 102491 136989 102507
rect 1809 102205 1843 102221
rect 1809 102155 1843 102171
rect 136955 102205 136989 102221
rect 136955 102155 136989 102171
rect 1809 101869 1843 101885
rect 1809 101819 1843 101835
rect 136955 101869 136989 101885
rect 136955 101819 136989 101835
rect 1809 101533 1843 101549
rect 1809 101483 1843 101499
rect 136955 101533 136989 101549
rect 136955 101483 136989 101499
rect 1809 101197 1843 101213
rect 1809 101147 1843 101163
rect 136955 101197 136989 101213
rect 136955 101147 136989 101163
rect 1809 100861 1843 100877
rect 1809 100811 1843 100827
rect 136955 100861 136989 100877
rect 136955 100811 136989 100827
rect 1809 100525 1843 100541
rect 1809 100475 1843 100491
rect 136955 100525 136989 100541
rect 136955 100475 136989 100491
rect 1809 100189 1843 100205
rect 1809 100139 1843 100155
rect 136955 100189 136989 100205
rect 136955 100139 136989 100155
rect 1809 99853 1843 99869
rect 1809 99803 1843 99819
rect 136955 99853 136989 99869
rect 136955 99803 136989 99819
rect 1809 99517 1843 99533
rect 1809 99467 1843 99483
rect 136955 99517 136989 99533
rect 136955 99467 136989 99483
rect 1809 99181 1843 99197
rect 1809 99131 1843 99147
rect 136955 99181 136989 99197
rect 136955 99131 136989 99147
rect 1809 98845 1843 98861
rect 1809 98795 1843 98811
rect 136955 98845 136989 98861
rect 136955 98795 136989 98811
rect 1809 98509 1843 98525
rect 1809 98459 1843 98475
rect 136955 98509 136989 98525
rect 136955 98459 136989 98475
rect 1809 98173 1843 98189
rect 1809 98123 1843 98139
rect 136955 98173 136989 98189
rect 136955 98123 136989 98139
rect 1809 97837 1843 97853
rect 1809 97787 1843 97803
rect 136955 97837 136989 97853
rect 136955 97787 136989 97803
rect 1809 97501 1843 97517
rect 1809 97451 1843 97467
rect 136955 97501 136989 97517
rect 136955 97451 136989 97467
rect 1809 97165 1843 97181
rect 1809 97115 1843 97131
rect 136955 97165 136989 97181
rect 136955 97115 136989 97131
rect 1809 96829 1843 96845
rect 1809 96779 1843 96795
rect 136955 96829 136989 96845
rect 136955 96779 136989 96795
rect 1809 96493 1843 96509
rect 1809 96443 1843 96459
rect 136955 96493 136989 96509
rect 136955 96443 136989 96459
rect 1809 96157 1843 96173
rect 1809 96107 1843 96123
rect 136955 96157 136989 96173
rect 136955 96107 136989 96123
rect 1809 95821 1843 95837
rect 1809 95771 1843 95787
rect 136955 95821 136989 95837
rect 136955 95771 136989 95787
rect 1809 95485 1843 95501
rect 1809 95435 1843 95451
rect 136955 95485 136989 95501
rect 136955 95435 136989 95451
rect 1809 95149 1843 95165
rect 1809 95099 1843 95115
rect 136955 95149 136989 95165
rect 136955 95099 136989 95115
rect 1809 94813 1843 94829
rect 1809 94763 1843 94779
rect 136955 94813 136989 94829
rect 136955 94763 136989 94779
rect 1809 94477 1843 94493
rect 1809 94427 1843 94443
rect 136955 94477 136989 94493
rect 136955 94427 136989 94443
rect 1809 94141 1843 94157
rect 1809 94091 1843 94107
rect 136955 94141 136989 94157
rect 136955 94091 136989 94107
rect 1809 93805 1843 93821
rect 1809 93755 1843 93771
rect 136955 93805 136989 93821
rect 136955 93755 136989 93771
rect 1809 93469 1843 93485
rect 1809 93419 1843 93435
rect 136955 93469 136989 93485
rect 136955 93419 136989 93435
rect 1809 93133 1843 93149
rect 1809 93083 1843 93099
rect 136955 93133 136989 93149
rect 136955 93083 136989 93099
rect 1809 92797 1843 92813
rect 1809 92747 1843 92763
rect 136955 92797 136989 92813
rect 136955 92747 136989 92763
rect 1809 92461 1843 92477
rect 1809 92411 1843 92427
rect 136955 92461 136989 92477
rect 136955 92411 136989 92427
rect 1809 92125 1843 92141
rect 1809 92075 1843 92091
rect 136955 92125 136989 92141
rect 136955 92075 136989 92091
rect 1809 91789 1843 91805
rect 1809 91739 1843 91755
rect 136955 91789 136989 91805
rect 136955 91739 136989 91755
rect 1809 91453 1843 91469
rect 1809 91403 1843 91419
rect 136955 91453 136989 91469
rect 136955 91403 136989 91419
rect 1809 91117 1843 91133
rect 1809 91067 1843 91083
rect 136955 91117 136989 91133
rect 136955 91067 136989 91083
rect 1809 90781 1843 90797
rect 1809 90731 1843 90747
rect 136955 90781 136989 90797
rect 136955 90731 136989 90747
rect 1809 90445 1843 90461
rect 1809 90395 1843 90411
rect 136955 90445 136989 90461
rect 136955 90395 136989 90411
rect 1809 90109 1843 90125
rect 1809 90059 1843 90075
rect 136955 90109 136989 90125
rect 136955 90059 136989 90075
rect 1809 89773 1843 89789
rect 1809 89723 1843 89739
rect 136955 89773 136989 89789
rect 136955 89723 136989 89739
rect 1809 89437 1843 89453
rect 1809 89387 1843 89403
rect 136955 89437 136989 89453
rect 136955 89387 136989 89403
rect 1809 89101 1843 89117
rect 1809 89051 1843 89067
rect 136955 89101 136989 89117
rect 136955 89051 136989 89067
rect 1809 88765 1843 88781
rect 1809 88715 1843 88731
rect 136955 88765 136989 88781
rect 136955 88715 136989 88731
rect 1809 88429 1843 88445
rect 1809 88379 1843 88395
rect 136955 88429 136989 88445
rect 136955 88379 136989 88395
rect 1809 88093 1843 88109
rect 1809 88043 1843 88059
rect 136955 88093 136989 88109
rect 136955 88043 136989 88059
rect 1809 87757 1843 87773
rect 1809 87707 1843 87723
rect 136955 87757 136989 87773
rect 136955 87707 136989 87723
rect 1809 87421 1843 87437
rect 1809 87371 1843 87387
rect 136955 87421 136989 87437
rect 136955 87371 136989 87387
rect 1809 87085 1843 87101
rect 1809 87035 1843 87051
rect 136955 87085 136989 87101
rect 136955 87035 136989 87051
rect 1809 86749 1843 86765
rect 1809 86699 1843 86715
rect 136955 86749 136989 86765
rect 136955 86699 136989 86715
rect 1809 86413 1843 86429
rect 1809 86363 1843 86379
rect 136955 86413 136989 86429
rect 136955 86363 136989 86379
rect 1809 86077 1843 86093
rect 1809 86027 1843 86043
rect 136955 86077 136989 86093
rect 136955 86027 136989 86043
rect 1809 85741 1843 85757
rect 1809 85691 1843 85707
rect 136955 85741 136989 85757
rect 136955 85691 136989 85707
rect 1809 85405 1843 85421
rect 1809 85355 1843 85371
rect 136955 85405 136989 85421
rect 136955 85355 136989 85371
rect 1809 85069 1843 85085
rect 1809 85019 1843 85035
rect 136955 85069 136989 85085
rect 136955 85019 136989 85035
rect 1809 84733 1843 84749
rect 1809 84683 1843 84699
rect 136955 84733 136989 84749
rect 136955 84683 136989 84699
rect 1809 84397 1843 84413
rect 1809 84347 1843 84363
rect 136955 84397 136989 84413
rect 136955 84347 136989 84363
rect 1809 84061 1843 84077
rect 1809 84011 1843 84027
rect 136955 84061 136989 84077
rect 136955 84011 136989 84027
rect 1809 83725 1843 83741
rect 1809 83675 1843 83691
rect 136955 83725 136989 83741
rect 136955 83675 136989 83691
rect 1809 83389 1843 83405
rect 1809 83339 1843 83355
rect 136955 83389 136989 83405
rect 136955 83339 136989 83355
rect 1809 83053 1843 83069
rect 1809 83003 1843 83019
rect 136955 83053 136989 83069
rect 136955 83003 136989 83019
rect 1809 82717 1843 82733
rect 1809 82667 1843 82683
rect 136955 82717 136989 82733
rect 136955 82667 136989 82683
rect 1809 82381 1843 82397
rect 1809 82331 1843 82347
rect 136955 82381 136989 82397
rect 136955 82331 136989 82347
rect 1809 82045 1843 82061
rect 1809 81995 1843 82011
rect 136955 82045 136989 82061
rect 136955 81995 136989 82011
rect 1809 81709 1843 81725
rect 1809 81659 1843 81675
rect 136955 81709 136989 81725
rect 136955 81659 136989 81675
rect 1809 81373 1843 81389
rect 1809 81323 1843 81339
rect 136955 81373 136989 81389
rect 136955 81323 136989 81339
rect 1809 81037 1843 81053
rect 1809 80987 1843 81003
rect 136955 81037 136989 81053
rect 136955 80987 136989 81003
rect 1809 80701 1843 80717
rect 1809 80651 1843 80667
rect 136955 80701 136989 80717
rect 136955 80651 136989 80667
rect 1809 80365 1843 80381
rect 1809 80315 1843 80331
rect 136955 80365 136989 80381
rect 136955 80315 136989 80331
rect 1809 80029 1843 80045
rect 1809 79979 1843 79995
rect 136955 80029 136989 80045
rect 136955 79979 136989 79995
rect 1809 79693 1843 79709
rect 1809 79643 1843 79659
rect 136955 79693 136989 79709
rect 136955 79643 136989 79659
rect 1809 79357 1843 79373
rect 1809 79307 1843 79323
rect 136955 79357 136989 79373
rect 136955 79307 136989 79323
rect 1809 79021 1843 79037
rect 1809 78971 1843 78987
rect 136955 79021 136989 79037
rect 136955 78971 136989 78987
rect 1809 78685 1843 78701
rect 1809 78635 1843 78651
rect 136955 78685 136989 78701
rect 136955 78635 136989 78651
rect 1809 78349 1843 78365
rect 1809 78299 1843 78315
rect 136955 78349 136989 78365
rect 136955 78299 136989 78315
rect 1809 78013 1843 78029
rect 1809 77963 1843 77979
rect 136955 78013 136989 78029
rect 136955 77963 136989 77979
rect 1809 77677 1843 77693
rect 1809 77627 1843 77643
rect 136955 77677 136989 77693
rect 136955 77627 136989 77643
rect 1809 77341 1843 77357
rect 1809 77291 1843 77307
rect 136955 77341 136989 77357
rect 136955 77291 136989 77307
rect 1809 77005 1843 77021
rect 1809 76955 1843 76971
rect 136955 77005 136989 77021
rect 136955 76955 136989 76971
rect 1809 76669 1843 76685
rect 1809 76619 1843 76635
rect 136955 76669 136989 76685
rect 136955 76619 136989 76635
rect 1809 76333 1843 76349
rect 1809 76283 1843 76299
rect 136955 76333 136989 76349
rect 136955 76283 136989 76299
rect 1809 75997 1843 76013
rect 1809 75947 1843 75963
rect 136955 75997 136989 76013
rect 136955 75947 136989 75963
rect 1809 75661 1843 75677
rect 1809 75611 1843 75627
rect 136955 75661 136989 75677
rect 136955 75611 136989 75627
rect 1809 75325 1843 75341
rect 1809 75275 1843 75291
rect 136955 75325 136989 75341
rect 136955 75275 136989 75291
rect 1809 74989 1843 75005
rect 1809 74939 1843 74955
rect 136955 74989 136989 75005
rect 136955 74939 136989 74955
rect 1809 74653 1843 74669
rect 1809 74603 1843 74619
rect 136955 74653 136989 74669
rect 136955 74603 136989 74619
rect 1809 74317 1843 74333
rect 1809 74267 1843 74283
rect 136955 74317 136989 74333
rect 136955 74267 136989 74283
rect 1809 73981 1843 73997
rect 1809 73931 1843 73947
rect 136955 73981 136989 73997
rect 136955 73931 136989 73947
rect 1809 73645 1843 73661
rect 1809 73595 1843 73611
rect 136955 73645 136989 73661
rect 136955 73595 136989 73611
rect 1809 73309 1843 73325
rect 1809 73259 1843 73275
rect 136955 73309 136989 73325
rect 136955 73259 136989 73275
rect 1809 72973 1843 72989
rect 1809 72923 1843 72939
rect 136955 72973 136989 72989
rect 136955 72923 136989 72939
rect 1809 72637 1843 72653
rect 1809 72587 1843 72603
rect 136955 72637 136989 72653
rect 136955 72587 136989 72603
rect 1809 72301 1843 72317
rect 1809 72251 1843 72267
rect 136955 72301 136989 72317
rect 136955 72251 136989 72267
rect 1809 71965 1843 71981
rect 1809 71915 1843 71931
rect 136955 71965 136989 71981
rect 136955 71915 136989 71931
rect 1809 71629 1843 71645
rect 1809 71579 1843 71595
rect 136955 71629 136989 71645
rect 136955 71579 136989 71595
rect 1809 71293 1843 71309
rect 1809 71243 1843 71259
rect 136955 71293 136989 71309
rect 136955 71243 136989 71259
rect 1809 70957 1843 70973
rect 1809 70907 1843 70923
rect 136955 70957 136989 70973
rect 136955 70907 136989 70923
rect 1809 70621 1843 70637
rect 1809 70571 1843 70587
rect 136955 70621 136989 70637
rect 136955 70571 136989 70587
rect 1809 70285 1843 70301
rect 1809 70235 1843 70251
rect 136955 70285 136989 70301
rect 136955 70235 136989 70251
rect 1809 69949 1843 69965
rect 1809 69899 1843 69915
rect 136955 69949 136989 69965
rect 136955 69899 136989 69915
rect 1809 69613 1843 69629
rect 1809 69563 1843 69579
rect 136955 69613 136989 69629
rect 136955 69563 136989 69579
rect 1809 69277 1843 69293
rect 1809 69227 1843 69243
rect 136955 69277 136989 69293
rect 136955 69227 136989 69243
rect 1809 68941 1843 68957
rect 1809 68891 1843 68907
rect 136955 68941 136989 68957
rect 136955 68891 136989 68907
rect 1809 68605 1843 68621
rect 1809 68555 1843 68571
rect 136955 68605 136989 68621
rect 136955 68555 136989 68571
rect 1809 68269 1843 68285
rect 1809 68219 1843 68235
rect 136955 68269 136989 68285
rect 136955 68219 136989 68235
rect 1809 67933 1843 67949
rect 1809 67883 1843 67899
rect 136955 67933 136989 67949
rect 136955 67883 136989 67899
rect 1809 67597 1843 67613
rect 1809 67547 1843 67563
rect 136955 67597 136989 67613
rect 136955 67547 136989 67563
rect 1809 67261 1843 67277
rect 1809 67211 1843 67227
rect 136955 67261 136989 67277
rect 136955 67211 136989 67227
rect 1809 66925 1843 66941
rect 1809 66875 1843 66891
rect 136955 66925 136989 66941
rect 136955 66875 136989 66891
rect 1809 66589 1843 66605
rect 1809 66539 1843 66555
rect 136955 66589 136989 66605
rect 136955 66539 136989 66555
rect 1809 66253 1843 66269
rect 1809 66203 1843 66219
rect 136955 66253 136989 66269
rect 136955 66203 136989 66219
rect 1809 65917 1843 65933
rect 1809 65867 1843 65883
rect 136955 65917 136989 65933
rect 136955 65867 136989 65883
rect 1809 65581 1843 65597
rect 1809 65531 1843 65547
rect 136955 65581 136989 65597
rect 136955 65531 136989 65547
rect 1809 65245 1843 65261
rect 1809 65195 1843 65211
rect 136955 65245 136989 65261
rect 136955 65195 136989 65211
rect 1809 64909 1843 64925
rect 1809 64859 1843 64875
rect 136955 64909 136989 64925
rect 136955 64859 136989 64875
rect 1809 64573 1843 64589
rect 1809 64523 1843 64539
rect 136955 64573 136989 64589
rect 136955 64523 136989 64539
rect 1809 64237 1843 64253
rect 1809 64187 1843 64203
rect 136955 64237 136989 64253
rect 136955 64187 136989 64203
rect 1809 63901 1843 63917
rect 1809 63851 1843 63867
rect 136955 63901 136989 63917
rect 136955 63851 136989 63867
rect 1809 63565 1843 63581
rect 1809 63515 1843 63531
rect 136955 63565 136989 63581
rect 136955 63515 136989 63531
rect 1809 63229 1843 63245
rect 1809 63179 1843 63195
rect 136955 63229 136989 63245
rect 136955 63179 136989 63195
rect 1809 62893 1843 62909
rect 1809 62843 1843 62859
rect 136955 62893 136989 62909
rect 136955 62843 136989 62859
rect 1809 62557 1843 62573
rect 1809 62507 1843 62523
rect 136955 62557 136989 62573
rect 136955 62507 136989 62523
rect 1809 62221 1843 62237
rect 1809 62171 1843 62187
rect 136955 62221 136989 62237
rect 136955 62171 136989 62187
rect 1809 61885 1843 61901
rect 1809 61835 1843 61851
rect 136955 61885 136989 61901
rect 136955 61835 136989 61851
rect 1809 61549 1843 61565
rect 1809 61499 1843 61515
rect 136955 61549 136989 61565
rect 136955 61499 136989 61515
rect 1809 61213 1843 61229
rect 1809 61163 1843 61179
rect 136955 61213 136989 61229
rect 136955 61163 136989 61179
rect 1809 60877 1843 60893
rect 1809 60827 1843 60843
rect 136955 60877 136989 60893
rect 136955 60827 136989 60843
rect 1809 60541 1843 60557
rect 1809 60491 1843 60507
rect 136955 60541 136989 60557
rect 136955 60491 136989 60507
rect 1809 60205 1843 60221
rect 1809 60155 1843 60171
rect 136955 60205 136989 60221
rect 136955 60155 136989 60171
rect 1809 59869 1843 59885
rect 1809 59819 1843 59835
rect 136955 59869 136989 59885
rect 136955 59819 136989 59835
rect 1809 59533 1843 59549
rect 1809 59483 1843 59499
rect 136955 59533 136989 59549
rect 136955 59483 136989 59499
rect 1809 59197 1843 59213
rect 1809 59147 1843 59163
rect 136955 59197 136989 59213
rect 136955 59147 136989 59163
rect 1809 58861 1843 58877
rect 1809 58811 1843 58827
rect 136955 58861 136989 58877
rect 136955 58811 136989 58827
rect 1809 58525 1843 58541
rect 1809 58475 1843 58491
rect 136955 58525 136989 58541
rect 136955 58475 136989 58491
rect 1809 58189 1843 58205
rect 1809 58139 1843 58155
rect 136955 58189 136989 58205
rect 136955 58139 136989 58155
rect 1809 57853 1843 57869
rect 1809 57803 1843 57819
rect 136955 57853 136989 57869
rect 136955 57803 136989 57819
rect 1809 57517 1843 57533
rect 1809 57467 1843 57483
rect 136955 57517 136989 57533
rect 136955 57467 136989 57483
rect 1809 57181 1843 57197
rect 1809 57131 1843 57147
rect 136955 57181 136989 57197
rect 136955 57131 136989 57147
rect 1809 56845 1843 56861
rect 1809 56795 1843 56811
rect 136955 56845 136989 56861
rect 136955 56795 136989 56811
rect 1809 56509 1843 56525
rect 1809 56459 1843 56475
rect 136955 56509 136989 56525
rect 136955 56459 136989 56475
rect 1809 56173 1843 56189
rect 1809 56123 1843 56139
rect 136955 56173 136989 56189
rect 136955 56123 136989 56139
rect 1809 55837 1843 55853
rect 1809 55787 1843 55803
rect 136955 55837 136989 55853
rect 136955 55787 136989 55803
rect 1809 55501 1843 55517
rect 1809 55451 1843 55467
rect 136955 55501 136989 55517
rect 136955 55451 136989 55467
rect 1809 55165 1843 55181
rect 1809 55115 1843 55131
rect 136955 55165 136989 55181
rect 136955 55115 136989 55131
rect 1809 54829 1843 54845
rect 1809 54779 1843 54795
rect 136955 54829 136989 54845
rect 136955 54779 136989 54795
rect 1809 54493 1843 54509
rect 1809 54443 1843 54459
rect 136955 54493 136989 54509
rect 136955 54443 136989 54459
rect 1809 54157 1843 54173
rect 1809 54107 1843 54123
rect 136955 54157 136989 54173
rect 136955 54107 136989 54123
rect 1809 53821 1843 53837
rect 1809 53771 1843 53787
rect 136955 53821 136989 53837
rect 136955 53771 136989 53787
rect 1809 53485 1843 53501
rect 1809 53435 1843 53451
rect 136955 53485 136989 53501
rect 136955 53435 136989 53451
rect 1809 53149 1843 53165
rect 1809 53099 1843 53115
rect 136955 53149 136989 53165
rect 136955 53099 136989 53115
rect 1809 52813 1843 52829
rect 1809 52763 1843 52779
rect 136955 52813 136989 52829
rect 136955 52763 136989 52779
rect 1809 52477 1843 52493
rect 1809 52427 1843 52443
rect 136955 52477 136989 52493
rect 136955 52427 136989 52443
rect 1809 52141 1843 52157
rect 1809 52091 1843 52107
rect 136955 52141 136989 52157
rect 136955 52091 136989 52107
rect 1809 51805 1843 51821
rect 1809 51755 1843 51771
rect 136955 51805 136989 51821
rect 136955 51755 136989 51771
rect 1809 51469 1843 51485
rect 1809 51419 1843 51435
rect 136955 51469 136989 51485
rect 136955 51419 136989 51435
rect 1809 51133 1843 51149
rect 1809 51083 1843 51099
rect 136955 51133 136989 51149
rect 136955 51083 136989 51099
rect 1809 50797 1843 50813
rect 1809 50747 1843 50763
rect 136955 50797 136989 50813
rect 136955 50747 136989 50763
rect 1809 50461 1843 50477
rect 1809 50411 1843 50427
rect 136955 50461 136989 50477
rect 136955 50411 136989 50427
rect 1809 50125 1843 50141
rect 1809 50075 1843 50091
rect 136955 50125 136989 50141
rect 136955 50075 136989 50091
rect 1809 49789 1843 49805
rect 1809 49739 1843 49755
rect 136955 49789 136989 49805
rect 136955 49739 136989 49755
rect 1809 49453 1843 49469
rect 1809 49403 1843 49419
rect 136955 49453 136989 49469
rect 136955 49403 136989 49419
rect 1809 49117 1843 49133
rect 1809 49067 1843 49083
rect 136955 49117 136989 49133
rect 136955 49067 136989 49083
rect 1809 48781 1843 48797
rect 1809 48731 1843 48747
rect 136955 48781 136989 48797
rect 136955 48731 136989 48747
rect 1809 48445 1843 48461
rect 1809 48395 1843 48411
rect 136955 48445 136989 48461
rect 136955 48395 136989 48411
rect 1809 48109 1843 48125
rect 1809 48059 1843 48075
rect 136955 48109 136989 48125
rect 136955 48059 136989 48075
rect 1809 47773 1843 47789
rect 1809 47723 1843 47739
rect 136955 47773 136989 47789
rect 136955 47723 136989 47739
rect 1809 47437 1843 47453
rect 1809 47387 1843 47403
rect 136955 47437 136989 47453
rect 136955 47387 136989 47403
rect 1809 47101 1843 47117
rect 1809 47051 1843 47067
rect 136955 47101 136989 47117
rect 136955 47051 136989 47067
rect 1809 46765 1843 46781
rect 1809 46715 1843 46731
rect 136955 46765 136989 46781
rect 136955 46715 136989 46731
rect 1809 46429 1843 46445
rect 1809 46379 1843 46395
rect 136955 46429 136989 46445
rect 136955 46379 136989 46395
rect 1809 46093 1843 46109
rect 1809 46043 1843 46059
rect 136955 46093 136989 46109
rect 136955 46043 136989 46059
rect 1809 45757 1843 45773
rect 1809 45707 1843 45723
rect 136955 45757 136989 45773
rect 136955 45707 136989 45723
rect 1809 45421 1843 45437
rect 1809 45371 1843 45387
rect 136955 45421 136989 45437
rect 136955 45371 136989 45387
rect 1809 45085 1843 45101
rect 1809 45035 1843 45051
rect 136955 45085 136989 45101
rect 136955 45035 136989 45051
rect 1809 44749 1843 44765
rect 1809 44699 1843 44715
rect 136955 44749 136989 44765
rect 136955 44699 136989 44715
rect 1809 44413 1843 44429
rect 1809 44363 1843 44379
rect 136955 44413 136989 44429
rect 136955 44363 136989 44379
rect 1809 44077 1843 44093
rect 1809 44027 1843 44043
rect 136955 44077 136989 44093
rect 136955 44027 136989 44043
rect 1809 43741 1843 43757
rect 1809 43691 1843 43707
rect 136955 43741 136989 43757
rect 136955 43691 136989 43707
rect 1809 43405 1843 43421
rect 1809 43355 1843 43371
rect 136955 43405 136989 43421
rect 136955 43355 136989 43371
rect 1809 43069 1843 43085
rect 1809 43019 1843 43035
rect 136955 43069 136989 43085
rect 136955 43019 136989 43035
rect 1809 42733 1843 42749
rect 1809 42683 1843 42699
rect 136955 42733 136989 42749
rect 136955 42683 136989 42699
rect 1809 42397 1843 42413
rect 1809 42347 1843 42363
rect 136955 42397 136989 42413
rect 136955 42347 136989 42363
rect 1809 42061 1843 42077
rect 1809 42011 1843 42027
rect 136955 42061 136989 42077
rect 136955 42011 136989 42027
rect 1809 41725 1843 41741
rect 1809 41675 1843 41691
rect 136955 41725 136989 41741
rect 136955 41675 136989 41691
rect 1809 41389 1843 41405
rect 1809 41339 1843 41355
rect 136955 41389 136989 41405
rect 136955 41339 136989 41355
rect 1809 41053 1843 41069
rect 1809 41003 1843 41019
rect 136955 41053 136989 41069
rect 136955 41003 136989 41019
rect 1809 40717 1843 40733
rect 1809 40667 1843 40683
rect 136955 40717 136989 40733
rect 136955 40667 136989 40683
rect 1809 40381 1843 40397
rect 1809 40331 1843 40347
rect 136955 40381 136989 40397
rect 136955 40331 136989 40347
rect 1809 40045 1843 40061
rect 1809 39995 1843 40011
rect 136955 40045 136989 40061
rect 136955 39995 136989 40011
rect 1809 39709 1843 39725
rect 1809 39659 1843 39675
rect 136955 39709 136989 39725
rect 136955 39659 136989 39675
rect 1809 39373 1843 39389
rect 1809 39323 1843 39339
rect 136955 39373 136989 39389
rect 136955 39323 136989 39339
rect 1809 39037 1843 39053
rect 1809 38987 1843 39003
rect 136955 39037 136989 39053
rect 136955 38987 136989 39003
rect 1809 38701 1843 38717
rect 1809 38651 1843 38667
rect 136955 38701 136989 38717
rect 136955 38651 136989 38667
rect 1809 38365 1843 38381
rect 1809 38315 1843 38331
rect 136955 38365 136989 38381
rect 136955 38315 136989 38331
rect 1809 38029 1843 38045
rect 1809 37979 1843 37995
rect 136955 38029 136989 38045
rect 136955 37979 136989 37995
rect 1809 37693 1843 37709
rect 1809 37643 1843 37659
rect 136955 37693 136989 37709
rect 136955 37643 136989 37659
rect 1809 37357 1843 37373
rect 1809 37307 1843 37323
rect 136955 37357 136989 37373
rect 136955 37307 136989 37323
rect 1809 37021 1843 37037
rect 1809 36971 1843 36987
rect 136955 37021 136989 37037
rect 136955 36971 136989 36987
rect 1809 36685 1843 36701
rect 1809 36635 1843 36651
rect 136955 36685 136989 36701
rect 136955 36635 136989 36651
rect 1809 36349 1843 36365
rect 1809 36299 1843 36315
rect 136955 36349 136989 36365
rect 136955 36299 136989 36315
rect 1809 36013 1843 36029
rect 1809 35963 1843 35979
rect 136955 36013 136989 36029
rect 136955 35963 136989 35979
rect 1809 35677 1843 35693
rect 1809 35627 1843 35643
rect 136955 35677 136989 35693
rect 136955 35627 136989 35643
rect 1809 35341 1843 35357
rect 1809 35291 1843 35307
rect 136955 35341 136989 35357
rect 136955 35291 136989 35307
rect 1809 35005 1843 35021
rect 1809 34955 1843 34971
rect 136955 35005 136989 35021
rect 136955 34955 136989 34971
rect 1809 34669 1843 34685
rect 1809 34619 1843 34635
rect 136955 34669 136989 34685
rect 136955 34619 136989 34635
rect 1809 34333 1843 34349
rect 1809 34283 1843 34299
rect 136955 34333 136989 34349
rect 136955 34283 136989 34299
rect 1809 33997 1843 34013
rect 1809 33947 1843 33963
rect 136955 33997 136989 34013
rect 136955 33947 136989 33963
rect 1809 33661 1843 33677
rect 1809 33611 1843 33627
rect 136955 33661 136989 33677
rect 136955 33611 136989 33627
rect 1809 33325 1843 33341
rect 1809 33275 1843 33291
rect 136955 33325 136989 33341
rect 136955 33275 136989 33291
rect 1809 32989 1843 33005
rect 1809 32939 1843 32955
rect 136955 32989 136989 33005
rect 136955 32939 136989 32955
rect 1809 32653 1843 32669
rect 1809 32603 1843 32619
rect 136955 32653 136989 32669
rect 136955 32603 136989 32619
rect 1809 32317 1843 32333
rect 1809 32267 1843 32283
rect 136955 32317 136989 32333
rect 136955 32267 136989 32283
rect 1809 31981 1843 31997
rect 1809 31931 1843 31947
rect 136955 31981 136989 31997
rect 136955 31931 136989 31947
rect 1809 31645 1843 31661
rect 1809 31595 1843 31611
rect 136955 31645 136989 31661
rect 136955 31595 136989 31611
rect 1809 31309 1843 31325
rect 1809 31259 1843 31275
rect 136955 31309 136989 31325
rect 136955 31259 136989 31275
rect 1809 30973 1843 30989
rect 1809 30923 1843 30939
rect 136955 30973 136989 30989
rect 136955 30923 136989 30939
rect 1809 30637 1843 30653
rect 1809 30587 1843 30603
rect 136955 30637 136989 30653
rect 136955 30587 136989 30603
rect 1809 30301 1843 30317
rect 1809 30251 1843 30267
rect 136955 30301 136989 30317
rect 136955 30251 136989 30267
rect 1809 29965 1843 29981
rect 1809 29915 1843 29931
rect 136955 29965 136989 29981
rect 136955 29915 136989 29931
rect 1809 29629 1843 29645
rect 1809 29579 1843 29595
rect 136955 29629 136989 29645
rect 136955 29579 136989 29595
rect 1809 29293 1843 29309
rect 1809 29243 1843 29259
rect 136955 29293 136989 29309
rect 136955 29243 136989 29259
rect 1809 28957 1843 28973
rect 1809 28907 1843 28923
rect 136955 28957 136989 28973
rect 136955 28907 136989 28923
rect 1809 28621 1843 28637
rect 1809 28571 1843 28587
rect 136955 28621 136989 28637
rect 136955 28571 136989 28587
rect 1809 28285 1843 28301
rect 1809 28235 1843 28251
rect 136955 28285 136989 28301
rect 136955 28235 136989 28251
rect 1809 27949 1843 27965
rect 1809 27899 1843 27915
rect 136955 27949 136989 27965
rect 136955 27899 136989 27915
rect 1809 27613 1843 27629
rect 1809 27563 1843 27579
rect 136955 27613 136989 27629
rect 136955 27563 136989 27579
rect 1809 27277 1843 27293
rect 1809 27227 1843 27243
rect 136955 27277 136989 27293
rect 136955 27227 136989 27243
rect 1809 26941 1843 26957
rect 1809 26891 1843 26907
rect 136955 26941 136989 26957
rect 136955 26891 136989 26907
rect 1809 26605 1843 26621
rect 1809 26555 1843 26571
rect 136955 26605 136989 26621
rect 136955 26555 136989 26571
rect 1809 26269 1843 26285
rect 1809 26219 1843 26235
rect 136955 26269 136989 26285
rect 136955 26219 136989 26235
rect 1809 25933 1843 25949
rect 1809 25883 1843 25899
rect 136955 25933 136989 25949
rect 136955 25883 136989 25899
rect 1809 25597 1843 25613
rect 1809 25547 1843 25563
rect 136955 25597 136989 25613
rect 136955 25547 136989 25563
rect 1809 25261 1843 25277
rect 1809 25211 1843 25227
rect 136955 25261 136989 25277
rect 136955 25211 136989 25227
rect 1809 24925 1843 24941
rect 1809 24875 1843 24891
rect 136955 24925 136989 24941
rect 136955 24875 136989 24891
rect 1809 24589 1843 24605
rect 1809 24539 1843 24555
rect 136955 24589 136989 24605
rect 136955 24539 136989 24555
rect 1809 24253 1843 24269
rect 1809 24203 1843 24219
rect 136955 24253 136989 24269
rect 136955 24203 136989 24219
rect 1809 23917 1843 23933
rect 1809 23867 1843 23883
rect 136955 23917 136989 23933
rect 136955 23867 136989 23883
rect 1809 23581 1843 23597
rect 1809 23531 1843 23547
rect 136955 23581 136989 23597
rect 136955 23531 136989 23547
rect 1809 23245 1843 23261
rect 1809 23195 1843 23211
rect 136955 23245 136989 23261
rect 136955 23195 136989 23211
rect 1809 22909 1843 22925
rect 1809 22859 1843 22875
rect 136955 22909 136989 22925
rect 136955 22859 136989 22875
rect 1809 22573 1843 22589
rect 1809 22523 1843 22539
rect 136955 22573 136989 22589
rect 136955 22523 136989 22539
rect 1809 22237 1843 22253
rect 1809 22187 1843 22203
rect 136955 22237 136989 22253
rect 136955 22187 136989 22203
rect 1809 21901 1843 21917
rect 1809 21851 1843 21867
rect 136955 21901 136989 21917
rect 136955 21851 136989 21867
rect 1809 21565 1843 21581
rect 1809 21515 1843 21531
rect 136955 21565 136989 21581
rect 136955 21515 136989 21531
rect 1809 21229 1843 21245
rect 1809 21179 1843 21195
rect 136955 21229 136989 21245
rect 136955 21179 136989 21195
rect 1809 20893 1843 20909
rect 1809 20843 1843 20859
rect 136955 20893 136989 20909
rect 136955 20843 136989 20859
rect 1809 20557 1843 20573
rect 1809 20507 1843 20523
rect 136955 20557 136989 20573
rect 136955 20507 136989 20523
rect 1809 20221 1843 20237
rect 1809 20171 1843 20187
rect 136955 20221 136989 20237
rect 136955 20171 136989 20187
rect 1809 19885 1843 19901
rect 1809 19835 1843 19851
rect 136955 19885 136989 19901
rect 136955 19835 136989 19851
rect 1809 19549 1843 19565
rect 1809 19499 1843 19515
rect 136955 19549 136989 19565
rect 136955 19499 136989 19515
rect 1809 19213 1843 19229
rect 1809 19163 1843 19179
rect 136955 19213 136989 19229
rect 136955 19163 136989 19179
rect 1809 18877 1843 18893
rect 1809 18827 1843 18843
rect 136955 18877 136989 18893
rect 136955 18827 136989 18843
rect 1809 18541 1843 18557
rect 1809 18491 1843 18507
rect 136955 18541 136989 18557
rect 136955 18491 136989 18507
rect 1809 18205 1843 18221
rect 1809 18155 1843 18171
rect 136955 18205 136989 18221
rect 136955 18155 136989 18171
rect 1809 17869 1843 17885
rect 1809 17819 1843 17835
rect 136955 17869 136989 17885
rect 136955 17819 136989 17835
rect 1809 17533 1843 17549
rect 1809 17483 1843 17499
rect 136955 17533 136989 17549
rect 136955 17483 136989 17499
rect 1809 17197 1843 17213
rect 1809 17147 1843 17163
rect 136955 17197 136989 17213
rect 136955 17147 136989 17163
rect 1809 16861 1843 16877
rect 1809 16811 1843 16827
rect 136955 16861 136989 16877
rect 136955 16811 136989 16827
rect 1809 16525 1843 16541
rect 1809 16475 1843 16491
rect 136955 16525 136989 16541
rect 136955 16475 136989 16491
rect 1809 16189 1843 16205
rect 1809 16139 1843 16155
rect 136955 16189 136989 16205
rect 136955 16139 136989 16155
rect 1809 15853 1843 15869
rect 1809 15803 1843 15819
rect 136955 15853 136989 15869
rect 136955 15803 136989 15819
rect 1809 15517 1843 15533
rect 1809 15467 1843 15483
rect 136955 15517 136989 15533
rect 136955 15467 136989 15483
rect 1809 15181 1843 15197
rect 1809 15131 1843 15147
rect 136955 15181 136989 15197
rect 136955 15131 136989 15147
rect 1809 14845 1843 14861
rect 1809 14795 1843 14811
rect 136955 14845 136989 14861
rect 136955 14795 136989 14811
rect 1809 14509 1843 14525
rect 1809 14459 1843 14475
rect 136955 14509 136989 14525
rect 136955 14459 136989 14475
rect 1809 14173 1843 14189
rect 1809 14123 1843 14139
rect 136955 14173 136989 14189
rect 136955 14123 136989 14139
rect 1809 13837 1843 13853
rect 1809 13787 1843 13803
rect 136955 13837 136989 13853
rect 136955 13787 136989 13803
rect 1809 13501 1843 13517
rect 1809 13451 1843 13467
rect 136955 13501 136989 13517
rect 136955 13451 136989 13467
rect 1809 13165 1843 13181
rect 1809 13115 1843 13131
rect 136955 13165 136989 13181
rect 136955 13115 136989 13131
rect 1809 12829 1843 12845
rect 1809 12779 1843 12795
rect 136955 12829 136989 12845
rect 136955 12779 136989 12795
rect 1809 12493 1843 12509
rect 1809 12443 1843 12459
rect 136955 12493 136989 12509
rect 136955 12443 136989 12459
rect 1809 12157 1843 12173
rect 1809 12107 1843 12123
rect 136955 12157 136989 12173
rect 136955 12107 136989 12123
rect 1809 11821 1843 11837
rect 1809 11771 1843 11787
rect 136955 11821 136989 11837
rect 136955 11771 136989 11787
rect 1809 11485 1843 11501
rect 1809 11435 1843 11451
rect 136955 11485 136989 11501
rect 136955 11435 136989 11451
rect 1809 11149 1843 11165
rect 1809 11099 1843 11115
rect 136955 11149 136989 11165
rect 136955 11099 136989 11115
rect 1809 10813 1843 10829
rect 1809 10763 1843 10779
rect 136955 10813 136989 10829
rect 136955 10763 136989 10779
rect 1809 10477 1843 10493
rect 1809 10427 1843 10443
rect 136955 10477 136989 10493
rect 136955 10427 136989 10443
rect 1809 10141 1843 10157
rect 1809 10091 1843 10107
rect 136955 10141 136989 10157
rect 136955 10091 136989 10107
rect 1809 9805 1843 9821
rect 1809 9755 1843 9771
rect 136955 9805 136989 9821
rect 136955 9755 136989 9771
rect 1809 9469 1843 9485
rect 1809 9419 1843 9435
rect 136955 9469 136989 9485
rect 136955 9419 136989 9435
rect 1809 9133 1843 9149
rect 1809 9083 1843 9099
rect 136955 9133 136989 9149
rect 136955 9083 136989 9099
rect 1809 8797 1843 8813
rect 1809 8747 1843 8763
rect 136955 8797 136989 8813
rect 136955 8747 136989 8763
rect 1809 8461 1843 8477
rect 1809 8411 1843 8427
rect 136955 8461 136989 8477
rect 136955 8411 136989 8427
rect 1809 8125 1843 8141
rect 1809 8075 1843 8091
rect 136955 8125 136989 8141
rect 136955 8075 136989 8091
rect 1809 7789 1843 7805
rect 1809 7739 1843 7755
rect 136955 7789 136989 7805
rect 136955 7739 136989 7755
rect 1809 7453 1843 7469
rect 1809 7403 1843 7419
rect 136955 7453 136989 7469
rect 136955 7403 136989 7419
rect 1809 7117 1843 7133
rect 1809 7067 1843 7083
rect 136955 7117 136989 7133
rect 136955 7067 136989 7083
rect 1809 6781 1843 6797
rect 1809 6731 1843 6747
rect 136955 6781 136989 6797
rect 136955 6731 136989 6747
rect 1809 6445 1843 6461
rect 1809 6395 1843 6411
rect 136955 6445 136989 6461
rect 136955 6395 136989 6411
rect 1809 6109 1843 6125
rect 1809 6059 1843 6075
rect 136955 6109 136989 6125
rect 136955 6059 136989 6075
rect 1809 5773 1843 5789
rect 1809 5723 1843 5739
rect 136955 5773 136989 5789
rect 136955 5723 136989 5739
rect 1809 5437 1843 5453
rect 1809 5387 1843 5403
rect 136955 5437 136989 5453
rect 136955 5387 136989 5403
rect 1809 5101 1843 5117
rect 1809 5051 1843 5067
rect 136955 5101 136989 5117
rect 136955 5051 136989 5067
rect 1809 4765 1843 4781
rect 1809 4715 1843 4731
rect 136955 4765 136989 4781
rect 136955 4715 136989 4731
rect 1809 4429 1843 4445
rect 1809 4379 1843 4395
rect 136955 4429 136989 4445
rect 136955 4379 136989 4395
rect 1809 4093 1843 4109
rect 1809 4043 1843 4059
rect 136955 4093 136989 4109
rect 136955 4043 136989 4059
rect 1809 3757 1843 3773
rect 1809 3707 1843 3723
rect 136955 3757 136989 3773
rect 136955 3707 136989 3723
rect 1809 3421 1843 3437
rect 1809 3371 1843 3387
rect 136955 3421 136989 3437
rect 136955 3371 136989 3387
rect 1809 3085 1843 3101
rect 1809 3035 1843 3051
rect 136955 3085 136989 3101
rect 136955 3035 136989 3051
rect 1809 2749 1843 2765
rect 1809 2699 1843 2715
rect 136955 2749 136989 2765
rect 136955 2699 136989 2715
rect 1809 2413 1843 2429
rect 1809 2363 1843 2379
rect 136955 2413 136989 2429
rect 136955 2363 136989 2379
rect 1809 2077 1843 2093
rect 1809 2027 1843 2043
rect 136955 2077 136989 2093
rect 136955 2027 136989 2043
rect 2145 1741 2179 1757
rect 2145 1691 2179 1707
rect 2481 1741 2515 1757
rect 2481 1691 2515 1707
rect 2817 1741 2851 1757
rect 2817 1691 2851 1707
rect 3153 1741 3187 1757
rect 3153 1691 3187 1707
rect 3489 1741 3523 1757
rect 3489 1691 3523 1707
rect 3825 1741 3859 1757
rect 3825 1691 3859 1707
rect 4161 1741 4195 1757
rect 4161 1691 4195 1707
rect 4497 1741 4531 1757
rect 4497 1691 4531 1707
rect 4833 1741 4867 1757
rect 4833 1691 4867 1707
rect 5169 1741 5203 1757
rect 5169 1691 5203 1707
rect 5505 1741 5539 1757
rect 5505 1691 5539 1707
rect 5841 1741 5875 1757
rect 5841 1691 5875 1707
rect 6177 1741 6211 1757
rect 6177 1691 6211 1707
rect 6513 1741 6547 1757
rect 6513 1691 6547 1707
rect 6849 1741 6883 1757
rect 6849 1691 6883 1707
rect 7185 1741 7219 1757
rect 7185 1691 7219 1707
rect 7521 1741 7555 1757
rect 7521 1691 7555 1707
rect 7857 1741 7891 1757
rect 7857 1691 7891 1707
rect 8193 1741 8227 1757
rect 8193 1691 8227 1707
rect 8529 1741 8563 1757
rect 8529 1691 8563 1707
rect 8865 1741 8899 1757
rect 8865 1691 8899 1707
rect 9201 1741 9235 1757
rect 9201 1691 9235 1707
rect 9537 1741 9571 1757
rect 9537 1691 9571 1707
rect 9873 1741 9907 1757
rect 9873 1691 9907 1707
rect 10209 1741 10243 1757
rect 10209 1691 10243 1707
rect 10545 1741 10579 1757
rect 10545 1691 10579 1707
rect 10881 1741 10915 1757
rect 10881 1691 10915 1707
rect 11217 1741 11251 1757
rect 11217 1691 11251 1707
rect 11553 1741 11587 1757
rect 11553 1691 11587 1707
rect 11889 1741 11923 1757
rect 11889 1691 11923 1707
rect 12225 1741 12259 1757
rect 12225 1691 12259 1707
rect 12561 1741 12595 1757
rect 12561 1691 12595 1707
rect 12897 1741 12931 1757
rect 12897 1691 12931 1707
rect 13233 1741 13267 1757
rect 13233 1691 13267 1707
rect 13569 1741 13603 1757
rect 13569 1691 13603 1707
rect 13905 1741 13939 1757
rect 13905 1691 13939 1707
rect 14241 1741 14275 1757
rect 14241 1691 14275 1707
rect 14577 1741 14611 1757
rect 14577 1691 14611 1707
rect 14913 1741 14947 1757
rect 14913 1691 14947 1707
rect 15249 1741 15283 1757
rect 15249 1691 15283 1707
rect 15585 1741 15619 1757
rect 15585 1691 15619 1707
rect 15921 1741 15955 1757
rect 15921 1691 15955 1707
rect 16257 1741 16291 1757
rect 16257 1691 16291 1707
rect 16593 1741 16627 1757
rect 16593 1691 16627 1707
rect 16929 1741 16963 1757
rect 16929 1691 16963 1707
rect 17265 1741 17299 1757
rect 17265 1691 17299 1707
rect 17601 1741 17635 1757
rect 17601 1691 17635 1707
rect 17937 1741 17971 1757
rect 17937 1691 17971 1707
rect 18273 1741 18307 1757
rect 18273 1691 18307 1707
rect 18609 1741 18643 1757
rect 18609 1691 18643 1707
rect 18945 1741 18979 1757
rect 18945 1691 18979 1707
rect 19281 1741 19315 1757
rect 19281 1691 19315 1707
rect 19617 1741 19651 1757
rect 19617 1691 19651 1707
rect 19953 1741 19987 1757
rect 19953 1691 19987 1707
rect 20289 1741 20323 1757
rect 20289 1691 20323 1707
rect 20625 1741 20659 1757
rect 20625 1691 20659 1707
rect 20961 1741 20995 1757
rect 20961 1691 20995 1707
rect 21297 1741 21331 1757
rect 21297 1691 21331 1707
rect 21633 1741 21667 1757
rect 21633 1691 21667 1707
rect 21969 1741 22003 1757
rect 21969 1691 22003 1707
rect 22305 1741 22339 1757
rect 22305 1691 22339 1707
rect 22641 1741 22675 1757
rect 22641 1691 22675 1707
rect 22977 1741 23011 1757
rect 22977 1691 23011 1707
rect 23313 1741 23347 1757
rect 23313 1691 23347 1707
rect 23649 1741 23683 1757
rect 23649 1691 23683 1707
rect 23985 1741 24019 1757
rect 23985 1691 24019 1707
rect 24321 1741 24355 1757
rect 24321 1691 24355 1707
rect 24657 1741 24691 1757
rect 24657 1691 24691 1707
rect 24993 1741 25027 1757
rect 24993 1691 25027 1707
rect 25329 1741 25363 1757
rect 25329 1691 25363 1707
rect 25665 1741 25699 1757
rect 25665 1691 25699 1707
rect 26001 1741 26035 1757
rect 26001 1691 26035 1707
rect 26337 1741 26371 1757
rect 26337 1691 26371 1707
rect 26673 1741 26707 1757
rect 26673 1691 26707 1707
rect 27009 1741 27043 1757
rect 27009 1691 27043 1707
rect 27345 1741 27379 1757
rect 27345 1691 27379 1707
rect 27681 1741 27715 1757
rect 27681 1691 27715 1707
rect 28017 1741 28051 1757
rect 28017 1691 28051 1707
rect 28353 1741 28387 1757
rect 28353 1691 28387 1707
rect 28689 1741 28723 1757
rect 28689 1691 28723 1707
rect 29025 1741 29059 1757
rect 29025 1691 29059 1707
rect 29361 1741 29395 1757
rect 29361 1691 29395 1707
rect 29697 1741 29731 1757
rect 29697 1691 29731 1707
rect 30033 1741 30067 1757
rect 30033 1691 30067 1707
rect 30369 1741 30403 1757
rect 30369 1691 30403 1707
rect 30705 1741 30739 1757
rect 30705 1691 30739 1707
rect 31041 1741 31075 1757
rect 31041 1691 31075 1707
rect 31377 1741 31411 1757
rect 31377 1691 31411 1707
rect 31713 1741 31747 1757
rect 31713 1691 31747 1707
rect 32049 1741 32083 1757
rect 32049 1691 32083 1707
rect 32385 1741 32419 1757
rect 32385 1691 32419 1707
rect 32721 1741 32755 1757
rect 32721 1691 32755 1707
rect 33057 1741 33091 1757
rect 33057 1691 33091 1707
rect 33393 1741 33427 1757
rect 33393 1691 33427 1707
rect 33729 1741 33763 1757
rect 33729 1691 33763 1707
rect 34065 1741 34099 1757
rect 34065 1691 34099 1707
rect 34401 1741 34435 1757
rect 34401 1691 34435 1707
rect 34737 1741 34771 1757
rect 34737 1691 34771 1707
rect 35073 1741 35107 1757
rect 35073 1691 35107 1707
rect 35409 1741 35443 1757
rect 35409 1691 35443 1707
rect 35745 1741 35779 1757
rect 35745 1691 35779 1707
rect 36081 1741 36115 1757
rect 36081 1691 36115 1707
rect 36417 1741 36451 1757
rect 36417 1691 36451 1707
rect 36753 1741 36787 1757
rect 36753 1691 36787 1707
rect 37089 1741 37123 1757
rect 37089 1691 37123 1707
rect 37425 1741 37459 1757
rect 37425 1691 37459 1707
rect 37761 1741 37795 1757
rect 37761 1691 37795 1707
rect 38097 1741 38131 1757
rect 38097 1691 38131 1707
rect 38433 1741 38467 1757
rect 38433 1691 38467 1707
rect 38769 1741 38803 1757
rect 38769 1691 38803 1707
rect 39105 1741 39139 1757
rect 39105 1691 39139 1707
rect 39441 1741 39475 1757
rect 39441 1691 39475 1707
rect 39777 1741 39811 1757
rect 39777 1691 39811 1707
rect 40113 1741 40147 1757
rect 40113 1691 40147 1707
rect 40449 1741 40483 1757
rect 40449 1691 40483 1707
rect 40785 1741 40819 1757
rect 40785 1691 40819 1707
rect 41121 1741 41155 1757
rect 41121 1691 41155 1707
rect 41457 1741 41491 1757
rect 41457 1691 41491 1707
rect 41793 1741 41827 1757
rect 41793 1691 41827 1707
rect 42129 1741 42163 1757
rect 42129 1691 42163 1707
rect 42465 1741 42499 1757
rect 42465 1691 42499 1707
rect 42801 1741 42835 1757
rect 42801 1691 42835 1707
rect 43137 1741 43171 1757
rect 43137 1691 43171 1707
rect 43473 1741 43507 1757
rect 43473 1691 43507 1707
rect 43809 1741 43843 1757
rect 43809 1691 43843 1707
rect 44145 1741 44179 1757
rect 44145 1691 44179 1707
rect 44481 1741 44515 1757
rect 44481 1691 44515 1707
rect 44817 1741 44851 1757
rect 44817 1691 44851 1707
rect 45153 1741 45187 1757
rect 45153 1691 45187 1707
rect 45489 1741 45523 1757
rect 45489 1691 45523 1707
rect 45825 1741 45859 1757
rect 45825 1691 45859 1707
rect 46161 1741 46195 1757
rect 46161 1691 46195 1707
rect 46497 1741 46531 1757
rect 46497 1691 46531 1707
rect 46833 1741 46867 1757
rect 46833 1691 46867 1707
rect 47169 1741 47203 1757
rect 47169 1691 47203 1707
rect 47505 1741 47539 1757
rect 47505 1691 47539 1707
rect 47841 1741 47875 1757
rect 47841 1691 47875 1707
rect 48177 1741 48211 1757
rect 48177 1691 48211 1707
rect 48513 1741 48547 1757
rect 48513 1691 48547 1707
rect 48849 1741 48883 1757
rect 48849 1691 48883 1707
rect 49185 1741 49219 1757
rect 49185 1691 49219 1707
rect 49521 1741 49555 1757
rect 49521 1691 49555 1707
rect 49857 1741 49891 1757
rect 49857 1691 49891 1707
rect 50193 1741 50227 1757
rect 50193 1691 50227 1707
rect 50529 1741 50563 1757
rect 50529 1691 50563 1707
rect 50865 1741 50899 1757
rect 50865 1691 50899 1707
rect 51201 1741 51235 1757
rect 51201 1691 51235 1707
rect 51537 1741 51571 1757
rect 51537 1691 51571 1707
rect 51873 1741 51907 1757
rect 51873 1691 51907 1707
rect 52209 1741 52243 1757
rect 52209 1691 52243 1707
rect 52545 1741 52579 1757
rect 52545 1691 52579 1707
rect 52881 1741 52915 1757
rect 52881 1691 52915 1707
rect 53217 1741 53251 1757
rect 53217 1691 53251 1707
rect 53553 1741 53587 1757
rect 53553 1691 53587 1707
rect 53889 1741 53923 1757
rect 53889 1691 53923 1707
rect 54225 1741 54259 1757
rect 54225 1691 54259 1707
rect 54561 1741 54595 1757
rect 54561 1691 54595 1707
rect 54897 1741 54931 1757
rect 54897 1691 54931 1707
rect 55233 1741 55267 1757
rect 55233 1691 55267 1707
rect 55569 1741 55603 1757
rect 55569 1691 55603 1707
rect 55905 1741 55939 1757
rect 55905 1691 55939 1707
rect 56241 1741 56275 1757
rect 56241 1691 56275 1707
rect 56577 1741 56611 1757
rect 56577 1691 56611 1707
rect 56913 1741 56947 1757
rect 56913 1691 56947 1707
rect 57249 1741 57283 1757
rect 57249 1691 57283 1707
rect 57585 1741 57619 1757
rect 57585 1691 57619 1707
rect 57921 1741 57955 1757
rect 57921 1691 57955 1707
rect 58257 1741 58291 1757
rect 58257 1691 58291 1707
rect 58593 1741 58627 1757
rect 58593 1691 58627 1707
rect 58929 1741 58963 1757
rect 58929 1691 58963 1707
rect 59265 1741 59299 1757
rect 59265 1691 59299 1707
rect 59601 1741 59635 1757
rect 59601 1691 59635 1707
rect 59937 1741 59971 1757
rect 59937 1691 59971 1707
rect 60273 1741 60307 1757
rect 60273 1691 60307 1707
rect 60609 1741 60643 1757
rect 60609 1691 60643 1707
rect 60945 1741 60979 1757
rect 60945 1691 60979 1707
rect 61281 1741 61315 1757
rect 61281 1691 61315 1707
rect 61617 1741 61651 1757
rect 61617 1691 61651 1707
rect 61953 1741 61987 1757
rect 61953 1691 61987 1707
rect 62289 1741 62323 1757
rect 62289 1691 62323 1707
rect 62625 1741 62659 1757
rect 62625 1691 62659 1707
rect 62961 1741 62995 1757
rect 62961 1691 62995 1707
rect 63297 1741 63331 1757
rect 63297 1691 63331 1707
rect 63633 1741 63667 1757
rect 63633 1691 63667 1707
rect 63969 1741 64003 1757
rect 63969 1691 64003 1707
rect 64305 1741 64339 1757
rect 64305 1691 64339 1707
rect 64641 1741 64675 1757
rect 64641 1691 64675 1707
rect 64977 1741 65011 1757
rect 64977 1691 65011 1707
rect 65313 1741 65347 1757
rect 65313 1691 65347 1707
rect 65649 1741 65683 1757
rect 65649 1691 65683 1707
rect 65985 1741 66019 1757
rect 65985 1691 66019 1707
rect 66321 1741 66355 1757
rect 66321 1691 66355 1707
rect 66657 1741 66691 1757
rect 66657 1691 66691 1707
rect 66993 1741 67027 1757
rect 66993 1691 67027 1707
rect 67329 1741 67363 1757
rect 67329 1691 67363 1707
rect 67665 1741 67699 1757
rect 67665 1691 67699 1707
rect 68001 1741 68035 1757
rect 68001 1691 68035 1707
rect 68337 1741 68371 1757
rect 68337 1691 68371 1707
rect 68673 1741 68707 1757
rect 68673 1691 68707 1707
rect 69009 1741 69043 1757
rect 69009 1691 69043 1707
rect 69345 1741 69379 1757
rect 69345 1691 69379 1707
rect 69681 1741 69715 1757
rect 69681 1691 69715 1707
rect 70017 1741 70051 1757
rect 70017 1691 70051 1707
rect 70353 1741 70387 1757
rect 70353 1691 70387 1707
rect 70689 1741 70723 1757
rect 70689 1691 70723 1707
rect 71025 1741 71059 1757
rect 71025 1691 71059 1707
rect 71361 1741 71395 1757
rect 71361 1691 71395 1707
rect 71697 1741 71731 1757
rect 71697 1691 71731 1707
rect 72033 1741 72067 1757
rect 72033 1691 72067 1707
rect 72369 1741 72403 1757
rect 72369 1691 72403 1707
rect 72705 1741 72739 1757
rect 72705 1691 72739 1707
rect 73041 1741 73075 1757
rect 73041 1691 73075 1707
rect 73377 1741 73411 1757
rect 73377 1691 73411 1707
rect 73713 1741 73747 1757
rect 73713 1691 73747 1707
rect 74049 1741 74083 1757
rect 74049 1691 74083 1707
rect 74385 1741 74419 1757
rect 74385 1691 74419 1707
rect 74721 1741 74755 1757
rect 74721 1691 74755 1707
rect 75057 1741 75091 1757
rect 75057 1691 75091 1707
rect 75393 1741 75427 1757
rect 75393 1691 75427 1707
rect 75729 1741 75763 1757
rect 75729 1691 75763 1707
rect 76065 1741 76099 1757
rect 76065 1691 76099 1707
rect 76401 1741 76435 1757
rect 76401 1691 76435 1707
rect 76737 1741 76771 1757
rect 76737 1691 76771 1707
rect 77073 1741 77107 1757
rect 77073 1691 77107 1707
rect 77409 1741 77443 1757
rect 77409 1691 77443 1707
rect 77745 1741 77779 1757
rect 77745 1691 77779 1707
rect 78081 1741 78115 1757
rect 78081 1691 78115 1707
rect 78417 1741 78451 1757
rect 78417 1691 78451 1707
rect 78753 1741 78787 1757
rect 78753 1691 78787 1707
rect 79089 1741 79123 1757
rect 79089 1691 79123 1707
rect 79425 1741 79459 1757
rect 79425 1691 79459 1707
rect 79761 1741 79795 1757
rect 79761 1691 79795 1707
rect 80097 1741 80131 1757
rect 80097 1691 80131 1707
rect 80433 1741 80467 1757
rect 80433 1691 80467 1707
rect 80769 1741 80803 1757
rect 80769 1691 80803 1707
rect 81105 1741 81139 1757
rect 81105 1691 81139 1707
rect 81441 1741 81475 1757
rect 81441 1691 81475 1707
rect 81777 1741 81811 1757
rect 81777 1691 81811 1707
rect 82113 1741 82147 1757
rect 82113 1691 82147 1707
rect 82449 1741 82483 1757
rect 82449 1691 82483 1707
rect 82785 1741 82819 1757
rect 82785 1691 82819 1707
rect 83121 1741 83155 1757
rect 83121 1691 83155 1707
rect 83457 1741 83491 1757
rect 83457 1691 83491 1707
rect 83793 1741 83827 1757
rect 83793 1691 83827 1707
rect 84129 1741 84163 1757
rect 84129 1691 84163 1707
rect 84465 1741 84499 1757
rect 84465 1691 84499 1707
rect 84801 1741 84835 1757
rect 84801 1691 84835 1707
rect 85137 1741 85171 1757
rect 85137 1691 85171 1707
rect 85473 1741 85507 1757
rect 85473 1691 85507 1707
rect 85809 1741 85843 1757
rect 85809 1691 85843 1707
rect 86145 1741 86179 1757
rect 86145 1691 86179 1707
rect 86481 1741 86515 1757
rect 86481 1691 86515 1707
rect 86817 1741 86851 1757
rect 86817 1691 86851 1707
rect 87153 1741 87187 1757
rect 87153 1691 87187 1707
rect 87489 1741 87523 1757
rect 87489 1691 87523 1707
rect 87825 1741 87859 1757
rect 87825 1691 87859 1707
rect 88161 1741 88195 1757
rect 88161 1691 88195 1707
rect 88497 1741 88531 1757
rect 88497 1691 88531 1707
rect 88833 1741 88867 1757
rect 88833 1691 88867 1707
rect 89169 1741 89203 1757
rect 89169 1691 89203 1707
rect 89505 1741 89539 1757
rect 89505 1691 89539 1707
rect 89841 1741 89875 1757
rect 89841 1691 89875 1707
rect 90177 1741 90211 1757
rect 90177 1691 90211 1707
rect 90513 1741 90547 1757
rect 90513 1691 90547 1707
rect 90849 1741 90883 1757
rect 90849 1691 90883 1707
rect 91185 1741 91219 1757
rect 91185 1691 91219 1707
rect 91521 1741 91555 1757
rect 91521 1691 91555 1707
rect 91857 1741 91891 1757
rect 91857 1691 91891 1707
rect 92193 1741 92227 1757
rect 92193 1691 92227 1707
rect 92529 1741 92563 1757
rect 92529 1691 92563 1707
rect 92865 1741 92899 1757
rect 92865 1691 92899 1707
rect 93201 1741 93235 1757
rect 93201 1691 93235 1707
rect 93537 1741 93571 1757
rect 93537 1691 93571 1707
rect 93873 1741 93907 1757
rect 93873 1691 93907 1707
rect 94209 1741 94243 1757
rect 94209 1691 94243 1707
rect 94545 1741 94579 1757
rect 94545 1691 94579 1707
rect 94881 1741 94915 1757
rect 94881 1691 94915 1707
rect 95217 1741 95251 1757
rect 95217 1691 95251 1707
rect 95553 1741 95587 1757
rect 95553 1691 95587 1707
rect 95889 1741 95923 1757
rect 95889 1691 95923 1707
rect 96225 1741 96259 1757
rect 96225 1691 96259 1707
rect 96561 1741 96595 1757
rect 96561 1691 96595 1707
rect 96897 1741 96931 1757
rect 96897 1691 96931 1707
rect 97233 1741 97267 1757
rect 97233 1691 97267 1707
rect 97569 1741 97603 1757
rect 97569 1691 97603 1707
rect 97905 1741 97939 1757
rect 97905 1691 97939 1707
rect 98241 1741 98275 1757
rect 98241 1691 98275 1707
rect 98577 1741 98611 1757
rect 98577 1691 98611 1707
rect 98913 1741 98947 1757
rect 98913 1691 98947 1707
rect 99249 1741 99283 1757
rect 99249 1691 99283 1707
rect 99585 1741 99619 1757
rect 99585 1691 99619 1707
rect 99921 1741 99955 1757
rect 99921 1691 99955 1707
rect 100257 1741 100291 1757
rect 100257 1691 100291 1707
rect 100593 1741 100627 1757
rect 100593 1691 100627 1707
rect 100929 1741 100963 1757
rect 100929 1691 100963 1707
rect 101265 1741 101299 1757
rect 101265 1691 101299 1707
rect 101601 1741 101635 1757
rect 101601 1691 101635 1707
rect 101937 1741 101971 1757
rect 101937 1691 101971 1707
rect 102273 1741 102307 1757
rect 102273 1691 102307 1707
rect 102609 1741 102643 1757
rect 102609 1691 102643 1707
rect 102945 1741 102979 1757
rect 102945 1691 102979 1707
rect 103281 1741 103315 1757
rect 103281 1691 103315 1707
rect 103617 1741 103651 1757
rect 103617 1691 103651 1707
rect 103953 1741 103987 1757
rect 103953 1691 103987 1707
rect 104289 1741 104323 1757
rect 104289 1691 104323 1707
rect 104625 1741 104659 1757
rect 104625 1691 104659 1707
rect 104961 1741 104995 1757
rect 104961 1691 104995 1707
rect 105297 1741 105331 1757
rect 105297 1691 105331 1707
rect 105633 1741 105667 1757
rect 105633 1691 105667 1707
rect 105969 1741 106003 1757
rect 105969 1691 106003 1707
rect 106305 1741 106339 1757
rect 106305 1691 106339 1707
rect 106641 1741 106675 1757
rect 106641 1691 106675 1707
rect 106977 1741 107011 1757
rect 106977 1691 107011 1707
rect 107313 1741 107347 1757
rect 107313 1691 107347 1707
rect 107649 1741 107683 1757
rect 107649 1691 107683 1707
rect 107985 1741 108019 1757
rect 107985 1691 108019 1707
rect 108321 1741 108355 1757
rect 108321 1691 108355 1707
rect 108657 1741 108691 1757
rect 108657 1691 108691 1707
rect 108993 1741 109027 1757
rect 108993 1691 109027 1707
rect 109329 1741 109363 1757
rect 109329 1691 109363 1707
rect 109665 1741 109699 1757
rect 109665 1691 109699 1707
rect 110001 1741 110035 1757
rect 110001 1691 110035 1707
rect 110337 1741 110371 1757
rect 110337 1691 110371 1707
rect 110673 1741 110707 1757
rect 110673 1691 110707 1707
rect 111009 1741 111043 1757
rect 111009 1691 111043 1707
rect 111345 1741 111379 1757
rect 111345 1691 111379 1707
rect 111681 1741 111715 1757
rect 111681 1691 111715 1707
rect 112017 1741 112051 1757
rect 112017 1691 112051 1707
rect 112353 1741 112387 1757
rect 112353 1691 112387 1707
rect 112689 1741 112723 1757
rect 112689 1691 112723 1707
rect 113025 1741 113059 1757
rect 113025 1691 113059 1707
rect 113361 1741 113395 1757
rect 113361 1691 113395 1707
rect 113697 1741 113731 1757
rect 113697 1691 113731 1707
rect 114033 1741 114067 1757
rect 114033 1691 114067 1707
rect 114369 1741 114403 1757
rect 114369 1691 114403 1707
rect 114705 1741 114739 1757
rect 114705 1691 114739 1707
rect 115041 1741 115075 1757
rect 115041 1691 115075 1707
rect 115377 1741 115411 1757
rect 115377 1691 115411 1707
rect 115713 1741 115747 1757
rect 115713 1691 115747 1707
rect 116049 1741 116083 1757
rect 116049 1691 116083 1707
rect 116385 1741 116419 1757
rect 116385 1691 116419 1707
rect 116721 1741 116755 1757
rect 116721 1691 116755 1707
rect 117057 1741 117091 1757
rect 117057 1691 117091 1707
rect 117393 1741 117427 1757
rect 117393 1691 117427 1707
rect 117729 1741 117763 1757
rect 117729 1691 117763 1707
rect 118065 1741 118099 1757
rect 118065 1691 118099 1707
rect 118401 1741 118435 1757
rect 118401 1691 118435 1707
rect 118737 1741 118771 1757
rect 118737 1691 118771 1707
rect 119073 1741 119107 1757
rect 119073 1691 119107 1707
rect 119409 1741 119443 1757
rect 119409 1691 119443 1707
rect 119745 1741 119779 1757
rect 119745 1691 119779 1707
rect 120081 1741 120115 1757
rect 120081 1691 120115 1707
rect 120417 1741 120451 1757
rect 120417 1691 120451 1707
rect 120753 1741 120787 1757
rect 120753 1691 120787 1707
rect 121089 1741 121123 1757
rect 121089 1691 121123 1707
rect 121425 1741 121459 1757
rect 121425 1691 121459 1707
rect 121761 1741 121795 1757
rect 121761 1691 121795 1707
rect 122097 1741 122131 1757
rect 122097 1691 122131 1707
rect 122433 1741 122467 1757
rect 122433 1691 122467 1707
rect 122769 1741 122803 1757
rect 122769 1691 122803 1707
rect 123105 1741 123139 1757
rect 123105 1691 123139 1707
rect 123441 1741 123475 1757
rect 123441 1691 123475 1707
rect 123777 1741 123811 1757
rect 123777 1691 123811 1707
rect 124113 1741 124147 1757
rect 124113 1691 124147 1707
rect 124449 1741 124483 1757
rect 124449 1691 124483 1707
rect 124785 1741 124819 1757
rect 124785 1691 124819 1707
rect 125121 1741 125155 1757
rect 125121 1691 125155 1707
rect 125457 1741 125491 1757
rect 125457 1691 125491 1707
rect 125793 1741 125827 1757
rect 125793 1691 125827 1707
rect 126129 1741 126163 1757
rect 126129 1691 126163 1707
rect 126465 1741 126499 1757
rect 126465 1691 126499 1707
rect 126801 1741 126835 1757
rect 126801 1691 126835 1707
rect 127137 1741 127171 1757
rect 127137 1691 127171 1707
rect 127473 1741 127507 1757
rect 127473 1691 127507 1707
rect 127809 1741 127843 1757
rect 127809 1691 127843 1707
rect 128145 1741 128179 1757
rect 128145 1691 128179 1707
rect 128481 1741 128515 1757
rect 128481 1691 128515 1707
rect 128817 1741 128851 1757
rect 128817 1691 128851 1707
rect 129153 1741 129187 1757
rect 129153 1691 129187 1707
rect 129489 1741 129523 1757
rect 129489 1691 129523 1707
rect 129825 1741 129859 1757
rect 129825 1691 129859 1707
rect 130161 1741 130195 1757
rect 130161 1691 130195 1707
rect 130497 1741 130531 1757
rect 130497 1691 130531 1707
rect 130833 1741 130867 1757
rect 130833 1691 130867 1707
rect 131169 1741 131203 1757
rect 131169 1691 131203 1707
rect 131505 1741 131539 1757
rect 131505 1691 131539 1707
rect 131841 1741 131875 1757
rect 131841 1691 131875 1707
rect 132177 1741 132211 1757
rect 132177 1691 132211 1707
rect 132513 1741 132547 1757
rect 132513 1691 132547 1707
rect 132849 1741 132883 1757
rect 132849 1691 132883 1707
rect 133185 1741 133219 1757
rect 133185 1691 133219 1707
rect 133521 1741 133555 1757
rect 133521 1691 133555 1707
rect 133857 1741 133891 1757
rect 133857 1691 133891 1707
rect 134193 1741 134227 1757
rect 134193 1691 134227 1707
rect 134529 1741 134563 1757
rect 134529 1691 134563 1707
rect 134865 1741 134899 1757
rect 134865 1691 134899 1707
rect 135201 1741 135235 1757
rect 135201 1691 135235 1707
rect 135537 1741 135571 1757
rect 135537 1691 135571 1707
rect 135873 1741 135907 1757
rect 135873 1691 135907 1707
rect 136209 1741 136243 1757
rect 136209 1691 136243 1707
rect 136545 1741 136579 1757
rect 136545 1691 136579 1707
<< viali >>
rect 2145 132016 2179 132050
rect 2481 132016 2515 132050
rect 2817 132016 2851 132050
rect 3153 132016 3187 132050
rect 3489 132016 3523 132050
rect 3825 132016 3859 132050
rect 4161 132016 4195 132050
rect 4497 132016 4531 132050
rect 4833 132016 4867 132050
rect 5169 132016 5203 132050
rect 5505 132016 5539 132050
rect 5841 132016 5875 132050
rect 6177 132016 6211 132050
rect 6513 132016 6547 132050
rect 6849 132016 6883 132050
rect 7185 132016 7219 132050
rect 7521 132016 7555 132050
rect 7857 132016 7891 132050
rect 8193 132016 8227 132050
rect 8529 132016 8563 132050
rect 8865 132016 8899 132050
rect 9201 132016 9235 132050
rect 9537 132016 9571 132050
rect 9873 132016 9907 132050
rect 10209 132016 10243 132050
rect 10545 132016 10579 132050
rect 10881 132016 10915 132050
rect 11217 132016 11251 132050
rect 11553 132016 11587 132050
rect 11889 132016 11923 132050
rect 12225 132016 12259 132050
rect 12561 132016 12595 132050
rect 12897 132016 12931 132050
rect 13233 132016 13267 132050
rect 13569 132016 13603 132050
rect 13905 132016 13939 132050
rect 14241 132016 14275 132050
rect 14577 132016 14611 132050
rect 14913 132016 14947 132050
rect 15249 132016 15283 132050
rect 15585 132016 15619 132050
rect 15921 132016 15955 132050
rect 16257 132016 16291 132050
rect 16593 132016 16627 132050
rect 16929 132016 16963 132050
rect 17265 132016 17299 132050
rect 17601 132016 17635 132050
rect 17937 132016 17971 132050
rect 18273 132016 18307 132050
rect 18609 132016 18643 132050
rect 18945 132016 18979 132050
rect 19281 132016 19315 132050
rect 19617 132016 19651 132050
rect 19953 132016 19987 132050
rect 20289 132016 20323 132050
rect 20625 132016 20659 132050
rect 20961 132016 20995 132050
rect 21297 132016 21331 132050
rect 21633 132016 21667 132050
rect 21969 132016 22003 132050
rect 22305 132016 22339 132050
rect 22641 132016 22675 132050
rect 22977 132016 23011 132050
rect 23313 132016 23347 132050
rect 23649 132016 23683 132050
rect 23985 132016 24019 132050
rect 24321 132016 24355 132050
rect 24657 132016 24691 132050
rect 24993 132016 25027 132050
rect 25329 132016 25363 132050
rect 25665 132016 25699 132050
rect 26001 132016 26035 132050
rect 26337 132016 26371 132050
rect 26673 132016 26707 132050
rect 27009 132016 27043 132050
rect 27345 132016 27379 132050
rect 27681 132016 27715 132050
rect 28017 132016 28051 132050
rect 28353 132016 28387 132050
rect 28689 132016 28723 132050
rect 29025 132016 29059 132050
rect 29361 132016 29395 132050
rect 29697 132016 29731 132050
rect 30033 132016 30067 132050
rect 30369 132016 30403 132050
rect 30705 132016 30739 132050
rect 31041 132016 31075 132050
rect 31377 132016 31411 132050
rect 31713 132016 31747 132050
rect 32049 132016 32083 132050
rect 32385 132016 32419 132050
rect 32721 132016 32755 132050
rect 33057 132016 33091 132050
rect 33393 132016 33427 132050
rect 33729 132016 33763 132050
rect 34065 132016 34099 132050
rect 34401 132016 34435 132050
rect 34737 132016 34771 132050
rect 35073 132016 35107 132050
rect 35409 132016 35443 132050
rect 35745 132016 35779 132050
rect 36081 132016 36115 132050
rect 36417 132016 36451 132050
rect 36753 132016 36787 132050
rect 37089 132016 37123 132050
rect 37425 132016 37459 132050
rect 37761 132016 37795 132050
rect 38097 132016 38131 132050
rect 38433 132016 38467 132050
rect 38769 132016 38803 132050
rect 39105 132016 39139 132050
rect 39441 132016 39475 132050
rect 39777 132016 39811 132050
rect 40113 132016 40147 132050
rect 40449 132016 40483 132050
rect 40785 132016 40819 132050
rect 41121 132016 41155 132050
rect 41457 132016 41491 132050
rect 41793 132016 41827 132050
rect 42129 132016 42163 132050
rect 42465 132016 42499 132050
rect 42801 132016 42835 132050
rect 43137 132016 43171 132050
rect 43473 132016 43507 132050
rect 43809 132016 43843 132050
rect 44145 132016 44179 132050
rect 44481 132016 44515 132050
rect 44817 132016 44851 132050
rect 45153 132016 45187 132050
rect 45489 132016 45523 132050
rect 45825 132016 45859 132050
rect 46161 132016 46195 132050
rect 46497 132016 46531 132050
rect 46833 132016 46867 132050
rect 47169 132016 47203 132050
rect 47505 132016 47539 132050
rect 47841 132016 47875 132050
rect 48177 132016 48211 132050
rect 48513 132016 48547 132050
rect 48849 132016 48883 132050
rect 49185 132016 49219 132050
rect 49521 132016 49555 132050
rect 49857 132016 49891 132050
rect 50193 132016 50227 132050
rect 50529 132016 50563 132050
rect 50865 132016 50899 132050
rect 51201 132016 51235 132050
rect 51537 132016 51571 132050
rect 51873 132016 51907 132050
rect 52209 132016 52243 132050
rect 52545 132016 52579 132050
rect 52881 132016 52915 132050
rect 53217 132016 53251 132050
rect 53553 132016 53587 132050
rect 53889 132016 53923 132050
rect 54225 132016 54259 132050
rect 54561 132016 54595 132050
rect 54897 132016 54931 132050
rect 55233 132016 55267 132050
rect 55569 132016 55603 132050
rect 55905 132016 55939 132050
rect 56241 132016 56275 132050
rect 56577 132016 56611 132050
rect 56913 132016 56947 132050
rect 57249 132016 57283 132050
rect 57585 132016 57619 132050
rect 57921 132016 57955 132050
rect 58257 132016 58291 132050
rect 58593 132016 58627 132050
rect 58929 132016 58963 132050
rect 59265 132016 59299 132050
rect 59601 132016 59635 132050
rect 59937 132016 59971 132050
rect 60273 132016 60307 132050
rect 60609 132016 60643 132050
rect 60945 132016 60979 132050
rect 61281 132016 61315 132050
rect 61617 132016 61651 132050
rect 61953 132016 61987 132050
rect 62289 132016 62323 132050
rect 62625 132016 62659 132050
rect 62961 132016 62995 132050
rect 63297 132016 63331 132050
rect 63633 132016 63667 132050
rect 63969 132016 64003 132050
rect 64305 132016 64339 132050
rect 64641 132016 64675 132050
rect 64977 132016 65011 132050
rect 65313 132016 65347 132050
rect 65649 132016 65683 132050
rect 65985 132016 66019 132050
rect 66321 132016 66355 132050
rect 66657 132016 66691 132050
rect 66993 132016 67027 132050
rect 67329 132016 67363 132050
rect 67665 132016 67699 132050
rect 68001 132016 68035 132050
rect 68337 132016 68371 132050
rect 68673 132016 68707 132050
rect 69009 132016 69043 132050
rect 69345 132016 69379 132050
rect 69681 132016 69715 132050
rect 70017 132016 70051 132050
rect 70353 132016 70387 132050
rect 70689 132016 70723 132050
rect 71025 132016 71059 132050
rect 71361 132016 71395 132050
rect 71697 132016 71731 132050
rect 72033 132016 72067 132050
rect 72369 132016 72403 132050
rect 72705 132016 72739 132050
rect 73041 132016 73075 132050
rect 73377 132016 73411 132050
rect 73713 132016 73747 132050
rect 74049 132016 74083 132050
rect 74385 132016 74419 132050
rect 74721 132016 74755 132050
rect 75057 132016 75091 132050
rect 75393 132016 75427 132050
rect 75729 132016 75763 132050
rect 76065 132016 76099 132050
rect 76401 132016 76435 132050
rect 76737 132016 76771 132050
rect 77073 132016 77107 132050
rect 77409 132016 77443 132050
rect 77745 132016 77779 132050
rect 78081 132016 78115 132050
rect 78417 132016 78451 132050
rect 78753 132016 78787 132050
rect 79089 132016 79123 132050
rect 79425 132016 79459 132050
rect 79761 132016 79795 132050
rect 80097 132016 80131 132050
rect 80433 132016 80467 132050
rect 80769 132016 80803 132050
rect 81105 132016 81139 132050
rect 81441 132016 81475 132050
rect 81777 132016 81811 132050
rect 82113 132016 82147 132050
rect 82449 132016 82483 132050
rect 82785 132016 82819 132050
rect 83121 132016 83155 132050
rect 83457 132016 83491 132050
rect 83793 132016 83827 132050
rect 84129 132016 84163 132050
rect 84465 132016 84499 132050
rect 84801 132016 84835 132050
rect 85137 132016 85171 132050
rect 85473 132016 85507 132050
rect 85809 132016 85843 132050
rect 86145 132016 86179 132050
rect 86481 132016 86515 132050
rect 86817 132016 86851 132050
rect 87153 132016 87187 132050
rect 87489 132016 87523 132050
rect 87825 132016 87859 132050
rect 88161 132016 88195 132050
rect 88497 132016 88531 132050
rect 88833 132016 88867 132050
rect 89169 132016 89203 132050
rect 89505 132016 89539 132050
rect 89841 132016 89875 132050
rect 90177 132016 90211 132050
rect 90513 132016 90547 132050
rect 90849 132016 90883 132050
rect 91185 132016 91219 132050
rect 91521 132016 91555 132050
rect 91857 132016 91891 132050
rect 92193 132016 92227 132050
rect 92529 132016 92563 132050
rect 92865 132016 92899 132050
rect 93201 132016 93235 132050
rect 93537 132016 93571 132050
rect 93873 132016 93907 132050
rect 94209 132016 94243 132050
rect 94545 132016 94579 132050
rect 94881 132016 94915 132050
rect 95217 132016 95251 132050
rect 95553 132016 95587 132050
rect 95889 132016 95923 132050
rect 96225 132016 96259 132050
rect 96561 132016 96595 132050
rect 96897 132016 96931 132050
rect 97233 132016 97267 132050
rect 97569 132016 97603 132050
rect 97905 132016 97939 132050
rect 98241 132016 98275 132050
rect 98577 132016 98611 132050
rect 98913 132016 98947 132050
rect 99249 132016 99283 132050
rect 99585 132016 99619 132050
rect 99921 132016 99955 132050
rect 100257 132016 100291 132050
rect 100593 132016 100627 132050
rect 100929 132016 100963 132050
rect 101265 132016 101299 132050
rect 101601 132016 101635 132050
rect 101937 132016 101971 132050
rect 102273 132016 102307 132050
rect 102609 132016 102643 132050
rect 102945 132016 102979 132050
rect 103281 132016 103315 132050
rect 103617 132016 103651 132050
rect 103953 132016 103987 132050
rect 104289 132016 104323 132050
rect 104625 132016 104659 132050
rect 104961 132016 104995 132050
rect 105297 132016 105331 132050
rect 105633 132016 105667 132050
rect 105969 132016 106003 132050
rect 106305 132016 106339 132050
rect 106641 132016 106675 132050
rect 106977 132016 107011 132050
rect 107313 132016 107347 132050
rect 107649 132016 107683 132050
rect 107985 132016 108019 132050
rect 108321 132016 108355 132050
rect 108657 132016 108691 132050
rect 108993 132016 109027 132050
rect 109329 132016 109363 132050
rect 109665 132016 109699 132050
rect 110001 132016 110035 132050
rect 110337 132016 110371 132050
rect 110673 132016 110707 132050
rect 111009 132016 111043 132050
rect 111345 132016 111379 132050
rect 111681 132016 111715 132050
rect 112017 132016 112051 132050
rect 112353 132016 112387 132050
rect 112689 132016 112723 132050
rect 113025 132016 113059 132050
rect 113361 132016 113395 132050
rect 113697 132016 113731 132050
rect 114033 132016 114067 132050
rect 114369 132016 114403 132050
rect 114705 132016 114739 132050
rect 115041 132016 115075 132050
rect 115377 132016 115411 132050
rect 115713 132016 115747 132050
rect 116049 132016 116083 132050
rect 116385 132016 116419 132050
rect 116721 132016 116755 132050
rect 117057 132016 117091 132050
rect 117393 132016 117427 132050
rect 117729 132016 117763 132050
rect 118065 132016 118099 132050
rect 118401 132016 118435 132050
rect 118737 132016 118771 132050
rect 119073 132016 119107 132050
rect 119409 132016 119443 132050
rect 119745 132016 119779 132050
rect 120081 132016 120115 132050
rect 120417 132016 120451 132050
rect 120753 132016 120787 132050
rect 121089 132016 121123 132050
rect 121425 132016 121459 132050
rect 121761 132016 121795 132050
rect 122097 132016 122131 132050
rect 122433 132016 122467 132050
rect 122769 132016 122803 132050
rect 123105 132016 123139 132050
rect 123441 132016 123475 132050
rect 123777 132016 123811 132050
rect 124113 132016 124147 132050
rect 124449 132016 124483 132050
rect 124785 132016 124819 132050
rect 125121 132016 125155 132050
rect 125457 132016 125491 132050
rect 125793 132016 125827 132050
rect 126129 132016 126163 132050
rect 126465 132016 126499 132050
rect 126801 132016 126835 132050
rect 127137 132016 127171 132050
rect 127473 132016 127507 132050
rect 127809 132016 127843 132050
rect 128145 132016 128179 132050
rect 128481 132016 128515 132050
rect 128817 132016 128851 132050
rect 129153 132016 129187 132050
rect 129489 132016 129523 132050
rect 129825 132016 129859 132050
rect 130161 132016 130195 132050
rect 130497 132016 130531 132050
rect 130833 132016 130867 132050
rect 131169 132016 131203 132050
rect 131505 132016 131539 132050
rect 131841 132016 131875 132050
rect 132177 132016 132211 132050
rect 132513 132016 132547 132050
rect 132849 132016 132883 132050
rect 133185 132016 133219 132050
rect 133521 132016 133555 132050
rect 133857 132016 133891 132050
rect 134193 132016 134227 132050
rect 134529 132016 134563 132050
rect 134865 132016 134899 132050
rect 135201 132016 135235 132050
rect 135537 132016 135571 132050
rect 135873 132016 135907 132050
rect 136209 132016 136243 132050
rect 136545 132016 136579 132050
rect 1809 131403 1843 131437
rect 136955 131403 136989 131437
rect 1809 131067 1843 131101
rect 136955 131067 136989 131101
rect 1809 130731 1843 130765
rect 136955 130731 136989 130765
rect 1809 130395 1843 130429
rect 136955 130395 136989 130429
rect 1809 130059 1843 130093
rect 136955 130059 136989 130093
rect 1809 129723 1843 129757
rect 136955 129723 136989 129757
rect 1809 129387 1843 129421
rect 136955 129387 136989 129421
rect 1809 129051 1843 129085
rect 136955 129051 136989 129085
rect 1809 128715 1843 128749
rect 136955 128715 136989 128749
rect 1809 128379 1843 128413
rect 136955 128379 136989 128413
rect 1809 128043 1843 128077
rect 136955 128043 136989 128077
rect 1809 127707 1843 127741
rect 136955 127707 136989 127741
rect 1809 127371 1843 127405
rect 136955 127371 136989 127405
rect 1809 127035 1843 127069
rect 136955 127035 136989 127069
rect 1809 126699 1843 126733
rect 136955 126699 136989 126733
rect 1809 126363 1843 126397
rect 136955 126363 136989 126397
rect 1809 126027 1843 126061
rect 136955 126027 136989 126061
rect 1809 125691 1843 125725
rect 136955 125691 136989 125725
rect 1809 125355 1843 125389
rect 136955 125355 136989 125389
rect 1809 125019 1843 125053
rect 136955 125019 136989 125053
rect 1809 124683 1843 124717
rect 136955 124683 136989 124717
rect 1809 124347 1843 124381
rect 136955 124347 136989 124381
rect 1809 124011 1843 124045
rect 136955 124011 136989 124045
rect 1809 123675 1843 123709
rect 136955 123675 136989 123709
rect 1809 123339 1843 123373
rect 136955 123339 136989 123373
rect 1809 123003 1843 123037
rect 136955 123003 136989 123037
rect 1809 122667 1843 122701
rect 136955 122667 136989 122701
rect 1809 122331 1843 122365
rect 136955 122331 136989 122365
rect 1809 121995 1843 122029
rect 136955 121995 136989 122029
rect 1809 121659 1843 121693
rect 136955 121659 136989 121693
rect 1809 121323 1843 121357
rect 136955 121323 136989 121357
rect 1809 120987 1843 121021
rect 136955 120987 136989 121021
rect 1809 120651 1843 120685
rect 136955 120651 136989 120685
rect 1809 120315 1843 120349
rect 136955 120315 136989 120349
rect 1809 119979 1843 120013
rect 136955 119979 136989 120013
rect 1809 119643 1843 119677
rect 136955 119643 136989 119677
rect 1809 119307 1843 119341
rect 136955 119307 136989 119341
rect 1809 118971 1843 119005
rect 136955 118971 136989 119005
rect 1809 118635 1843 118669
rect 136955 118635 136989 118669
rect 1809 118299 1843 118333
rect 136955 118299 136989 118333
rect 1809 117963 1843 117997
rect 136955 117963 136989 117997
rect 1809 117627 1843 117661
rect 136955 117627 136989 117661
rect 1809 117291 1843 117325
rect 136955 117291 136989 117325
rect 1809 116955 1843 116989
rect 136955 116955 136989 116989
rect 1809 116619 1843 116653
rect 136955 116619 136989 116653
rect 1809 116283 1843 116317
rect 136955 116283 136989 116317
rect 1809 115947 1843 115981
rect 136955 115947 136989 115981
rect 1809 115611 1843 115645
rect 136955 115611 136989 115645
rect 1809 115275 1843 115309
rect 136955 115275 136989 115309
rect 1809 114939 1843 114973
rect 136955 114939 136989 114973
rect 1809 114603 1843 114637
rect 136955 114603 136989 114637
rect 1809 114267 1843 114301
rect 136955 114267 136989 114301
rect 1809 113931 1843 113965
rect 136955 113931 136989 113965
rect 1809 113595 1843 113629
rect 136955 113595 136989 113629
rect 1809 113259 1843 113293
rect 136955 113259 136989 113293
rect 1809 112923 1843 112957
rect 136955 112923 136989 112957
rect 1809 112587 1843 112621
rect 136955 112587 136989 112621
rect 1809 112251 1843 112285
rect 136955 112251 136989 112285
rect 1809 111915 1843 111949
rect 136955 111915 136989 111949
rect 1809 111579 1843 111613
rect 136955 111579 136989 111613
rect 1809 111243 1843 111277
rect 136955 111243 136989 111277
rect 1809 110907 1843 110941
rect 136955 110907 136989 110941
rect 1809 110571 1843 110605
rect 136955 110571 136989 110605
rect 1809 110235 1843 110269
rect 136955 110235 136989 110269
rect 1809 109899 1843 109933
rect 136955 109899 136989 109933
rect 1809 109563 1843 109597
rect 136955 109563 136989 109597
rect 1809 109227 1843 109261
rect 136955 109227 136989 109261
rect 1809 108891 1843 108925
rect 136955 108891 136989 108925
rect 1809 108555 1843 108589
rect 136955 108555 136989 108589
rect 1809 108219 1843 108253
rect 136955 108219 136989 108253
rect 1809 107883 1843 107917
rect 136955 107883 136989 107917
rect 1809 107547 1843 107581
rect 136955 107547 136989 107581
rect 1809 107211 1843 107245
rect 136955 107211 136989 107245
rect 1809 106875 1843 106909
rect 136955 106875 136989 106909
rect 1809 106539 1843 106573
rect 136955 106539 136989 106573
rect 1809 106203 1843 106237
rect 136955 106203 136989 106237
rect 1809 105867 1843 105901
rect 136955 105867 136989 105901
rect 1809 105531 1843 105565
rect 136955 105531 136989 105565
rect 1809 105195 1843 105229
rect 136955 105195 136989 105229
rect 1809 104859 1843 104893
rect 136955 104859 136989 104893
rect 1809 104523 1843 104557
rect 136955 104523 136989 104557
rect 1809 104187 1843 104221
rect 136955 104187 136989 104221
rect 1809 103851 1843 103885
rect 136955 103851 136989 103885
rect 1809 103515 1843 103549
rect 136955 103515 136989 103549
rect 1809 103179 1843 103213
rect 136955 103179 136989 103213
rect 1809 102843 1843 102877
rect 136955 102843 136989 102877
rect 1809 102507 1843 102541
rect 136955 102507 136989 102541
rect 1809 102171 1843 102205
rect 136955 102171 136989 102205
rect 1809 101835 1843 101869
rect 136955 101835 136989 101869
rect 1809 101499 1843 101533
rect 136955 101499 136989 101533
rect 1809 101163 1843 101197
rect 136955 101163 136989 101197
rect 1809 100827 1843 100861
rect 136955 100827 136989 100861
rect 1809 100491 1843 100525
rect 136955 100491 136989 100525
rect 1809 100155 1843 100189
rect 136955 100155 136989 100189
rect 1809 99819 1843 99853
rect 136955 99819 136989 99853
rect 1809 99483 1843 99517
rect 136955 99483 136989 99517
rect 1809 99147 1843 99181
rect 136955 99147 136989 99181
rect 1809 98811 1843 98845
rect 136955 98811 136989 98845
rect 1809 98475 1843 98509
rect 136955 98475 136989 98509
rect 1809 98139 1843 98173
rect 136955 98139 136989 98173
rect 1809 97803 1843 97837
rect 136955 97803 136989 97837
rect 1809 97467 1843 97501
rect 136955 97467 136989 97501
rect 1809 97131 1843 97165
rect 136955 97131 136989 97165
rect 1809 96795 1843 96829
rect 136955 96795 136989 96829
rect 1809 96459 1843 96493
rect 136955 96459 136989 96493
rect 1809 96123 1843 96157
rect 136955 96123 136989 96157
rect 1809 95787 1843 95821
rect 136955 95787 136989 95821
rect 1809 95451 1843 95485
rect 136955 95451 136989 95485
rect 1809 95115 1843 95149
rect 136955 95115 136989 95149
rect 1809 94779 1843 94813
rect 136955 94779 136989 94813
rect 1809 94443 1843 94477
rect 136955 94443 136989 94477
rect 1809 94107 1843 94141
rect 136955 94107 136989 94141
rect 1809 93771 1843 93805
rect 136955 93771 136989 93805
rect 1809 93435 1843 93469
rect 136955 93435 136989 93469
rect 1809 93099 1843 93133
rect 136955 93099 136989 93133
rect 1809 92763 1843 92797
rect 136955 92763 136989 92797
rect 1809 92427 1843 92461
rect 136955 92427 136989 92461
rect 1809 92091 1843 92125
rect 136955 92091 136989 92125
rect 1809 91755 1843 91789
rect 136955 91755 136989 91789
rect 1809 91419 1843 91453
rect 136955 91419 136989 91453
rect 1809 91083 1843 91117
rect 136955 91083 136989 91117
rect 1809 90747 1843 90781
rect 136955 90747 136989 90781
rect 1809 90411 1843 90445
rect 136955 90411 136989 90445
rect 1809 90075 1843 90109
rect 136955 90075 136989 90109
rect 1809 89739 1843 89773
rect 136955 89739 136989 89773
rect 1809 89403 1843 89437
rect 136955 89403 136989 89437
rect 1809 89067 1843 89101
rect 136955 89067 136989 89101
rect 1809 88731 1843 88765
rect 136955 88731 136989 88765
rect 1809 88395 1843 88429
rect 136955 88395 136989 88429
rect 1809 88059 1843 88093
rect 136955 88059 136989 88093
rect 1809 87723 1843 87757
rect 136955 87723 136989 87757
rect 1809 87387 1843 87421
rect 136955 87387 136989 87421
rect 1809 87051 1843 87085
rect 136955 87051 136989 87085
rect 1809 86715 1843 86749
rect 136955 86715 136989 86749
rect 1809 86379 1843 86413
rect 136955 86379 136989 86413
rect 1809 86043 1843 86077
rect 136955 86043 136989 86077
rect 1809 85707 1843 85741
rect 136955 85707 136989 85741
rect 1809 85371 1843 85405
rect 136955 85371 136989 85405
rect 1809 85035 1843 85069
rect 136955 85035 136989 85069
rect 1809 84699 1843 84733
rect 136955 84699 136989 84733
rect 1809 84363 1843 84397
rect 136955 84363 136989 84397
rect 1809 84027 1843 84061
rect 136955 84027 136989 84061
rect 1809 83691 1843 83725
rect 136955 83691 136989 83725
rect 1809 83355 1843 83389
rect 136955 83355 136989 83389
rect 1809 83019 1843 83053
rect 136955 83019 136989 83053
rect 1809 82683 1843 82717
rect 136955 82683 136989 82717
rect 1809 82347 1843 82381
rect 136955 82347 136989 82381
rect 1809 82011 1843 82045
rect 136955 82011 136989 82045
rect 1809 81675 1843 81709
rect 136955 81675 136989 81709
rect 1809 81339 1843 81373
rect 136955 81339 136989 81373
rect 1809 81003 1843 81037
rect 136955 81003 136989 81037
rect 1809 80667 1843 80701
rect 136955 80667 136989 80701
rect 1809 80331 1843 80365
rect 136955 80331 136989 80365
rect 1809 79995 1843 80029
rect 136955 79995 136989 80029
rect 1809 79659 1843 79693
rect 136955 79659 136989 79693
rect 1809 79323 1843 79357
rect 136955 79323 136989 79357
rect 1809 78987 1843 79021
rect 136955 78987 136989 79021
rect 1809 78651 1843 78685
rect 136955 78651 136989 78685
rect 1809 78315 1843 78349
rect 136955 78315 136989 78349
rect 1809 77979 1843 78013
rect 136955 77979 136989 78013
rect 1809 77643 1843 77677
rect 136955 77643 136989 77677
rect 1809 77307 1843 77341
rect 136955 77307 136989 77341
rect 1809 76971 1843 77005
rect 136955 76971 136989 77005
rect 1809 76635 1843 76669
rect 136955 76635 136989 76669
rect 1809 76299 1843 76333
rect 136955 76299 136989 76333
rect 1809 75963 1843 75997
rect 136955 75963 136989 75997
rect 1809 75627 1843 75661
rect 136955 75627 136989 75661
rect 1809 75291 1843 75325
rect 136955 75291 136989 75325
rect 1809 74955 1843 74989
rect 136955 74955 136989 74989
rect 1809 74619 1843 74653
rect 136955 74619 136989 74653
rect 1809 74283 1843 74317
rect 136955 74283 136989 74317
rect 1809 73947 1843 73981
rect 136955 73947 136989 73981
rect 1809 73611 1843 73645
rect 136955 73611 136989 73645
rect 1809 73275 1843 73309
rect 136955 73275 136989 73309
rect 1809 72939 1843 72973
rect 136955 72939 136989 72973
rect 1809 72603 1843 72637
rect 136955 72603 136989 72637
rect 1809 72267 1843 72301
rect 136955 72267 136989 72301
rect 1809 71931 1843 71965
rect 136955 71931 136989 71965
rect 1809 71595 1843 71629
rect 136955 71595 136989 71629
rect 1809 71259 1843 71293
rect 136955 71259 136989 71293
rect 1809 70923 1843 70957
rect 136955 70923 136989 70957
rect 1809 70587 1843 70621
rect 136955 70587 136989 70621
rect 1809 70251 1843 70285
rect 136955 70251 136989 70285
rect 1809 69915 1843 69949
rect 136955 69915 136989 69949
rect 1809 69579 1843 69613
rect 136955 69579 136989 69613
rect 1809 69243 1843 69277
rect 136955 69243 136989 69277
rect 1809 68907 1843 68941
rect 136955 68907 136989 68941
rect 1809 68571 1843 68605
rect 136955 68571 136989 68605
rect 1809 68235 1843 68269
rect 136955 68235 136989 68269
rect 1809 67899 1843 67933
rect 136955 67899 136989 67933
rect 1809 67563 1843 67597
rect 136955 67563 136989 67597
rect 1809 67227 1843 67261
rect 136955 67227 136989 67261
rect 1809 66891 1843 66925
rect 136955 66891 136989 66925
rect 1809 66555 1843 66589
rect 136955 66555 136989 66589
rect 1809 66219 1843 66253
rect 136955 66219 136989 66253
rect 1809 65883 1843 65917
rect 136955 65883 136989 65917
rect 1809 65547 1843 65581
rect 136955 65547 136989 65581
rect 1809 65211 1843 65245
rect 136955 65211 136989 65245
rect 1809 64875 1843 64909
rect 136955 64875 136989 64909
rect 1809 64539 1843 64573
rect 136955 64539 136989 64573
rect 1809 64203 1843 64237
rect 136955 64203 136989 64237
rect 1809 63867 1843 63901
rect 136955 63867 136989 63901
rect 1809 63531 1843 63565
rect 136955 63531 136989 63565
rect 1809 63195 1843 63229
rect 136955 63195 136989 63229
rect 1809 62859 1843 62893
rect 136955 62859 136989 62893
rect 1809 62523 1843 62557
rect 136955 62523 136989 62557
rect 1809 62187 1843 62221
rect 136955 62187 136989 62221
rect 1809 61851 1843 61885
rect 136955 61851 136989 61885
rect 1809 61515 1843 61549
rect 136955 61515 136989 61549
rect 1809 61179 1843 61213
rect 136955 61179 136989 61213
rect 1809 60843 1843 60877
rect 136955 60843 136989 60877
rect 1809 60507 1843 60541
rect 136955 60507 136989 60541
rect 1809 60171 1843 60205
rect 136955 60171 136989 60205
rect 1809 59835 1843 59869
rect 136955 59835 136989 59869
rect 1809 59499 1843 59533
rect 136955 59499 136989 59533
rect 1809 59163 1843 59197
rect 136955 59163 136989 59197
rect 1809 58827 1843 58861
rect 136955 58827 136989 58861
rect 1809 58491 1843 58525
rect 136955 58491 136989 58525
rect 1809 58155 1843 58189
rect 136955 58155 136989 58189
rect 1809 57819 1843 57853
rect 136955 57819 136989 57853
rect 1809 57483 1843 57517
rect 136955 57483 136989 57517
rect 1809 57147 1843 57181
rect 136955 57147 136989 57181
rect 1809 56811 1843 56845
rect 136955 56811 136989 56845
rect 1809 56475 1843 56509
rect 136955 56475 136989 56509
rect 1809 56139 1843 56173
rect 136955 56139 136989 56173
rect 1809 55803 1843 55837
rect 136955 55803 136989 55837
rect 1809 55467 1843 55501
rect 136955 55467 136989 55501
rect 1809 55131 1843 55165
rect 136955 55131 136989 55165
rect 1809 54795 1843 54829
rect 136955 54795 136989 54829
rect 1809 54459 1843 54493
rect 136955 54459 136989 54493
rect 1809 54123 1843 54157
rect 136955 54123 136989 54157
rect 1809 53787 1843 53821
rect 136955 53787 136989 53821
rect 1809 53451 1843 53485
rect 136955 53451 136989 53485
rect 1809 53115 1843 53149
rect 136955 53115 136989 53149
rect 1809 52779 1843 52813
rect 136955 52779 136989 52813
rect 1809 52443 1843 52477
rect 136955 52443 136989 52477
rect 1809 52107 1843 52141
rect 136955 52107 136989 52141
rect 1809 51771 1843 51805
rect 136955 51771 136989 51805
rect 1809 51435 1843 51469
rect 136955 51435 136989 51469
rect 1809 51099 1843 51133
rect 136955 51099 136989 51133
rect 1809 50763 1843 50797
rect 136955 50763 136989 50797
rect 1809 50427 1843 50461
rect 136955 50427 136989 50461
rect 1809 50091 1843 50125
rect 136955 50091 136989 50125
rect 1809 49755 1843 49789
rect 136955 49755 136989 49789
rect 1809 49419 1843 49453
rect 136955 49419 136989 49453
rect 1809 49083 1843 49117
rect 136955 49083 136989 49117
rect 1809 48747 1843 48781
rect 136955 48747 136989 48781
rect 1809 48411 1843 48445
rect 136955 48411 136989 48445
rect 1809 48075 1843 48109
rect 136955 48075 136989 48109
rect 1809 47739 1843 47773
rect 136955 47739 136989 47773
rect 1809 47403 1843 47437
rect 136955 47403 136989 47437
rect 1809 47067 1843 47101
rect 136955 47067 136989 47101
rect 1809 46731 1843 46765
rect 136955 46731 136989 46765
rect 1809 46395 1843 46429
rect 136955 46395 136989 46429
rect 1809 46059 1843 46093
rect 136955 46059 136989 46093
rect 1809 45723 1843 45757
rect 136955 45723 136989 45757
rect 1809 45387 1843 45421
rect 136955 45387 136989 45421
rect 1809 45051 1843 45085
rect 136955 45051 136989 45085
rect 1809 44715 1843 44749
rect 136955 44715 136989 44749
rect 1809 44379 1843 44413
rect 136955 44379 136989 44413
rect 1809 44043 1843 44077
rect 136955 44043 136989 44077
rect 1809 43707 1843 43741
rect 136955 43707 136989 43741
rect 1809 43371 1843 43405
rect 136955 43371 136989 43405
rect 1809 43035 1843 43069
rect 136955 43035 136989 43069
rect 1809 42699 1843 42733
rect 136955 42699 136989 42733
rect 1809 42363 1843 42397
rect 136955 42363 136989 42397
rect 1809 42027 1843 42061
rect 136955 42027 136989 42061
rect 1809 41691 1843 41725
rect 136955 41691 136989 41725
rect 1809 41355 1843 41389
rect 136955 41355 136989 41389
rect 1809 41019 1843 41053
rect 136955 41019 136989 41053
rect 1809 40683 1843 40717
rect 136955 40683 136989 40717
rect 1809 40347 1843 40381
rect 136955 40347 136989 40381
rect 1809 40011 1843 40045
rect 136955 40011 136989 40045
rect 1809 39675 1843 39709
rect 136955 39675 136989 39709
rect 1809 39339 1843 39373
rect 136955 39339 136989 39373
rect 1809 39003 1843 39037
rect 136955 39003 136989 39037
rect 1809 38667 1843 38701
rect 136955 38667 136989 38701
rect 1809 38331 1843 38365
rect 136955 38331 136989 38365
rect 1809 37995 1843 38029
rect 136955 37995 136989 38029
rect 1809 37659 1843 37693
rect 136955 37659 136989 37693
rect 1809 37323 1843 37357
rect 136955 37323 136989 37357
rect 1809 36987 1843 37021
rect 136955 36987 136989 37021
rect 1809 36651 1843 36685
rect 136955 36651 136989 36685
rect 1809 36315 1843 36349
rect 136955 36315 136989 36349
rect 1809 35979 1843 36013
rect 136955 35979 136989 36013
rect 1809 35643 1843 35677
rect 136955 35643 136989 35677
rect 1809 35307 1843 35341
rect 136955 35307 136989 35341
rect 1809 34971 1843 35005
rect 136955 34971 136989 35005
rect 1809 34635 1843 34669
rect 136955 34635 136989 34669
rect 1809 34299 1843 34333
rect 136955 34299 136989 34333
rect 1809 33963 1843 33997
rect 136955 33963 136989 33997
rect 1809 33627 1843 33661
rect 136955 33627 136989 33661
rect 1809 33291 1843 33325
rect 136955 33291 136989 33325
rect 1809 32955 1843 32989
rect 136955 32955 136989 32989
rect 1809 32619 1843 32653
rect 136955 32619 136989 32653
rect 1809 32283 1843 32317
rect 136955 32283 136989 32317
rect 1809 31947 1843 31981
rect 136955 31947 136989 31981
rect 1809 31611 1843 31645
rect 136955 31611 136989 31645
rect 1809 31275 1843 31309
rect 136955 31275 136989 31309
rect 1809 30939 1843 30973
rect 136955 30939 136989 30973
rect 1809 30603 1843 30637
rect 136955 30603 136989 30637
rect 1809 30267 1843 30301
rect 136955 30267 136989 30301
rect 1809 29931 1843 29965
rect 136955 29931 136989 29965
rect 1809 29595 1843 29629
rect 136955 29595 136989 29629
rect 1809 29259 1843 29293
rect 136955 29259 136989 29293
rect 1809 28923 1843 28957
rect 136955 28923 136989 28957
rect 1809 28587 1843 28621
rect 136955 28587 136989 28621
rect 1809 28251 1843 28285
rect 136955 28251 136989 28285
rect 1809 27915 1843 27949
rect 136955 27915 136989 27949
rect 1809 27579 1843 27613
rect 136955 27579 136989 27613
rect 1809 27243 1843 27277
rect 136955 27243 136989 27277
rect 1809 26907 1843 26941
rect 136955 26907 136989 26941
rect 1809 26571 1843 26605
rect 136955 26571 136989 26605
rect 1809 26235 1843 26269
rect 136955 26235 136989 26269
rect 1809 25899 1843 25933
rect 136955 25899 136989 25933
rect 1809 25563 1843 25597
rect 136955 25563 136989 25597
rect 1809 25227 1843 25261
rect 136955 25227 136989 25261
rect 1809 24891 1843 24925
rect 136955 24891 136989 24925
rect 1809 24555 1843 24589
rect 136955 24555 136989 24589
rect 1809 24219 1843 24253
rect 136955 24219 136989 24253
rect 1809 23883 1843 23917
rect 136955 23883 136989 23917
rect 1809 23547 1843 23581
rect 136955 23547 136989 23581
rect 1809 23211 1843 23245
rect 136955 23211 136989 23245
rect 1809 22875 1843 22909
rect 136955 22875 136989 22909
rect 1809 22539 1843 22573
rect 136955 22539 136989 22573
rect 1809 22203 1843 22237
rect 136955 22203 136989 22237
rect 1809 21867 1843 21901
rect 136955 21867 136989 21901
rect 1809 21531 1843 21565
rect 136955 21531 136989 21565
rect 1809 21195 1843 21229
rect 136955 21195 136989 21229
rect 1809 20859 1843 20893
rect 136955 20859 136989 20893
rect 1809 20523 1843 20557
rect 136955 20523 136989 20557
rect 1809 20187 1843 20221
rect 136955 20187 136989 20221
rect 1809 19851 1843 19885
rect 136955 19851 136989 19885
rect 1809 19515 1843 19549
rect 136955 19515 136989 19549
rect 1809 19179 1843 19213
rect 136955 19179 136989 19213
rect 1809 18843 1843 18877
rect 136955 18843 136989 18877
rect 1809 18507 1843 18541
rect 136955 18507 136989 18541
rect 1809 18171 1843 18205
rect 136955 18171 136989 18205
rect 1809 17835 1843 17869
rect 136955 17835 136989 17869
rect 1809 17499 1843 17533
rect 136955 17499 136989 17533
rect 1809 17163 1843 17197
rect 136955 17163 136989 17197
rect 1809 16827 1843 16861
rect 136955 16827 136989 16861
rect 1809 16491 1843 16525
rect 136955 16491 136989 16525
rect 1809 16155 1843 16189
rect 136955 16155 136989 16189
rect 1809 15819 1843 15853
rect 136955 15819 136989 15853
rect 1809 15483 1843 15517
rect 136955 15483 136989 15517
rect 1809 15147 1843 15181
rect 136955 15147 136989 15181
rect 1809 14811 1843 14845
rect 136955 14811 136989 14845
rect 1809 14475 1843 14509
rect 136955 14475 136989 14509
rect 1809 14139 1843 14173
rect 136955 14139 136989 14173
rect 1809 13803 1843 13837
rect 136955 13803 136989 13837
rect 1809 13467 1843 13501
rect 136955 13467 136989 13501
rect 1809 13131 1843 13165
rect 136955 13131 136989 13165
rect 1809 12795 1843 12829
rect 136955 12795 136989 12829
rect 1809 12459 1843 12493
rect 136955 12459 136989 12493
rect 1809 12123 1843 12157
rect 136955 12123 136989 12157
rect 1809 11787 1843 11821
rect 136955 11787 136989 11821
rect 1809 11451 1843 11485
rect 136955 11451 136989 11485
rect 1809 11115 1843 11149
rect 136955 11115 136989 11149
rect 1809 10779 1843 10813
rect 136955 10779 136989 10813
rect 1809 10443 1843 10477
rect 136955 10443 136989 10477
rect 1809 10107 1843 10141
rect 136955 10107 136989 10141
rect 1809 9771 1843 9805
rect 136955 9771 136989 9805
rect 1809 9435 1843 9469
rect 136955 9435 136989 9469
rect 1809 9099 1843 9133
rect 136955 9099 136989 9133
rect 1809 8763 1843 8797
rect 136955 8763 136989 8797
rect 1809 8427 1843 8461
rect 136955 8427 136989 8461
rect 1809 8091 1843 8125
rect 136955 8091 136989 8125
rect 1809 7755 1843 7789
rect 136955 7755 136989 7789
rect 1809 7419 1843 7453
rect 136955 7419 136989 7453
rect 1809 7083 1843 7117
rect 136955 7083 136989 7117
rect 1809 6747 1843 6781
rect 136955 6747 136989 6781
rect 1809 6411 1843 6445
rect 136955 6411 136989 6445
rect 1809 6075 1843 6109
rect 136955 6075 136989 6109
rect 1809 5739 1843 5773
rect 136955 5739 136989 5773
rect 1809 5403 1843 5437
rect 136955 5403 136989 5437
rect 1809 5067 1843 5101
rect 136955 5067 136989 5101
rect 1809 4731 1843 4765
rect 136955 4731 136989 4765
rect 1809 4395 1843 4429
rect 136955 4395 136989 4429
rect 1809 4059 1843 4093
rect 136955 4059 136989 4093
rect 1809 3723 1843 3757
rect 136955 3723 136989 3757
rect 1809 3387 1843 3421
rect 136955 3387 136989 3421
rect 1809 3051 1843 3085
rect 136955 3051 136989 3085
rect 1809 2715 1843 2749
rect 136955 2715 136989 2749
rect 1809 2379 1843 2413
rect 136955 2379 136989 2413
rect 1809 2043 1843 2077
rect 136955 2043 136989 2077
rect 2145 1707 2179 1741
rect 2481 1707 2515 1741
rect 2817 1707 2851 1741
rect 3153 1707 3187 1741
rect 3489 1707 3523 1741
rect 3825 1707 3859 1741
rect 4161 1707 4195 1741
rect 4497 1707 4531 1741
rect 4833 1707 4867 1741
rect 5169 1707 5203 1741
rect 5505 1707 5539 1741
rect 5841 1707 5875 1741
rect 6177 1707 6211 1741
rect 6513 1707 6547 1741
rect 6849 1707 6883 1741
rect 7185 1707 7219 1741
rect 7521 1707 7555 1741
rect 7857 1707 7891 1741
rect 8193 1707 8227 1741
rect 8529 1707 8563 1741
rect 8865 1707 8899 1741
rect 9201 1707 9235 1741
rect 9537 1707 9571 1741
rect 9873 1707 9907 1741
rect 10209 1707 10243 1741
rect 10545 1707 10579 1741
rect 10881 1707 10915 1741
rect 11217 1707 11251 1741
rect 11553 1707 11587 1741
rect 11889 1707 11923 1741
rect 12225 1707 12259 1741
rect 12561 1707 12595 1741
rect 12897 1707 12931 1741
rect 13233 1707 13267 1741
rect 13569 1707 13603 1741
rect 13905 1707 13939 1741
rect 14241 1707 14275 1741
rect 14577 1707 14611 1741
rect 14913 1707 14947 1741
rect 15249 1707 15283 1741
rect 15585 1707 15619 1741
rect 15921 1707 15955 1741
rect 16257 1707 16291 1741
rect 16593 1707 16627 1741
rect 16929 1707 16963 1741
rect 17265 1707 17299 1741
rect 17601 1707 17635 1741
rect 17937 1707 17971 1741
rect 18273 1707 18307 1741
rect 18609 1707 18643 1741
rect 18945 1707 18979 1741
rect 19281 1707 19315 1741
rect 19617 1707 19651 1741
rect 19953 1707 19987 1741
rect 20289 1707 20323 1741
rect 20625 1707 20659 1741
rect 20961 1707 20995 1741
rect 21297 1707 21331 1741
rect 21633 1707 21667 1741
rect 21969 1707 22003 1741
rect 22305 1707 22339 1741
rect 22641 1707 22675 1741
rect 22977 1707 23011 1741
rect 23313 1707 23347 1741
rect 23649 1707 23683 1741
rect 23985 1707 24019 1741
rect 24321 1707 24355 1741
rect 24657 1707 24691 1741
rect 24993 1707 25027 1741
rect 25329 1707 25363 1741
rect 25665 1707 25699 1741
rect 26001 1707 26035 1741
rect 26337 1707 26371 1741
rect 26673 1707 26707 1741
rect 27009 1707 27043 1741
rect 27345 1707 27379 1741
rect 27681 1707 27715 1741
rect 28017 1707 28051 1741
rect 28353 1707 28387 1741
rect 28689 1707 28723 1741
rect 29025 1707 29059 1741
rect 29361 1707 29395 1741
rect 29697 1707 29731 1741
rect 30033 1707 30067 1741
rect 30369 1707 30403 1741
rect 30705 1707 30739 1741
rect 31041 1707 31075 1741
rect 31377 1707 31411 1741
rect 31713 1707 31747 1741
rect 32049 1707 32083 1741
rect 32385 1707 32419 1741
rect 32721 1707 32755 1741
rect 33057 1707 33091 1741
rect 33393 1707 33427 1741
rect 33729 1707 33763 1741
rect 34065 1707 34099 1741
rect 34401 1707 34435 1741
rect 34737 1707 34771 1741
rect 35073 1707 35107 1741
rect 35409 1707 35443 1741
rect 35745 1707 35779 1741
rect 36081 1707 36115 1741
rect 36417 1707 36451 1741
rect 36753 1707 36787 1741
rect 37089 1707 37123 1741
rect 37425 1707 37459 1741
rect 37761 1707 37795 1741
rect 38097 1707 38131 1741
rect 38433 1707 38467 1741
rect 38769 1707 38803 1741
rect 39105 1707 39139 1741
rect 39441 1707 39475 1741
rect 39777 1707 39811 1741
rect 40113 1707 40147 1741
rect 40449 1707 40483 1741
rect 40785 1707 40819 1741
rect 41121 1707 41155 1741
rect 41457 1707 41491 1741
rect 41793 1707 41827 1741
rect 42129 1707 42163 1741
rect 42465 1707 42499 1741
rect 42801 1707 42835 1741
rect 43137 1707 43171 1741
rect 43473 1707 43507 1741
rect 43809 1707 43843 1741
rect 44145 1707 44179 1741
rect 44481 1707 44515 1741
rect 44817 1707 44851 1741
rect 45153 1707 45187 1741
rect 45489 1707 45523 1741
rect 45825 1707 45859 1741
rect 46161 1707 46195 1741
rect 46497 1707 46531 1741
rect 46833 1707 46867 1741
rect 47169 1707 47203 1741
rect 47505 1707 47539 1741
rect 47841 1707 47875 1741
rect 48177 1707 48211 1741
rect 48513 1707 48547 1741
rect 48849 1707 48883 1741
rect 49185 1707 49219 1741
rect 49521 1707 49555 1741
rect 49857 1707 49891 1741
rect 50193 1707 50227 1741
rect 50529 1707 50563 1741
rect 50865 1707 50899 1741
rect 51201 1707 51235 1741
rect 51537 1707 51571 1741
rect 51873 1707 51907 1741
rect 52209 1707 52243 1741
rect 52545 1707 52579 1741
rect 52881 1707 52915 1741
rect 53217 1707 53251 1741
rect 53553 1707 53587 1741
rect 53889 1707 53923 1741
rect 54225 1707 54259 1741
rect 54561 1707 54595 1741
rect 54897 1707 54931 1741
rect 55233 1707 55267 1741
rect 55569 1707 55603 1741
rect 55905 1707 55939 1741
rect 56241 1707 56275 1741
rect 56577 1707 56611 1741
rect 56913 1707 56947 1741
rect 57249 1707 57283 1741
rect 57585 1707 57619 1741
rect 57921 1707 57955 1741
rect 58257 1707 58291 1741
rect 58593 1707 58627 1741
rect 58929 1707 58963 1741
rect 59265 1707 59299 1741
rect 59601 1707 59635 1741
rect 59937 1707 59971 1741
rect 60273 1707 60307 1741
rect 60609 1707 60643 1741
rect 60945 1707 60979 1741
rect 61281 1707 61315 1741
rect 61617 1707 61651 1741
rect 61953 1707 61987 1741
rect 62289 1707 62323 1741
rect 62625 1707 62659 1741
rect 62961 1707 62995 1741
rect 63297 1707 63331 1741
rect 63633 1707 63667 1741
rect 63969 1707 64003 1741
rect 64305 1707 64339 1741
rect 64641 1707 64675 1741
rect 64977 1707 65011 1741
rect 65313 1707 65347 1741
rect 65649 1707 65683 1741
rect 65985 1707 66019 1741
rect 66321 1707 66355 1741
rect 66657 1707 66691 1741
rect 66993 1707 67027 1741
rect 67329 1707 67363 1741
rect 67665 1707 67699 1741
rect 68001 1707 68035 1741
rect 68337 1707 68371 1741
rect 68673 1707 68707 1741
rect 69009 1707 69043 1741
rect 69345 1707 69379 1741
rect 69681 1707 69715 1741
rect 70017 1707 70051 1741
rect 70353 1707 70387 1741
rect 70689 1707 70723 1741
rect 71025 1707 71059 1741
rect 71361 1707 71395 1741
rect 71697 1707 71731 1741
rect 72033 1707 72067 1741
rect 72369 1707 72403 1741
rect 72705 1707 72739 1741
rect 73041 1707 73075 1741
rect 73377 1707 73411 1741
rect 73713 1707 73747 1741
rect 74049 1707 74083 1741
rect 74385 1707 74419 1741
rect 74721 1707 74755 1741
rect 75057 1707 75091 1741
rect 75393 1707 75427 1741
rect 75729 1707 75763 1741
rect 76065 1707 76099 1741
rect 76401 1707 76435 1741
rect 76737 1707 76771 1741
rect 77073 1707 77107 1741
rect 77409 1707 77443 1741
rect 77745 1707 77779 1741
rect 78081 1707 78115 1741
rect 78417 1707 78451 1741
rect 78753 1707 78787 1741
rect 79089 1707 79123 1741
rect 79425 1707 79459 1741
rect 79761 1707 79795 1741
rect 80097 1707 80131 1741
rect 80433 1707 80467 1741
rect 80769 1707 80803 1741
rect 81105 1707 81139 1741
rect 81441 1707 81475 1741
rect 81777 1707 81811 1741
rect 82113 1707 82147 1741
rect 82449 1707 82483 1741
rect 82785 1707 82819 1741
rect 83121 1707 83155 1741
rect 83457 1707 83491 1741
rect 83793 1707 83827 1741
rect 84129 1707 84163 1741
rect 84465 1707 84499 1741
rect 84801 1707 84835 1741
rect 85137 1707 85171 1741
rect 85473 1707 85507 1741
rect 85809 1707 85843 1741
rect 86145 1707 86179 1741
rect 86481 1707 86515 1741
rect 86817 1707 86851 1741
rect 87153 1707 87187 1741
rect 87489 1707 87523 1741
rect 87825 1707 87859 1741
rect 88161 1707 88195 1741
rect 88497 1707 88531 1741
rect 88833 1707 88867 1741
rect 89169 1707 89203 1741
rect 89505 1707 89539 1741
rect 89841 1707 89875 1741
rect 90177 1707 90211 1741
rect 90513 1707 90547 1741
rect 90849 1707 90883 1741
rect 91185 1707 91219 1741
rect 91521 1707 91555 1741
rect 91857 1707 91891 1741
rect 92193 1707 92227 1741
rect 92529 1707 92563 1741
rect 92865 1707 92899 1741
rect 93201 1707 93235 1741
rect 93537 1707 93571 1741
rect 93873 1707 93907 1741
rect 94209 1707 94243 1741
rect 94545 1707 94579 1741
rect 94881 1707 94915 1741
rect 95217 1707 95251 1741
rect 95553 1707 95587 1741
rect 95889 1707 95923 1741
rect 96225 1707 96259 1741
rect 96561 1707 96595 1741
rect 96897 1707 96931 1741
rect 97233 1707 97267 1741
rect 97569 1707 97603 1741
rect 97905 1707 97939 1741
rect 98241 1707 98275 1741
rect 98577 1707 98611 1741
rect 98913 1707 98947 1741
rect 99249 1707 99283 1741
rect 99585 1707 99619 1741
rect 99921 1707 99955 1741
rect 100257 1707 100291 1741
rect 100593 1707 100627 1741
rect 100929 1707 100963 1741
rect 101265 1707 101299 1741
rect 101601 1707 101635 1741
rect 101937 1707 101971 1741
rect 102273 1707 102307 1741
rect 102609 1707 102643 1741
rect 102945 1707 102979 1741
rect 103281 1707 103315 1741
rect 103617 1707 103651 1741
rect 103953 1707 103987 1741
rect 104289 1707 104323 1741
rect 104625 1707 104659 1741
rect 104961 1707 104995 1741
rect 105297 1707 105331 1741
rect 105633 1707 105667 1741
rect 105969 1707 106003 1741
rect 106305 1707 106339 1741
rect 106641 1707 106675 1741
rect 106977 1707 107011 1741
rect 107313 1707 107347 1741
rect 107649 1707 107683 1741
rect 107985 1707 108019 1741
rect 108321 1707 108355 1741
rect 108657 1707 108691 1741
rect 108993 1707 109027 1741
rect 109329 1707 109363 1741
rect 109665 1707 109699 1741
rect 110001 1707 110035 1741
rect 110337 1707 110371 1741
rect 110673 1707 110707 1741
rect 111009 1707 111043 1741
rect 111345 1707 111379 1741
rect 111681 1707 111715 1741
rect 112017 1707 112051 1741
rect 112353 1707 112387 1741
rect 112689 1707 112723 1741
rect 113025 1707 113059 1741
rect 113361 1707 113395 1741
rect 113697 1707 113731 1741
rect 114033 1707 114067 1741
rect 114369 1707 114403 1741
rect 114705 1707 114739 1741
rect 115041 1707 115075 1741
rect 115377 1707 115411 1741
rect 115713 1707 115747 1741
rect 116049 1707 116083 1741
rect 116385 1707 116419 1741
rect 116721 1707 116755 1741
rect 117057 1707 117091 1741
rect 117393 1707 117427 1741
rect 117729 1707 117763 1741
rect 118065 1707 118099 1741
rect 118401 1707 118435 1741
rect 118737 1707 118771 1741
rect 119073 1707 119107 1741
rect 119409 1707 119443 1741
rect 119745 1707 119779 1741
rect 120081 1707 120115 1741
rect 120417 1707 120451 1741
rect 120753 1707 120787 1741
rect 121089 1707 121123 1741
rect 121425 1707 121459 1741
rect 121761 1707 121795 1741
rect 122097 1707 122131 1741
rect 122433 1707 122467 1741
rect 122769 1707 122803 1741
rect 123105 1707 123139 1741
rect 123441 1707 123475 1741
rect 123777 1707 123811 1741
rect 124113 1707 124147 1741
rect 124449 1707 124483 1741
rect 124785 1707 124819 1741
rect 125121 1707 125155 1741
rect 125457 1707 125491 1741
rect 125793 1707 125827 1741
rect 126129 1707 126163 1741
rect 126465 1707 126499 1741
rect 126801 1707 126835 1741
rect 127137 1707 127171 1741
rect 127473 1707 127507 1741
rect 127809 1707 127843 1741
rect 128145 1707 128179 1741
rect 128481 1707 128515 1741
rect 128817 1707 128851 1741
rect 129153 1707 129187 1741
rect 129489 1707 129523 1741
rect 129825 1707 129859 1741
rect 130161 1707 130195 1741
rect 130497 1707 130531 1741
rect 130833 1707 130867 1741
rect 131169 1707 131203 1741
rect 131505 1707 131539 1741
rect 131841 1707 131875 1741
rect 132177 1707 132211 1741
rect 132513 1707 132547 1741
rect 132849 1707 132883 1741
rect 133185 1707 133219 1741
rect 133521 1707 133555 1741
rect 133857 1707 133891 1741
rect 134193 1707 134227 1741
rect 134529 1707 134563 1741
rect 134865 1707 134899 1741
rect 135201 1707 135235 1741
rect 135537 1707 135571 1741
rect 135873 1707 135907 1741
rect 136209 1707 136243 1741
rect 136545 1707 136579 1741
<< metal1 >>
rect 1714 132059 137084 132145
rect 1714 132007 2136 132059
rect 2188 132050 3816 132059
rect 3868 132050 5496 132059
rect 5548 132050 7176 132059
rect 7228 132050 8856 132059
rect 8908 132050 10536 132059
rect 10588 132050 12216 132059
rect 12268 132050 13896 132059
rect 13948 132050 15576 132059
rect 15628 132050 17256 132059
rect 17308 132050 18936 132059
rect 18988 132050 20616 132059
rect 20668 132050 22296 132059
rect 22348 132050 23976 132059
rect 24028 132050 25656 132059
rect 25708 132050 27336 132059
rect 27388 132050 29016 132059
rect 29068 132050 30696 132059
rect 30748 132050 32376 132059
rect 32428 132050 34056 132059
rect 34108 132050 35736 132059
rect 35788 132050 37416 132059
rect 37468 132050 39096 132059
rect 39148 132050 40776 132059
rect 40828 132050 42456 132059
rect 42508 132050 44136 132059
rect 44188 132050 45816 132059
rect 45868 132050 47496 132059
rect 47548 132050 49176 132059
rect 49228 132050 50856 132059
rect 50908 132050 52536 132059
rect 52588 132050 54216 132059
rect 54268 132050 55896 132059
rect 55948 132050 57576 132059
rect 57628 132050 59256 132059
rect 59308 132050 60936 132059
rect 60988 132050 62616 132059
rect 62668 132050 64296 132059
rect 64348 132050 65976 132059
rect 66028 132050 67656 132059
rect 67708 132050 69336 132059
rect 69388 132050 71016 132059
rect 71068 132050 72696 132059
rect 72748 132050 74376 132059
rect 74428 132050 76056 132059
rect 76108 132050 77736 132059
rect 77788 132050 79416 132059
rect 79468 132050 81096 132059
rect 81148 132050 82776 132059
rect 82828 132050 84456 132059
rect 84508 132050 86136 132059
rect 86188 132050 87816 132059
rect 87868 132050 89496 132059
rect 89548 132050 91176 132059
rect 91228 132050 92856 132059
rect 92908 132050 94536 132059
rect 94588 132050 96216 132059
rect 96268 132050 97896 132059
rect 97948 132050 99576 132059
rect 99628 132050 101256 132059
rect 101308 132050 102936 132059
rect 102988 132050 104616 132059
rect 104668 132050 106296 132059
rect 106348 132050 107976 132059
rect 108028 132050 109656 132059
rect 109708 132050 111336 132059
rect 111388 132050 113016 132059
rect 113068 132050 114696 132059
rect 114748 132050 116376 132059
rect 116428 132050 118056 132059
rect 118108 132050 119736 132059
rect 119788 132050 121416 132059
rect 121468 132050 123096 132059
rect 123148 132050 124776 132059
rect 124828 132050 126456 132059
rect 126508 132050 128136 132059
rect 128188 132050 129816 132059
rect 129868 132050 131496 132059
rect 131548 132050 133176 132059
rect 133228 132050 134856 132059
rect 134908 132050 136536 132059
rect 2188 132016 2481 132050
rect 2515 132016 2817 132050
rect 2851 132016 3153 132050
rect 3187 132016 3489 132050
rect 3523 132016 3816 132050
rect 3868 132016 4161 132050
rect 4195 132016 4497 132050
rect 4531 132016 4833 132050
rect 4867 132016 5169 132050
rect 5203 132016 5496 132050
rect 5548 132016 5841 132050
rect 5875 132016 6177 132050
rect 6211 132016 6513 132050
rect 6547 132016 6849 132050
rect 6883 132016 7176 132050
rect 7228 132016 7521 132050
rect 7555 132016 7857 132050
rect 7891 132016 8193 132050
rect 8227 132016 8529 132050
rect 8563 132016 8856 132050
rect 8908 132016 9201 132050
rect 9235 132016 9537 132050
rect 9571 132016 9873 132050
rect 9907 132016 10209 132050
rect 10243 132016 10536 132050
rect 10588 132016 10881 132050
rect 10915 132016 11217 132050
rect 11251 132016 11553 132050
rect 11587 132016 11889 132050
rect 11923 132016 12216 132050
rect 12268 132016 12561 132050
rect 12595 132016 12897 132050
rect 12931 132016 13233 132050
rect 13267 132016 13569 132050
rect 13603 132016 13896 132050
rect 13948 132016 14241 132050
rect 14275 132016 14577 132050
rect 14611 132016 14913 132050
rect 14947 132016 15249 132050
rect 15283 132016 15576 132050
rect 15628 132016 15921 132050
rect 15955 132016 16257 132050
rect 16291 132016 16593 132050
rect 16627 132016 16929 132050
rect 16963 132016 17256 132050
rect 17308 132016 17601 132050
rect 17635 132016 17937 132050
rect 17971 132016 18273 132050
rect 18307 132016 18609 132050
rect 18643 132016 18936 132050
rect 18988 132016 19281 132050
rect 19315 132016 19617 132050
rect 19651 132016 19953 132050
rect 19987 132016 20289 132050
rect 20323 132016 20616 132050
rect 20668 132016 20961 132050
rect 20995 132016 21297 132050
rect 21331 132016 21633 132050
rect 21667 132016 21969 132050
rect 22003 132016 22296 132050
rect 22348 132016 22641 132050
rect 22675 132016 22977 132050
rect 23011 132016 23313 132050
rect 23347 132016 23649 132050
rect 23683 132016 23976 132050
rect 24028 132016 24321 132050
rect 24355 132016 24657 132050
rect 24691 132016 24993 132050
rect 25027 132016 25329 132050
rect 25363 132016 25656 132050
rect 25708 132016 26001 132050
rect 26035 132016 26337 132050
rect 26371 132016 26673 132050
rect 26707 132016 27009 132050
rect 27043 132016 27336 132050
rect 27388 132016 27681 132050
rect 27715 132016 28017 132050
rect 28051 132016 28353 132050
rect 28387 132016 28689 132050
rect 28723 132016 29016 132050
rect 29068 132016 29361 132050
rect 29395 132016 29697 132050
rect 29731 132016 30033 132050
rect 30067 132016 30369 132050
rect 30403 132016 30696 132050
rect 30748 132016 31041 132050
rect 31075 132016 31377 132050
rect 31411 132016 31713 132050
rect 31747 132016 32049 132050
rect 32083 132016 32376 132050
rect 32428 132016 32721 132050
rect 32755 132016 33057 132050
rect 33091 132016 33393 132050
rect 33427 132016 33729 132050
rect 33763 132016 34056 132050
rect 34108 132016 34401 132050
rect 34435 132016 34737 132050
rect 34771 132016 35073 132050
rect 35107 132016 35409 132050
rect 35443 132016 35736 132050
rect 35788 132016 36081 132050
rect 36115 132016 36417 132050
rect 36451 132016 36753 132050
rect 36787 132016 37089 132050
rect 37123 132016 37416 132050
rect 37468 132016 37761 132050
rect 37795 132016 38097 132050
rect 38131 132016 38433 132050
rect 38467 132016 38769 132050
rect 38803 132016 39096 132050
rect 39148 132016 39441 132050
rect 39475 132016 39777 132050
rect 39811 132016 40113 132050
rect 40147 132016 40449 132050
rect 40483 132016 40776 132050
rect 40828 132016 41121 132050
rect 41155 132016 41457 132050
rect 41491 132016 41793 132050
rect 41827 132016 42129 132050
rect 42163 132016 42456 132050
rect 42508 132016 42801 132050
rect 42835 132016 43137 132050
rect 43171 132016 43473 132050
rect 43507 132016 43809 132050
rect 43843 132016 44136 132050
rect 44188 132016 44481 132050
rect 44515 132016 44817 132050
rect 44851 132016 45153 132050
rect 45187 132016 45489 132050
rect 45523 132016 45816 132050
rect 45868 132016 46161 132050
rect 46195 132016 46497 132050
rect 46531 132016 46833 132050
rect 46867 132016 47169 132050
rect 47203 132016 47496 132050
rect 47548 132016 47841 132050
rect 47875 132016 48177 132050
rect 48211 132016 48513 132050
rect 48547 132016 48849 132050
rect 48883 132016 49176 132050
rect 49228 132016 49521 132050
rect 49555 132016 49857 132050
rect 49891 132016 50193 132050
rect 50227 132016 50529 132050
rect 50563 132016 50856 132050
rect 50908 132016 51201 132050
rect 51235 132016 51537 132050
rect 51571 132016 51873 132050
rect 51907 132016 52209 132050
rect 52243 132016 52536 132050
rect 52588 132016 52881 132050
rect 52915 132016 53217 132050
rect 53251 132016 53553 132050
rect 53587 132016 53889 132050
rect 53923 132016 54216 132050
rect 54268 132016 54561 132050
rect 54595 132016 54897 132050
rect 54931 132016 55233 132050
rect 55267 132016 55569 132050
rect 55603 132016 55896 132050
rect 55948 132016 56241 132050
rect 56275 132016 56577 132050
rect 56611 132016 56913 132050
rect 56947 132016 57249 132050
rect 57283 132016 57576 132050
rect 57628 132016 57921 132050
rect 57955 132016 58257 132050
rect 58291 132016 58593 132050
rect 58627 132016 58929 132050
rect 58963 132016 59256 132050
rect 59308 132016 59601 132050
rect 59635 132016 59937 132050
rect 59971 132016 60273 132050
rect 60307 132016 60609 132050
rect 60643 132016 60936 132050
rect 60988 132016 61281 132050
rect 61315 132016 61617 132050
rect 61651 132016 61953 132050
rect 61987 132016 62289 132050
rect 62323 132016 62616 132050
rect 62668 132016 62961 132050
rect 62995 132016 63297 132050
rect 63331 132016 63633 132050
rect 63667 132016 63969 132050
rect 64003 132016 64296 132050
rect 64348 132016 64641 132050
rect 64675 132016 64977 132050
rect 65011 132016 65313 132050
rect 65347 132016 65649 132050
rect 65683 132016 65976 132050
rect 66028 132016 66321 132050
rect 66355 132016 66657 132050
rect 66691 132016 66993 132050
rect 67027 132016 67329 132050
rect 67363 132016 67656 132050
rect 67708 132016 68001 132050
rect 68035 132016 68337 132050
rect 68371 132016 68673 132050
rect 68707 132016 69009 132050
rect 69043 132016 69336 132050
rect 69388 132016 69681 132050
rect 69715 132016 70017 132050
rect 70051 132016 70353 132050
rect 70387 132016 70689 132050
rect 70723 132016 71016 132050
rect 71068 132016 71361 132050
rect 71395 132016 71697 132050
rect 71731 132016 72033 132050
rect 72067 132016 72369 132050
rect 72403 132016 72696 132050
rect 72748 132016 73041 132050
rect 73075 132016 73377 132050
rect 73411 132016 73713 132050
rect 73747 132016 74049 132050
rect 74083 132016 74376 132050
rect 74428 132016 74721 132050
rect 74755 132016 75057 132050
rect 75091 132016 75393 132050
rect 75427 132016 75729 132050
rect 75763 132016 76056 132050
rect 76108 132016 76401 132050
rect 76435 132016 76737 132050
rect 76771 132016 77073 132050
rect 77107 132016 77409 132050
rect 77443 132016 77736 132050
rect 77788 132016 78081 132050
rect 78115 132016 78417 132050
rect 78451 132016 78753 132050
rect 78787 132016 79089 132050
rect 79123 132016 79416 132050
rect 79468 132016 79761 132050
rect 79795 132016 80097 132050
rect 80131 132016 80433 132050
rect 80467 132016 80769 132050
rect 80803 132016 81096 132050
rect 81148 132016 81441 132050
rect 81475 132016 81777 132050
rect 81811 132016 82113 132050
rect 82147 132016 82449 132050
rect 82483 132016 82776 132050
rect 82828 132016 83121 132050
rect 83155 132016 83457 132050
rect 83491 132016 83793 132050
rect 83827 132016 84129 132050
rect 84163 132016 84456 132050
rect 84508 132016 84801 132050
rect 84835 132016 85137 132050
rect 85171 132016 85473 132050
rect 85507 132016 85809 132050
rect 85843 132016 86136 132050
rect 86188 132016 86481 132050
rect 86515 132016 86817 132050
rect 86851 132016 87153 132050
rect 87187 132016 87489 132050
rect 87523 132016 87816 132050
rect 87868 132016 88161 132050
rect 88195 132016 88497 132050
rect 88531 132016 88833 132050
rect 88867 132016 89169 132050
rect 89203 132016 89496 132050
rect 89548 132016 89841 132050
rect 89875 132016 90177 132050
rect 90211 132016 90513 132050
rect 90547 132016 90849 132050
rect 90883 132016 91176 132050
rect 91228 132016 91521 132050
rect 91555 132016 91857 132050
rect 91891 132016 92193 132050
rect 92227 132016 92529 132050
rect 92563 132016 92856 132050
rect 92908 132016 93201 132050
rect 93235 132016 93537 132050
rect 93571 132016 93873 132050
rect 93907 132016 94209 132050
rect 94243 132016 94536 132050
rect 94588 132016 94881 132050
rect 94915 132016 95217 132050
rect 95251 132016 95553 132050
rect 95587 132016 95889 132050
rect 95923 132016 96216 132050
rect 96268 132016 96561 132050
rect 96595 132016 96897 132050
rect 96931 132016 97233 132050
rect 97267 132016 97569 132050
rect 97603 132016 97896 132050
rect 97948 132016 98241 132050
rect 98275 132016 98577 132050
rect 98611 132016 98913 132050
rect 98947 132016 99249 132050
rect 99283 132016 99576 132050
rect 99628 132016 99921 132050
rect 99955 132016 100257 132050
rect 100291 132016 100593 132050
rect 100627 132016 100929 132050
rect 100963 132016 101256 132050
rect 101308 132016 101601 132050
rect 101635 132016 101937 132050
rect 101971 132016 102273 132050
rect 102307 132016 102609 132050
rect 102643 132016 102936 132050
rect 102988 132016 103281 132050
rect 103315 132016 103617 132050
rect 103651 132016 103953 132050
rect 103987 132016 104289 132050
rect 104323 132016 104616 132050
rect 104668 132016 104961 132050
rect 104995 132016 105297 132050
rect 105331 132016 105633 132050
rect 105667 132016 105969 132050
rect 106003 132016 106296 132050
rect 106348 132016 106641 132050
rect 106675 132016 106977 132050
rect 107011 132016 107313 132050
rect 107347 132016 107649 132050
rect 107683 132016 107976 132050
rect 108028 132016 108321 132050
rect 108355 132016 108657 132050
rect 108691 132016 108993 132050
rect 109027 132016 109329 132050
rect 109363 132016 109656 132050
rect 109708 132016 110001 132050
rect 110035 132016 110337 132050
rect 110371 132016 110673 132050
rect 110707 132016 111009 132050
rect 111043 132016 111336 132050
rect 111388 132016 111681 132050
rect 111715 132016 112017 132050
rect 112051 132016 112353 132050
rect 112387 132016 112689 132050
rect 112723 132016 113016 132050
rect 113068 132016 113361 132050
rect 113395 132016 113697 132050
rect 113731 132016 114033 132050
rect 114067 132016 114369 132050
rect 114403 132016 114696 132050
rect 114748 132016 115041 132050
rect 115075 132016 115377 132050
rect 115411 132016 115713 132050
rect 115747 132016 116049 132050
rect 116083 132016 116376 132050
rect 116428 132016 116721 132050
rect 116755 132016 117057 132050
rect 117091 132016 117393 132050
rect 117427 132016 117729 132050
rect 117763 132016 118056 132050
rect 118108 132016 118401 132050
rect 118435 132016 118737 132050
rect 118771 132016 119073 132050
rect 119107 132016 119409 132050
rect 119443 132016 119736 132050
rect 119788 132016 120081 132050
rect 120115 132016 120417 132050
rect 120451 132016 120753 132050
rect 120787 132016 121089 132050
rect 121123 132016 121416 132050
rect 121468 132016 121761 132050
rect 121795 132016 122097 132050
rect 122131 132016 122433 132050
rect 122467 132016 122769 132050
rect 122803 132016 123096 132050
rect 123148 132016 123441 132050
rect 123475 132016 123777 132050
rect 123811 132016 124113 132050
rect 124147 132016 124449 132050
rect 124483 132016 124776 132050
rect 124828 132016 125121 132050
rect 125155 132016 125457 132050
rect 125491 132016 125793 132050
rect 125827 132016 126129 132050
rect 126163 132016 126456 132050
rect 126508 132016 126801 132050
rect 126835 132016 127137 132050
rect 127171 132016 127473 132050
rect 127507 132016 127809 132050
rect 127843 132016 128136 132050
rect 128188 132016 128481 132050
rect 128515 132016 128817 132050
rect 128851 132016 129153 132050
rect 129187 132016 129489 132050
rect 129523 132016 129816 132050
rect 129868 132016 130161 132050
rect 130195 132016 130497 132050
rect 130531 132016 130833 132050
rect 130867 132016 131169 132050
rect 131203 132016 131496 132050
rect 131548 132016 131841 132050
rect 131875 132016 132177 132050
rect 132211 132016 132513 132050
rect 132547 132016 132849 132050
rect 132883 132016 133176 132050
rect 133228 132016 133521 132050
rect 133555 132016 133857 132050
rect 133891 132016 134193 132050
rect 134227 132016 134529 132050
rect 134563 132016 134856 132050
rect 134908 132016 135201 132050
rect 135235 132016 135537 132050
rect 135571 132016 135873 132050
rect 135907 132016 136209 132050
rect 136243 132016 136536 132050
rect 2188 132007 3816 132016
rect 3868 132007 5496 132016
rect 5548 132007 7176 132016
rect 7228 132007 8856 132016
rect 8908 132007 10536 132016
rect 10588 132007 12216 132016
rect 12268 132007 13896 132016
rect 13948 132007 15576 132016
rect 15628 132007 17256 132016
rect 17308 132007 18936 132016
rect 18988 132007 20616 132016
rect 20668 132007 22296 132016
rect 22348 132007 23976 132016
rect 24028 132007 25656 132016
rect 25708 132007 27336 132016
rect 27388 132007 29016 132016
rect 29068 132007 30696 132016
rect 30748 132007 32376 132016
rect 32428 132007 34056 132016
rect 34108 132007 35736 132016
rect 35788 132007 37416 132016
rect 37468 132007 39096 132016
rect 39148 132007 40776 132016
rect 40828 132007 42456 132016
rect 42508 132007 44136 132016
rect 44188 132007 45816 132016
rect 45868 132007 47496 132016
rect 47548 132007 49176 132016
rect 49228 132007 50856 132016
rect 50908 132007 52536 132016
rect 52588 132007 54216 132016
rect 54268 132007 55896 132016
rect 55948 132007 57576 132016
rect 57628 132007 59256 132016
rect 59308 132007 60936 132016
rect 60988 132007 62616 132016
rect 62668 132007 64296 132016
rect 64348 132007 65976 132016
rect 66028 132007 67656 132016
rect 67708 132007 69336 132016
rect 69388 132007 71016 132016
rect 71068 132007 72696 132016
rect 72748 132007 74376 132016
rect 74428 132007 76056 132016
rect 76108 132007 77736 132016
rect 77788 132007 79416 132016
rect 79468 132007 81096 132016
rect 81148 132007 82776 132016
rect 82828 132007 84456 132016
rect 84508 132007 86136 132016
rect 86188 132007 87816 132016
rect 87868 132007 89496 132016
rect 89548 132007 91176 132016
rect 91228 132007 92856 132016
rect 92908 132007 94536 132016
rect 94588 132007 96216 132016
rect 96268 132007 97896 132016
rect 97948 132007 99576 132016
rect 99628 132007 101256 132016
rect 101308 132007 102936 132016
rect 102988 132007 104616 132016
rect 104668 132007 106296 132016
rect 106348 132007 107976 132016
rect 108028 132007 109656 132016
rect 109708 132007 111336 132016
rect 111388 132007 113016 132016
rect 113068 132007 114696 132016
rect 114748 132007 116376 132016
rect 116428 132007 118056 132016
rect 118108 132007 119736 132016
rect 119788 132007 121416 132016
rect 121468 132007 123096 132016
rect 123148 132007 124776 132016
rect 124828 132007 126456 132016
rect 126508 132007 128136 132016
rect 128188 132007 129816 132016
rect 129868 132007 131496 132016
rect 131548 132007 133176 132016
rect 133228 132007 134856 132016
rect 134908 132007 136536 132016
rect 136588 132007 137084 132059
rect 1714 131921 137084 132007
rect 1794 131394 1800 131446
rect 1852 131394 1858 131446
rect 136940 131394 136946 131446
rect 136998 131394 137004 131446
rect 1794 131058 1800 131110
rect 1852 131058 1858 131110
rect 136940 131058 136946 131110
rect 136998 131058 137004 131110
rect 1794 130722 1800 130774
rect 1852 130722 1858 130774
rect 136940 130722 136946 130774
rect 136998 130722 137004 130774
rect 1794 130386 1800 130438
rect 1852 130386 1858 130438
rect 136940 130386 136946 130438
rect 136998 130386 137004 130438
rect 1794 130050 1800 130102
rect 1852 130050 1858 130102
rect 136940 130050 136946 130102
rect 136998 130050 137004 130102
rect 1794 129714 1800 129766
rect 1852 129714 1858 129766
rect 136940 129714 136946 129766
rect 136998 129714 137004 129766
rect 1794 129378 1800 129430
rect 1852 129378 1858 129430
rect 136940 129378 136946 129430
rect 136998 129378 137004 129430
rect 1794 129042 1800 129094
rect 1852 129042 1858 129094
rect 136940 129042 136946 129094
rect 136998 129042 137004 129094
rect 1794 128706 1800 128758
rect 1852 128706 1858 128758
rect 136940 128706 136946 128758
rect 136998 128706 137004 128758
rect 1794 128370 1800 128422
rect 1852 128370 1858 128422
rect 136940 128370 136946 128422
rect 136998 128370 137004 128422
rect 1794 128034 1800 128086
rect 1852 128034 1858 128086
rect 136940 128034 136946 128086
rect 136998 128034 137004 128086
rect 1794 127698 1800 127750
rect 1852 127698 1858 127750
rect 136940 127698 136946 127750
rect 136998 127698 137004 127750
rect 29558 127553 29564 127605
rect 29616 127553 29622 127605
rect 32054 127553 32060 127605
rect 32112 127553 32118 127605
rect 34550 127553 34556 127605
rect 34608 127553 34614 127605
rect 37046 127553 37052 127605
rect 37104 127553 37110 127605
rect 39542 127553 39548 127605
rect 39600 127553 39606 127605
rect 42038 127553 42044 127605
rect 42096 127553 42102 127605
rect 44534 127553 44540 127605
rect 44592 127553 44598 127605
rect 47030 127553 47036 127605
rect 47088 127553 47094 127605
rect 49526 127553 49532 127605
rect 49584 127553 49590 127605
rect 52022 127553 52028 127605
rect 52080 127553 52086 127605
rect 54518 127553 54524 127605
rect 54576 127553 54582 127605
rect 57014 127553 57020 127605
rect 57072 127553 57078 127605
rect 59510 127553 59516 127605
rect 59568 127553 59574 127605
rect 62006 127553 62012 127605
rect 62064 127553 62070 127605
rect 64502 127553 64508 127605
rect 64560 127553 64566 127605
rect 66998 127553 67004 127605
rect 67056 127553 67062 127605
rect 69494 127553 69500 127605
rect 69552 127553 69558 127605
rect 71990 127553 71996 127605
rect 72048 127553 72054 127605
rect 74486 127553 74492 127605
rect 74544 127553 74550 127605
rect 76982 127553 76988 127605
rect 77040 127553 77046 127605
rect 79478 127553 79484 127605
rect 79536 127553 79542 127605
rect 81974 127553 81980 127605
rect 82032 127553 82038 127605
rect 84470 127553 84476 127605
rect 84528 127553 84534 127605
rect 86966 127553 86972 127605
rect 87024 127553 87030 127605
rect 89462 127553 89468 127605
rect 89520 127553 89526 127605
rect 91958 127553 91964 127605
rect 92016 127553 92022 127605
rect 94454 127553 94460 127605
rect 94512 127553 94518 127605
rect 96950 127553 96956 127605
rect 97008 127553 97014 127605
rect 99446 127553 99452 127605
rect 99504 127553 99510 127605
rect 101942 127553 101948 127605
rect 102000 127553 102006 127605
rect 104438 127553 104444 127605
rect 104496 127553 104502 127605
rect 106934 127553 106940 127605
rect 106992 127553 106998 127605
rect 1794 127362 1800 127414
rect 1852 127362 1858 127414
rect 136940 127362 136946 127414
rect 136998 127362 137004 127414
rect 1794 127026 1800 127078
rect 1852 127026 1858 127078
rect 136940 127026 136946 127078
rect 136998 127026 137004 127078
rect 1794 126690 1800 126742
rect 1852 126690 1858 126742
rect 136940 126690 136946 126742
rect 136998 126690 137004 126742
rect 1794 126354 1800 126406
rect 1852 126354 1858 126406
rect 136940 126354 136946 126406
rect 136998 126354 137004 126406
rect 1794 126018 1800 126070
rect 1852 126018 1858 126070
rect 136940 126018 136946 126070
rect 136998 126018 137004 126070
rect 1794 125682 1800 125734
rect 1852 125682 1858 125734
rect 136940 125682 136946 125734
rect 136998 125682 137004 125734
rect 1794 125346 1800 125398
rect 1852 125346 1858 125398
rect 136940 125346 136946 125398
rect 136998 125346 137004 125398
rect 1794 125010 1800 125062
rect 1852 125010 1858 125062
rect 136940 125010 136946 125062
rect 136998 125010 137004 125062
rect 1794 124674 1800 124726
rect 1852 124674 1858 124726
rect 136940 124674 136946 124726
rect 136998 124674 137004 124726
rect 1794 124338 1800 124390
rect 1852 124338 1858 124390
rect 136940 124338 136946 124390
rect 136998 124338 137004 124390
rect 1794 124002 1800 124054
rect 1852 124002 1858 124054
rect 136940 124002 136946 124054
rect 136998 124002 137004 124054
rect 1794 123666 1800 123718
rect 1852 123666 1858 123718
rect 136940 123666 136946 123718
rect 136998 123666 137004 123718
rect 1794 123330 1800 123382
rect 1852 123330 1858 123382
rect 136940 123330 136946 123382
rect 136998 123330 137004 123382
rect 1794 122994 1800 123046
rect 1852 122994 1858 123046
rect 136940 122994 136946 123046
rect 136998 122994 137004 123046
rect 1794 122658 1800 122710
rect 1852 122658 1858 122710
rect 136940 122658 136946 122710
rect 136998 122658 137004 122710
rect 1794 122322 1800 122374
rect 1852 122322 1858 122374
rect 136940 122322 136946 122374
rect 136998 122322 137004 122374
rect 1794 121986 1800 122038
rect 1852 121986 1858 122038
rect 136940 121986 136946 122038
rect 136998 121986 137004 122038
rect 1794 121650 1800 121702
rect 1852 121650 1858 121702
rect 136940 121650 136946 121702
rect 136998 121650 137004 121702
rect 1794 121314 1800 121366
rect 1852 121314 1858 121366
rect 136940 121314 136946 121366
rect 136998 121314 137004 121366
rect 1794 120978 1800 121030
rect 1852 120978 1858 121030
rect 136940 120978 136946 121030
rect 136998 120978 137004 121030
rect 1794 120642 1800 120694
rect 1852 120642 1858 120694
rect 136940 120642 136946 120694
rect 136998 120642 137004 120694
rect 1794 120306 1800 120358
rect 1852 120306 1858 120358
rect 136940 120306 136946 120358
rect 136998 120306 137004 120358
rect 1794 119970 1800 120022
rect 1852 119970 1858 120022
rect 136940 119970 136946 120022
rect 136998 119970 137004 120022
rect 1794 119634 1800 119686
rect 1852 119634 1858 119686
rect 136940 119634 136946 119686
rect 136998 119634 137004 119686
rect 1794 119298 1800 119350
rect 1852 119298 1858 119350
rect 136940 119298 136946 119350
rect 136998 119298 137004 119350
rect 1794 118962 1800 119014
rect 1852 118962 1858 119014
rect 136940 118962 136946 119014
rect 136998 118962 137004 119014
rect 1794 118626 1800 118678
rect 1852 118626 1858 118678
rect 136940 118626 136946 118678
rect 136998 118626 137004 118678
rect 1794 118290 1800 118342
rect 1852 118290 1858 118342
rect 136940 118290 136946 118342
rect 136998 118290 137004 118342
rect 1794 117954 1800 118006
rect 1852 117954 1858 118006
rect 136940 117954 136946 118006
rect 136998 117954 137004 118006
rect 1794 117618 1800 117670
rect 1852 117618 1858 117670
rect 136940 117618 136946 117670
rect 136998 117618 137004 117670
rect 1794 117282 1800 117334
rect 1852 117282 1858 117334
rect 136940 117282 136946 117334
rect 136998 117282 137004 117334
rect 1794 116946 1800 116998
rect 1852 116946 1858 116998
rect 136940 116946 136946 116998
rect 136998 116946 137004 116998
rect 1794 116610 1800 116662
rect 1852 116610 1858 116662
rect 136940 116610 136946 116662
rect 136998 116610 137004 116662
rect 1794 116274 1800 116326
rect 1852 116274 1858 116326
rect 136940 116274 136946 116326
rect 136998 116274 137004 116326
rect 1794 115938 1800 115990
rect 1852 115938 1858 115990
rect 136940 115938 136946 115990
rect 136998 115938 137004 115990
rect 1794 115602 1800 115654
rect 1852 115602 1858 115654
rect 136940 115602 136946 115654
rect 136998 115602 137004 115654
rect 1794 115266 1800 115318
rect 1852 115266 1858 115318
rect 136940 115266 136946 115318
rect 136998 115266 137004 115318
rect 1794 114930 1800 114982
rect 1852 114930 1858 114982
rect 136940 114930 136946 114982
rect 136998 114930 137004 114982
rect 1794 114594 1800 114646
rect 1852 114594 1858 114646
rect 136940 114594 136946 114646
rect 136998 114594 137004 114646
rect 1794 114258 1800 114310
rect 1852 114258 1858 114310
rect 136940 114258 136946 114310
rect 136998 114258 137004 114310
rect 1794 113922 1800 113974
rect 1852 113922 1858 113974
rect 136940 113922 136946 113974
rect 136998 113922 137004 113974
rect 1794 113586 1800 113638
rect 1852 113586 1858 113638
rect 136940 113586 136946 113638
rect 136998 113586 137004 113638
rect 1794 113250 1800 113302
rect 1852 113250 1858 113302
rect 136940 113250 136946 113302
rect 136998 113250 137004 113302
rect 1794 112914 1800 112966
rect 1852 112914 1858 112966
rect 136940 112914 136946 112966
rect 136998 112914 137004 112966
rect 1794 112578 1800 112630
rect 1852 112578 1858 112630
rect 136940 112578 136946 112630
rect 136998 112578 137004 112630
rect 1794 112242 1800 112294
rect 1852 112242 1858 112294
rect 136940 112242 136946 112294
rect 136998 112242 137004 112294
rect 1794 111906 1800 111958
rect 1852 111906 1858 111958
rect 136940 111906 136946 111958
rect 136998 111906 137004 111958
rect 1794 111570 1800 111622
rect 1852 111570 1858 111622
rect 136940 111570 136946 111622
rect 136998 111570 137004 111622
rect 1794 111234 1800 111286
rect 1852 111234 1858 111286
rect 136940 111234 136946 111286
rect 136998 111234 137004 111286
rect 1794 110898 1800 110950
rect 1852 110898 1858 110950
rect 136940 110898 136946 110950
rect 136998 110898 137004 110950
rect 1794 110562 1800 110614
rect 1852 110562 1858 110614
rect 136940 110562 136946 110614
rect 136998 110562 137004 110614
rect 1794 110226 1800 110278
rect 1852 110226 1858 110278
rect 136940 110226 136946 110278
rect 136998 110226 137004 110278
rect 1794 109890 1800 109942
rect 1852 109890 1858 109942
rect 136940 109890 136946 109942
rect 136998 109890 137004 109942
rect 1794 109554 1800 109606
rect 1852 109554 1858 109606
rect 136940 109554 136946 109606
rect 136998 109554 137004 109606
rect 1794 109218 1800 109270
rect 1852 109218 1858 109270
rect 136940 109218 136946 109270
rect 136998 109218 137004 109270
rect 1794 108882 1800 108934
rect 1852 108882 1858 108934
rect 136940 108882 136946 108934
rect 136998 108882 137004 108934
rect 1794 108546 1800 108598
rect 1852 108546 1858 108598
rect 136940 108546 136946 108598
rect 136998 108546 137004 108598
rect 1794 108210 1800 108262
rect 1852 108210 1858 108262
rect 136940 108210 136946 108262
rect 136998 108210 137004 108262
rect 1794 107874 1800 107926
rect 1852 107874 1858 107926
rect 136940 107874 136946 107926
rect 136998 107874 137004 107926
rect 1794 107538 1800 107590
rect 1852 107538 1858 107590
rect 136940 107538 136946 107590
rect 136998 107538 137004 107590
rect 1794 107202 1800 107254
rect 1852 107202 1858 107254
rect 136940 107202 136946 107254
rect 136998 107202 137004 107254
rect 1794 106866 1800 106918
rect 1852 106866 1858 106918
rect 136940 106866 136946 106918
rect 136998 106866 137004 106918
rect 1794 106530 1800 106582
rect 1852 106530 1858 106582
rect 136940 106530 136946 106582
rect 136998 106530 137004 106582
rect 1794 106194 1800 106246
rect 1852 106194 1858 106246
rect 136940 106194 136946 106246
rect 136998 106194 137004 106246
rect 1794 105858 1800 105910
rect 1852 105858 1858 105910
rect 136940 105858 136946 105910
rect 136998 105858 137004 105910
rect 1794 105522 1800 105574
rect 1852 105522 1858 105574
rect 136940 105522 136946 105574
rect 136998 105522 137004 105574
rect 1794 105186 1800 105238
rect 1852 105186 1858 105238
rect 136940 105186 136946 105238
rect 136998 105186 137004 105238
rect 1794 104850 1800 104902
rect 1852 104850 1858 104902
rect 136940 104850 136946 104902
rect 136998 104850 137004 104902
rect 1794 104514 1800 104566
rect 1852 104514 1858 104566
rect 136940 104514 136946 104566
rect 136998 104514 137004 104566
rect 1794 104178 1800 104230
rect 1852 104178 1858 104230
rect 136940 104178 136946 104230
rect 136998 104178 137004 104230
rect 1794 103842 1800 103894
rect 1852 103842 1858 103894
rect 136940 103842 136946 103894
rect 136998 103842 137004 103894
rect 1794 103506 1800 103558
rect 1852 103506 1858 103558
rect 136940 103506 136946 103558
rect 136998 103506 137004 103558
rect 1794 103170 1800 103222
rect 1852 103170 1858 103222
rect 136940 103170 136946 103222
rect 136998 103170 137004 103222
rect 1794 102834 1800 102886
rect 1852 102834 1858 102886
rect 136940 102834 136946 102886
rect 136998 102834 137004 102886
rect 1794 102498 1800 102550
rect 1852 102498 1858 102550
rect 136940 102498 136946 102550
rect 136998 102498 137004 102550
rect 1794 102162 1800 102214
rect 1852 102162 1858 102214
rect 136940 102162 136946 102214
rect 136998 102162 137004 102214
rect 1794 101826 1800 101878
rect 1852 101826 1858 101878
rect 136940 101826 136946 101878
rect 136998 101826 137004 101878
rect 1794 101490 1800 101542
rect 1852 101490 1858 101542
rect 136940 101490 136946 101542
rect 136998 101490 137004 101542
rect 1794 101154 1800 101206
rect 1852 101154 1858 101206
rect 136940 101154 136946 101206
rect 136998 101154 137004 101206
rect 1794 100818 1800 100870
rect 1852 100818 1858 100870
rect 136940 100818 136946 100870
rect 136998 100818 137004 100870
rect 1794 100482 1800 100534
rect 1852 100482 1858 100534
rect 136940 100482 136946 100534
rect 136998 100482 137004 100534
rect 1794 100146 1800 100198
rect 1852 100146 1858 100198
rect 136940 100146 136946 100198
rect 136998 100146 137004 100198
rect 1794 99810 1800 99862
rect 1852 99810 1858 99862
rect 136940 99810 136946 99862
rect 136998 99810 137004 99862
rect 1794 99474 1800 99526
rect 1852 99474 1858 99526
rect 136940 99474 136946 99526
rect 136998 99474 137004 99526
rect 1794 99138 1800 99190
rect 1852 99138 1858 99190
rect 136940 99138 136946 99190
rect 136998 99138 137004 99190
rect 1794 98802 1800 98854
rect 1852 98802 1858 98854
rect 136940 98802 136946 98854
rect 136998 98802 137004 98854
rect 1794 98466 1800 98518
rect 1852 98466 1858 98518
rect 136940 98466 136946 98518
rect 136998 98466 137004 98518
rect 1794 98130 1800 98182
rect 1852 98130 1858 98182
rect 136940 98130 136946 98182
rect 136998 98130 137004 98182
rect 1794 97794 1800 97846
rect 1852 97794 1858 97846
rect 136940 97794 136946 97846
rect 136998 97794 137004 97846
rect 1794 97458 1800 97510
rect 1852 97458 1858 97510
rect 136940 97458 136946 97510
rect 136998 97458 137004 97510
rect 1794 97122 1800 97174
rect 1852 97122 1858 97174
rect 136940 97122 136946 97174
rect 136998 97122 137004 97174
rect 1794 96786 1800 96838
rect 1852 96786 1858 96838
rect 136940 96786 136946 96838
rect 136998 96786 137004 96838
rect 1794 96450 1800 96502
rect 1852 96450 1858 96502
rect 136940 96450 136946 96502
rect 136998 96450 137004 96502
rect 1794 96114 1800 96166
rect 1852 96114 1858 96166
rect 136940 96114 136946 96166
rect 136998 96114 137004 96166
rect 1794 95778 1800 95830
rect 1852 95778 1858 95830
rect 136940 95778 136946 95830
rect 136998 95778 137004 95830
rect 1794 95442 1800 95494
rect 1852 95442 1858 95494
rect 136940 95442 136946 95494
rect 136998 95442 137004 95494
rect 1794 95106 1800 95158
rect 1852 95106 1858 95158
rect 136940 95106 136946 95158
rect 136998 95106 137004 95158
rect 1794 94770 1800 94822
rect 1852 94770 1858 94822
rect 136940 94770 136946 94822
rect 136998 94770 137004 94822
rect 1794 94434 1800 94486
rect 1852 94434 1858 94486
rect 136940 94434 136946 94486
rect 136998 94434 137004 94486
rect 1794 94098 1800 94150
rect 1852 94098 1858 94150
rect 136940 94098 136946 94150
rect 136998 94098 137004 94150
rect 1794 93762 1800 93814
rect 1852 93762 1858 93814
rect 136940 93762 136946 93814
rect 136998 93762 137004 93814
rect 1794 93426 1800 93478
rect 1852 93426 1858 93478
rect 136940 93426 136946 93478
rect 136998 93426 137004 93478
rect 1794 93090 1800 93142
rect 1852 93090 1858 93142
rect 136940 93090 136946 93142
rect 136998 93090 137004 93142
rect 1794 92754 1800 92806
rect 1852 92754 1858 92806
rect 136940 92754 136946 92806
rect 136998 92754 137004 92806
rect 1794 92418 1800 92470
rect 1852 92418 1858 92470
rect 136940 92418 136946 92470
rect 136998 92418 137004 92470
rect 1794 92082 1800 92134
rect 1852 92082 1858 92134
rect 136940 92082 136946 92134
rect 136998 92082 137004 92134
rect 1794 91746 1800 91798
rect 1852 91746 1858 91798
rect 136940 91746 136946 91798
rect 136998 91746 137004 91798
rect 1794 91410 1800 91462
rect 1852 91410 1858 91462
rect 136940 91410 136946 91462
rect 136998 91410 137004 91462
rect 1794 91074 1800 91126
rect 1852 91074 1858 91126
rect 136940 91074 136946 91126
rect 136998 91074 137004 91126
rect 1794 90738 1800 90790
rect 1852 90738 1858 90790
rect 136940 90738 136946 90790
rect 136998 90738 137004 90790
rect 1794 90402 1800 90454
rect 1852 90402 1858 90454
rect 136940 90402 136946 90454
rect 136998 90402 137004 90454
rect 1794 90066 1800 90118
rect 1852 90066 1858 90118
rect 136940 90066 136946 90118
rect 136998 90066 137004 90118
rect 1794 89730 1800 89782
rect 1852 89730 1858 89782
rect 136940 89730 136946 89782
rect 136998 89730 137004 89782
rect 1794 89394 1800 89446
rect 1852 89394 1858 89446
rect 136940 89394 136946 89446
rect 136998 89394 137004 89446
rect 1794 89058 1800 89110
rect 1852 89058 1858 89110
rect 136940 89058 136946 89110
rect 136998 89058 137004 89110
rect 1794 88722 1800 88774
rect 1852 88722 1858 88774
rect 136940 88722 136946 88774
rect 136998 88722 137004 88774
rect 1794 88386 1800 88438
rect 1852 88386 1858 88438
rect 136940 88386 136946 88438
rect 136998 88386 137004 88438
rect 1794 88050 1800 88102
rect 1852 88050 1858 88102
rect 136940 88050 136946 88102
rect 136998 88050 137004 88102
rect 1794 87714 1800 87766
rect 1852 87714 1858 87766
rect 136940 87714 136946 87766
rect 136998 87714 137004 87766
rect 1794 87378 1800 87430
rect 1852 87378 1858 87430
rect 136940 87378 136946 87430
rect 136998 87378 137004 87430
rect 1794 87042 1800 87094
rect 1852 87042 1858 87094
rect 136940 87042 136946 87094
rect 136998 87042 137004 87094
rect 1794 86706 1800 86758
rect 1852 86706 1858 86758
rect 136940 86706 136946 86758
rect 136998 86706 137004 86758
rect 1794 86370 1800 86422
rect 1852 86370 1858 86422
rect 136940 86370 136946 86422
rect 136998 86370 137004 86422
rect 1794 86034 1800 86086
rect 1852 86034 1858 86086
rect 136940 86034 136946 86086
rect 136998 86034 137004 86086
rect 1794 85698 1800 85750
rect 1852 85698 1858 85750
rect 136940 85698 136946 85750
rect 136998 85698 137004 85750
rect 1794 85362 1800 85414
rect 1852 85362 1858 85414
rect 136940 85362 136946 85414
rect 136998 85362 137004 85414
rect 1794 85026 1800 85078
rect 1852 85026 1858 85078
rect 136940 85026 136946 85078
rect 136998 85026 137004 85078
rect 1794 84690 1800 84742
rect 1852 84690 1858 84742
rect 136940 84690 136946 84742
rect 136998 84690 137004 84742
rect 1794 84354 1800 84406
rect 1852 84354 1858 84406
rect 136940 84354 136946 84406
rect 136998 84354 137004 84406
rect 1794 84018 1800 84070
rect 1852 84018 1858 84070
rect 136940 84018 136946 84070
rect 136998 84018 137004 84070
rect 1794 83682 1800 83734
rect 1852 83682 1858 83734
rect 136940 83682 136946 83734
rect 136998 83682 137004 83734
rect 1794 83346 1800 83398
rect 1852 83346 1858 83398
rect 136940 83346 136946 83398
rect 136998 83346 137004 83398
rect 1794 83010 1800 83062
rect 1852 83010 1858 83062
rect 136940 83010 136946 83062
rect 136998 83010 137004 83062
rect 1794 82674 1800 82726
rect 1852 82674 1858 82726
rect 136940 82674 136946 82726
rect 136998 82674 137004 82726
rect 1794 82338 1800 82390
rect 1852 82338 1858 82390
rect 136940 82338 136946 82390
rect 136998 82338 137004 82390
rect 1794 82002 1800 82054
rect 1852 82002 1858 82054
rect 136940 82002 136946 82054
rect 136998 82002 137004 82054
rect 1794 81666 1800 81718
rect 1852 81666 1858 81718
rect 136940 81666 136946 81718
rect 136998 81666 137004 81718
rect 1794 81330 1800 81382
rect 1852 81330 1858 81382
rect 136940 81330 136946 81382
rect 136998 81330 137004 81382
rect 1794 80994 1800 81046
rect 1852 80994 1858 81046
rect 136940 80994 136946 81046
rect 136998 80994 137004 81046
rect 1794 80658 1800 80710
rect 1852 80658 1858 80710
rect 136940 80658 136946 80710
rect 136998 80658 137004 80710
rect 1794 80322 1800 80374
rect 1852 80322 1858 80374
rect 136940 80322 136946 80374
rect 136998 80322 137004 80374
rect 1794 79986 1800 80038
rect 1852 79986 1858 80038
rect 136940 79986 136946 80038
rect 136998 79986 137004 80038
rect 1794 79650 1800 79702
rect 1852 79650 1858 79702
rect 136940 79650 136946 79702
rect 136998 79650 137004 79702
rect 1794 79314 1800 79366
rect 1852 79314 1858 79366
rect 136940 79314 136946 79366
rect 136998 79314 137004 79366
rect 1794 78978 1800 79030
rect 1852 78978 1858 79030
rect 136940 78978 136946 79030
rect 136998 78978 137004 79030
rect 1794 78642 1800 78694
rect 1852 78642 1858 78694
rect 136940 78642 136946 78694
rect 136998 78642 137004 78694
rect 1794 78306 1800 78358
rect 1852 78306 1858 78358
rect 136940 78306 136946 78358
rect 136998 78306 137004 78358
rect 1794 77970 1800 78022
rect 1852 77970 1858 78022
rect 136940 77970 136946 78022
rect 136998 77970 137004 78022
rect 1794 77634 1800 77686
rect 1852 77634 1858 77686
rect 136940 77634 136946 77686
rect 136998 77634 137004 77686
rect 1794 77298 1800 77350
rect 1852 77298 1858 77350
rect 136940 77298 136946 77350
rect 136998 77298 137004 77350
rect 1794 76962 1800 77014
rect 1852 76962 1858 77014
rect 136940 76962 136946 77014
rect 136998 76962 137004 77014
rect 1794 76626 1800 76678
rect 1852 76626 1858 76678
rect 136940 76626 136946 76678
rect 136998 76626 137004 76678
rect 1794 76290 1800 76342
rect 1852 76290 1858 76342
rect 136940 76290 136946 76342
rect 136998 76290 137004 76342
rect 1794 75954 1800 76006
rect 1852 75954 1858 76006
rect 136940 75954 136946 76006
rect 136998 75954 137004 76006
rect 1794 75618 1800 75670
rect 1852 75618 1858 75670
rect 136940 75618 136946 75670
rect 136998 75618 137004 75670
rect 1794 75282 1800 75334
rect 1852 75282 1858 75334
rect 136940 75282 136946 75334
rect 136998 75282 137004 75334
rect 1794 74946 1800 74998
rect 1852 74946 1858 74998
rect 136940 74946 136946 74998
rect 136998 74946 137004 74998
rect 1794 74610 1800 74662
rect 1852 74610 1858 74662
rect 136940 74610 136946 74662
rect 136998 74610 137004 74662
rect 1794 74274 1800 74326
rect 1852 74274 1858 74326
rect 136940 74274 136946 74326
rect 136998 74274 137004 74326
rect 1794 73938 1800 73990
rect 1852 73938 1858 73990
rect 136940 73938 136946 73990
rect 136998 73938 137004 73990
rect 1794 73602 1800 73654
rect 1852 73602 1858 73654
rect 136940 73602 136946 73654
rect 136998 73602 137004 73654
rect 1794 73266 1800 73318
rect 1852 73266 1858 73318
rect 136940 73266 136946 73318
rect 136998 73266 137004 73318
rect 1794 72930 1800 72982
rect 1852 72930 1858 72982
rect 136940 72930 136946 72982
rect 136998 72930 137004 72982
rect 1794 72594 1800 72646
rect 1852 72594 1858 72646
rect 136940 72594 136946 72646
rect 136998 72594 137004 72646
rect 1794 72258 1800 72310
rect 1852 72258 1858 72310
rect 136940 72258 136946 72310
rect 136998 72258 137004 72310
rect 1794 71922 1800 71974
rect 1852 71922 1858 71974
rect 136940 71922 136946 71974
rect 136998 71922 137004 71974
rect 1794 71586 1800 71638
rect 1852 71586 1858 71638
rect 136940 71586 136946 71638
rect 136998 71586 137004 71638
rect 1794 71250 1800 71302
rect 1852 71250 1858 71302
rect 136940 71250 136946 71302
rect 136998 71250 137004 71302
rect 1794 70914 1800 70966
rect 1852 70914 1858 70966
rect 136940 70914 136946 70966
rect 136998 70914 137004 70966
rect 1794 70578 1800 70630
rect 1852 70578 1858 70630
rect 136940 70578 136946 70630
rect 136998 70578 137004 70630
rect 1794 70242 1800 70294
rect 1852 70242 1858 70294
rect 136940 70242 136946 70294
rect 136998 70242 137004 70294
rect 1794 69906 1800 69958
rect 1852 69906 1858 69958
rect 136940 69906 136946 69958
rect 136998 69906 137004 69958
rect 1794 69570 1800 69622
rect 1852 69570 1858 69622
rect 136940 69570 136946 69622
rect 136998 69570 137004 69622
rect 1794 69234 1800 69286
rect 1852 69234 1858 69286
rect 136940 69234 136946 69286
rect 136998 69234 137004 69286
rect 1794 68898 1800 68950
rect 1852 68898 1858 68950
rect 136940 68898 136946 68950
rect 136998 68898 137004 68950
rect 1794 68562 1800 68614
rect 1852 68562 1858 68614
rect 136940 68562 136946 68614
rect 136998 68562 137004 68614
rect 1794 68226 1800 68278
rect 1852 68226 1858 68278
rect 136940 68226 136946 68278
rect 136998 68226 137004 68278
rect 1794 67890 1800 67942
rect 1852 67890 1858 67942
rect 136940 67890 136946 67942
rect 136998 67890 137004 67942
rect 1794 67554 1800 67606
rect 1852 67554 1858 67606
rect 136940 67554 136946 67606
rect 136998 67554 137004 67606
rect 1794 67218 1800 67270
rect 1852 67218 1858 67270
rect 136940 67218 136946 67270
rect 136998 67218 137004 67270
rect 1794 66882 1800 66934
rect 1852 66882 1858 66934
rect 136940 66882 136946 66934
rect 136998 66882 137004 66934
rect 1794 66546 1800 66598
rect 1852 66546 1858 66598
rect 136940 66546 136946 66598
rect 136998 66546 137004 66598
rect 1794 66210 1800 66262
rect 1852 66210 1858 66262
rect 136940 66210 136946 66262
rect 136998 66210 137004 66262
rect 1794 65874 1800 65926
rect 1852 65874 1858 65926
rect 136940 65874 136946 65926
rect 136998 65874 137004 65926
rect 1794 65538 1800 65590
rect 1852 65538 1858 65590
rect 136940 65538 136946 65590
rect 136998 65538 137004 65590
rect 1794 65202 1800 65254
rect 1852 65202 1858 65254
rect 136940 65202 136946 65254
rect 136998 65202 137004 65254
rect 1794 64866 1800 64918
rect 1852 64866 1858 64918
rect 136940 64866 136946 64918
rect 136998 64866 137004 64918
rect 1794 64530 1800 64582
rect 1852 64530 1858 64582
rect 136940 64530 136946 64582
rect 136998 64530 137004 64582
rect 1794 64194 1800 64246
rect 1852 64194 1858 64246
rect 136940 64194 136946 64246
rect 136998 64194 137004 64246
rect 1794 63858 1800 63910
rect 1852 63858 1858 63910
rect 136940 63858 136946 63910
rect 136998 63858 137004 63910
rect 1794 63522 1800 63574
rect 1852 63522 1858 63574
rect 136940 63522 136946 63574
rect 136998 63522 137004 63574
rect 1794 63186 1800 63238
rect 1852 63186 1858 63238
rect 136940 63186 136946 63238
rect 136998 63186 137004 63238
rect 1794 62850 1800 62902
rect 1852 62850 1858 62902
rect 136940 62850 136946 62902
rect 136998 62850 137004 62902
rect 1794 62514 1800 62566
rect 1852 62514 1858 62566
rect 136940 62514 136946 62566
rect 136998 62514 137004 62566
rect 1794 62178 1800 62230
rect 1852 62178 1858 62230
rect 136940 62178 136946 62230
rect 136998 62178 137004 62230
rect 1794 61842 1800 61894
rect 1852 61842 1858 61894
rect 136940 61842 136946 61894
rect 136998 61842 137004 61894
rect 1794 61506 1800 61558
rect 1852 61506 1858 61558
rect 136940 61506 136946 61558
rect 136998 61506 137004 61558
rect 1794 61170 1800 61222
rect 1852 61170 1858 61222
rect 136940 61170 136946 61222
rect 136998 61170 137004 61222
rect 1794 60834 1800 60886
rect 1852 60834 1858 60886
rect 136940 60834 136946 60886
rect 136998 60834 137004 60886
rect 1794 60498 1800 60550
rect 1852 60498 1858 60550
rect 136940 60498 136946 60550
rect 136998 60498 137004 60550
rect 1794 60162 1800 60214
rect 1852 60162 1858 60214
rect 136940 60162 136946 60214
rect 136998 60162 137004 60214
rect 1794 59826 1800 59878
rect 1852 59826 1858 59878
rect 136940 59826 136946 59878
rect 136998 59826 137004 59878
rect 1794 59490 1800 59542
rect 1852 59490 1858 59542
rect 136940 59490 136946 59542
rect 136998 59490 137004 59542
rect 1794 59154 1800 59206
rect 1852 59154 1858 59206
rect 136940 59154 136946 59206
rect 136998 59154 137004 59206
rect 1794 58818 1800 58870
rect 1852 58818 1858 58870
rect 136940 58818 136946 58870
rect 136998 58818 137004 58870
rect 1794 58482 1800 58534
rect 1852 58482 1858 58534
rect 136940 58482 136946 58534
rect 136998 58482 137004 58534
rect 1794 58146 1800 58198
rect 1852 58146 1858 58198
rect 136940 58146 136946 58198
rect 136998 58146 137004 58198
rect 1794 57810 1800 57862
rect 1852 57810 1858 57862
rect 136940 57810 136946 57862
rect 136998 57810 137004 57862
rect 1794 57474 1800 57526
rect 1852 57474 1858 57526
rect 136940 57474 136946 57526
rect 136998 57474 137004 57526
rect 1794 57138 1800 57190
rect 1852 57138 1858 57190
rect 136940 57138 136946 57190
rect 136998 57138 137004 57190
rect 1794 56802 1800 56854
rect 1852 56802 1858 56854
rect 136940 56802 136946 56854
rect 136998 56802 137004 56854
rect 1794 56466 1800 56518
rect 1852 56466 1858 56518
rect 136940 56466 136946 56518
rect 136998 56466 137004 56518
rect 1794 56130 1800 56182
rect 1852 56130 1858 56182
rect 136940 56130 136946 56182
rect 136998 56130 137004 56182
rect 1794 55794 1800 55846
rect 1852 55794 1858 55846
rect 136940 55794 136946 55846
rect 136998 55794 137004 55846
rect 1794 55458 1800 55510
rect 1852 55458 1858 55510
rect 136940 55458 136946 55510
rect 136998 55458 137004 55510
rect 1794 55122 1800 55174
rect 1852 55122 1858 55174
rect 136940 55122 136946 55174
rect 136998 55122 137004 55174
rect 1794 54786 1800 54838
rect 1852 54786 1858 54838
rect 136940 54786 136946 54838
rect 136998 54786 137004 54838
rect 1794 54450 1800 54502
rect 1852 54450 1858 54502
rect 136940 54450 136946 54502
rect 136998 54450 137004 54502
rect 1794 54114 1800 54166
rect 1852 54114 1858 54166
rect 136940 54114 136946 54166
rect 136998 54114 137004 54166
rect 1794 53778 1800 53830
rect 1852 53778 1858 53830
rect 136940 53778 136946 53830
rect 136998 53778 137004 53830
rect 1794 53442 1800 53494
rect 1852 53442 1858 53494
rect 136940 53442 136946 53494
rect 136998 53442 137004 53494
rect 1794 53106 1800 53158
rect 1852 53106 1858 53158
rect 136940 53106 136946 53158
rect 136998 53106 137004 53158
rect 1794 52770 1800 52822
rect 1852 52770 1858 52822
rect 136940 52770 136946 52822
rect 136998 52770 137004 52822
rect 1794 52434 1800 52486
rect 1852 52434 1858 52486
rect 136940 52434 136946 52486
rect 136998 52434 137004 52486
rect 1794 52098 1800 52150
rect 1852 52098 1858 52150
rect 136940 52098 136946 52150
rect 136998 52098 137004 52150
rect 1794 51762 1800 51814
rect 1852 51762 1858 51814
rect 136940 51762 136946 51814
rect 136998 51762 137004 51814
rect 1794 51426 1800 51478
rect 1852 51426 1858 51478
rect 136940 51426 136946 51478
rect 136998 51426 137004 51478
rect 1794 51090 1800 51142
rect 1852 51090 1858 51142
rect 136940 51090 136946 51142
rect 136998 51090 137004 51142
rect 1794 50754 1800 50806
rect 1852 50754 1858 50806
rect 136940 50754 136946 50806
rect 136998 50754 137004 50806
rect 1794 50418 1800 50470
rect 1852 50418 1858 50470
rect 136940 50418 136946 50470
rect 136998 50418 137004 50470
rect 1794 50082 1800 50134
rect 1852 50082 1858 50134
rect 136940 50082 136946 50134
rect 136998 50082 137004 50134
rect 1794 49746 1800 49798
rect 1852 49746 1858 49798
rect 136940 49746 136946 49798
rect 136998 49746 137004 49798
rect 1794 49410 1800 49462
rect 1852 49410 1858 49462
rect 136940 49410 136946 49462
rect 136998 49410 137004 49462
rect 1794 49074 1800 49126
rect 1852 49074 1858 49126
rect 136940 49074 136946 49126
rect 136998 49074 137004 49126
rect 1794 48738 1800 48790
rect 1852 48738 1858 48790
rect 136940 48738 136946 48790
rect 136998 48738 137004 48790
rect 1794 48402 1800 48454
rect 1852 48402 1858 48454
rect 136940 48402 136946 48454
rect 136998 48402 137004 48454
rect 1794 48066 1800 48118
rect 1852 48066 1858 48118
rect 136940 48066 136946 48118
rect 136998 48066 137004 48118
rect 1794 47730 1800 47782
rect 1852 47730 1858 47782
rect 136940 47730 136946 47782
rect 136998 47730 137004 47782
rect 1794 47394 1800 47446
rect 1852 47394 1858 47446
rect 136940 47394 136946 47446
rect 136998 47394 137004 47446
rect 1794 47058 1800 47110
rect 1852 47058 1858 47110
rect 136940 47058 136946 47110
rect 136998 47058 137004 47110
rect 1794 46722 1800 46774
rect 1852 46722 1858 46774
rect 136940 46722 136946 46774
rect 136998 46722 137004 46774
rect 1794 46386 1800 46438
rect 1852 46386 1858 46438
rect 136940 46386 136946 46438
rect 136998 46386 137004 46438
rect 1794 46050 1800 46102
rect 1852 46050 1858 46102
rect 136940 46050 136946 46102
rect 136998 46050 137004 46102
rect 1794 45714 1800 45766
rect 1852 45714 1858 45766
rect 136940 45714 136946 45766
rect 136998 45714 137004 45766
rect 1794 45378 1800 45430
rect 1852 45378 1858 45430
rect 136940 45378 136946 45430
rect 136998 45378 137004 45430
rect 1794 45042 1800 45094
rect 1852 45042 1858 45094
rect 136940 45042 136946 45094
rect 136998 45042 137004 45094
rect 1794 44706 1800 44758
rect 1852 44706 1858 44758
rect 136940 44706 136946 44758
rect 136998 44706 137004 44758
rect 1794 44370 1800 44422
rect 1852 44370 1858 44422
rect 136940 44370 136946 44422
rect 136998 44370 137004 44422
rect 1794 44034 1800 44086
rect 1852 44034 1858 44086
rect 136940 44034 136946 44086
rect 136998 44034 137004 44086
rect 1794 43698 1800 43750
rect 1852 43698 1858 43750
rect 136940 43698 136946 43750
rect 136998 43698 137004 43750
rect 1794 43362 1800 43414
rect 1852 43362 1858 43414
rect 136940 43362 136946 43414
rect 136998 43362 137004 43414
rect 1794 43026 1800 43078
rect 1852 43026 1858 43078
rect 136940 43026 136946 43078
rect 136998 43026 137004 43078
rect 1794 42690 1800 42742
rect 1852 42690 1858 42742
rect 136940 42690 136946 42742
rect 136998 42690 137004 42742
rect 1794 42354 1800 42406
rect 1852 42354 1858 42406
rect 136940 42354 136946 42406
rect 136998 42354 137004 42406
rect 1794 42018 1800 42070
rect 1852 42018 1858 42070
rect 136940 42018 136946 42070
rect 136998 42018 137004 42070
rect 1794 41682 1800 41734
rect 1852 41682 1858 41734
rect 136940 41682 136946 41734
rect 136998 41682 137004 41734
rect 1794 41346 1800 41398
rect 1852 41346 1858 41398
rect 136940 41346 136946 41398
rect 136998 41346 137004 41398
rect 1794 41010 1800 41062
rect 1852 41010 1858 41062
rect 136940 41010 136946 41062
rect 136998 41010 137004 41062
rect 1794 40674 1800 40726
rect 1852 40674 1858 40726
rect 136940 40674 136946 40726
rect 136998 40674 137004 40726
rect 1794 40338 1800 40390
rect 1852 40338 1858 40390
rect 136940 40338 136946 40390
rect 136998 40338 137004 40390
rect 1794 40002 1800 40054
rect 1852 40002 1858 40054
rect 15967 39977 15973 40029
rect 16025 39977 16031 40029
rect 136940 40002 136946 40054
rect 136998 40002 137004 40054
rect 1794 39666 1800 39718
rect 1852 39666 1858 39718
rect 1794 39330 1800 39382
rect 1852 39330 1858 39382
rect 1794 38994 1800 39046
rect 1852 38994 1858 39046
rect 1794 38658 1800 38710
rect 1852 38658 1858 38710
rect 15887 38419 15893 38471
rect 15945 38419 15951 38471
rect 1794 38322 1800 38374
rect 1852 38322 1858 38374
rect 1794 37986 1800 38038
rect 1852 37986 1858 38038
rect 1794 37650 1800 37702
rect 1852 37650 1858 37702
rect 1794 37314 1800 37366
rect 1852 37314 1858 37366
rect 15807 37149 15813 37201
rect 15865 37149 15871 37201
rect 1794 36978 1800 37030
rect 1852 36978 1858 37030
rect 1794 36642 1800 36694
rect 1852 36642 1858 36694
rect 1794 36306 1800 36358
rect 1852 36306 1858 36358
rect 1794 35970 1800 36022
rect 1852 35970 1858 36022
rect 1794 35634 1800 35686
rect 1852 35634 1858 35686
rect 15727 35591 15733 35643
rect 15785 35591 15791 35643
rect 1794 35298 1800 35350
rect 1852 35298 1858 35350
rect 1794 34962 1800 35014
rect 1852 34962 1858 35014
rect 1794 34626 1800 34678
rect 1852 34626 1858 34678
rect 1794 34290 1800 34342
rect 1852 34290 1858 34342
rect 15647 34321 15653 34373
rect 15705 34321 15711 34373
rect 1794 33954 1800 34006
rect 1852 33954 1858 34006
rect 1794 33618 1800 33670
rect 1852 33618 1858 33670
rect 1794 33282 1800 33334
rect 1852 33282 1858 33334
rect 1794 32946 1800 32998
rect 1852 32946 1858 32998
rect 15567 32763 15573 32815
rect 15625 32763 15631 32815
rect 1794 32610 1800 32662
rect 1852 32610 1858 32662
rect 1794 32274 1800 32326
rect 1852 32274 1858 32326
rect 1794 31938 1800 31990
rect 1852 31938 1858 31990
rect 1794 31602 1800 31654
rect 1852 31602 1858 31654
rect 15487 31493 15493 31545
rect 15545 31493 15551 31545
rect 1794 31266 1800 31318
rect 1852 31266 1858 31318
rect 1794 30930 1800 30982
rect 1852 30930 1858 30982
rect 1794 30594 1800 30646
rect 1852 30594 1858 30646
rect 1794 30258 1800 30310
rect 1852 30258 1858 30310
rect 1794 29922 1800 29974
rect 1852 29922 1858 29974
rect 15407 29935 15413 29987
rect 15465 29935 15471 29987
rect 1794 29586 1800 29638
rect 1852 29586 1858 29638
rect 1794 29250 1800 29302
rect 1852 29250 1858 29302
rect 1794 28914 1800 28966
rect 1852 28914 1858 28966
rect 1794 28578 1800 28630
rect 1852 28578 1858 28630
rect 1794 28242 1800 28294
rect 1852 28242 1858 28294
rect 1794 27906 1800 27958
rect 1852 27906 1858 27958
rect 1794 27570 1800 27622
rect 1852 27570 1858 27622
rect 1794 27234 1800 27286
rect 1852 27234 1858 27286
rect 1794 26898 1800 26950
rect 1852 26898 1858 26950
rect 1794 26562 1800 26614
rect 1852 26562 1858 26614
rect 1794 26226 1800 26278
rect 1852 26226 1858 26278
rect 1794 25890 1800 25942
rect 1852 25890 1858 25942
rect 1794 25554 1800 25606
rect 1852 25554 1858 25606
rect 1794 25218 1800 25270
rect 1852 25218 1858 25270
rect 1794 24882 1800 24934
rect 1852 24882 1858 24934
rect 1794 24546 1800 24598
rect 1852 24546 1858 24598
rect 15425 24586 15453 29935
rect 15505 24586 15533 31493
rect 15585 24586 15613 32763
rect 15665 24586 15693 34321
rect 15745 24586 15773 35591
rect 15825 24586 15853 37149
rect 15905 24586 15933 38419
rect 15985 24586 16013 39977
rect 136940 39666 136946 39718
rect 136998 39666 137004 39718
rect 136940 39330 136946 39382
rect 136998 39330 137004 39382
rect 136940 38994 136946 39046
rect 136998 38994 137004 39046
rect 136940 38658 136946 38710
rect 136998 38658 137004 38710
rect 136940 38322 136946 38374
rect 136998 38322 137004 38374
rect 136940 37986 136946 38038
rect 136998 37986 137004 38038
rect 136940 37650 136946 37702
rect 136998 37650 137004 37702
rect 136940 37314 136946 37366
rect 136998 37314 137004 37366
rect 136940 36978 136946 37030
rect 136998 36978 137004 37030
rect 136940 36642 136946 36694
rect 136998 36642 137004 36694
rect 136940 36306 136946 36358
rect 136998 36306 137004 36358
rect 136940 35970 136946 36022
rect 136998 35970 137004 36022
rect 136940 35634 136946 35686
rect 136998 35634 137004 35686
rect 136940 35298 136946 35350
rect 136998 35298 137004 35350
rect 136940 34962 136946 35014
rect 136998 34962 137004 35014
rect 136940 34626 136946 34678
rect 136998 34626 137004 34678
rect 136940 34290 136946 34342
rect 136998 34290 137004 34342
rect 136940 33954 136946 34006
rect 136998 33954 137004 34006
rect 136940 33618 136946 33670
rect 136998 33618 137004 33670
rect 136940 33282 136946 33334
rect 136998 33282 137004 33334
rect 136940 32946 136946 32998
rect 136998 32946 137004 32998
rect 136940 32610 136946 32662
rect 136998 32610 137004 32662
rect 136940 32274 136946 32326
rect 136998 32274 137004 32326
rect 136940 31938 136946 31990
rect 136998 31938 137004 31990
rect 136940 31602 136946 31654
rect 136998 31602 137004 31654
rect 136940 31266 136946 31318
rect 136998 31266 137004 31318
rect 136940 30930 136946 30982
rect 136998 30930 137004 30982
rect 136940 30594 136946 30646
rect 136998 30594 137004 30646
rect 136940 30258 136946 30310
rect 136998 30258 137004 30310
rect 136940 29922 136946 29974
rect 136998 29922 137004 29974
rect 136940 29586 136946 29638
rect 136998 29586 137004 29638
rect 136940 29250 136946 29302
rect 136998 29250 137004 29302
rect 136940 28914 136946 28966
rect 136998 28914 137004 28966
rect 136940 28578 136946 28630
rect 136998 28578 137004 28630
rect 136940 28242 136946 28294
rect 136998 28242 137004 28294
rect 136940 27906 136946 27958
rect 136998 27906 137004 27958
rect 136940 27570 136946 27622
rect 136998 27570 137004 27622
rect 136940 27234 136946 27286
rect 136998 27234 137004 27286
rect 136940 26898 136946 26950
rect 136998 26898 137004 26950
rect 136940 26562 136946 26614
rect 136998 26562 137004 26614
rect 136940 26226 136946 26278
rect 136998 26226 137004 26278
rect 136940 25890 136946 25942
rect 136998 25890 137004 25942
rect 136940 25554 136946 25606
rect 136998 25554 137004 25606
rect 136940 25218 136946 25270
rect 136998 25218 137004 25270
rect 136940 24882 136946 24934
rect 136998 24882 137004 24934
rect 1794 24210 1800 24262
rect 1852 24210 1858 24262
rect 1794 23874 1800 23926
rect 1852 23874 1858 23926
rect 1794 23538 1800 23590
rect 1852 23538 1858 23590
rect 1794 23202 1800 23254
rect 1852 23202 1858 23254
rect 1794 22866 1800 22918
rect 1852 22866 1858 22918
rect 1794 22530 1800 22582
rect 1852 22530 1858 22582
rect 1794 22194 1800 22246
rect 1852 22194 1858 22246
rect 1794 21858 1800 21910
rect 1852 21858 1858 21910
rect 1794 21522 1800 21574
rect 1852 21522 1858 21574
rect 1794 21186 1800 21238
rect 1852 21186 1858 21238
rect 1794 20850 1800 20902
rect 1852 20850 1858 20902
rect 1794 20514 1800 20566
rect 1852 20514 1858 20566
rect 1794 20178 1800 20230
rect 1852 20178 1858 20230
rect 1794 19842 1800 19894
rect 1852 19842 1858 19894
rect 1794 19506 1800 19558
rect 1852 19506 1858 19558
rect 1794 19170 1800 19222
rect 1852 19170 1858 19222
rect 1794 18834 1800 18886
rect 1852 18834 1858 18886
rect 1794 18498 1800 18550
rect 1852 18498 1858 18550
rect 1794 18162 1800 18214
rect 1852 18162 1858 18214
rect 1794 17826 1800 17878
rect 1852 17826 1858 17878
rect 1794 17490 1800 17542
rect 1852 17490 1858 17542
rect 1794 17154 1800 17206
rect 1852 17154 1858 17206
rect 1794 16818 1800 16870
rect 1852 16818 1858 16870
rect 1794 16482 1800 16534
rect 1852 16482 1858 16534
rect 1794 16146 1800 16198
rect 1852 16146 1858 16198
rect 1794 15810 1800 15862
rect 1852 15810 1858 15862
rect 1794 15474 1800 15526
rect 1852 15474 1858 15526
rect 1794 15138 1800 15190
rect 1852 15138 1858 15190
rect 1794 14802 1800 14854
rect 1852 14802 1858 14854
rect 1794 14466 1800 14518
rect 1852 14466 1858 14518
rect 1794 14130 1800 14182
rect 1852 14130 1858 14182
rect 1794 13794 1800 13846
rect 1852 13794 1858 13846
rect 1794 13458 1800 13510
rect 1852 13458 1858 13510
rect 29558 13207 29564 13259
rect 29616 13207 29622 13259
rect 32054 13207 32060 13259
rect 32112 13207 32118 13259
rect 34550 13207 34556 13259
rect 34608 13207 34614 13259
rect 37046 13207 37052 13259
rect 37104 13207 37110 13259
rect 39542 13207 39548 13259
rect 39600 13207 39606 13259
rect 42038 13207 42044 13259
rect 42096 13207 42102 13259
rect 44534 13207 44540 13259
rect 44592 13207 44598 13259
rect 47030 13207 47036 13259
rect 47088 13207 47094 13259
rect 49526 13207 49532 13259
rect 49584 13207 49590 13259
rect 52022 13207 52028 13259
rect 52080 13207 52086 13259
rect 54518 13207 54524 13259
rect 54576 13207 54582 13259
rect 57014 13207 57020 13259
rect 57072 13207 57078 13259
rect 59510 13207 59516 13259
rect 59568 13207 59574 13259
rect 62006 13207 62012 13259
rect 62064 13207 62070 13259
rect 64502 13207 64508 13259
rect 64560 13207 64566 13259
rect 66998 13207 67004 13259
rect 67056 13207 67062 13259
rect 69494 13207 69500 13259
rect 69552 13207 69558 13259
rect 71990 13207 71996 13259
rect 72048 13207 72054 13259
rect 74486 13207 74492 13259
rect 74544 13207 74550 13259
rect 76982 13207 76988 13259
rect 77040 13207 77046 13259
rect 79478 13207 79484 13259
rect 79536 13207 79542 13259
rect 81974 13207 81980 13259
rect 82032 13207 82038 13259
rect 84470 13207 84476 13259
rect 84528 13207 84534 13259
rect 86966 13207 86972 13259
rect 87024 13207 87030 13259
rect 89462 13207 89468 13259
rect 89520 13207 89526 13259
rect 91958 13207 91964 13259
rect 92016 13207 92022 13259
rect 94454 13207 94460 13259
rect 94512 13207 94518 13259
rect 96950 13207 96956 13259
rect 97008 13207 97014 13259
rect 99446 13207 99452 13259
rect 99504 13207 99510 13259
rect 101942 13207 101948 13259
rect 102000 13207 102006 13259
rect 104438 13207 104444 13259
rect 104496 13207 104502 13259
rect 106934 13207 106940 13259
rect 106992 13207 106998 13259
rect 1794 13122 1800 13174
rect 1852 13122 1858 13174
rect 1794 12786 1800 12838
rect 1852 12786 1858 12838
rect 1794 12450 1800 12502
rect 1852 12450 1858 12502
rect 1794 12114 1800 12166
rect 1852 12114 1858 12166
rect 1794 11778 1800 11830
rect 1852 11778 1858 11830
rect 1794 11442 1800 11494
rect 1852 11442 1858 11494
rect 1794 11106 1800 11158
rect 1852 11106 1858 11158
rect 1794 10770 1800 10822
rect 1852 10770 1858 10822
rect 1794 10434 1800 10486
rect 1852 10434 1858 10486
rect 1794 10098 1800 10150
rect 1852 10098 1858 10150
rect 1794 9762 1800 9814
rect 1852 9762 1858 9814
rect 1794 9426 1800 9478
rect 1852 9426 1858 9478
rect 122785 9195 122813 24586
rect 122865 10753 122893 24586
rect 122945 12023 122973 24586
rect 123025 13581 123053 24586
rect 123105 14851 123133 24586
rect 123185 16409 123213 24586
rect 123265 17679 123293 24586
rect 123345 19237 123373 24586
rect 136940 24546 136946 24598
rect 136998 24546 137004 24598
rect 136940 24210 136946 24262
rect 136998 24210 137004 24262
rect 136940 23874 136946 23926
rect 136998 23874 137004 23926
rect 136940 23538 136946 23590
rect 136998 23538 137004 23590
rect 136940 23202 136946 23254
rect 136998 23202 137004 23254
rect 136940 22866 136946 22918
rect 136998 22866 137004 22918
rect 136940 22530 136946 22582
rect 136998 22530 137004 22582
rect 136940 22194 136946 22246
rect 136998 22194 137004 22246
rect 136940 21858 136946 21910
rect 136998 21858 137004 21910
rect 136940 21522 136946 21574
rect 136998 21522 137004 21574
rect 136940 21186 136946 21238
rect 136998 21186 137004 21238
rect 136940 20850 136946 20902
rect 136998 20850 137004 20902
rect 136940 20514 136946 20566
rect 136998 20514 137004 20566
rect 136940 20178 136946 20230
rect 136998 20178 137004 20230
rect 136940 19842 136946 19894
rect 136998 19842 137004 19894
rect 136940 19506 136946 19558
rect 136998 19506 137004 19558
rect 123327 19185 123333 19237
rect 123385 19185 123391 19237
rect 136940 19170 136946 19222
rect 136998 19170 137004 19222
rect 136940 18834 136946 18886
rect 136998 18834 137004 18886
rect 136940 18498 136946 18550
rect 136998 18498 137004 18550
rect 136940 18162 136946 18214
rect 136998 18162 137004 18214
rect 136940 17826 136946 17878
rect 136998 17826 137004 17878
rect 123247 17627 123253 17679
rect 123305 17627 123311 17679
rect 136940 17490 136946 17542
rect 136998 17490 137004 17542
rect 136940 17154 136946 17206
rect 136998 17154 137004 17206
rect 136940 16818 136946 16870
rect 136998 16818 137004 16870
rect 136940 16482 136946 16534
rect 136998 16482 137004 16534
rect 123167 16357 123173 16409
rect 123225 16357 123231 16409
rect 136940 16146 136946 16198
rect 136998 16146 137004 16198
rect 136940 15810 136946 15862
rect 136998 15810 137004 15862
rect 136940 15474 136946 15526
rect 136998 15474 137004 15526
rect 136940 15138 136946 15190
rect 136998 15138 137004 15190
rect 123087 14799 123093 14851
rect 123145 14799 123151 14851
rect 136940 14802 136946 14854
rect 136998 14802 137004 14854
rect 136940 14466 136946 14518
rect 136998 14466 137004 14518
rect 136940 14130 136946 14182
rect 136998 14130 137004 14182
rect 136940 13794 136946 13846
rect 136998 13794 137004 13846
rect 123007 13529 123013 13581
rect 123065 13529 123071 13581
rect 136940 13458 136946 13510
rect 136998 13458 137004 13510
rect 136940 13122 136946 13174
rect 136998 13122 137004 13174
rect 136940 12786 136946 12838
rect 136998 12786 137004 12838
rect 136940 12450 136946 12502
rect 136998 12450 137004 12502
rect 136940 12114 136946 12166
rect 136998 12114 137004 12166
rect 122927 11971 122933 12023
rect 122985 11971 122991 12023
rect 136940 11778 136946 11830
rect 136998 11778 137004 11830
rect 136940 11442 136946 11494
rect 136998 11442 137004 11494
rect 136940 11106 136946 11158
rect 136998 11106 137004 11158
rect 136940 10770 136946 10822
rect 136998 10770 137004 10822
rect 122847 10701 122853 10753
rect 122905 10701 122911 10753
rect 136940 10434 136946 10486
rect 136998 10434 137004 10486
rect 136940 10098 136946 10150
rect 136998 10098 137004 10150
rect 136940 9762 136946 9814
rect 136998 9762 137004 9814
rect 136940 9426 136946 9478
rect 136998 9426 137004 9478
rect 122767 9143 122773 9195
rect 122825 9143 122831 9195
rect 1794 9090 1800 9142
rect 1852 9090 1858 9142
rect 136940 9090 136946 9142
rect 136998 9090 137004 9142
rect 1794 8754 1800 8806
rect 1852 8754 1858 8806
rect 136940 8754 136946 8806
rect 136998 8754 137004 8806
rect 1794 8418 1800 8470
rect 1852 8418 1858 8470
rect 136940 8418 136946 8470
rect 136998 8418 137004 8470
rect 1794 8082 1800 8134
rect 1852 8082 1858 8134
rect 136940 8082 136946 8134
rect 136998 8082 137004 8134
rect 1794 7746 1800 7798
rect 1852 7746 1858 7798
rect 136940 7746 136946 7798
rect 136998 7746 137004 7798
rect 1794 7410 1800 7462
rect 1852 7410 1858 7462
rect 136940 7410 136946 7462
rect 136998 7410 137004 7462
rect 1794 7074 1800 7126
rect 1852 7074 1858 7126
rect 136940 7074 136946 7126
rect 136998 7074 137004 7126
rect 1794 6738 1800 6790
rect 1852 6738 1858 6790
rect 136940 6738 136946 6790
rect 136998 6738 137004 6790
rect 1794 6402 1800 6454
rect 1852 6402 1858 6454
rect 136940 6402 136946 6454
rect 136998 6402 137004 6454
rect 1794 6066 1800 6118
rect 1852 6066 1858 6118
rect 136940 6066 136946 6118
rect 136998 6066 137004 6118
rect 1794 5730 1800 5782
rect 1852 5730 1858 5782
rect 136940 5730 136946 5782
rect 136998 5730 137004 5782
rect 1794 5394 1800 5446
rect 1852 5394 1858 5446
rect 136940 5394 136946 5446
rect 136998 5394 137004 5446
rect 1794 5058 1800 5110
rect 1852 5058 1858 5110
rect 136940 5058 136946 5110
rect 136998 5058 137004 5110
rect 1794 4722 1800 4774
rect 1852 4722 1858 4774
rect 136940 4722 136946 4774
rect 136998 4722 137004 4774
rect 1794 4386 1800 4438
rect 1852 4386 1858 4438
rect 136940 4386 136946 4438
rect 136998 4386 137004 4438
rect 1794 4050 1800 4102
rect 1852 4050 1858 4102
rect 136940 4050 136946 4102
rect 136998 4050 137004 4102
rect 1794 3714 1800 3766
rect 1852 3714 1858 3766
rect 136940 3714 136946 3766
rect 136998 3714 137004 3766
rect 1794 3378 1800 3430
rect 1852 3378 1858 3430
rect 136940 3378 136946 3430
rect 136998 3378 137004 3430
rect 1794 3042 1800 3094
rect 1852 3042 1858 3094
rect 136940 3042 136946 3094
rect 136998 3042 137004 3094
rect 1794 2706 1800 2758
rect 1852 2706 1858 2758
rect 136940 2706 136946 2758
rect 136998 2706 137004 2758
rect 1794 2370 1800 2422
rect 1852 2370 1858 2422
rect 136940 2370 136946 2422
rect 136998 2370 137004 2422
rect 1794 2034 1800 2086
rect 1852 2034 1858 2086
rect 136940 2034 136946 2086
rect 136998 2034 137004 2086
rect 1714 1750 137084 1836
rect 1714 1698 2136 1750
rect 2188 1741 3816 1750
rect 3868 1741 5496 1750
rect 5548 1741 7176 1750
rect 7228 1741 8856 1750
rect 8908 1741 10536 1750
rect 10588 1741 12216 1750
rect 12268 1741 13896 1750
rect 13948 1741 15576 1750
rect 15628 1741 17256 1750
rect 17308 1741 18936 1750
rect 18988 1741 20616 1750
rect 20668 1741 22296 1750
rect 22348 1741 23976 1750
rect 24028 1741 25656 1750
rect 25708 1741 27336 1750
rect 27388 1741 29016 1750
rect 29068 1741 30696 1750
rect 30748 1741 32376 1750
rect 32428 1741 34056 1750
rect 34108 1741 35736 1750
rect 35788 1741 37416 1750
rect 37468 1741 39096 1750
rect 39148 1741 40776 1750
rect 40828 1741 42456 1750
rect 42508 1741 44136 1750
rect 44188 1741 45816 1750
rect 45868 1741 47496 1750
rect 47548 1741 49176 1750
rect 49228 1741 50856 1750
rect 50908 1741 52536 1750
rect 52588 1741 54216 1750
rect 54268 1741 55896 1750
rect 55948 1741 57576 1750
rect 57628 1741 59256 1750
rect 59308 1741 60936 1750
rect 60988 1741 62616 1750
rect 62668 1741 64296 1750
rect 64348 1741 65976 1750
rect 66028 1741 67656 1750
rect 67708 1741 69336 1750
rect 69388 1741 71016 1750
rect 71068 1741 72696 1750
rect 72748 1741 74376 1750
rect 74428 1741 76056 1750
rect 76108 1741 77736 1750
rect 77788 1741 79416 1750
rect 79468 1741 81096 1750
rect 81148 1741 82776 1750
rect 82828 1741 84456 1750
rect 84508 1741 86136 1750
rect 86188 1741 87816 1750
rect 87868 1741 89496 1750
rect 89548 1741 91176 1750
rect 91228 1741 92856 1750
rect 92908 1741 94536 1750
rect 94588 1741 96216 1750
rect 96268 1741 97896 1750
rect 97948 1741 99576 1750
rect 99628 1741 101256 1750
rect 101308 1741 102936 1750
rect 102988 1741 104616 1750
rect 104668 1741 106296 1750
rect 106348 1741 107976 1750
rect 108028 1741 109656 1750
rect 109708 1741 111336 1750
rect 111388 1741 113016 1750
rect 113068 1741 114696 1750
rect 114748 1741 116376 1750
rect 116428 1741 118056 1750
rect 118108 1741 119736 1750
rect 119788 1741 121416 1750
rect 121468 1741 123096 1750
rect 123148 1741 124776 1750
rect 124828 1741 126456 1750
rect 126508 1741 128136 1750
rect 128188 1741 129816 1750
rect 129868 1741 131496 1750
rect 131548 1741 133176 1750
rect 133228 1741 134856 1750
rect 134908 1741 136536 1750
rect 2188 1707 2481 1741
rect 2515 1707 2817 1741
rect 2851 1707 3153 1741
rect 3187 1707 3489 1741
rect 3523 1707 3816 1741
rect 3868 1707 4161 1741
rect 4195 1707 4497 1741
rect 4531 1707 4833 1741
rect 4867 1707 5169 1741
rect 5203 1707 5496 1741
rect 5548 1707 5841 1741
rect 5875 1707 6177 1741
rect 6211 1707 6513 1741
rect 6547 1707 6849 1741
rect 6883 1707 7176 1741
rect 7228 1707 7521 1741
rect 7555 1707 7857 1741
rect 7891 1707 8193 1741
rect 8227 1707 8529 1741
rect 8563 1707 8856 1741
rect 8908 1707 9201 1741
rect 9235 1707 9537 1741
rect 9571 1707 9873 1741
rect 9907 1707 10209 1741
rect 10243 1707 10536 1741
rect 10588 1707 10881 1741
rect 10915 1707 11217 1741
rect 11251 1707 11553 1741
rect 11587 1707 11889 1741
rect 11923 1707 12216 1741
rect 12268 1707 12561 1741
rect 12595 1707 12897 1741
rect 12931 1707 13233 1741
rect 13267 1707 13569 1741
rect 13603 1707 13896 1741
rect 13948 1707 14241 1741
rect 14275 1707 14577 1741
rect 14611 1707 14913 1741
rect 14947 1707 15249 1741
rect 15283 1707 15576 1741
rect 15628 1707 15921 1741
rect 15955 1707 16257 1741
rect 16291 1707 16593 1741
rect 16627 1707 16929 1741
rect 16963 1707 17256 1741
rect 17308 1707 17601 1741
rect 17635 1707 17937 1741
rect 17971 1707 18273 1741
rect 18307 1707 18609 1741
rect 18643 1707 18936 1741
rect 18988 1707 19281 1741
rect 19315 1707 19617 1741
rect 19651 1707 19953 1741
rect 19987 1707 20289 1741
rect 20323 1707 20616 1741
rect 20668 1707 20961 1741
rect 20995 1707 21297 1741
rect 21331 1707 21633 1741
rect 21667 1707 21969 1741
rect 22003 1707 22296 1741
rect 22348 1707 22641 1741
rect 22675 1707 22977 1741
rect 23011 1707 23313 1741
rect 23347 1707 23649 1741
rect 23683 1707 23976 1741
rect 24028 1707 24321 1741
rect 24355 1707 24657 1741
rect 24691 1707 24993 1741
rect 25027 1707 25329 1741
rect 25363 1707 25656 1741
rect 25708 1707 26001 1741
rect 26035 1707 26337 1741
rect 26371 1707 26673 1741
rect 26707 1707 27009 1741
rect 27043 1707 27336 1741
rect 27388 1707 27681 1741
rect 27715 1707 28017 1741
rect 28051 1707 28353 1741
rect 28387 1707 28689 1741
rect 28723 1707 29016 1741
rect 29068 1707 29361 1741
rect 29395 1707 29697 1741
rect 29731 1707 30033 1741
rect 30067 1707 30369 1741
rect 30403 1707 30696 1741
rect 30748 1707 31041 1741
rect 31075 1707 31377 1741
rect 31411 1707 31713 1741
rect 31747 1707 32049 1741
rect 32083 1707 32376 1741
rect 32428 1707 32721 1741
rect 32755 1707 33057 1741
rect 33091 1707 33393 1741
rect 33427 1707 33729 1741
rect 33763 1707 34056 1741
rect 34108 1707 34401 1741
rect 34435 1707 34737 1741
rect 34771 1707 35073 1741
rect 35107 1707 35409 1741
rect 35443 1707 35736 1741
rect 35788 1707 36081 1741
rect 36115 1707 36417 1741
rect 36451 1707 36753 1741
rect 36787 1707 37089 1741
rect 37123 1707 37416 1741
rect 37468 1707 37761 1741
rect 37795 1707 38097 1741
rect 38131 1707 38433 1741
rect 38467 1707 38769 1741
rect 38803 1707 39096 1741
rect 39148 1707 39441 1741
rect 39475 1707 39777 1741
rect 39811 1707 40113 1741
rect 40147 1707 40449 1741
rect 40483 1707 40776 1741
rect 40828 1707 41121 1741
rect 41155 1707 41457 1741
rect 41491 1707 41793 1741
rect 41827 1707 42129 1741
rect 42163 1707 42456 1741
rect 42508 1707 42801 1741
rect 42835 1707 43137 1741
rect 43171 1707 43473 1741
rect 43507 1707 43809 1741
rect 43843 1707 44136 1741
rect 44188 1707 44481 1741
rect 44515 1707 44817 1741
rect 44851 1707 45153 1741
rect 45187 1707 45489 1741
rect 45523 1707 45816 1741
rect 45868 1707 46161 1741
rect 46195 1707 46497 1741
rect 46531 1707 46833 1741
rect 46867 1707 47169 1741
rect 47203 1707 47496 1741
rect 47548 1707 47841 1741
rect 47875 1707 48177 1741
rect 48211 1707 48513 1741
rect 48547 1707 48849 1741
rect 48883 1707 49176 1741
rect 49228 1707 49521 1741
rect 49555 1707 49857 1741
rect 49891 1707 50193 1741
rect 50227 1707 50529 1741
rect 50563 1707 50856 1741
rect 50908 1707 51201 1741
rect 51235 1707 51537 1741
rect 51571 1707 51873 1741
rect 51907 1707 52209 1741
rect 52243 1707 52536 1741
rect 52588 1707 52881 1741
rect 52915 1707 53217 1741
rect 53251 1707 53553 1741
rect 53587 1707 53889 1741
rect 53923 1707 54216 1741
rect 54268 1707 54561 1741
rect 54595 1707 54897 1741
rect 54931 1707 55233 1741
rect 55267 1707 55569 1741
rect 55603 1707 55896 1741
rect 55948 1707 56241 1741
rect 56275 1707 56577 1741
rect 56611 1707 56913 1741
rect 56947 1707 57249 1741
rect 57283 1707 57576 1741
rect 57628 1707 57921 1741
rect 57955 1707 58257 1741
rect 58291 1707 58593 1741
rect 58627 1707 58929 1741
rect 58963 1707 59256 1741
rect 59308 1707 59601 1741
rect 59635 1707 59937 1741
rect 59971 1707 60273 1741
rect 60307 1707 60609 1741
rect 60643 1707 60936 1741
rect 60988 1707 61281 1741
rect 61315 1707 61617 1741
rect 61651 1707 61953 1741
rect 61987 1707 62289 1741
rect 62323 1707 62616 1741
rect 62668 1707 62961 1741
rect 62995 1707 63297 1741
rect 63331 1707 63633 1741
rect 63667 1707 63969 1741
rect 64003 1707 64296 1741
rect 64348 1707 64641 1741
rect 64675 1707 64977 1741
rect 65011 1707 65313 1741
rect 65347 1707 65649 1741
rect 65683 1707 65976 1741
rect 66028 1707 66321 1741
rect 66355 1707 66657 1741
rect 66691 1707 66993 1741
rect 67027 1707 67329 1741
rect 67363 1707 67656 1741
rect 67708 1707 68001 1741
rect 68035 1707 68337 1741
rect 68371 1707 68673 1741
rect 68707 1707 69009 1741
rect 69043 1707 69336 1741
rect 69388 1707 69681 1741
rect 69715 1707 70017 1741
rect 70051 1707 70353 1741
rect 70387 1707 70689 1741
rect 70723 1707 71016 1741
rect 71068 1707 71361 1741
rect 71395 1707 71697 1741
rect 71731 1707 72033 1741
rect 72067 1707 72369 1741
rect 72403 1707 72696 1741
rect 72748 1707 73041 1741
rect 73075 1707 73377 1741
rect 73411 1707 73713 1741
rect 73747 1707 74049 1741
rect 74083 1707 74376 1741
rect 74428 1707 74721 1741
rect 74755 1707 75057 1741
rect 75091 1707 75393 1741
rect 75427 1707 75729 1741
rect 75763 1707 76056 1741
rect 76108 1707 76401 1741
rect 76435 1707 76737 1741
rect 76771 1707 77073 1741
rect 77107 1707 77409 1741
rect 77443 1707 77736 1741
rect 77788 1707 78081 1741
rect 78115 1707 78417 1741
rect 78451 1707 78753 1741
rect 78787 1707 79089 1741
rect 79123 1707 79416 1741
rect 79468 1707 79761 1741
rect 79795 1707 80097 1741
rect 80131 1707 80433 1741
rect 80467 1707 80769 1741
rect 80803 1707 81096 1741
rect 81148 1707 81441 1741
rect 81475 1707 81777 1741
rect 81811 1707 82113 1741
rect 82147 1707 82449 1741
rect 82483 1707 82776 1741
rect 82828 1707 83121 1741
rect 83155 1707 83457 1741
rect 83491 1707 83793 1741
rect 83827 1707 84129 1741
rect 84163 1707 84456 1741
rect 84508 1707 84801 1741
rect 84835 1707 85137 1741
rect 85171 1707 85473 1741
rect 85507 1707 85809 1741
rect 85843 1707 86136 1741
rect 86188 1707 86481 1741
rect 86515 1707 86817 1741
rect 86851 1707 87153 1741
rect 87187 1707 87489 1741
rect 87523 1707 87816 1741
rect 87868 1707 88161 1741
rect 88195 1707 88497 1741
rect 88531 1707 88833 1741
rect 88867 1707 89169 1741
rect 89203 1707 89496 1741
rect 89548 1707 89841 1741
rect 89875 1707 90177 1741
rect 90211 1707 90513 1741
rect 90547 1707 90849 1741
rect 90883 1707 91176 1741
rect 91228 1707 91521 1741
rect 91555 1707 91857 1741
rect 91891 1707 92193 1741
rect 92227 1707 92529 1741
rect 92563 1707 92856 1741
rect 92908 1707 93201 1741
rect 93235 1707 93537 1741
rect 93571 1707 93873 1741
rect 93907 1707 94209 1741
rect 94243 1707 94536 1741
rect 94588 1707 94881 1741
rect 94915 1707 95217 1741
rect 95251 1707 95553 1741
rect 95587 1707 95889 1741
rect 95923 1707 96216 1741
rect 96268 1707 96561 1741
rect 96595 1707 96897 1741
rect 96931 1707 97233 1741
rect 97267 1707 97569 1741
rect 97603 1707 97896 1741
rect 97948 1707 98241 1741
rect 98275 1707 98577 1741
rect 98611 1707 98913 1741
rect 98947 1707 99249 1741
rect 99283 1707 99576 1741
rect 99628 1707 99921 1741
rect 99955 1707 100257 1741
rect 100291 1707 100593 1741
rect 100627 1707 100929 1741
rect 100963 1707 101256 1741
rect 101308 1707 101601 1741
rect 101635 1707 101937 1741
rect 101971 1707 102273 1741
rect 102307 1707 102609 1741
rect 102643 1707 102936 1741
rect 102988 1707 103281 1741
rect 103315 1707 103617 1741
rect 103651 1707 103953 1741
rect 103987 1707 104289 1741
rect 104323 1707 104616 1741
rect 104668 1707 104961 1741
rect 104995 1707 105297 1741
rect 105331 1707 105633 1741
rect 105667 1707 105969 1741
rect 106003 1707 106296 1741
rect 106348 1707 106641 1741
rect 106675 1707 106977 1741
rect 107011 1707 107313 1741
rect 107347 1707 107649 1741
rect 107683 1707 107976 1741
rect 108028 1707 108321 1741
rect 108355 1707 108657 1741
rect 108691 1707 108993 1741
rect 109027 1707 109329 1741
rect 109363 1707 109656 1741
rect 109708 1707 110001 1741
rect 110035 1707 110337 1741
rect 110371 1707 110673 1741
rect 110707 1707 111009 1741
rect 111043 1707 111336 1741
rect 111388 1707 111681 1741
rect 111715 1707 112017 1741
rect 112051 1707 112353 1741
rect 112387 1707 112689 1741
rect 112723 1707 113016 1741
rect 113068 1707 113361 1741
rect 113395 1707 113697 1741
rect 113731 1707 114033 1741
rect 114067 1707 114369 1741
rect 114403 1707 114696 1741
rect 114748 1707 115041 1741
rect 115075 1707 115377 1741
rect 115411 1707 115713 1741
rect 115747 1707 116049 1741
rect 116083 1707 116376 1741
rect 116428 1707 116721 1741
rect 116755 1707 117057 1741
rect 117091 1707 117393 1741
rect 117427 1707 117729 1741
rect 117763 1707 118056 1741
rect 118108 1707 118401 1741
rect 118435 1707 118737 1741
rect 118771 1707 119073 1741
rect 119107 1707 119409 1741
rect 119443 1707 119736 1741
rect 119788 1707 120081 1741
rect 120115 1707 120417 1741
rect 120451 1707 120753 1741
rect 120787 1707 121089 1741
rect 121123 1707 121416 1741
rect 121468 1707 121761 1741
rect 121795 1707 122097 1741
rect 122131 1707 122433 1741
rect 122467 1707 122769 1741
rect 122803 1707 123096 1741
rect 123148 1707 123441 1741
rect 123475 1707 123777 1741
rect 123811 1707 124113 1741
rect 124147 1707 124449 1741
rect 124483 1707 124776 1741
rect 124828 1707 125121 1741
rect 125155 1707 125457 1741
rect 125491 1707 125793 1741
rect 125827 1707 126129 1741
rect 126163 1707 126456 1741
rect 126508 1707 126801 1741
rect 126835 1707 127137 1741
rect 127171 1707 127473 1741
rect 127507 1707 127809 1741
rect 127843 1707 128136 1741
rect 128188 1707 128481 1741
rect 128515 1707 128817 1741
rect 128851 1707 129153 1741
rect 129187 1707 129489 1741
rect 129523 1707 129816 1741
rect 129868 1707 130161 1741
rect 130195 1707 130497 1741
rect 130531 1707 130833 1741
rect 130867 1707 131169 1741
rect 131203 1707 131496 1741
rect 131548 1707 131841 1741
rect 131875 1707 132177 1741
rect 132211 1707 132513 1741
rect 132547 1707 132849 1741
rect 132883 1707 133176 1741
rect 133228 1707 133521 1741
rect 133555 1707 133857 1741
rect 133891 1707 134193 1741
rect 134227 1707 134529 1741
rect 134563 1707 134856 1741
rect 134908 1707 135201 1741
rect 135235 1707 135537 1741
rect 135571 1707 135873 1741
rect 135907 1707 136209 1741
rect 136243 1707 136536 1741
rect 2188 1698 3816 1707
rect 3868 1698 5496 1707
rect 5548 1698 7176 1707
rect 7228 1698 8856 1707
rect 8908 1698 10536 1707
rect 10588 1698 12216 1707
rect 12268 1698 13896 1707
rect 13948 1698 15576 1707
rect 15628 1698 17256 1707
rect 17308 1698 18936 1707
rect 18988 1698 20616 1707
rect 20668 1698 22296 1707
rect 22348 1698 23976 1707
rect 24028 1698 25656 1707
rect 25708 1698 27336 1707
rect 27388 1698 29016 1707
rect 29068 1698 30696 1707
rect 30748 1698 32376 1707
rect 32428 1698 34056 1707
rect 34108 1698 35736 1707
rect 35788 1698 37416 1707
rect 37468 1698 39096 1707
rect 39148 1698 40776 1707
rect 40828 1698 42456 1707
rect 42508 1698 44136 1707
rect 44188 1698 45816 1707
rect 45868 1698 47496 1707
rect 47548 1698 49176 1707
rect 49228 1698 50856 1707
rect 50908 1698 52536 1707
rect 52588 1698 54216 1707
rect 54268 1698 55896 1707
rect 55948 1698 57576 1707
rect 57628 1698 59256 1707
rect 59308 1698 60936 1707
rect 60988 1698 62616 1707
rect 62668 1698 64296 1707
rect 64348 1698 65976 1707
rect 66028 1698 67656 1707
rect 67708 1698 69336 1707
rect 69388 1698 71016 1707
rect 71068 1698 72696 1707
rect 72748 1698 74376 1707
rect 74428 1698 76056 1707
rect 76108 1698 77736 1707
rect 77788 1698 79416 1707
rect 79468 1698 81096 1707
rect 81148 1698 82776 1707
rect 82828 1698 84456 1707
rect 84508 1698 86136 1707
rect 86188 1698 87816 1707
rect 87868 1698 89496 1707
rect 89548 1698 91176 1707
rect 91228 1698 92856 1707
rect 92908 1698 94536 1707
rect 94588 1698 96216 1707
rect 96268 1698 97896 1707
rect 97948 1698 99576 1707
rect 99628 1698 101256 1707
rect 101308 1698 102936 1707
rect 102988 1698 104616 1707
rect 104668 1698 106296 1707
rect 106348 1698 107976 1707
rect 108028 1698 109656 1707
rect 109708 1698 111336 1707
rect 111388 1698 113016 1707
rect 113068 1698 114696 1707
rect 114748 1698 116376 1707
rect 116428 1698 118056 1707
rect 118108 1698 119736 1707
rect 119788 1698 121416 1707
rect 121468 1698 123096 1707
rect 123148 1698 124776 1707
rect 124828 1698 126456 1707
rect 126508 1698 128136 1707
rect 128188 1698 129816 1707
rect 129868 1698 131496 1707
rect 131548 1698 133176 1707
rect 133228 1698 134856 1707
rect 134908 1698 136536 1707
rect 136588 1698 137084 1750
rect 1714 1612 137084 1698
<< via1 >>
rect 2136 132050 2188 132059
rect 3816 132050 3868 132059
rect 5496 132050 5548 132059
rect 7176 132050 7228 132059
rect 8856 132050 8908 132059
rect 10536 132050 10588 132059
rect 12216 132050 12268 132059
rect 13896 132050 13948 132059
rect 15576 132050 15628 132059
rect 17256 132050 17308 132059
rect 18936 132050 18988 132059
rect 20616 132050 20668 132059
rect 22296 132050 22348 132059
rect 23976 132050 24028 132059
rect 25656 132050 25708 132059
rect 27336 132050 27388 132059
rect 29016 132050 29068 132059
rect 30696 132050 30748 132059
rect 32376 132050 32428 132059
rect 34056 132050 34108 132059
rect 35736 132050 35788 132059
rect 37416 132050 37468 132059
rect 39096 132050 39148 132059
rect 40776 132050 40828 132059
rect 42456 132050 42508 132059
rect 44136 132050 44188 132059
rect 45816 132050 45868 132059
rect 47496 132050 47548 132059
rect 49176 132050 49228 132059
rect 50856 132050 50908 132059
rect 52536 132050 52588 132059
rect 54216 132050 54268 132059
rect 55896 132050 55948 132059
rect 57576 132050 57628 132059
rect 59256 132050 59308 132059
rect 60936 132050 60988 132059
rect 62616 132050 62668 132059
rect 64296 132050 64348 132059
rect 65976 132050 66028 132059
rect 67656 132050 67708 132059
rect 69336 132050 69388 132059
rect 71016 132050 71068 132059
rect 72696 132050 72748 132059
rect 74376 132050 74428 132059
rect 76056 132050 76108 132059
rect 77736 132050 77788 132059
rect 79416 132050 79468 132059
rect 81096 132050 81148 132059
rect 82776 132050 82828 132059
rect 84456 132050 84508 132059
rect 86136 132050 86188 132059
rect 87816 132050 87868 132059
rect 89496 132050 89548 132059
rect 91176 132050 91228 132059
rect 92856 132050 92908 132059
rect 94536 132050 94588 132059
rect 96216 132050 96268 132059
rect 97896 132050 97948 132059
rect 99576 132050 99628 132059
rect 101256 132050 101308 132059
rect 102936 132050 102988 132059
rect 104616 132050 104668 132059
rect 106296 132050 106348 132059
rect 107976 132050 108028 132059
rect 109656 132050 109708 132059
rect 111336 132050 111388 132059
rect 113016 132050 113068 132059
rect 114696 132050 114748 132059
rect 116376 132050 116428 132059
rect 118056 132050 118108 132059
rect 119736 132050 119788 132059
rect 121416 132050 121468 132059
rect 123096 132050 123148 132059
rect 124776 132050 124828 132059
rect 126456 132050 126508 132059
rect 128136 132050 128188 132059
rect 129816 132050 129868 132059
rect 131496 132050 131548 132059
rect 133176 132050 133228 132059
rect 134856 132050 134908 132059
rect 136536 132050 136588 132059
rect 2136 132016 2145 132050
rect 2145 132016 2179 132050
rect 2179 132016 2188 132050
rect 3816 132016 3825 132050
rect 3825 132016 3859 132050
rect 3859 132016 3868 132050
rect 5496 132016 5505 132050
rect 5505 132016 5539 132050
rect 5539 132016 5548 132050
rect 7176 132016 7185 132050
rect 7185 132016 7219 132050
rect 7219 132016 7228 132050
rect 8856 132016 8865 132050
rect 8865 132016 8899 132050
rect 8899 132016 8908 132050
rect 10536 132016 10545 132050
rect 10545 132016 10579 132050
rect 10579 132016 10588 132050
rect 12216 132016 12225 132050
rect 12225 132016 12259 132050
rect 12259 132016 12268 132050
rect 13896 132016 13905 132050
rect 13905 132016 13939 132050
rect 13939 132016 13948 132050
rect 15576 132016 15585 132050
rect 15585 132016 15619 132050
rect 15619 132016 15628 132050
rect 17256 132016 17265 132050
rect 17265 132016 17299 132050
rect 17299 132016 17308 132050
rect 18936 132016 18945 132050
rect 18945 132016 18979 132050
rect 18979 132016 18988 132050
rect 20616 132016 20625 132050
rect 20625 132016 20659 132050
rect 20659 132016 20668 132050
rect 22296 132016 22305 132050
rect 22305 132016 22339 132050
rect 22339 132016 22348 132050
rect 23976 132016 23985 132050
rect 23985 132016 24019 132050
rect 24019 132016 24028 132050
rect 25656 132016 25665 132050
rect 25665 132016 25699 132050
rect 25699 132016 25708 132050
rect 27336 132016 27345 132050
rect 27345 132016 27379 132050
rect 27379 132016 27388 132050
rect 29016 132016 29025 132050
rect 29025 132016 29059 132050
rect 29059 132016 29068 132050
rect 30696 132016 30705 132050
rect 30705 132016 30739 132050
rect 30739 132016 30748 132050
rect 32376 132016 32385 132050
rect 32385 132016 32419 132050
rect 32419 132016 32428 132050
rect 34056 132016 34065 132050
rect 34065 132016 34099 132050
rect 34099 132016 34108 132050
rect 35736 132016 35745 132050
rect 35745 132016 35779 132050
rect 35779 132016 35788 132050
rect 37416 132016 37425 132050
rect 37425 132016 37459 132050
rect 37459 132016 37468 132050
rect 39096 132016 39105 132050
rect 39105 132016 39139 132050
rect 39139 132016 39148 132050
rect 40776 132016 40785 132050
rect 40785 132016 40819 132050
rect 40819 132016 40828 132050
rect 42456 132016 42465 132050
rect 42465 132016 42499 132050
rect 42499 132016 42508 132050
rect 44136 132016 44145 132050
rect 44145 132016 44179 132050
rect 44179 132016 44188 132050
rect 45816 132016 45825 132050
rect 45825 132016 45859 132050
rect 45859 132016 45868 132050
rect 47496 132016 47505 132050
rect 47505 132016 47539 132050
rect 47539 132016 47548 132050
rect 49176 132016 49185 132050
rect 49185 132016 49219 132050
rect 49219 132016 49228 132050
rect 50856 132016 50865 132050
rect 50865 132016 50899 132050
rect 50899 132016 50908 132050
rect 52536 132016 52545 132050
rect 52545 132016 52579 132050
rect 52579 132016 52588 132050
rect 54216 132016 54225 132050
rect 54225 132016 54259 132050
rect 54259 132016 54268 132050
rect 55896 132016 55905 132050
rect 55905 132016 55939 132050
rect 55939 132016 55948 132050
rect 57576 132016 57585 132050
rect 57585 132016 57619 132050
rect 57619 132016 57628 132050
rect 59256 132016 59265 132050
rect 59265 132016 59299 132050
rect 59299 132016 59308 132050
rect 60936 132016 60945 132050
rect 60945 132016 60979 132050
rect 60979 132016 60988 132050
rect 62616 132016 62625 132050
rect 62625 132016 62659 132050
rect 62659 132016 62668 132050
rect 64296 132016 64305 132050
rect 64305 132016 64339 132050
rect 64339 132016 64348 132050
rect 65976 132016 65985 132050
rect 65985 132016 66019 132050
rect 66019 132016 66028 132050
rect 67656 132016 67665 132050
rect 67665 132016 67699 132050
rect 67699 132016 67708 132050
rect 69336 132016 69345 132050
rect 69345 132016 69379 132050
rect 69379 132016 69388 132050
rect 71016 132016 71025 132050
rect 71025 132016 71059 132050
rect 71059 132016 71068 132050
rect 72696 132016 72705 132050
rect 72705 132016 72739 132050
rect 72739 132016 72748 132050
rect 74376 132016 74385 132050
rect 74385 132016 74419 132050
rect 74419 132016 74428 132050
rect 76056 132016 76065 132050
rect 76065 132016 76099 132050
rect 76099 132016 76108 132050
rect 77736 132016 77745 132050
rect 77745 132016 77779 132050
rect 77779 132016 77788 132050
rect 79416 132016 79425 132050
rect 79425 132016 79459 132050
rect 79459 132016 79468 132050
rect 81096 132016 81105 132050
rect 81105 132016 81139 132050
rect 81139 132016 81148 132050
rect 82776 132016 82785 132050
rect 82785 132016 82819 132050
rect 82819 132016 82828 132050
rect 84456 132016 84465 132050
rect 84465 132016 84499 132050
rect 84499 132016 84508 132050
rect 86136 132016 86145 132050
rect 86145 132016 86179 132050
rect 86179 132016 86188 132050
rect 87816 132016 87825 132050
rect 87825 132016 87859 132050
rect 87859 132016 87868 132050
rect 89496 132016 89505 132050
rect 89505 132016 89539 132050
rect 89539 132016 89548 132050
rect 91176 132016 91185 132050
rect 91185 132016 91219 132050
rect 91219 132016 91228 132050
rect 92856 132016 92865 132050
rect 92865 132016 92899 132050
rect 92899 132016 92908 132050
rect 94536 132016 94545 132050
rect 94545 132016 94579 132050
rect 94579 132016 94588 132050
rect 96216 132016 96225 132050
rect 96225 132016 96259 132050
rect 96259 132016 96268 132050
rect 97896 132016 97905 132050
rect 97905 132016 97939 132050
rect 97939 132016 97948 132050
rect 99576 132016 99585 132050
rect 99585 132016 99619 132050
rect 99619 132016 99628 132050
rect 101256 132016 101265 132050
rect 101265 132016 101299 132050
rect 101299 132016 101308 132050
rect 102936 132016 102945 132050
rect 102945 132016 102979 132050
rect 102979 132016 102988 132050
rect 104616 132016 104625 132050
rect 104625 132016 104659 132050
rect 104659 132016 104668 132050
rect 106296 132016 106305 132050
rect 106305 132016 106339 132050
rect 106339 132016 106348 132050
rect 107976 132016 107985 132050
rect 107985 132016 108019 132050
rect 108019 132016 108028 132050
rect 109656 132016 109665 132050
rect 109665 132016 109699 132050
rect 109699 132016 109708 132050
rect 111336 132016 111345 132050
rect 111345 132016 111379 132050
rect 111379 132016 111388 132050
rect 113016 132016 113025 132050
rect 113025 132016 113059 132050
rect 113059 132016 113068 132050
rect 114696 132016 114705 132050
rect 114705 132016 114739 132050
rect 114739 132016 114748 132050
rect 116376 132016 116385 132050
rect 116385 132016 116419 132050
rect 116419 132016 116428 132050
rect 118056 132016 118065 132050
rect 118065 132016 118099 132050
rect 118099 132016 118108 132050
rect 119736 132016 119745 132050
rect 119745 132016 119779 132050
rect 119779 132016 119788 132050
rect 121416 132016 121425 132050
rect 121425 132016 121459 132050
rect 121459 132016 121468 132050
rect 123096 132016 123105 132050
rect 123105 132016 123139 132050
rect 123139 132016 123148 132050
rect 124776 132016 124785 132050
rect 124785 132016 124819 132050
rect 124819 132016 124828 132050
rect 126456 132016 126465 132050
rect 126465 132016 126499 132050
rect 126499 132016 126508 132050
rect 128136 132016 128145 132050
rect 128145 132016 128179 132050
rect 128179 132016 128188 132050
rect 129816 132016 129825 132050
rect 129825 132016 129859 132050
rect 129859 132016 129868 132050
rect 131496 132016 131505 132050
rect 131505 132016 131539 132050
rect 131539 132016 131548 132050
rect 133176 132016 133185 132050
rect 133185 132016 133219 132050
rect 133219 132016 133228 132050
rect 134856 132016 134865 132050
rect 134865 132016 134899 132050
rect 134899 132016 134908 132050
rect 136536 132016 136545 132050
rect 136545 132016 136579 132050
rect 136579 132016 136588 132050
rect 2136 132007 2188 132016
rect 3816 132007 3868 132016
rect 5496 132007 5548 132016
rect 7176 132007 7228 132016
rect 8856 132007 8908 132016
rect 10536 132007 10588 132016
rect 12216 132007 12268 132016
rect 13896 132007 13948 132016
rect 15576 132007 15628 132016
rect 17256 132007 17308 132016
rect 18936 132007 18988 132016
rect 20616 132007 20668 132016
rect 22296 132007 22348 132016
rect 23976 132007 24028 132016
rect 25656 132007 25708 132016
rect 27336 132007 27388 132016
rect 29016 132007 29068 132016
rect 30696 132007 30748 132016
rect 32376 132007 32428 132016
rect 34056 132007 34108 132016
rect 35736 132007 35788 132016
rect 37416 132007 37468 132016
rect 39096 132007 39148 132016
rect 40776 132007 40828 132016
rect 42456 132007 42508 132016
rect 44136 132007 44188 132016
rect 45816 132007 45868 132016
rect 47496 132007 47548 132016
rect 49176 132007 49228 132016
rect 50856 132007 50908 132016
rect 52536 132007 52588 132016
rect 54216 132007 54268 132016
rect 55896 132007 55948 132016
rect 57576 132007 57628 132016
rect 59256 132007 59308 132016
rect 60936 132007 60988 132016
rect 62616 132007 62668 132016
rect 64296 132007 64348 132016
rect 65976 132007 66028 132016
rect 67656 132007 67708 132016
rect 69336 132007 69388 132016
rect 71016 132007 71068 132016
rect 72696 132007 72748 132016
rect 74376 132007 74428 132016
rect 76056 132007 76108 132016
rect 77736 132007 77788 132016
rect 79416 132007 79468 132016
rect 81096 132007 81148 132016
rect 82776 132007 82828 132016
rect 84456 132007 84508 132016
rect 86136 132007 86188 132016
rect 87816 132007 87868 132016
rect 89496 132007 89548 132016
rect 91176 132007 91228 132016
rect 92856 132007 92908 132016
rect 94536 132007 94588 132016
rect 96216 132007 96268 132016
rect 97896 132007 97948 132016
rect 99576 132007 99628 132016
rect 101256 132007 101308 132016
rect 102936 132007 102988 132016
rect 104616 132007 104668 132016
rect 106296 132007 106348 132016
rect 107976 132007 108028 132016
rect 109656 132007 109708 132016
rect 111336 132007 111388 132016
rect 113016 132007 113068 132016
rect 114696 132007 114748 132016
rect 116376 132007 116428 132016
rect 118056 132007 118108 132016
rect 119736 132007 119788 132016
rect 121416 132007 121468 132016
rect 123096 132007 123148 132016
rect 124776 132007 124828 132016
rect 126456 132007 126508 132016
rect 128136 132007 128188 132016
rect 129816 132007 129868 132016
rect 131496 132007 131548 132016
rect 133176 132007 133228 132016
rect 134856 132007 134908 132016
rect 136536 132007 136588 132016
rect 1800 131437 1852 131446
rect 1800 131403 1809 131437
rect 1809 131403 1843 131437
rect 1843 131403 1852 131437
rect 1800 131394 1852 131403
rect 136946 131437 136998 131446
rect 136946 131403 136955 131437
rect 136955 131403 136989 131437
rect 136989 131403 136998 131437
rect 136946 131394 136998 131403
rect 1800 131101 1852 131110
rect 1800 131067 1809 131101
rect 1809 131067 1843 131101
rect 1843 131067 1852 131101
rect 1800 131058 1852 131067
rect 136946 131101 136998 131110
rect 136946 131067 136955 131101
rect 136955 131067 136989 131101
rect 136989 131067 136998 131101
rect 136946 131058 136998 131067
rect 1800 130765 1852 130774
rect 1800 130731 1809 130765
rect 1809 130731 1843 130765
rect 1843 130731 1852 130765
rect 1800 130722 1852 130731
rect 136946 130765 136998 130774
rect 136946 130731 136955 130765
rect 136955 130731 136989 130765
rect 136989 130731 136998 130765
rect 136946 130722 136998 130731
rect 1800 130429 1852 130438
rect 1800 130395 1809 130429
rect 1809 130395 1843 130429
rect 1843 130395 1852 130429
rect 1800 130386 1852 130395
rect 136946 130429 136998 130438
rect 136946 130395 136955 130429
rect 136955 130395 136989 130429
rect 136989 130395 136998 130429
rect 136946 130386 136998 130395
rect 1800 130093 1852 130102
rect 1800 130059 1809 130093
rect 1809 130059 1843 130093
rect 1843 130059 1852 130093
rect 1800 130050 1852 130059
rect 136946 130093 136998 130102
rect 136946 130059 136955 130093
rect 136955 130059 136989 130093
rect 136989 130059 136998 130093
rect 136946 130050 136998 130059
rect 1800 129757 1852 129766
rect 1800 129723 1809 129757
rect 1809 129723 1843 129757
rect 1843 129723 1852 129757
rect 1800 129714 1852 129723
rect 136946 129757 136998 129766
rect 136946 129723 136955 129757
rect 136955 129723 136989 129757
rect 136989 129723 136998 129757
rect 136946 129714 136998 129723
rect 1800 129421 1852 129430
rect 1800 129387 1809 129421
rect 1809 129387 1843 129421
rect 1843 129387 1852 129421
rect 1800 129378 1852 129387
rect 136946 129421 136998 129430
rect 136946 129387 136955 129421
rect 136955 129387 136989 129421
rect 136989 129387 136998 129421
rect 136946 129378 136998 129387
rect 1800 129085 1852 129094
rect 1800 129051 1809 129085
rect 1809 129051 1843 129085
rect 1843 129051 1852 129085
rect 1800 129042 1852 129051
rect 136946 129085 136998 129094
rect 136946 129051 136955 129085
rect 136955 129051 136989 129085
rect 136989 129051 136998 129085
rect 136946 129042 136998 129051
rect 1800 128749 1852 128758
rect 1800 128715 1809 128749
rect 1809 128715 1843 128749
rect 1843 128715 1852 128749
rect 1800 128706 1852 128715
rect 136946 128749 136998 128758
rect 136946 128715 136955 128749
rect 136955 128715 136989 128749
rect 136989 128715 136998 128749
rect 136946 128706 136998 128715
rect 1800 128413 1852 128422
rect 1800 128379 1809 128413
rect 1809 128379 1843 128413
rect 1843 128379 1852 128413
rect 1800 128370 1852 128379
rect 136946 128413 136998 128422
rect 136946 128379 136955 128413
rect 136955 128379 136989 128413
rect 136989 128379 136998 128413
rect 136946 128370 136998 128379
rect 1800 128077 1852 128086
rect 1800 128043 1809 128077
rect 1809 128043 1843 128077
rect 1843 128043 1852 128077
rect 1800 128034 1852 128043
rect 136946 128077 136998 128086
rect 136946 128043 136955 128077
rect 136955 128043 136989 128077
rect 136989 128043 136998 128077
rect 136946 128034 136998 128043
rect 1800 127741 1852 127750
rect 1800 127707 1809 127741
rect 1809 127707 1843 127741
rect 1843 127707 1852 127741
rect 1800 127698 1852 127707
rect 136946 127741 136998 127750
rect 136946 127707 136955 127741
rect 136955 127707 136989 127741
rect 136989 127707 136998 127741
rect 136946 127698 136998 127707
rect 29564 127553 29616 127605
rect 32060 127553 32112 127605
rect 34556 127553 34608 127605
rect 37052 127553 37104 127605
rect 39548 127553 39600 127605
rect 42044 127553 42096 127605
rect 44540 127553 44592 127605
rect 47036 127553 47088 127605
rect 49532 127553 49584 127605
rect 52028 127553 52080 127605
rect 54524 127553 54576 127605
rect 57020 127553 57072 127605
rect 59516 127553 59568 127605
rect 62012 127553 62064 127605
rect 64508 127553 64560 127605
rect 67004 127553 67056 127605
rect 69500 127553 69552 127605
rect 71996 127553 72048 127605
rect 74492 127553 74544 127605
rect 76988 127553 77040 127605
rect 79484 127553 79536 127605
rect 81980 127553 82032 127605
rect 84476 127553 84528 127605
rect 86972 127553 87024 127605
rect 89468 127553 89520 127605
rect 91964 127553 92016 127605
rect 94460 127553 94512 127605
rect 96956 127553 97008 127605
rect 99452 127553 99504 127605
rect 101948 127553 102000 127605
rect 104444 127553 104496 127605
rect 106940 127553 106992 127605
rect 1800 127405 1852 127414
rect 1800 127371 1809 127405
rect 1809 127371 1843 127405
rect 1843 127371 1852 127405
rect 1800 127362 1852 127371
rect 136946 127405 136998 127414
rect 136946 127371 136955 127405
rect 136955 127371 136989 127405
rect 136989 127371 136998 127405
rect 136946 127362 136998 127371
rect 1800 127069 1852 127078
rect 1800 127035 1809 127069
rect 1809 127035 1843 127069
rect 1843 127035 1852 127069
rect 1800 127026 1852 127035
rect 136946 127069 136998 127078
rect 136946 127035 136955 127069
rect 136955 127035 136989 127069
rect 136989 127035 136998 127069
rect 136946 127026 136998 127035
rect 1800 126733 1852 126742
rect 1800 126699 1809 126733
rect 1809 126699 1843 126733
rect 1843 126699 1852 126733
rect 1800 126690 1852 126699
rect 136946 126733 136998 126742
rect 136946 126699 136955 126733
rect 136955 126699 136989 126733
rect 136989 126699 136998 126733
rect 136946 126690 136998 126699
rect 1800 126397 1852 126406
rect 1800 126363 1809 126397
rect 1809 126363 1843 126397
rect 1843 126363 1852 126397
rect 1800 126354 1852 126363
rect 136946 126397 136998 126406
rect 136946 126363 136955 126397
rect 136955 126363 136989 126397
rect 136989 126363 136998 126397
rect 136946 126354 136998 126363
rect 1800 126061 1852 126070
rect 1800 126027 1809 126061
rect 1809 126027 1843 126061
rect 1843 126027 1852 126061
rect 1800 126018 1852 126027
rect 136946 126061 136998 126070
rect 136946 126027 136955 126061
rect 136955 126027 136989 126061
rect 136989 126027 136998 126061
rect 136946 126018 136998 126027
rect 1800 125725 1852 125734
rect 1800 125691 1809 125725
rect 1809 125691 1843 125725
rect 1843 125691 1852 125725
rect 1800 125682 1852 125691
rect 136946 125725 136998 125734
rect 136946 125691 136955 125725
rect 136955 125691 136989 125725
rect 136989 125691 136998 125725
rect 136946 125682 136998 125691
rect 1800 125389 1852 125398
rect 1800 125355 1809 125389
rect 1809 125355 1843 125389
rect 1843 125355 1852 125389
rect 1800 125346 1852 125355
rect 136946 125389 136998 125398
rect 136946 125355 136955 125389
rect 136955 125355 136989 125389
rect 136989 125355 136998 125389
rect 136946 125346 136998 125355
rect 1800 125053 1852 125062
rect 1800 125019 1809 125053
rect 1809 125019 1843 125053
rect 1843 125019 1852 125053
rect 1800 125010 1852 125019
rect 136946 125053 136998 125062
rect 136946 125019 136955 125053
rect 136955 125019 136989 125053
rect 136989 125019 136998 125053
rect 136946 125010 136998 125019
rect 1800 124717 1852 124726
rect 1800 124683 1809 124717
rect 1809 124683 1843 124717
rect 1843 124683 1852 124717
rect 1800 124674 1852 124683
rect 136946 124717 136998 124726
rect 136946 124683 136955 124717
rect 136955 124683 136989 124717
rect 136989 124683 136998 124717
rect 136946 124674 136998 124683
rect 1800 124381 1852 124390
rect 1800 124347 1809 124381
rect 1809 124347 1843 124381
rect 1843 124347 1852 124381
rect 1800 124338 1852 124347
rect 136946 124381 136998 124390
rect 136946 124347 136955 124381
rect 136955 124347 136989 124381
rect 136989 124347 136998 124381
rect 136946 124338 136998 124347
rect 1800 124045 1852 124054
rect 1800 124011 1809 124045
rect 1809 124011 1843 124045
rect 1843 124011 1852 124045
rect 1800 124002 1852 124011
rect 136946 124045 136998 124054
rect 136946 124011 136955 124045
rect 136955 124011 136989 124045
rect 136989 124011 136998 124045
rect 136946 124002 136998 124011
rect 1800 123709 1852 123718
rect 1800 123675 1809 123709
rect 1809 123675 1843 123709
rect 1843 123675 1852 123709
rect 1800 123666 1852 123675
rect 136946 123709 136998 123718
rect 136946 123675 136955 123709
rect 136955 123675 136989 123709
rect 136989 123675 136998 123709
rect 136946 123666 136998 123675
rect 1800 123373 1852 123382
rect 1800 123339 1809 123373
rect 1809 123339 1843 123373
rect 1843 123339 1852 123373
rect 1800 123330 1852 123339
rect 136946 123373 136998 123382
rect 136946 123339 136955 123373
rect 136955 123339 136989 123373
rect 136989 123339 136998 123373
rect 136946 123330 136998 123339
rect 1800 123037 1852 123046
rect 1800 123003 1809 123037
rect 1809 123003 1843 123037
rect 1843 123003 1852 123037
rect 1800 122994 1852 123003
rect 136946 123037 136998 123046
rect 136946 123003 136955 123037
rect 136955 123003 136989 123037
rect 136989 123003 136998 123037
rect 136946 122994 136998 123003
rect 1800 122701 1852 122710
rect 1800 122667 1809 122701
rect 1809 122667 1843 122701
rect 1843 122667 1852 122701
rect 1800 122658 1852 122667
rect 136946 122701 136998 122710
rect 136946 122667 136955 122701
rect 136955 122667 136989 122701
rect 136989 122667 136998 122701
rect 136946 122658 136998 122667
rect 1800 122365 1852 122374
rect 1800 122331 1809 122365
rect 1809 122331 1843 122365
rect 1843 122331 1852 122365
rect 1800 122322 1852 122331
rect 136946 122365 136998 122374
rect 136946 122331 136955 122365
rect 136955 122331 136989 122365
rect 136989 122331 136998 122365
rect 136946 122322 136998 122331
rect 1800 122029 1852 122038
rect 1800 121995 1809 122029
rect 1809 121995 1843 122029
rect 1843 121995 1852 122029
rect 1800 121986 1852 121995
rect 136946 122029 136998 122038
rect 136946 121995 136955 122029
rect 136955 121995 136989 122029
rect 136989 121995 136998 122029
rect 136946 121986 136998 121995
rect 1800 121693 1852 121702
rect 1800 121659 1809 121693
rect 1809 121659 1843 121693
rect 1843 121659 1852 121693
rect 1800 121650 1852 121659
rect 136946 121693 136998 121702
rect 136946 121659 136955 121693
rect 136955 121659 136989 121693
rect 136989 121659 136998 121693
rect 136946 121650 136998 121659
rect 1800 121357 1852 121366
rect 1800 121323 1809 121357
rect 1809 121323 1843 121357
rect 1843 121323 1852 121357
rect 1800 121314 1852 121323
rect 136946 121357 136998 121366
rect 136946 121323 136955 121357
rect 136955 121323 136989 121357
rect 136989 121323 136998 121357
rect 136946 121314 136998 121323
rect 1800 121021 1852 121030
rect 1800 120987 1809 121021
rect 1809 120987 1843 121021
rect 1843 120987 1852 121021
rect 1800 120978 1852 120987
rect 136946 121021 136998 121030
rect 136946 120987 136955 121021
rect 136955 120987 136989 121021
rect 136989 120987 136998 121021
rect 136946 120978 136998 120987
rect 1800 120685 1852 120694
rect 1800 120651 1809 120685
rect 1809 120651 1843 120685
rect 1843 120651 1852 120685
rect 1800 120642 1852 120651
rect 136946 120685 136998 120694
rect 136946 120651 136955 120685
rect 136955 120651 136989 120685
rect 136989 120651 136998 120685
rect 136946 120642 136998 120651
rect 1800 120349 1852 120358
rect 1800 120315 1809 120349
rect 1809 120315 1843 120349
rect 1843 120315 1852 120349
rect 1800 120306 1852 120315
rect 136946 120349 136998 120358
rect 136946 120315 136955 120349
rect 136955 120315 136989 120349
rect 136989 120315 136998 120349
rect 136946 120306 136998 120315
rect 1800 120013 1852 120022
rect 1800 119979 1809 120013
rect 1809 119979 1843 120013
rect 1843 119979 1852 120013
rect 1800 119970 1852 119979
rect 136946 120013 136998 120022
rect 136946 119979 136955 120013
rect 136955 119979 136989 120013
rect 136989 119979 136998 120013
rect 136946 119970 136998 119979
rect 1800 119677 1852 119686
rect 1800 119643 1809 119677
rect 1809 119643 1843 119677
rect 1843 119643 1852 119677
rect 1800 119634 1852 119643
rect 136946 119677 136998 119686
rect 136946 119643 136955 119677
rect 136955 119643 136989 119677
rect 136989 119643 136998 119677
rect 136946 119634 136998 119643
rect 1800 119341 1852 119350
rect 1800 119307 1809 119341
rect 1809 119307 1843 119341
rect 1843 119307 1852 119341
rect 1800 119298 1852 119307
rect 136946 119341 136998 119350
rect 136946 119307 136955 119341
rect 136955 119307 136989 119341
rect 136989 119307 136998 119341
rect 136946 119298 136998 119307
rect 1800 119005 1852 119014
rect 1800 118971 1809 119005
rect 1809 118971 1843 119005
rect 1843 118971 1852 119005
rect 1800 118962 1852 118971
rect 136946 119005 136998 119014
rect 136946 118971 136955 119005
rect 136955 118971 136989 119005
rect 136989 118971 136998 119005
rect 136946 118962 136998 118971
rect 1800 118669 1852 118678
rect 1800 118635 1809 118669
rect 1809 118635 1843 118669
rect 1843 118635 1852 118669
rect 1800 118626 1852 118635
rect 136946 118669 136998 118678
rect 136946 118635 136955 118669
rect 136955 118635 136989 118669
rect 136989 118635 136998 118669
rect 136946 118626 136998 118635
rect 1800 118333 1852 118342
rect 1800 118299 1809 118333
rect 1809 118299 1843 118333
rect 1843 118299 1852 118333
rect 1800 118290 1852 118299
rect 136946 118333 136998 118342
rect 136946 118299 136955 118333
rect 136955 118299 136989 118333
rect 136989 118299 136998 118333
rect 136946 118290 136998 118299
rect 1800 117997 1852 118006
rect 1800 117963 1809 117997
rect 1809 117963 1843 117997
rect 1843 117963 1852 117997
rect 1800 117954 1852 117963
rect 136946 117997 136998 118006
rect 136946 117963 136955 117997
rect 136955 117963 136989 117997
rect 136989 117963 136998 117997
rect 136946 117954 136998 117963
rect 1800 117661 1852 117670
rect 1800 117627 1809 117661
rect 1809 117627 1843 117661
rect 1843 117627 1852 117661
rect 1800 117618 1852 117627
rect 136946 117661 136998 117670
rect 136946 117627 136955 117661
rect 136955 117627 136989 117661
rect 136989 117627 136998 117661
rect 136946 117618 136998 117627
rect 1800 117325 1852 117334
rect 1800 117291 1809 117325
rect 1809 117291 1843 117325
rect 1843 117291 1852 117325
rect 1800 117282 1852 117291
rect 136946 117325 136998 117334
rect 136946 117291 136955 117325
rect 136955 117291 136989 117325
rect 136989 117291 136998 117325
rect 136946 117282 136998 117291
rect 1800 116989 1852 116998
rect 1800 116955 1809 116989
rect 1809 116955 1843 116989
rect 1843 116955 1852 116989
rect 1800 116946 1852 116955
rect 136946 116989 136998 116998
rect 136946 116955 136955 116989
rect 136955 116955 136989 116989
rect 136989 116955 136998 116989
rect 136946 116946 136998 116955
rect 1800 116653 1852 116662
rect 1800 116619 1809 116653
rect 1809 116619 1843 116653
rect 1843 116619 1852 116653
rect 1800 116610 1852 116619
rect 136946 116653 136998 116662
rect 136946 116619 136955 116653
rect 136955 116619 136989 116653
rect 136989 116619 136998 116653
rect 136946 116610 136998 116619
rect 1800 116317 1852 116326
rect 1800 116283 1809 116317
rect 1809 116283 1843 116317
rect 1843 116283 1852 116317
rect 1800 116274 1852 116283
rect 136946 116317 136998 116326
rect 136946 116283 136955 116317
rect 136955 116283 136989 116317
rect 136989 116283 136998 116317
rect 136946 116274 136998 116283
rect 1800 115981 1852 115990
rect 1800 115947 1809 115981
rect 1809 115947 1843 115981
rect 1843 115947 1852 115981
rect 1800 115938 1852 115947
rect 136946 115981 136998 115990
rect 136946 115947 136955 115981
rect 136955 115947 136989 115981
rect 136989 115947 136998 115981
rect 136946 115938 136998 115947
rect 1800 115645 1852 115654
rect 1800 115611 1809 115645
rect 1809 115611 1843 115645
rect 1843 115611 1852 115645
rect 1800 115602 1852 115611
rect 136946 115645 136998 115654
rect 136946 115611 136955 115645
rect 136955 115611 136989 115645
rect 136989 115611 136998 115645
rect 136946 115602 136998 115611
rect 1800 115309 1852 115318
rect 1800 115275 1809 115309
rect 1809 115275 1843 115309
rect 1843 115275 1852 115309
rect 1800 115266 1852 115275
rect 136946 115309 136998 115318
rect 136946 115275 136955 115309
rect 136955 115275 136989 115309
rect 136989 115275 136998 115309
rect 136946 115266 136998 115275
rect 1800 114973 1852 114982
rect 1800 114939 1809 114973
rect 1809 114939 1843 114973
rect 1843 114939 1852 114973
rect 1800 114930 1852 114939
rect 136946 114973 136998 114982
rect 136946 114939 136955 114973
rect 136955 114939 136989 114973
rect 136989 114939 136998 114973
rect 136946 114930 136998 114939
rect 1800 114637 1852 114646
rect 1800 114603 1809 114637
rect 1809 114603 1843 114637
rect 1843 114603 1852 114637
rect 1800 114594 1852 114603
rect 136946 114637 136998 114646
rect 136946 114603 136955 114637
rect 136955 114603 136989 114637
rect 136989 114603 136998 114637
rect 136946 114594 136998 114603
rect 1800 114301 1852 114310
rect 1800 114267 1809 114301
rect 1809 114267 1843 114301
rect 1843 114267 1852 114301
rect 1800 114258 1852 114267
rect 136946 114301 136998 114310
rect 136946 114267 136955 114301
rect 136955 114267 136989 114301
rect 136989 114267 136998 114301
rect 136946 114258 136998 114267
rect 1800 113965 1852 113974
rect 1800 113931 1809 113965
rect 1809 113931 1843 113965
rect 1843 113931 1852 113965
rect 1800 113922 1852 113931
rect 136946 113965 136998 113974
rect 136946 113931 136955 113965
rect 136955 113931 136989 113965
rect 136989 113931 136998 113965
rect 136946 113922 136998 113931
rect 1800 113629 1852 113638
rect 1800 113595 1809 113629
rect 1809 113595 1843 113629
rect 1843 113595 1852 113629
rect 1800 113586 1852 113595
rect 136946 113629 136998 113638
rect 136946 113595 136955 113629
rect 136955 113595 136989 113629
rect 136989 113595 136998 113629
rect 136946 113586 136998 113595
rect 1800 113293 1852 113302
rect 1800 113259 1809 113293
rect 1809 113259 1843 113293
rect 1843 113259 1852 113293
rect 1800 113250 1852 113259
rect 136946 113293 136998 113302
rect 136946 113259 136955 113293
rect 136955 113259 136989 113293
rect 136989 113259 136998 113293
rect 136946 113250 136998 113259
rect 1800 112957 1852 112966
rect 1800 112923 1809 112957
rect 1809 112923 1843 112957
rect 1843 112923 1852 112957
rect 1800 112914 1852 112923
rect 136946 112957 136998 112966
rect 136946 112923 136955 112957
rect 136955 112923 136989 112957
rect 136989 112923 136998 112957
rect 136946 112914 136998 112923
rect 1800 112621 1852 112630
rect 1800 112587 1809 112621
rect 1809 112587 1843 112621
rect 1843 112587 1852 112621
rect 1800 112578 1852 112587
rect 136946 112621 136998 112630
rect 136946 112587 136955 112621
rect 136955 112587 136989 112621
rect 136989 112587 136998 112621
rect 136946 112578 136998 112587
rect 1800 112285 1852 112294
rect 1800 112251 1809 112285
rect 1809 112251 1843 112285
rect 1843 112251 1852 112285
rect 1800 112242 1852 112251
rect 136946 112285 136998 112294
rect 136946 112251 136955 112285
rect 136955 112251 136989 112285
rect 136989 112251 136998 112285
rect 136946 112242 136998 112251
rect 1800 111949 1852 111958
rect 1800 111915 1809 111949
rect 1809 111915 1843 111949
rect 1843 111915 1852 111949
rect 1800 111906 1852 111915
rect 136946 111949 136998 111958
rect 136946 111915 136955 111949
rect 136955 111915 136989 111949
rect 136989 111915 136998 111949
rect 136946 111906 136998 111915
rect 1800 111613 1852 111622
rect 1800 111579 1809 111613
rect 1809 111579 1843 111613
rect 1843 111579 1852 111613
rect 1800 111570 1852 111579
rect 136946 111613 136998 111622
rect 136946 111579 136955 111613
rect 136955 111579 136989 111613
rect 136989 111579 136998 111613
rect 136946 111570 136998 111579
rect 1800 111277 1852 111286
rect 1800 111243 1809 111277
rect 1809 111243 1843 111277
rect 1843 111243 1852 111277
rect 1800 111234 1852 111243
rect 136946 111277 136998 111286
rect 136946 111243 136955 111277
rect 136955 111243 136989 111277
rect 136989 111243 136998 111277
rect 136946 111234 136998 111243
rect 1800 110941 1852 110950
rect 1800 110907 1809 110941
rect 1809 110907 1843 110941
rect 1843 110907 1852 110941
rect 1800 110898 1852 110907
rect 136946 110941 136998 110950
rect 136946 110907 136955 110941
rect 136955 110907 136989 110941
rect 136989 110907 136998 110941
rect 136946 110898 136998 110907
rect 1800 110605 1852 110614
rect 1800 110571 1809 110605
rect 1809 110571 1843 110605
rect 1843 110571 1852 110605
rect 1800 110562 1852 110571
rect 136946 110605 136998 110614
rect 136946 110571 136955 110605
rect 136955 110571 136989 110605
rect 136989 110571 136998 110605
rect 136946 110562 136998 110571
rect 1800 110269 1852 110278
rect 1800 110235 1809 110269
rect 1809 110235 1843 110269
rect 1843 110235 1852 110269
rect 1800 110226 1852 110235
rect 136946 110269 136998 110278
rect 136946 110235 136955 110269
rect 136955 110235 136989 110269
rect 136989 110235 136998 110269
rect 136946 110226 136998 110235
rect 1800 109933 1852 109942
rect 1800 109899 1809 109933
rect 1809 109899 1843 109933
rect 1843 109899 1852 109933
rect 1800 109890 1852 109899
rect 136946 109933 136998 109942
rect 136946 109899 136955 109933
rect 136955 109899 136989 109933
rect 136989 109899 136998 109933
rect 136946 109890 136998 109899
rect 1800 109597 1852 109606
rect 1800 109563 1809 109597
rect 1809 109563 1843 109597
rect 1843 109563 1852 109597
rect 1800 109554 1852 109563
rect 136946 109597 136998 109606
rect 136946 109563 136955 109597
rect 136955 109563 136989 109597
rect 136989 109563 136998 109597
rect 136946 109554 136998 109563
rect 1800 109261 1852 109270
rect 1800 109227 1809 109261
rect 1809 109227 1843 109261
rect 1843 109227 1852 109261
rect 1800 109218 1852 109227
rect 136946 109261 136998 109270
rect 136946 109227 136955 109261
rect 136955 109227 136989 109261
rect 136989 109227 136998 109261
rect 136946 109218 136998 109227
rect 1800 108925 1852 108934
rect 1800 108891 1809 108925
rect 1809 108891 1843 108925
rect 1843 108891 1852 108925
rect 1800 108882 1852 108891
rect 136946 108925 136998 108934
rect 136946 108891 136955 108925
rect 136955 108891 136989 108925
rect 136989 108891 136998 108925
rect 136946 108882 136998 108891
rect 1800 108589 1852 108598
rect 1800 108555 1809 108589
rect 1809 108555 1843 108589
rect 1843 108555 1852 108589
rect 1800 108546 1852 108555
rect 136946 108589 136998 108598
rect 136946 108555 136955 108589
rect 136955 108555 136989 108589
rect 136989 108555 136998 108589
rect 136946 108546 136998 108555
rect 1800 108253 1852 108262
rect 1800 108219 1809 108253
rect 1809 108219 1843 108253
rect 1843 108219 1852 108253
rect 1800 108210 1852 108219
rect 136946 108253 136998 108262
rect 136946 108219 136955 108253
rect 136955 108219 136989 108253
rect 136989 108219 136998 108253
rect 136946 108210 136998 108219
rect 1800 107917 1852 107926
rect 1800 107883 1809 107917
rect 1809 107883 1843 107917
rect 1843 107883 1852 107917
rect 1800 107874 1852 107883
rect 136946 107917 136998 107926
rect 136946 107883 136955 107917
rect 136955 107883 136989 107917
rect 136989 107883 136998 107917
rect 136946 107874 136998 107883
rect 1800 107581 1852 107590
rect 1800 107547 1809 107581
rect 1809 107547 1843 107581
rect 1843 107547 1852 107581
rect 1800 107538 1852 107547
rect 136946 107581 136998 107590
rect 136946 107547 136955 107581
rect 136955 107547 136989 107581
rect 136989 107547 136998 107581
rect 136946 107538 136998 107547
rect 1800 107245 1852 107254
rect 1800 107211 1809 107245
rect 1809 107211 1843 107245
rect 1843 107211 1852 107245
rect 1800 107202 1852 107211
rect 136946 107245 136998 107254
rect 136946 107211 136955 107245
rect 136955 107211 136989 107245
rect 136989 107211 136998 107245
rect 136946 107202 136998 107211
rect 1800 106909 1852 106918
rect 1800 106875 1809 106909
rect 1809 106875 1843 106909
rect 1843 106875 1852 106909
rect 1800 106866 1852 106875
rect 136946 106909 136998 106918
rect 136946 106875 136955 106909
rect 136955 106875 136989 106909
rect 136989 106875 136998 106909
rect 136946 106866 136998 106875
rect 1800 106573 1852 106582
rect 1800 106539 1809 106573
rect 1809 106539 1843 106573
rect 1843 106539 1852 106573
rect 1800 106530 1852 106539
rect 136946 106573 136998 106582
rect 136946 106539 136955 106573
rect 136955 106539 136989 106573
rect 136989 106539 136998 106573
rect 136946 106530 136998 106539
rect 1800 106237 1852 106246
rect 1800 106203 1809 106237
rect 1809 106203 1843 106237
rect 1843 106203 1852 106237
rect 1800 106194 1852 106203
rect 136946 106237 136998 106246
rect 136946 106203 136955 106237
rect 136955 106203 136989 106237
rect 136989 106203 136998 106237
rect 136946 106194 136998 106203
rect 1800 105901 1852 105910
rect 1800 105867 1809 105901
rect 1809 105867 1843 105901
rect 1843 105867 1852 105901
rect 1800 105858 1852 105867
rect 136946 105901 136998 105910
rect 136946 105867 136955 105901
rect 136955 105867 136989 105901
rect 136989 105867 136998 105901
rect 136946 105858 136998 105867
rect 1800 105565 1852 105574
rect 1800 105531 1809 105565
rect 1809 105531 1843 105565
rect 1843 105531 1852 105565
rect 1800 105522 1852 105531
rect 136946 105565 136998 105574
rect 136946 105531 136955 105565
rect 136955 105531 136989 105565
rect 136989 105531 136998 105565
rect 136946 105522 136998 105531
rect 1800 105229 1852 105238
rect 1800 105195 1809 105229
rect 1809 105195 1843 105229
rect 1843 105195 1852 105229
rect 1800 105186 1852 105195
rect 136946 105229 136998 105238
rect 136946 105195 136955 105229
rect 136955 105195 136989 105229
rect 136989 105195 136998 105229
rect 136946 105186 136998 105195
rect 1800 104893 1852 104902
rect 1800 104859 1809 104893
rect 1809 104859 1843 104893
rect 1843 104859 1852 104893
rect 1800 104850 1852 104859
rect 136946 104893 136998 104902
rect 136946 104859 136955 104893
rect 136955 104859 136989 104893
rect 136989 104859 136998 104893
rect 136946 104850 136998 104859
rect 1800 104557 1852 104566
rect 1800 104523 1809 104557
rect 1809 104523 1843 104557
rect 1843 104523 1852 104557
rect 1800 104514 1852 104523
rect 136946 104557 136998 104566
rect 136946 104523 136955 104557
rect 136955 104523 136989 104557
rect 136989 104523 136998 104557
rect 136946 104514 136998 104523
rect 1800 104221 1852 104230
rect 1800 104187 1809 104221
rect 1809 104187 1843 104221
rect 1843 104187 1852 104221
rect 1800 104178 1852 104187
rect 136946 104221 136998 104230
rect 136946 104187 136955 104221
rect 136955 104187 136989 104221
rect 136989 104187 136998 104221
rect 136946 104178 136998 104187
rect 1800 103885 1852 103894
rect 1800 103851 1809 103885
rect 1809 103851 1843 103885
rect 1843 103851 1852 103885
rect 1800 103842 1852 103851
rect 136946 103885 136998 103894
rect 136946 103851 136955 103885
rect 136955 103851 136989 103885
rect 136989 103851 136998 103885
rect 136946 103842 136998 103851
rect 1800 103549 1852 103558
rect 1800 103515 1809 103549
rect 1809 103515 1843 103549
rect 1843 103515 1852 103549
rect 1800 103506 1852 103515
rect 136946 103549 136998 103558
rect 136946 103515 136955 103549
rect 136955 103515 136989 103549
rect 136989 103515 136998 103549
rect 136946 103506 136998 103515
rect 1800 103213 1852 103222
rect 1800 103179 1809 103213
rect 1809 103179 1843 103213
rect 1843 103179 1852 103213
rect 1800 103170 1852 103179
rect 136946 103213 136998 103222
rect 136946 103179 136955 103213
rect 136955 103179 136989 103213
rect 136989 103179 136998 103213
rect 136946 103170 136998 103179
rect 1800 102877 1852 102886
rect 1800 102843 1809 102877
rect 1809 102843 1843 102877
rect 1843 102843 1852 102877
rect 1800 102834 1852 102843
rect 136946 102877 136998 102886
rect 136946 102843 136955 102877
rect 136955 102843 136989 102877
rect 136989 102843 136998 102877
rect 136946 102834 136998 102843
rect 1800 102541 1852 102550
rect 1800 102507 1809 102541
rect 1809 102507 1843 102541
rect 1843 102507 1852 102541
rect 1800 102498 1852 102507
rect 136946 102541 136998 102550
rect 136946 102507 136955 102541
rect 136955 102507 136989 102541
rect 136989 102507 136998 102541
rect 136946 102498 136998 102507
rect 1800 102205 1852 102214
rect 1800 102171 1809 102205
rect 1809 102171 1843 102205
rect 1843 102171 1852 102205
rect 1800 102162 1852 102171
rect 136946 102205 136998 102214
rect 136946 102171 136955 102205
rect 136955 102171 136989 102205
rect 136989 102171 136998 102205
rect 136946 102162 136998 102171
rect 1800 101869 1852 101878
rect 1800 101835 1809 101869
rect 1809 101835 1843 101869
rect 1843 101835 1852 101869
rect 1800 101826 1852 101835
rect 136946 101869 136998 101878
rect 136946 101835 136955 101869
rect 136955 101835 136989 101869
rect 136989 101835 136998 101869
rect 136946 101826 136998 101835
rect 1800 101533 1852 101542
rect 1800 101499 1809 101533
rect 1809 101499 1843 101533
rect 1843 101499 1852 101533
rect 1800 101490 1852 101499
rect 136946 101533 136998 101542
rect 136946 101499 136955 101533
rect 136955 101499 136989 101533
rect 136989 101499 136998 101533
rect 136946 101490 136998 101499
rect 1800 101197 1852 101206
rect 1800 101163 1809 101197
rect 1809 101163 1843 101197
rect 1843 101163 1852 101197
rect 1800 101154 1852 101163
rect 136946 101197 136998 101206
rect 136946 101163 136955 101197
rect 136955 101163 136989 101197
rect 136989 101163 136998 101197
rect 136946 101154 136998 101163
rect 1800 100861 1852 100870
rect 1800 100827 1809 100861
rect 1809 100827 1843 100861
rect 1843 100827 1852 100861
rect 1800 100818 1852 100827
rect 136946 100861 136998 100870
rect 136946 100827 136955 100861
rect 136955 100827 136989 100861
rect 136989 100827 136998 100861
rect 136946 100818 136998 100827
rect 1800 100525 1852 100534
rect 1800 100491 1809 100525
rect 1809 100491 1843 100525
rect 1843 100491 1852 100525
rect 1800 100482 1852 100491
rect 136946 100525 136998 100534
rect 136946 100491 136955 100525
rect 136955 100491 136989 100525
rect 136989 100491 136998 100525
rect 136946 100482 136998 100491
rect 1800 100189 1852 100198
rect 1800 100155 1809 100189
rect 1809 100155 1843 100189
rect 1843 100155 1852 100189
rect 1800 100146 1852 100155
rect 136946 100189 136998 100198
rect 136946 100155 136955 100189
rect 136955 100155 136989 100189
rect 136989 100155 136998 100189
rect 136946 100146 136998 100155
rect 1800 99853 1852 99862
rect 1800 99819 1809 99853
rect 1809 99819 1843 99853
rect 1843 99819 1852 99853
rect 1800 99810 1852 99819
rect 136946 99853 136998 99862
rect 136946 99819 136955 99853
rect 136955 99819 136989 99853
rect 136989 99819 136998 99853
rect 136946 99810 136998 99819
rect 1800 99517 1852 99526
rect 1800 99483 1809 99517
rect 1809 99483 1843 99517
rect 1843 99483 1852 99517
rect 1800 99474 1852 99483
rect 136946 99517 136998 99526
rect 136946 99483 136955 99517
rect 136955 99483 136989 99517
rect 136989 99483 136998 99517
rect 136946 99474 136998 99483
rect 1800 99181 1852 99190
rect 1800 99147 1809 99181
rect 1809 99147 1843 99181
rect 1843 99147 1852 99181
rect 1800 99138 1852 99147
rect 136946 99181 136998 99190
rect 136946 99147 136955 99181
rect 136955 99147 136989 99181
rect 136989 99147 136998 99181
rect 136946 99138 136998 99147
rect 1800 98845 1852 98854
rect 1800 98811 1809 98845
rect 1809 98811 1843 98845
rect 1843 98811 1852 98845
rect 1800 98802 1852 98811
rect 136946 98845 136998 98854
rect 136946 98811 136955 98845
rect 136955 98811 136989 98845
rect 136989 98811 136998 98845
rect 136946 98802 136998 98811
rect 1800 98509 1852 98518
rect 1800 98475 1809 98509
rect 1809 98475 1843 98509
rect 1843 98475 1852 98509
rect 1800 98466 1852 98475
rect 136946 98509 136998 98518
rect 136946 98475 136955 98509
rect 136955 98475 136989 98509
rect 136989 98475 136998 98509
rect 136946 98466 136998 98475
rect 1800 98173 1852 98182
rect 1800 98139 1809 98173
rect 1809 98139 1843 98173
rect 1843 98139 1852 98173
rect 1800 98130 1852 98139
rect 136946 98173 136998 98182
rect 136946 98139 136955 98173
rect 136955 98139 136989 98173
rect 136989 98139 136998 98173
rect 136946 98130 136998 98139
rect 1800 97837 1852 97846
rect 1800 97803 1809 97837
rect 1809 97803 1843 97837
rect 1843 97803 1852 97837
rect 1800 97794 1852 97803
rect 136946 97837 136998 97846
rect 136946 97803 136955 97837
rect 136955 97803 136989 97837
rect 136989 97803 136998 97837
rect 136946 97794 136998 97803
rect 1800 97501 1852 97510
rect 1800 97467 1809 97501
rect 1809 97467 1843 97501
rect 1843 97467 1852 97501
rect 1800 97458 1852 97467
rect 136946 97501 136998 97510
rect 136946 97467 136955 97501
rect 136955 97467 136989 97501
rect 136989 97467 136998 97501
rect 136946 97458 136998 97467
rect 1800 97165 1852 97174
rect 1800 97131 1809 97165
rect 1809 97131 1843 97165
rect 1843 97131 1852 97165
rect 1800 97122 1852 97131
rect 136946 97165 136998 97174
rect 136946 97131 136955 97165
rect 136955 97131 136989 97165
rect 136989 97131 136998 97165
rect 136946 97122 136998 97131
rect 1800 96829 1852 96838
rect 1800 96795 1809 96829
rect 1809 96795 1843 96829
rect 1843 96795 1852 96829
rect 1800 96786 1852 96795
rect 136946 96829 136998 96838
rect 136946 96795 136955 96829
rect 136955 96795 136989 96829
rect 136989 96795 136998 96829
rect 136946 96786 136998 96795
rect 1800 96493 1852 96502
rect 1800 96459 1809 96493
rect 1809 96459 1843 96493
rect 1843 96459 1852 96493
rect 1800 96450 1852 96459
rect 136946 96493 136998 96502
rect 136946 96459 136955 96493
rect 136955 96459 136989 96493
rect 136989 96459 136998 96493
rect 136946 96450 136998 96459
rect 1800 96157 1852 96166
rect 1800 96123 1809 96157
rect 1809 96123 1843 96157
rect 1843 96123 1852 96157
rect 1800 96114 1852 96123
rect 136946 96157 136998 96166
rect 136946 96123 136955 96157
rect 136955 96123 136989 96157
rect 136989 96123 136998 96157
rect 136946 96114 136998 96123
rect 1800 95821 1852 95830
rect 1800 95787 1809 95821
rect 1809 95787 1843 95821
rect 1843 95787 1852 95821
rect 1800 95778 1852 95787
rect 136946 95821 136998 95830
rect 136946 95787 136955 95821
rect 136955 95787 136989 95821
rect 136989 95787 136998 95821
rect 136946 95778 136998 95787
rect 1800 95485 1852 95494
rect 1800 95451 1809 95485
rect 1809 95451 1843 95485
rect 1843 95451 1852 95485
rect 1800 95442 1852 95451
rect 136946 95485 136998 95494
rect 136946 95451 136955 95485
rect 136955 95451 136989 95485
rect 136989 95451 136998 95485
rect 136946 95442 136998 95451
rect 1800 95149 1852 95158
rect 1800 95115 1809 95149
rect 1809 95115 1843 95149
rect 1843 95115 1852 95149
rect 1800 95106 1852 95115
rect 136946 95149 136998 95158
rect 136946 95115 136955 95149
rect 136955 95115 136989 95149
rect 136989 95115 136998 95149
rect 136946 95106 136998 95115
rect 1800 94813 1852 94822
rect 1800 94779 1809 94813
rect 1809 94779 1843 94813
rect 1843 94779 1852 94813
rect 1800 94770 1852 94779
rect 136946 94813 136998 94822
rect 136946 94779 136955 94813
rect 136955 94779 136989 94813
rect 136989 94779 136998 94813
rect 136946 94770 136998 94779
rect 1800 94477 1852 94486
rect 1800 94443 1809 94477
rect 1809 94443 1843 94477
rect 1843 94443 1852 94477
rect 1800 94434 1852 94443
rect 136946 94477 136998 94486
rect 136946 94443 136955 94477
rect 136955 94443 136989 94477
rect 136989 94443 136998 94477
rect 136946 94434 136998 94443
rect 1800 94141 1852 94150
rect 1800 94107 1809 94141
rect 1809 94107 1843 94141
rect 1843 94107 1852 94141
rect 1800 94098 1852 94107
rect 136946 94141 136998 94150
rect 136946 94107 136955 94141
rect 136955 94107 136989 94141
rect 136989 94107 136998 94141
rect 136946 94098 136998 94107
rect 1800 93805 1852 93814
rect 1800 93771 1809 93805
rect 1809 93771 1843 93805
rect 1843 93771 1852 93805
rect 1800 93762 1852 93771
rect 136946 93805 136998 93814
rect 136946 93771 136955 93805
rect 136955 93771 136989 93805
rect 136989 93771 136998 93805
rect 136946 93762 136998 93771
rect 1800 93469 1852 93478
rect 1800 93435 1809 93469
rect 1809 93435 1843 93469
rect 1843 93435 1852 93469
rect 1800 93426 1852 93435
rect 136946 93469 136998 93478
rect 136946 93435 136955 93469
rect 136955 93435 136989 93469
rect 136989 93435 136998 93469
rect 136946 93426 136998 93435
rect 1800 93133 1852 93142
rect 1800 93099 1809 93133
rect 1809 93099 1843 93133
rect 1843 93099 1852 93133
rect 1800 93090 1852 93099
rect 136946 93133 136998 93142
rect 136946 93099 136955 93133
rect 136955 93099 136989 93133
rect 136989 93099 136998 93133
rect 136946 93090 136998 93099
rect 1800 92797 1852 92806
rect 1800 92763 1809 92797
rect 1809 92763 1843 92797
rect 1843 92763 1852 92797
rect 1800 92754 1852 92763
rect 136946 92797 136998 92806
rect 136946 92763 136955 92797
rect 136955 92763 136989 92797
rect 136989 92763 136998 92797
rect 136946 92754 136998 92763
rect 1800 92461 1852 92470
rect 1800 92427 1809 92461
rect 1809 92427 1843 92461
rect 1843 92427 1852 92461
rect 1800 92418 1852 92427
rect 136946 92461 136998 92470
rect 136946 92427 136955 92461
rect 136955 92427 136989 92461
rect 136989 92427 136998 92461
rect 136946 92418 136998 92427
rect 1800 92125 1852 92134
rect 1800 92091 1809 92125
rect 1809 92091 1843 92125
rect 1843 92091 1852 92125
rect 1800 92082 1852 92091
rect 136946 92125 136998 92134
rect 136946 92091 136955 92125
rect 136955 92091 136989 92125
rect 136989 92091 136998 92125
rect 136946 92082 136998 92091
rect 1800 91789 1852 91798
rect 1800 91755 1809 91789
rect 1809 91755 1843 91789
rect 1843 91755 1852 91789
rect 1800 91746 1852 91755
rect 136946 91789 136998 91798
rect 136946 91755 136955 91789
rect 136955 91755 136989 91789
rect 136989 91755 136998 91789
rect 136946 91746 136998 91755
rect 1800 91453 1852 91462
rect 1800 91419 1809 91453
rect 1809 91419 1843 91453
rect 1843 91419 1852 91453
rect 1800 91410 1852 91419
rect 136946 91453 136998 91462
rect 136946 91419 136955 91453
rect 136955 91419 136989 91453
rect 136989 91419 136998 91453
rect 136946 91410 136998 91419
rect 1800 91117 1852 91126
rect 1800 91083 1809 91117
rect 1809 91083 1843 91117
rect 1843 91083 1852 91117
rect 1800 91074 1852 91083
rect 136946 91117 136998 91126
rect 136946 91083 136955 91117
rect 136955 91083 136989 91117
rect 136989 91083 136998 91117
rect 136946 91074 136998 91083
rect 1800 90781 1852 90790
rect 1800 90747 1809 90781
rect 1809 90747 1843 90781
rect 1843 90747 1852 90781
rect 1800 90738 1852 90747
rect 136946 90781 136998 90790
rect 136946 90747 136955 90781
rect 136955 90747 136989 90781
rect 136989 90747 136998 90781
rect 136946 90738 136998 90747
rect 1800 90445 1852 90454
rect 1800 90411 1809 90445
rect 1809 90411 1843 90445
rect 1843 90411 1852 90445
rect 1800 90402 1852 90411
rect 136946 90445 136998 90454
rect 136946 90411 136955 90445
rect 136955 90411 136989 90445
rect 136989 90411 136998 90445
rect 136946 90402 136998 90411
rect 1800 90109 1852 90118
rect 1800 90075 1809 90109
rect 1809 90075 1843 90109
rect 1843 90075 1852 90109
rect 1800 90066 1852 90075
rect 136946 90109 136998 90118
rect 136946 90075 136955 90109
rect 136955 90075 136989 90109
rect 136989 90075 136998 90109
rect 136946 90066 136998 90075
rect 1800 89773 1852 89782
rect 1800 89739 1809 89773
rect 1809 89739 1843 89773
rect 1843 89739 1852 89773
rect 1800 89730 1852 89739
rect 136946 89773 136998 89782
rect 136946 89739 136955 89773
rect 136955 89739 136989 89773
rect 136989 89739 136998 89773
rect 136946 89730 136998 89739
rect 1800 89437 1852 89446
rect 1800 89403 1809 89437
rect 1809 89403 1843 89437
rect 1843 89403 1852 89437
rect 1800 89394 1852 89403
rect 136946 89437 136998 89446
rect 136946 89403 136955 89437
rect 136955 89403 136989 89437
rect 136989 89403 136998 89437
rect 136946 89394 136998 89403
rect 1800 89101 1852 89110
rect 1800 89067 1809 89101
rect 1809 89067 1843 89101
rect 1843 89067 1852 89101
rect 1800 89058 1852 89067
rect 136946 89101 136998 89110
rect 136946 89067 136955 89101
rect 136955 89067 136989 89101
rect 136989 89067 136998 89101
rect 136946 89058 136998 89067
rect 1800 88765 1852 88774
rect 1800 88731 1809 88765
rect 1809 88731 1843 88765
rect 1843 88731 1852 88765
rect 1800 88722 1852 88731
rect 136946 88765 136998 88774
rect 136946 88731 136955 88765
rect 136955 88731 136989 88765
rect 136989 88731 136998 88765
rect 136946 88722 136998 88731
rect 1800 88429 1852 88438
rect 1800 88395 1809 88429
rect 1809 88395 1843 88429
rect 1843 88395 1852 88429
rect 1800 88386 1852 88395
rect 136946 88429 136998 88438
rect 136946 88395 136955 88429
rect 136955 88395 136989 88429
rect 136989 88395 136998 88429
rect 136946 88386 136998 88395
rect 1800 88093 1852 88102
rect 1800 88059 1809 88093
rect 1809 88059 1843 88093
rect 1843 88059 1852 88093
rect 1800 88050 1852 88059
rect 136946 88093 136998 88102
rect 136946 88059 136955 88093
rect 136955 88059 136989 88093
rect 136989 88059 136998 88093
rect 136946 88050 136998 88059
rect 1800 87757 1852 87766
rect 1800 87723 1809 87757
rect 1809 87723 1843 87757
rect 1843 87723 1852 87757
rect 1800 87714 1852 87723
rect 136946 87757 136998 87766
rect 136946 87723 136955 87757
rect 136955 87723 136989 87757
rect 136989 87723 136998 87757
rect 136946 87714 136998 87723
rect 1800 87421 1852 87430
rect 1800 87387 1809 87421
rect 1809 87387 1843 87421
rect 1843 87387 1852 87421
rect 1800 87378 1852 87387
rect 136946 87421 136998 87430
rect 136946 87387 136955 87421
rect 136955 87387 136989 87421
rect 136989 87387 136998 87421
rect 136946 87378 136998 87387
rect 1800 87085 1852 87094
rect 1800 87051 1809 87085
rect 1809 87051 1843 87085
rect 1843 87051 1852 87085
rect 1800 87042 1852 87051
rect 136946 87085 136998 87094
rect 136946 87051 136955 87085
rect 136955 87051 136989 87085
rect 136989 87051 136998 87085
rect 136946 87042 136998 87051
rect 1800 86749 1852 86758
rect 1800 86715 1809 86749
rect 1809 86715 1843 86749
rect 1843 86715 1852 86749
rect 1800 86706 1852 86715
rect 136946 86749 136998 86758
rect 136946 86715 136955 86749
rect 136955 86715 136989 86749
rect 136989 86715 136998 86749
rect 136946 86706 136998 86715
rect 1800 86413 1852 86422
rect 1800 86379 1809 86413
rect 1809 86379 1843 86413
rect 1843 86379 1852 86413
rect 1800 86370 1852 86379
rect 136946 86413 136998 86422
rect 136946 86379 136955 86413
rect 136955 86379 136989 86413
rect 136989 86379 136998 86413
rect 136946 86370 136998 86379
rect 1800 86077 1852 86086
rect 1800 86043 1809 86077
rect 1809 86043 1843 86077
rect 1843 86043 1852 86077
rect 1800 86034 1852 86043
rect 136946 86077 136998 86086
rect 136946 86043 136955 86077
rect 136955 86043 136989 86077
rect 136989 86043 136998 86077
rect 136946 86034 136998 86043
rect 1800 85741 1852 85750
rect 1800 85707 1809 85741
rect 1809 85707 1843 85741
rect 1843 85707 1852 85741
rect 1800 85698 1852 85707
rect 136946 85741 136998 85750
rect 136946 85707 136955 85741
rect 136955 85707 136989 85741
rect 136989 85707 136998 85741
rect 136946 85698 136998 85707
rect 1800 85405 1852 85414
rect 1800 85371 1809 85405
rect 1809 85371 1843 85405
rect 1843 85371 1852 85405
rect 1800 85362 1852 85371
rect 136946 85405 136998 85414
rect 136946 85371 136955 85405
rect 136955 85371 136989 85405
rect 136989 85371 136998 85405
rect 136946 85362 136998 85371
rect 1800 85069 1852 85078
rect 1800 85035 1809 85069
rect 1809 85035 1843 85069
rect 1843 85035 1852 85069
rect 1800 85026 1852 85035
rect 136946 85069 136998 85078
rect 136946 85035 136955 85069
rect 136955 85035 136989 85069
rect 136989 85035 136998 85069
rect 136946 85026 136998 85035
rect 1800 84733 1852 84742
rect 1800 84699 1809 84733
rect 1809 84699 1843 84733
rect 1843 84699 1852 84733
rect 1800 84690 1852 84699
rect 136946 84733 136998 84742
rect 136946 84699 136955 84733
rect 136955 84699 136989 84733
rect 136989 84699 136998 84733
rect 136946 84690 136998 84699
rect 1800 84397 1852 84406
rect 1800 84363 1809 84397
rect 1809 84363 1843 84397
rect 1843 84363 1852 84397
rect 1800 84354 1852 84363
rect 136946 84397 136998 84406
rect 136946 84363 136955 84397
rect 136955 84363 136989 84397
rect 136989 84363 136998 84397
rect 136946 84354 136998 84363
rect 1800 84061 1852 84070
rect 1800 84027 1809 84061
rect 1809 84027 1843 84061
rect 1843 84027 1852 84061
rect 1800 84018 1852 84027
rect 136946 84061 136998 84070
rect 136946 84027 136955 84061
rect 136955 84027 136989 84061
rect 136989 84027 136998 84061
rect 136946 84018 136998 84027
rect 1800 83725 1852 83734
rect 1800 83691 1809 83725
rect 1809 83691 1843 83725
rect 1843 83691 1852 83725
rect 1800 83682 1852 83691
rect 136946 83725 136998 83734
rect 136946 83691 136955 83725
rect 136955 83691 136989 83725
rect 136989 83691 136998 83725
rect 136946 83682 136998 83691
rect 1800 83389 1852 83398
rect 1800 83355 1809 83389
rect 1809 83355 1843 83389
rect 1843 83355 1852 83389
rect 1800 83346 1852 83355
rect 136946 83389 136998 83398
rect 136946 83355 136955 83389
rect 136955 83355 136989 83389
rect 136989 83355 136998 83389
rect 136946 83346 136998 83355
rect 1800 83053 1852 83062
rect 1800 83019 1809 83053
rect 1809 83019 1843 83053
rect 1843 83019 1852 83053
rect 1800 83010 1852 83019
rect 136946 83053 136998 83062
rect 136946 83019 136955 83053
rect 136955 83019 136989 83053
rect 136989 83019 136998 83053
rect 136946 83010 136998 83019
rect 1800 82717 1852 82726
rect 1800 82683 1809 82717
rect 1809 82683 1843 82717
rect 1843 82683 1852 82717
rect 1800 82674 1852 82683
rect 136946 82717 136998 82726
rect 136946 82683 136955 82717
rect 136955 82683 136989 82717
rect 136989 82683 136998 82717
rect 136946 82674 136998 82683
rect 1800 82381 1852 82390
rect 1800 82347 1809 82381
rect 1809 82347 1843 82381
rect 1843 82347 1852 82381
rect 1800 82338 1852 82347
rect 136946 82381 136998 82390
rect 136946 82347 136955 82381
rect 136955 82347 136989 82381
rect 136989 82347 136998 82381
rect 136946 82338 136998 82347
rect 1800 82045 1852 82054
rect 1800 82011 1809 82045
rect 1809 82011 1843 82045
rect 1843 82011 1852 82045
rect 1800 82002 1852 82011
rect 136946 82045 136998 82054
rect 136946 82011 136955 82045
rect 136955 82011 136989 82045
rect 136989 82011 136998 82045
rect 136946 82002 136998 82011
rect 1800 81709 1852 81718
rect 1800 81675 1809 81709
rect 1809 81675 1843 81709
rect 1843 81675 1852 81709
rect 1800 81666 1852 81675
rect 136946 81709 136998 81718
rect 136946 81675 136955 81709
rect 136955 81675 136989 81709
rect 136989 81675 136998 81709
rect 136946 81666 136998 81675
rect 1800 81373 1852 81382
rect 1800 81339 1809 81373
rect 1809 81339 1843 81373
rect 1843 81339 1852 81373
rect 1800 81330 1852 81339
rect 136946 81373 136998 81382
rect 136946 81339 136955 81373
rect 136955 81339 136989 81373
rect 136989 81339 136998 81373
rect 136946 81330 136998 81339
rect 1800 81037 1852 81046
rect 1800 81003 1809 81037
rect 1809 81003 1843 81037
rect 1843 81003 1852 81037
rect 1800 80994 1852 81003
rect 136946 81037 136998 81046
rect 136946 81003 136955 81037
rect 136955 81003 136989 81037
rect 136989 81003 136998 81037
rect 136946 80994 136998 81003
rect 1800 80701 1852 80710
rect 1800 80667 1809 80701
rect 1809 80667 1843 80701
rect 1843 80667 1852 80701
rect 1800 80658 1852 80667
rect 136946 80701 136998 80710
rect 136946 80667 136955 80701
rect 136955 80667 136989 80701
rect 136989 80667 136998 80701
rect 136946 80658 136998 80667
rect 1800 80365 1852 80374
rect 1800 80331 1809 80365
rect 1809 80331 1843 80365
rect 1843 80331 1852 80365
rect 1800 80322 1852 80331
rect 136946 80365 136998 80374
rect 136946 80331 136955 80365
rect 136955 80331 136989 80365
rect 136989 80331 136998 80365
rect 136946 80322 136998 80331
rect 1800 80029 1852 80038
rect 1800 79995 1809 80029
rect 1809 79995 1843 80029
rect 1843 79995 1852 80029
rect 1800 79986 1852 79995
rect 136946 80029 136998 80038
rect 136946 79995 136955 80029
rect 136955 79995 136989 80029
rect 136989 79995 136998 80029
rect 136946 79986 136998 79995
rect 1800 79693 1852 79702
rect 1800 79659 1809 79693
rect 1809 79659 1843 79693
rect 1843 79659 1852 79693
rect 1800 79650 1852 79659
rect 136946 79693 136998 79702
rect 136946 79659 136955 79693
rect 136955 79659 136989 79693
rect 136989 79659 136998 79693
rect 136946 79650 136998 79659
rect 1800 79357 1852 79366
rect 1800 79323 1809 79357
rect 1809 79323 1843 79357
rect 1843 79323 1852 79357
rect 1800 79314 1852 79323
rect 136946 79357 136998 79366
rect 136946 79323 136955 79357
rect 136955 79323 136989 79357
rect 136989 79323 136998 79357
rect 136946 79314 136998 79323
rect 1800 79021 1852 79030
rect 1800 78987 1809 79021
rect 1809 78987 1843 79021
rect 1843 78987 1852 79021
rect 1800 78978 1852 78987
rect 136946 79021 136998 79030
rect 136946 78987 136955 79021
rect 136955 78987 136989 79021
rect 136989 78987 136998 79021
rect 136946 78978 136998 78987
rect 1800 78685 1852 78694
rect 1800 78651 1809 78685
rect 1809 78651 1843 78685
rect 1843 78651 1852 78685
rect 1800 78642 1852 78651
rect 136946 78685 136998 78694
rect 136946 78651 136955 78685
rect 136955 78651 136989 78685
rect 136989 78651 136998 78685
rect 136946 78642 136998 78651
rect 1800 78349 1852 78358
rect 1800 78315 1809 78349
rect 1809 78315 1843 78349
rect 1843 78315 1852 78349
rect 1800 78306 1852 78315
rect 136946 78349 136998 78358
rect 136946 78315 136955 78349
rect 136955 78315 136989 78349
rect 136989 78315 136998 78349
rect 136946 78306 136998 78315
rect 1800 78013 1852 78022
rect 1800 77979 1809 78013
rect 1809 77979 1843 78013
rect 1843 77979 1852 78013
rect 1800 77970 1852 77979
rect 136946 78013 136998 78022
rect 136946 77979 136955 78013
rect 136955 77979 136989 78013
rect 136989 77979 136998 78013
rect 136946 77970 136998 77979
rect 1800 77677 1852 77686
rect 1800 77643 1809 77677
rect 1809 77643 1843 77677
rect 1843 77643 1852 77677
rect 1800 77634 1852 77643
rect 136946 77677 136998 77686
rect 136946 77643 136955 77677
rect 136955 77643 136989 77677
rect 136989 77643 136998 77677
rect 136946 77634 136998 77643
rect 1800 77341 1852 77350
rect 1800 77307 1809 77341
rect 1809 77307 1843 77341
rect 1843 77307 1852 77341
rect 1800 77298 1852 77307
rect 136946 77341 136998 77350
rect 136946 77307 136955 77341
rect 136955 77307 136989 77341
rect 136989 77307 136998 77341
rect 136946 77298 136998 77307
rect 1800 77005 1852 77014
rect 1800 76971 1809 77005
rect 1809 76971 1843 77005
rect 1843 76971 1852 77005
rect 1800 76962 1852 76971
rect 136946 77005 136998 77014
rect 136946 76971 136955 77005
rect 136955 76971 136989 77005
rect 136989 76971 136998 77005
rect 136946 76962 136998 76971
rect 1800 76669 1852 76678
rect 1800 76635 1809 76669
rect 1809 76635 1843 76669
rect 1843 76635 1852 76669
rect 1800 76626 1852 76635
rect 136946 76669 136998 76678
rect 136946 76635 136955 76669
rect 136955 76635 136989 76669
rect 136989 76635 136998 76669
rect 136946 76626 136998 76635
rect 1800 76333 1852 76342
rect 1800 76299 1809 76333
rect 1809 76299 1843 76333
rect 1843 76299 1852 76333
rect 1800 76290 1852 76299
rect 136946 76333 136998 76342
rect 136946 76299 136955 76333
rect 136955 76299 136989 76333
rect 136989 76299 136998 76333
rect 136946 76290 136998 76299
rect 1800 75997 1852 76006
rect 1800 75963 1809 75997
rect 1809 75963 1843 75997
rect 1843 75963 1852 75997
rect 1800 75954 1852 75963
rect 136946 75997 136998 76006
rect 136946 75963 136955 75997
rect 136955 75963 136989 75997
rect 136989 75963 136998 75997
rect 136946 75954 136998 75963
rect 1800 75661 1852 75670
rect 1800 75627 1809 75661
rect 1809 75627 1843 75661
rect 1843 75627 1852 75661
rect 1800 75618 1852 75627
rect 136946 75661 136998 75670
rect 136946 75627 136955 75661
rect 136955 75627 136989 75661
rect 136989 75627 136998 75661
rect 136946 75618 136998 75627
rect 1800 75325 1852 75334
rect 1800 75291 1809 75325
rect 1809 75291 1843 75325
rect 1843 75291 1852 75325
rect 1800 75282 1852 75291
rect 136946 75325 136998 75334
rect 136946 75291 136955 75325
rect 136955 75291 136989 75325
rect 136989 75291 136998 75325
rect 136946 75282 136998 75291
rect 1800 74989 1852 74998
rect 1800 74955 1809 74989
rect 1809 74955 1843 74989
rect 1843 74955 1852 74989
rect 1800 74946 1852 74955
rect 136946 74989 136998 74998
rect 136946 74955 136955 74989
rect 136955 74955 136989 74989
rect 136989 74955 136998 74989
rect 136946 74946 136998 74955
rect 1800 74653 1852 74662
rect 1800 74619 1809 74653
rect 1809 74619 1843 74653
rect 1843 74619 1852 74653
rect 1800 74610 1852 74619
rect 136946 74653 136998 74662
rect 136946 74619 136955 74653
rect 136955 74619 136989 74653
rect 136989 74619 136998 74653
rect 136946 74610 136998 74619
rect 1800 74317 1852 74326
rect 1800 74283 1809 74317
rect 1809 74283 1843 74317
rect 1843 74283 1852 74317
rect 1800 74274 1852 74283
rect 136946 74317 136998 74326
rect 136946 74283 136955 74317
rect 136955 74283 136989 74317
rect 136989 74283 136998 74317
rect 136946 74274 136998 74283
rect 1800 73981 1852 73990
rect 1800 73947 1809 73981
rect 1809 73947 1843 73981
rect 1843 73947 1852 73981
rect 1800 73938 1852 73947
rect 136946 73981 136998 73990
rect 136946 73947 136955 73981
rect 136955 73947 136989 73981
rect 136989 73947 136998 73981
rect 136946 73938 136998 73947
rect 1800 73645 1852 73654
rect 1800 73611 1809 73645
rect 1809 73611 1843 73645
rect 1843 73611 1852 73645
rect 1800 73602 1852 73611
rect 136946 73645 136998 73654
rect 136946 73611 136955 73645
rect 136955 73611 136989 73645
rect 136989 73611 136998 73645
rect 136946 73602 136998 73611
rect 1800 73309 1852 73318
rect 1800 73275 1809 73309
rect 1809 73275 1843 73309
rect 1843 73275 1852 73309
rect 1800 73266 1852 73275
rect 136946 73309 136998 73318
rect 136946 73275 136955 73309
rect 136955 73275 136989 73309
rect 136989 73275 136998 73309
rect 136946 73266 136998 73275
rect 1800 72973 1852 72982
rect 1800 72939 1809 72973
rect 1809 72939 1843 72973
rect 1843 72939 1852 72973
rect 1800 72930 1852 72939
rect 136946 72973 136998 72982
rect 136946 72939 136955 72973
rect 136955 72939 136989 72973
rect 136989 72939 136998 72973
rect 136946 72930 136998 72939
rect 1800 72637 1852 72646
rect 1800 72603 1809 72637
rect 1809 72603 1843 72637
rect 1843 72603 1852 72637
rect 1800 72594 1852 72603
rect 136946 72637 136998 72646
rect 136946 72603 136955 72637
rect 136955 72603 136989 72637
rect 136989 72603 136998 72637
rect 136946 72594 136998 72603
rect 1800 72301 1852 72310
rect 1800 72267 1809 72301
rect 1809 72267 1843 72301
rect 1843 72267 1852 72301
rect 1800 72258 1852 72267
rect 136946 72301 136998 72310
rect 136946 72267 136955 72301
rect 136955 72267 136989 72301
rect 136989 72267 136998 72301
rect 136946 72258 136998 72267
rect 1800 71965 1852 71974
rect 1800 71931 1809 71965
rect 1809 71931 1843 71965
rect 1843 71931 1852 71965
rect 1800 71922 1852 71931
rect 136946 71965 136998 71974
rect 136946 71931 136955 71965
rect 136955 71931 136989 71965
rect 136989 71931 136998 71965
rect 136946 71922 136998 71931
rect 1800 71629 1852 71638
rect 1800 71595 1809 71629
rect 1809 71595 1843 71629
rect 1843 71595 1852 71629
rect 1800 71586 1852 71595
rect 136946 71629 136998 71638
rect 136946 71595 136955 71629
rect 136955 71595 136989 71629
rect 136989 71595 136998 71629
rect 136946 71586 136998 71595
rect 1800 71293 1852 71302
rect 1800 71259 1809 71293
rect 1809 71259 1843 71293
rect 1843 71259 1852 71293
rect 1800 71250 1852 71259
rect 136946 71293 136998 71302
rect 136946 71259 136955 71293
rect 136955 71259 136989 71293
rect 136989 71259 136998 71293
rect 136946 71250 136998 71259
rect 1800 70957 1852 70966
rect 1800 70923 1809 70957
rect 1809 70923 1843 70957
rect 1843 70923 1852 70957
rect 1800 70914 1852 70923
rect 136946 70957 136998 70966
rect 136946 70923 136955 70957
rect 136955 70923 136989 70957
rect 136989 70923 136998 70957
rect 136946 70914 136998 70923
rect 1800 70621 1852 70630
rect 1800 70587 1809 70621
rect 1809 70587 1843 70621
rect 1843 70587 1852 70621
rect 1800 70578 1852 70587
rect 136946 70621 136998 70630
rect 136946 70587 136955 70621
rect 136955 70587 136989 70621
rect 136989 70587 136998 70621
rect 136946 70578 136998 70587
rect 1800 70285 1852 70294
rect 1800 70251 1809 70285
rect 1809 70251 1843 70285
rect 1843 70251 1852 70285
rect 1800 70242 1852 70251
rect 136946 70285 136998 70294
rect 136946 70251 136955 70285
rect 136955 70251 136989 70285
rect 136989 70251 136998 70285
rect 136946 70242 136998 70251
rect 1800 69949 1852 69958
rect 1800 69915 1809 69949
rect 1809 69915 1843 69949
rect 1843 69915 1852 69949
rect 1800 69906 1852 69915
rect 136946 69949 136998 69958
rect 136946 69915 136955 69949
rect 136955 69915 136989 69949
rect 136989 69915 136998 69949
rect 136946 69906 136998 69915
rect 1800 69613 1852 69622
rect 1800 69579 1809 69613
rect 1809 69579 1843 69613
rect 1843 69579 1852 69613
rect 1800 69570 1852 69579
rect 136946 69613 136998 69622
rect 136946 69579 136955 69613
rect 136955 69579 136989 69613
rect 136989 69579 136998 69613
rect 136946 69570 136998 69579
rect 1800 69277 1852 69286
rect 1800 69243 1809 69277
rect 1809 69243 1843 69277
rect 1843 69243 1852 69277
rect 1800 69234 1852 69243
rect 136946 69277 136998 69286
rect 136946 69243 136955 69277
rect 136955 69243 136989 69277
rect 136989 69243 136998 69277
rect 136946 69234 136998 69243
rect 1800 68941 1852 68950
rect 1800 68907 1809 68941
rect 1809 68907 1843 68941
rect 1843 68907 1852 68941
rect 1800 68898 1852 68907
rect 136946 68941 136998 68950
rect 136946 68907 136955 68941
rect 136955 68907 136989 68941
rect 136989 68907 136998 68941
rect 136946 68898 136998 68907
rect 1800 68605 1852 68614
rect 1800 68571 1809 68605
rect 1809 68571 1843 68605
rect 1843 68571 1852 68605
rect 1800 68562 1852 68571
rect 136946 68605 136998 68614
rect 136946 68571 136955 68605
rect 136955 68571 136989 68605
rect 136989 68571 136998 68605
rect 136946 68562 136998 68571
rect 1800 68269 1852 68278
rect 1800 68235 1809 68269
rect 1809 68235 1843 68269
rect 1843 68235 1852 68269
rect 1800 68226 1852 68235
rect 136946 68269 136998 68278
rect 136946 68235 136955 68269
rect 136955 68235 136989 68269
rect 136989 68235 136998 68269
rect 136946 68226 136998 68235
rect 1800 67933 1852 67942
rect 1800 67899 1809 67933
rect 1809 67899 1843 67933
rect 1843 67899 1852 67933
rect 1800 67890 1852 67899
rect 136946 67933 136998 67942
rect 136946 67899 136955 67933
rect 136955 67899 136989 67933
rect 136989 67899 136998 67933
rect 136946 67890 136998 67899
rect 1800 67597 1852 67606
rect 1800 67563 1809 67597
rect 1809 67563 1843 67597
rect 1843 67563 1852 67597
rect 1800 67554 1852 67563
rect 136946 67597 136998 67606
rect 136946 67563 136955 67597
rect 136955 67563 136989 67597
rect 136989 67563 136998 67597
rect 136946 67554 136998 67563
rect 1800 67261 1852 67270
rect 1800 67227 1809 67261
rect 1809 67227 1843 67261
rect 1843 67227 1852 67261
rect 1800 67218 1852 67227
rect 136946 67261 136998 67270
rect 136946 67227 136955 67261
rect 136955 67227 136989 67261
rect 136989 67227 136998 67261
rect 136946 67218 136998 67227
rect 1800 66925 1852 66934
rect 1800 66891 1809 66925
rect 1809 66891 1843 66925
rect 1843 66891 1852 66925
rect 1800 66882 1852 66891
rect 136946 66925 136998 66934
rect 136946 66891 136955 66925
rect 136955 66891 136989 66925
rect 136989 66891 136998 66925
rect 136946 66882 136998 66891
rect 1800 66589 1852 66598
rect 1800 66555 1809 66589
rect 1809 66555 1843 66589
rect 1843 66555 1852 66589
rect 1800 66546 1852 66555
rect 136946 66589 136998 66598
rect 136946 66555 136955 66589
rect 136955 66555 136989 66589
rect 136989 66555 136998 66589
rect 136946 66546 136998 66555
rect 1800 66253 1852 66262
rect 1800 66219 1809 66253
rect 1809 66219 1843 66253
rect 1843 66219 1852 66253
rect 1800 66210 1852 66219
rect 136946 66253 136998 66262
rect 136946 66219 136955 66253
rect 136955 66219 136989 66253
rect 136989 66219 136998 66253
rect 136946 66210 136998 66219
rect 1800 65917 1852 65926
rect 1800 65883 1809 65917
rect 1809 65883 1843 65917
rect 1843 65883 1852 65917
rect 1800 65874 1852 65883
rect 136946 65917 136998 65926
rect 136946 65883 136955 65917
rect 136955 65883 136989 65917
rect 136989 65883 136998 65917
rect 136946 65874 136998 65883
rect 1800 65581 1852 65590
rect 1800 65547 1809 65581
rect 1809 65547 1843 65581
rect 1843 65547 1852 65581
rect 1800 65538 1852 65547
rect 136946 65581 136998 65590
rect 136946 65547 136955 65581
rect 136955 65547 136989 65581
rect 136989 65547 136998 65581
rect 136946 65538 136998 65547
rect 1800 65245 1852 65254
rect 1800 65211 1809 65245
rect 1809 65211 1843 65245
rect 1843 65211 1852 65245
rect 1800 65202 1852 65211
rect 136946 65245 136998 65254
rect 136946 65211 136955 65245
rect 136955 65211 136989 65245
rect 136989 65211 136998 65245
rect 136946 65202 136998 65211
rect 1800 64909 1852 64918
rect 1800 64875 1809 64909
rect 1809 64875 1843 64909
rect 1843 64875 1852 64909
rect 1800 64866 1852 64875
rect 136946 64909 136998 64918
rect 136946 64875 136955 64909
rect 136955 64875 136989 64909
rect 136989 64875 136998 64909
rect 136946 64866 136998 64875
rect 1800 64573 1852 64582
rect 1800 64539 1809 64573
rect 1809 64539 1843 64573
rect 1843 64539 1852 64573
rect 1800 64530 1852 64539
rect 136946 64573 136998 64582
rect 136946 64539 136955 64573
rect 136955 64539 136989 64573
rect 136989 64539 136998 64573
rect 136946 64530 136998 64539
rect 1800 64237 1852 64246
rect 1800 64203 1809 64237
rect 1809 64203 1843 64237
rect 1843 64203 1852 64237
rect 1800 64194 1852 64203
rect 136946 64237 136998 64246
rect 136946 64203 136955 64237
rect 136955 64203 136989 64237
rect 136989 64203 136998 64237
rect 136946 64194 136998 64203
rect 1800 63901 1852 63910
rect 1800 63867 1809 63901
rect 1809 63867 1843 63901
rect 1843 63867 1852 63901
rect 1800 63858 1852 63867
rect 136946 63901 136998 63910
rect 136946 63867 136955 63901
rect 136955 63867 136989 63901
rect 136989 63867 136998 63901
rect 136946 63858 136998 63867
rect 1800 63565 1852 63574
rect 1800 63531 1809 63565
rect 1809 63531 1843 63565
rect 1843 63531 1852 63565
rect 1800 63522 1852 63531
rect 136946 63565 136998 63574
rect 136946 63531 136955 63565
rect 136955 63531 136989 63565
rect 136989 63531 136998 63565
rect 136946 63522 136998 63531
rect 1800 63229 1852 63238
rect 1800 63195 1809 63229
rect 1809 63195 1843 63229
rect 1843 63195 1852 63229
rect 1800 63186 1852 63195
rect 136946 63229 136998 63238
rect 136946 63195 136955 63229
rect 136955 63195 136989 63229
rect 136989 63195 136998 63229
rect 136946 63186 136998 63195
rect 1800 62893 1852 62902
rect 1800 62859 1809 62893
rect 1809 62859 1843 62893
rect 1843 62859 1852 62893
rect 1800 62850 1852 62859
rect 136946 62893 136998 62902
rect 136946 62859 136955 62893
rect 136955 62859 136989 62893
rect 136989 62859 136998 62893
rect 136946 62850 136998 62859
rect 1800 62557 1852 62566
rect 1800 62523 1809 62557
rect 1809 62523 1843 62557
rect 1843 62523 1852 62557
rect 1800 62514 1852 62523
rect 136946 62557 136998 62566
rect 136946 62523 136955 62557
rect 136955 62523 136989 62557
rect 136989 62523 136998 62557
rect 136946 62514 136998 62523
rect 1800 62221 1852 62230
rect 1800 62187 1809 62221
rect 1809 62187 1843 62221
rect 1843 62187 1852 62221
rect 1800 62178 1852 62187
rect 136946 62221 136998 62230
rect 136946 62187 136955 62221
rect 136955 62187 136989 62221
rect 136989 62187 136998 62221
rect 136946 62178 136998 62187
rect 1800 61885 1852 61894
rect 1800 61851 1809 61885
rect 1809 61851 1843 61885
rect 1843 61851 1852 61885
rect 1800 61842 1852 61851
rect 136946 61885 136998 61894
rect 136946 61851 136955 61885
rect 136955 61851 136989 61885
rect 136989 61851 136998 61885
rect 136946 61842 136998 61851
rect 1800 61549 1852 61558
rect 1800 61515 1809 61549
rect 1809 61515 1843 61549
rect 1843 61515 1852 61549
rect 1800 61506 1852 61515
rect 136946 61549 136998 61558
rect 136946 61515 136955 61549
rect 136955 61515 136989 61549
rect 136989 61515 136998 61549
rect 136946 61506 136998 61515
rect 1800 61213 1852 61222
rect 1800 61179 1809 61213
rect 1809 61179 1843 61213
rect 1843 61179 1852 61213
rect 1800 61170 1852 61179
rect 136946 61213 136998 61222
rect 136946 61179 136955 61213
rect 136955 61179 136989 61213
rect 136989 61179 136998 61213
rect 136946 61170 136998 61179
rect 1800 60877 1852 60886
rect 1800 60843 1809 60877
rect 1809 60843 1843 60877
rect 1843 60843 1852 60877
rect 1800 60834 1852 60843
rect 136946 60877 136998 60886
rect 136946 60843 136955 60877
rect 136955 60843 136989 60877
rect 136989 60843 136998 60877
rect 136946 60834 136998 60843
rect 1800 60541 1852 60550
rect 1800 60507 1809 60541
rect 1809 60507 1843 60541
rect 1843 60507 1852 60541
rect 1800 60498 1852 60507
rect 136946 60541 136998 60550
rect 136946 60507 136955 60541
rect 136955 60507 136989 60541
rect 136989 60507 136998 60541
rect 136946 60498 136998 60507
rect 1800 60205 1852 60214
rect 1800 60171 1809 60205
rect 1809 60171 1843 60205
rect 1843 60171 1852 60205
rect 1800 60162 1852 60171
rect 136946 60205 136998 60214
rect 136946 60171 136955 60205
rect 136955 60171 136989 60205
rect 136989 60171 136998 60205
rect 136946 60162 136998 60171
rect 1800 59869 1852 59878
rect 1800 59835 1809 59869
rect 1809 59835 1843 59869
rect 1843 59835 1852 59869
rect 1800 59826 1852 59835
rect 136946 59869 136998 59878
rect 136946 59835 136955 59869
rect 136955 59835 136989 59869
rect 136989 59835 136998 59869
rect 136946 59826 136998 59835
rect 1800 59533 1852 59542
rect 1800 59499 1809 59533
rect 1809 59499 1843 59533
rect 1843 59499 1852 59533
rect 1800 59490 1852 59499
rect 136946 59533 136998 59542
rect 136946 59499 136955 59533
rect 136955 59499 136989 59533
rect 136989 59499 136998 59533
rect 136946 59490 136998 59499
rect 1800 59197 1852 59206
rect 1800 59163 1809 59197
rect 1809 59163 1843 59197
rect 1843 59163 1852 59197
rect 1800 59154 1852 59163
rect 136946 59197 136998 59206
rect 136946 59163 136955 59197
rect 136955 59163 136989 59197
rect 136989 59163 136998 59197
rect 136946 59154 136998 59163
rect 1800 58861 1852 58870
rect 1800 58827 1809 58861
rect 1809 58827 1843 58861
rect 1843 58827 1852 58861
rect 1800 58818 1852 58827
rect 136946 58861 136998 58870
rect 136946 58827 136955 58861
rect 136955 58827 136989 58861
rect 136989 58827 136998 58861
rect 136946 58818 136998 58827
rect 1800 58525 1852 58534
rect 1800 58491 1809 58525
rect 1809 58491 1843 58525
rect 1843 58491 1852 58525
rect 1800 58482 1852 58491
rect 136946 58525 136998 58534
rect 136946 58491 136955 58525
rect 136955 58491 136989 58525
rect 136989 58491 136998 58525
rect 136946 58482 136998 58491
rect 1800 58189 1852 58198
rect 1800 58155 1809 58189
rect 1809 58155 1843 58189
rect 1843 58155 1852 58189
rect 1800 58146 1852 58155
rect 136946 58189 136998 58198
rect 136946 58155 136955 58189
rect 136955 58155 136989 58189
rect 136989 58155 136998 58189
rect 136946 58146 136998 58155
rect 1800 57853 1852 57862
rect 1800 57819 1809 57853
rect 1809 57819 1843 57853
rect 1843 57819 1852 57853
rect 1800 57810 1852 57819
rect 136946 57853 136998 57862
rect 136946 57819 136955 57853
rect 136955 57819 136989 57853
rect 136989 57819 136998 57853
rect 136946 57810 136998 57819
rect 1800 57517 1852 57526
rect 1800 57483 1809 57517
rect 1809 57483 1843 57517
rect 1843 57483 1852 57517
rect 1800 57474 1852 57483
rect 136946 57517 136998 57526
rect 136946 57483 136955 57517
rect 136955 57483 136989 57517
rect 136989 57483 136998 57517
rect 136946 57474 136998 57483
rect 1800 57181 1852 57190
rect 1800 57147 1809 57181
rect 1809 57147 1843 57181
rect 1843 57147 1852 57181
rect 1800 57138 1852 57147
rect 136946 57181 136998 57190
rect 136946 57147 136955 57181
rect 136955 57147 136989 57181
rect 136989 57147 136998 57181
rect 136946 57138 136998 57147
rect 1800 56845 1852 56854
rect 1800 56811 1809 56845
rect 1809 56811 1843 56845
rect 1843 56811 1852 56845
rect 1800 56802 1852 56811
rect 136946 56845 136998 56854
rect 136946 56811 136955 56845
rect 136955 56811 136989 56845
rect 136989 56811 136998 56845
rect 136946 56802 136998 56811
rect 1800 56509 1852 56518
rect 1800 56475 1809 56509
rect 1809 56475 1843 56509
rect 1843 56475 1852 56509
rect 1800 56466 1852 56475
rect 136946 56509 136998 56518
rect 136946 56475 136955 56509
rect 136955 56475 136989 56509
rect 136989 56475 136998 56509
rect 136946 56466 136998 56475
rect 1800 56173 1852 56182
rect 1800 56139 1809 56173
rect 1809 56139 1843 56173
rect 1843 56139 1852 56173
rect 1800 56130 1852 56139
rect 136946 56173 136998 56182
rect 136946 56139 136955 56173
rect 136955 56139 136989 56173
rect 136989 56139 136998 56173
rect 136946 56130 136998 56139
rect 1800 55837 1852 55846
rect 1800 55803 1809 55837
rect 1809 55803 1843 55837
rect 1843 55803 1852 55837
rect 1800 55794 1852 55803
rect 136946 55837 136998 55846
rect 136946 55803 136955 55837
rect 136955 55803 136989 55837
rect 136989 55803 136998 55837
rect 136946 55794 136998 55803
rect 1800 55501 1852 55510
rect 1800 55467 1809 55501
rect 1809 55467 1843 55501
rect 1843 55467 1852 55501
rect 1800 55458 1852 55467
rect 136946 55501 136998 55510
rect 136946 55467 136955 55501
rect 136955 55467 136989 55501
rect 136989 55467 136998 55501
rect 136946 55458 136998 55467
rect 1800 55165 1852 55174
rect 1800 55131 1809 55165
rect 1809 55131 1843 55165
rect 1843 55131 1852 55165
rect 1800 55122 1852 55131
rect 136946 55165 136998 55174
rect 136946 55131 136955 55165
rect 136955 55131 136989 55165
rect 136989 55131 136998 55165
rect 136946 55122 136998 55131
rect 1800 54829 1852 54838
rect 1800 54795 1809 54829
rect 1809 54795 1843 54829
rect 1843 54795 1852 54829
rect 1800 54786 1852 54795
rect 136946 54829 136998 54838
rect 136946 54795 136955 54829
rect 136955 54795 136989 54829
rect 136989 54795 136998 54829
rect 136946 54786 136998 54795
rect 1800 54493 1852 54502
rect 1800 54459 1809 54493
rect 1809 54459 1843 54493
rect 1843 54459 1852 54493
rect 1800 54450 1852 54459
rect 136946 54493 136998 54502
rect 136946 54459 136955 54493
rect 136955 54459 136989 54493
rect 136989 54459 136998 54493
rect 136946 54450 136998 54459
rect 1800 54157 1852 54166
rect 1800 54123 1809 54157
rect 1809 54123 1843 54157
rect 1843 54123 1852 54157
rect 1800 54114 1852 54123
rect 136946 54157 136998 54166
rect 136946 54123 136955 54157
rect 136955 54123 136989 54157
rect 136989 54123 136998 54157
rect 136946 54114 136998 54123
rect 1800 53821 1852 53830
rect 1800 53787 1809 53821
rect 1809 53787 1843 53821
rect 1843 53787 1852 53821
rect 1800 53778 1852 53787
rect 136946 53821 136998 53830
rect 136946 53787 136955 53821
rect 136955 53787 136989 53821
rect 136989 53787 136998 53821
rect 136946 53778 136998 53787
rect 1800 53485 1852 53494
rect 1800 53451 1809 53485
rect 1809 53451 1843 53485
rect 1843 53451 1852 53485
rect 1800 53442 1852 53451
rect 136946 53485 136998 53494
rect 136946 53451 136955 53485
rect 136955 53451 136989 53485
rect 136989 53451 136998 53485
rect 136946 53442 136998 53451
rect 1800 53149 1852 53158
rect 1800 53115 1809 53149
rect 1809 53115 1843 53149
rect 1843 53115 1852 53149
rect 1800 53106 1852 53115
rect 136946 53149 136998 53158
rect 136946 53115 136955 53149
rect 136955 53115 136989 53149
rect 136989 53115 136998 53149
rect 136946 53106 136998 53115
rect 1800 52813 1852 52822
rect 1800 52779 1809 52813
rect 1809 52779 1843 52813
rect 1843 52779 1852 52813
rect 1800 52770 1852 52779
rect 136946 52813 136998 52822
rect 136946 52779 136955 52813
rect 136955 52779 136989 52813
rect 136989 52779 136998 52813
rect 136946 52770 136998 52779
rect 1800 52477 1852 52486
rect 1800 52443 1809 52477
rect 1809 52443 1843 52477
rect 1843 52443 1852 52477
rect 1800 52434 1852 52443
rect 136946 52477 136998 52486
rect 136946 52443 136955 52477
rect 136955 52443 136989 52477
rect 136989 52443 136998 52477
rect 136946 52434 136998 52443
rect 1800 52141 1852 52150
rect 1800 52107 1809 52141
rect 1809 52107 1843 52141
rect 1843 52107 1852 52141
rect 1800 52098 1852 52107
rect 136946 52141 136998 52150
rect 136946 52107 136955 52141
rect 136955 52107 136989 52141
rect 136989 52107 136998 52141
rect 136946 52098 136998 52107
rect 1800 51805 1852 51814
rect 1800 51771 1809 51805
rect 1809 51771 1843 51805
rect 1843 51771 1852 51805
rect 1800 51762 1852 51771
rect 136946 51805 136998 51814
rect 136946 51771 136955 51805
rect 136955 51771 136989 51805
rect 136989 51771 136998 51805
rect 136946 51762 136998 51771
rect 1800 51469 1852 51478
rect 1800 51435 1809 51469
rect 1809 51435 1843 51469
rect 1843 51435 1852 51469
rect 1800 51426 1852 51435
rect 136946 51469 136998 51478
rect 136946 51435 136955 51469
rect 136955 51435 136989 51469
rect 136989 51435 136998 51469
rect 136946 51426 136998 51435
rect 1800 51133 1852 51142
rect 1800 51099 1809 51133
rect 1809 51099 1843 51133
rect 1843 51099 1852 51133
rect 1800 51090 1852 51099
rect 136946 51133 136998 51142
rect 136946 51099 136955 51133
rect 136955 51099 136989 51133
rect 136989 51099 136998 51133
rect 136946 51090 136998 51099
rect 1800 50797 1852 50806
rect 1800 50763 1809 50797
rect 1809 50763 1843 50797
rect 1843 50763 1852 50797
rect 1800 50754 1852 50763
rect 136946 50797 136998 50806
rect 136946 50763 136955 50797
rect 136955 50763 136989 50797
rect 136989 50763 136998 50797
rect 136946 50754 136998 50763
rect 1800 50461 1852 50470
rect 1800 50427 1809 50461
rect 1809 50427 1843 50461
rect 1843 50427 1852 50461
rect 1800 50418 1852 50427
rect 136946 50461 136998 50470
rect 136946 50427 136955 50461
rect 136955 50427 136989 50461
rect 136989 50427 136998 50461
rect 136946 50418 136998 50427
rect 1800 50125 1852 50134
rect 1800 50091 1809 50125
rect 1809 50091 1843 50125
rect 1843 50091 1852 50125
rect 1800 50082 1852 50091
rect 136946 50125 136998 50134
rect 136946 50091 136955 50125
rect 136955 50091 136989 50125
rect 136989 50091 136998 50125
rect 136946 50082 136998 50091
rect 1800 49789 1852 49798
rect 1800 49755 1809 49789
rect 1809 49755 1843 49789
rect 1843 49755 1852 49789
rect 1800 49746 1852 49755
rect 136946 49789 136998 49798
rect 136946 49755 136955 49789
rect 136955 49755 136989 49789
rect 136989 49755 136998 49789
rect 136946 49746 136998 49755
rect 1800 49453 1852 49462
rect 1800 49419 1809 49453
rect 1809 49419 1843 49453
rect 1843 49419 1852 49453
rect 1800 49410 1852 49419
rect 136946 49453 136998 49462
rect 136946 49419 136955 49453
rect 136955 49419 136989 49453
rect 136989 49419 136998 49453
rect 136946 49410 136998 49419
rect 1800 49117 1852 49126
rect 1800 49083 1809 49117
rect 1809 49083 1843 49117
rect 1843 49083 1852 49117
rect 1800 49074 1852 49083
rect 136946 49117 136998 49126
rect 136946 49083 136955 49117
rect 136955 49083 136989 49117
rect 136989 49083 136998 49117
rect 136946 49074 136998 49083
rect 1800 48781 1852 48790
rect 1800 48747 1809 48781
rect 1809 48747 1843 48781
rect 1843 48747 1852 48781
rect 1800 48738 1852 48747
rect 136946 48781 136998 48790
rect 136946 48747 136955 48781
rect 136955 48747 136989 48781
rect 136989 48747 136998 48781
rect 136946 48738 136998 48747
rect 1800 48445 1852 48454
rect 1800 48411 1809 48445
rect 1809 48411 1843 48445
rect 1843 48411 1852 48445
rect 1800 48402 1852 48411
rect 136946 48445 136998 48454
rect 136946 48411 136955 48445
rect 136955 48411 136989 48445
rect 136989 48411 136998 48445
rect 136946 48402 136998 48411
rect 1800 48109 1852 48118
rect 1800 48075 1809 48109
rect 1809 48075 1843 48109
rect 1843 48075 1852 48109
rect 1800 48066 1852 48075
rect 136946 48109 136998 48118
rect 136946 48075 136955 48109
rect 136955 48075 136989 48109
rect 136989 48075 136998 48109
rect 136946 48066 136998 48075
rect 1800 47773 1852 47782
rect 1800 47739 1809 47773
rect 1809 47739 1843 47773
rect 1843 47739 1852 47773
rect 1800 47730 1852 47739
rect 136946 47773 136998 47782
rect 136946 47739 136955 47773
rect 136955 47739 136989 47773
rect 136989 47739 136998 47773
rect 136946 47730 136998 47739
rect 1800 47437 1852 47446
rect 1800 47403 1809 47437
rect 1809 47403 1843 47437
rect 1843 47403 1852 47437
rect 1800 47394 1852 47403
rect 136946 47437 136998 47446
rect 136946 47403 136955 47437
rect 136955 47403 136989 47437
rect 136989 47403 136998 47437
rect 136946 47394 136998 47403
rect 1800 47101 1852 47110
rect 1800 47067 1809 47101
rect 1809 47067 1843 47101
rect 1843 47067 1852 47101
rect 1800 47058 1852 47067
rect 136946 47101 136998 47110
rect 136946 47067 136955 47101
rect 136955 47067 136989 47101
rect 136989 47067 136998 47101
rect 136946 47058 136998 47067
rect 1800 46765 1852 46774
rect 1800 46731 1809 46765
rect 1809 46731 1843 46765
rect 1843 46731 1852 46765
rect 1800 46722 1852 46731
rect 136946 46765 136998 46774
rect 136946 46731 136955 46765
rect 136955 46731 136989 46765
rect 136989 46731 136998 46765
rect 136946 46722 136998 46731
rect 1800 46429 1852 46438
rect 1800 46395 1809 46429
rect 1809 46395 1843 46429
rect 1843 46395 1852 46429
rect 1800 46386 1852 46395
rect 136946 46429 136998 46438
rect 136946 46395 136955 46429
rect 136955 46395 136989 46429
rect 136989 46395 136998 46429
rect 136946 46386 136998 46395
rect 1800 46093 1852 46102
rect 1800 46059 1809 46093
rect 1809 46059 1843 46093
rect 1843 46059 1852 46093
rect 1800 46050 1852 46059
rect 136946 46093 136998 46102
rect 136946 46059 136955 46093
rect 136955 46059 136989 46093
rect 136989 46059 136998 46093
rect 136946 46050 136998 46059
rect 1800 45757 1852 45766
rect 1800 45723 1809 45757
rect 1809 45723 1843 45757
rect 1843 45723 1852 45757
rect 1800 45714 1852 45723
rect 136946 45757 136998 45766
rect 136946 45723 136955 45757
rect 136955 45723 136989 45757
rect 136989 45723 136998 45757
rect 136946 45714 136998 45723
rect 1800 45421 1852 45430
rect 1800 45387 1809 45421
rect 1809 45387 1843 45421
rect 1843 45387 1852 45421
rect 1800 45378 1852 45387
rect 136946 45421 136998 45430
rect 136946 45387 136955 45421
rect 136955 45387 136989 45421
rect 136989 45387 136998 45421
rect 136946 45378 136998 45387
rect 1800 45085 1852 45094
rect 1800 45051 1809 45085
rect 1809 45051 1843 45085
rect 1843 45051 1852 45085
rect 1800 45042 1852 45051
rect 136946 45085 136998 45094
rect 136946 45051 136955 45085
rect 136955 45051 136989 45085
rect 136989 45051 136998 45085
rect 136946 45042 136998 45051
rect 1800 44749 1852 44758
rect 1800 44715 1809 44749
rect 1809 44715 1843 44749
rect 1843 44715 1852 44749
rect 1800 44706 1852 44715
rect 136946 44749 136998 44758
rect 136946 44715 136955 44749
rect 136955 44715 136989 44749
rect 136989 44715 136998 44749
rect 136946 44706 136998 44715
rect 1800 44413 1852 44422
rect 1800 44379 1809 44413
rect 1809 44379 1843 44413
rect 1843 44379 1852 44413
rect 1800 44370 1852 44379
rect 136946 44413 136998 44422
rect 136946 44379 136955 44413
rect 136955 44379 136989 44413
rect 136989 44379 136998 44413
rect 136946 44370 136998 44379
rect 1800 44077 1852 44086
rect 1800 44043 1809 44077
rect 1809 44043 1843 44077
rect 1843 44043 1852 44077
rect 1800 44034 1852 44043
rect 136946 44077 136998 44086
rect 136946 44043 136955 44077
rect 136955 44043 136989 44077
rect 136989 44043 136998 44077
rect 136946 44034 136998 44043
rect 1800 43741 1852 43750
rect 1800 43707 1809 43741
rect 1809 43707 1843 43741
rect 1843 43707 1852 43741
rect 1800 43698 1852 43707
rect 136946 43741 136998 43750
rect 136946 43707 136955 43741
rect 136955 43707 136989 43741
rect 136989 43707 136998 43741
rect 136946 43698 136998 43707
rect 1800 43405 1852 43414
rect 1800 43371 1809 43405
rect 1809 43371 1843 43405
rect 1843 43371 1852 43405
rect 1800 43362 1852 43371
rect 136946 43405 136998 43414
rect 136946 43371 136955 43405
rect 136955 43371 136989 43405
rect 136989 43371 136998 43405
rect 136946 43362 136998 43371
rect 1800 43069 1852 43078
rect 1800 43035 1809 43069
rect 1809 43035 1843 43069
rect 1843 43035 1852 43069
rect 1800 43026 1852 43035
rect 136946 43069 136998 43078
rect 136946 43035 136955 43069
rect 136955 43035 136989 43069
rect 136989 43035 136998 43069
rect 136946 43026 136998 43035
rect 1800 42733 1852 42742
rect 1800 42699 1809 42733
rect 1809 42699 1843 42733
rect 1843 42699 1852 42733
rect 1800 42690 1852 42699
rect 136946 42733 136998 42742
rect 136946 42699 136955 42733
rect 136955 42699 136989 42733
rect 136989 42699 136998 42733
rect 136946 42690 136998 42699
rect 1800 42397 1852 42406
rect 1800 42363 1809 42397
rect 1809 42363 1843 42397
rect 1843 42363 1852 42397
rect 1800 42354 1852 42363
rect 136946 42397 136998 42406
rect 136946 42363 136955 42397
rect 136955 42363 136989 42397
rect 136989 42363 136998 42397
rect 136946 42354 136998 42363
rect 1800 42061 1852 42070
rect 1800 42027 1809 42061
rect 1809 42027 1843 42061
rect 1843 42027 1852 42061
rect 1800 42018 1852 42027
rect 136946 42061 136998 42070
rect 136946 42027 136955 42061
rect 136955 42027 136989 42061
rect 136989 42027 136998 42061
rect 136946 42018 136998 42027
rect 1800 41725 1852 41734
rect 1800 41691 1809 41725
rect 1809 41691 1843 41725
rect 1843 41691 1852 41725
rect 1800 41682 1852 41691
rect 136946 41725 136998 41734
rect 136946 41691 136955 41725
rect 136955 41691 136989 41725
rect 136989 41691 136998 41725
rect 136946 41682 136998 41691
rect 1800 41389 1852 41398
rect 1800 41355 1809 41389
rect 1809 41355 1843 41389
rect 1843 41355 1852 41389
rect 1800 41346 1852 41355
rect 136946 41389 136998 41398
rect 136946 41355 136955 41389
rect 136955 41355 136989 41389
rect 136989 41355 136998 41389
rect 136946 41346 136998 41355
rect 1800 41053 1852 41062
rect 1800 41019 1809 41053
rect 1809 41019 1843 41053
rect 1843 41019 1852 41053
rect 1800 41010 1852 41019
rect 136946 41053 136998 41062
rect 136946 41019 136955 41053
rect 136955 41019 136989 41053
rect 136989 41019 136998 41053
rect 136946 41010 136998 41019
rect 1800 40717 1852 40726
rect 1800 40683 1809 40717
rect 1809 40683 1843 40717
rect 1843 40683 1852 40717
rect 1800 40674 1852 40683
rect 136946 40717 136998 40726
rect 136946 40683 136955 40717
rect 136955 40683 136989 40717
rect 136989 40683 136998 40717
rect 136946 40674 136998 40683
rect 1800 40381 1852 40390
rect 1800 40347 1809 40381
rect 1809 40347 1843 40381
rect 1843 40347 1852 40381
rect 1800 40338 1852 40347
rect 136946 40381 136998 40390
rect 136946 40347 136955 40381
rect 136955 40347 136989 40381
rect 136989 40347 136998 40381
rect 136946 40338 136998 40347
rect 1800 40045 1852 40054
rect 1800 40011 1809 40045
rect 1809 40011 1843 40045
rect 1843 40011 1852 40045
rect 1800 40002 1852 40011
rect 15973 39977 16025 40029
rect 136946 40045 136998 40054
rect 136946 40011 136955 40045
rect 136955 40011 136989 40045
rect 136989 40011 136998 40045
rect 136946 40002 136998 40011
rect 1800 39709 1852 39718
rect 1800 39675 1809 39709
rect 1809 39675 1843 39709
rect 1843 39675 1852 39709
rect 1800 39666 1852 39675
rect 1800 39373 1852 39382
rect 1800 39339 1809 39373
rect 1809 39339 1843 39373
rect 1843 39339 1852 39373
rect 1800 39330 1852 39339
rect 1800 39037 1852 39046
rect 1800 39003 1809 39037
rect 1809 39003 1843 39037
rect 1843 39003 1852 39037
rect 1800 38994 1852 39003
rect 1800 38701 1852 38710
rect 1800 38667 1809 38701
rect 1809 38667 1843 38701
rect 1843 38667 1852 38701
rect 1800 38658 1852 38667
rect 15893 38419 15945 38471
rect 1800 38365 1852 38374
rect 1800 38331 1809 38365
rect 1809 38331 1843 38365
rect 1843 38331 1852 38365
rect 1800 38322 1852 38331
rect 1800 38029 1852 38038
rect 1800 37995 1809 38029
rect 1809 37995 1843 38029
rect 1843 37995 1852 38029
rect 1800 37986 1852 37995
rect 1800 37693 1852 37702
rect 1800 37659 1809 37693
rect 1809 37659 1843 37693
rect 1843 37659 1852 37693
rect 1800 37650 1852 37659
rect 1800 37357 1852 37366
rect 1800 37323 1809 37357
rect 1809 37323 1843 37357
rect 1843 37323 1852 37357
rect 1800 37314 1852 37323
rect 15813 37149 15865 37201
rect 1800 37021 1852 37030
rect 1800 36987 1809 37021
rect 1809 36987 1843 37021
rect 1843 36987 1852 37021
rect 1800 36978 1852 36987
rect 1800 36685 1852 36694
rect 1800 36651 1809 36685
rect 1809 36651 1843 36685
rect 1843 36651 1852 36685
rect 1800 36642 1852 36651
rect 1800 36349 1852 36358
rect 1800 36315 1809 36349
rect 1809 36315 1843 36349
rect 1843 36315 1852 36349
rect 1800 36306 1852 36315
rect 1800 36013 1852 36022
rect 1800 35979 1809 36013
rect 1809 35979 1843 36013
rect 1843 35979 1852 36013
rect 1800 35970 1852 35979
rect 1800 35677 1852 35686
rect 1800 35643 1809 35677
rect 1809 35643 1843 35677
rect 1843 35643 1852 35677
rect 1800 35634 1852 35643
rect 15733 35591 15785 35643
rect 1800 35341 1852 35350
rect 1800 35307 1809 35341
rect 1809 35307 1843 35341
rect 1843 35307 1852 35341
rect 1800 35298 1852 35307
rect 1800 35005 1852 35014
rect 1800 34971 1809 35005
rect 1809 34971 1843 35005
rect 1843 34971 1852 35005
rect 1800 34962 1852 34971
rect 1800 34669 1852 34678
rect 1800 34635 1809 34669
rect 1809 34635 1843 34669
rect 1843 34635 1852 34669
rect 1800 34626 1852 34635
rect 1800 34333 1852 34342
rect 1800 34299 1809 34333
rect 1809 34299 1843 34333
rect 1843 34299 1852 34333
rect 1800 34290 1852 34299
rect 15653 34321 15705 34373
rect 1800 33997 1852 34006
rect 1800 33963 1809 33997
rect 1809 33963 1843 33997
rect 1843 33963 1852 33997
rect 1800 33954 1852 33963
rect 1800 33661 1852 33670
rect 1800 33627 1809 33661
rect 1809 33627 1843 33661
rect 1843 33627 1852 33661
rect 1800 33618 1852 33627
rect 1800 33325 1852 33334
rect 1800 33291 1809 33325
rect 1809 33291 1843 33325
rect 1843 33291 1852 33325
rect 1800 33282 1852 33291
rect 1800 32989 1852 32998
rect 1800 32955 1809 32989
rect 1809 32955 1843 32989
rect 1843 32955 1852 32989
rect 1800 32946 1852 32955
rect 15573 32763 15625 32815
rect 1800 32653 1852 32662
rect 1800 32619 1809 32653
rect 1809 32619 1843 32653
rect 1843 32619 1852 32653
rect 1800 32610 1852 32619
rect 1800 32317 1852 32326
rect 1800 32283 1809 32317
rect 1809 32283 1843 32317
rect 1843 32283 1852 32317
rect 1800 32274 1852 32283
rect 1800 31981 1852 31990
rect 1800 31947 1809 31981
rect 1809 31947 1843 31981
rect 1843 31947 1852 31981
rect 1800 31938 1852 31947
rect 1800 31645 1852 31654
rect 1800 31611 1809 31645
rect 1809 31611 1843 31645
rect 1843 31611 1852 31645
rect 1800 31602 1852 31611
rect 15493 31493 15545 31545
rect 1800 31309 1852 31318
rect 1800 31275 1809 31309
rect 1809 31275 1843 31309
rect 1843 31275 1852 31309
rect 1800 31266 1852 31275
rect 1800 30973 1852 30982
rect 1800 30939 1809 30973
rect 1809 30939 1843 30973
rect 1843 30939 1852 30973
rect 1800 30930 1852 30939
rect 1800 30637 1852 30646
rect 1800 30603 1809 30637
rect 1809 30603 1843 30637
rect 1843 30603 1852 30637
rect 1800 30594 1852 30603
rect 1800 30301 1852 30310
rect 1800 30267 1809 30301
rect 1809 30267 1843 30301
rect 1843 30267 1852 30301
rect 1800 30258 1852 30267
rect 1800 29965 1852 29974
rect 1800 29931 1809 29965
rect 1809 29931 1843 29965
rect 1843 29931 1852 29965
rect 1800 29922 1852 29931
rect 15413 29935 15465 29987
rect 1800 29629 1852 29638
rect 1800 29595 1809 29629
rect 1809 29595 1843 29629
rect 1843 29595 1852 29629
rect 1800 29586 1852 29595
rect 1800 29293 1852 29302
rect 1800 29259 1809 29293
rect 1809 29259 1843 29293
rect 1843 29259 1852 29293
rect 1800 29250 1852 29259
rect 1800 28957 1852 28966
rect 1800 28923 1809 28957
rect 1809 28923 1843 28957
rect 1843 28923 1852 28957
rect 1800 28914 1852 28923
rect 1800 28621 1852 28630
rect 1800 28587 1809 28621
rect 1809 28587 1843 28621
rect 1843 28587 1852 28621
rect 1800 28578 1852 28587
rect 1800 28285 1852 28294
rect 1800 28251 1809 28285
rect 1809 28251 1843 28285
rect 1843 28251 1852 28285
rect 1800 28242 1852 28251
rect 1800 27949 1852 27958
rect 1800 27915 1809 27949
rect 1809 27915 1843 27949
rect 1843 27915 1852 27949
rect 1800 27906 1852 27915
rect 1800 27613 1852 27622
rect 1800 27579 1809 27613
rect 1809 27579 1843 27613
rect 1843 27579 1852 27613
rect 1800 27570 1852 27579
rect 1800 27277 1852 27286
rect 1800 27243 1809 27277
rect 1809 27243 1843 27277
rect 1843 27243 1852 27277
rect 1800 27234 1852 27243
rect 1800 26941 1852 26950
rect 1800 26907 1809 26941
rect 1809 26907 1843 26941
rect 1843 26907 1852 26941
rect 1800 26898 1852 26907
rect 1800 26605 1852 26614
rect 1800 26571 1809 26605
rect 1809 26571 1843 26605
rect 1843 26571 1852 26605
rect 1800 26562 1852 26571
rect 1800 26269 1852 26278
rect 1800 26235 1809 26269
rect 1809 26235 1843 26269
rect 1843 26235 1852 26269
rect 1800 26226 1852 26235
rect 1800 25933 1852 25942
rect 1800 25899 1809 25933
rect 1809 25899 1843 25933
rect 1843 25899 1852 25933
rect 1800 25890 1852 25899
rect 1800 25597 1852 25606
rect 1800 25563 1809 25597
rect 1809 25563 1843 25597
rect 1843 25563 1852 25597
rect 1800 25554 1852 25563
rect 1800 25261 1852 25270
rect 1800 25227 1809 25261
rect 1809 25227 1843 25261
rect 1843 25227 1852 25261
rect 1800 25218 1852 25227
rect 1800 24925 1852 24934
rect 1800 24891 1809 24925
rect 1809 24891 1843 24925
rect 1843 24891 1852 24925
rect 1800 24882 1852 24891
rect 1800 24589 1852 24598
rect 1800 24555 1809 24589
rect 1809 24555 1843 24589
rect 1843 24555 1852 24589
rect 1800 24546 1852 24555
rect 136946 39709 136998 39718
rect 136946 39675 136955 39709
rect 136955 39675 136989 39709
rect 136989 39675 136998 39709
rect 136946 39666 136998 39675
rect 136946 39373 136998 39382
rect 136946 39339 136955 39373
rect 136955 39339 136989 39373
rect 136989 39339 136998 39373
rect 136946 39330 136998 39339
rect 136946 39037 136998 39046
rect 136946 39003 136955 39037
rect 136955 39003 136989 39037
rect 136989 39003 136998 39037
rect 136946 38994 136998 39003
rect 136946 38701 136998 38710
rect 136946 38667 136955 38701
rect 136955 38667 136989 38701
rect 136989 38667 136998 38701
rect 136946 38658 136998 38667
rect 136946 38365 136998 38374
rect 136946 38331 136955 38365
rect 136955 38331 136989 38365
rect 136989 38331 136998 38365
rect 136946 38322 136998 38331
rect 136946 38029 136998 38038
rect 136946 37995 136955 38029
rect 136955 37995 136989 38029
rect 136989 37995 136998 38029
rect 136946 37986 136998 37995
rect 136946 37693 136998 37702
rect 136946 37659 136955 37693
rect 136955 37659 136989 37693
rect 136989 37659 136998 37693
rect 136946 37650 136998 37659
rect 136946 37357 136998 37366
rect 136946 37323 136955 37357
rect 136955 37323 136989 37357
rect 136989 37323 136998 37357
rect 136946 37314 136998 37323
rect 136946 37021 136998 37030
rect 136946 36987 136955 37021
rect 136955 36987 136989 37021
rect 136989 36987 136998 37021
rect 136946 36978 136998 36987
rect 136946 36685 136998 36694
rect 136946 36651 136955 36685
rect 136955 36651 136989 36685
rect 136989 36651 136998 36685
rect 136946 36642 136998 36651
rect 136946 36349 136998 36358
rect 136946 36315 136955 36349
rect 136955 36315 136989 36349
rect 136989 36315 136998 36349
rect 136946 36306 136998 36315
rect 136946 36013 136998 36022
rect 136946 35979 136955 36013
rect 136955 35979 136989 36013
rect 136989 35979 136998 36013
rect 136946 35970 136998 35979
rect 136946 35677 136998 35686
rect 136946 35643 136955 35677
rect 136955 35643 136989 35677
rect 136989 35643 136998 35677
rect 136946 35634 136998 35643
rect 136946 35341 136998 35350
rect 136946 35307 136955 35341
rect 136955 35307 136989 35341
rect 136989 35307 136998 35341
rect 136946 35298 136998 35307
rect 136946 35005 136998 35014
rect 136946 34971 136955 35005
rect 136955 34971 136989 35005
rect 136989 34971 136998 35005
rect 136946 34962 136998 34971
rect 136946 34669 136998 34678
rect 136946 34635 136955 34669
rect 136955 34635 136989 34669
rect 136989 34635 136998 34669
rect 136946 34626 136998 34635
rect 136946 34333 136998 34342
rect 136946 34299 136955 34333
rect 136955 34299 136989 34333
rect 136989 34299 136998 34333
rect 136946 34290 136998 34299
rect 136946 33997 136998 34006
rect 136946 33963 136955 33997
rect 136955 33963 136989 33997
rect 136989 33963 136998 33997
rect 136946 33954 136998 33963
rect 136946 33661 136998 33670
rect 136946 33627 136955 33661
rect 136955 33627 136989 33661
rect 136989 33627 136998 33661
rect 136946 33618 136998 33627
rect 136946 33325 136998 33334
rect 136946 33291 136955 33325
rect 136955 33291 136989 33325
rect 136989 33291 136998 33325
rect 136946 33282 136998 33291
rect 136946 32989 136998 32998
rect 136946 32955 136955 32989
rect 136955 32955 136989 32989
rect 136989 32955 136998 32989
rect 136946 32946 136998 32955
rect 136946 32653 136998 32662
rect 136946 32619 136955 32653
rect 136955 32619 136989 32653
rect 136989 32619 136998 32653
rect 136946 32610 136998 32619
rect 136946 32317 136998 32326
rect 136946 32283 136955 32317
rect 136955 32283 136989 32317
rect 136989 32283 136998 32317
rect 136946 32274 136998 32283
rect 136946 31981 136998 31990
rect 136946 31947 136955 31981
rect 136955 31947 136989 31981
rect 136989 31947 136998 31981
rect 136946 31938 136998 31947
rect 136946 31645 136998 31654
rect 136946 31611 136955 31645
rect 136955 31611 136989 31645
rect 136989 31611 136998 31645
rect 136946 31602 136998 31611
rect 136946 31309 136998 31318
rect 136946 31275 136955 31309
rect 136955 31275 136989 31309
rect 136989 31275 136998 31309
rect 136946 31266 136998 31275
rect 136946 30973 136998 30982
rect 136946 30939 136955 30973
rect 136955 30939 136989 30973
rect 136989 30939 136998 30973
rect 136946 30930 136998 30939
rect 136946 30637 136998 30646
rect 136946 30603 136955 30637
rect 136955 30603 136989 30637
rect 136989 30603 136998 30637
rect 136946 30594 136998 30603
rect 136946 30301 136998 30310
rect 136946 30267 136955 30301
rect 136955 30267 136989 30301
rect 136989 30267 136998 30301
rect 136946 30258 136998 30267
rect 136946 29965 136998 29974
rect 136946 29931 136955 29965
rect 136955 29931 136989 29965
rect 136989 29931 136998 29965
rect 136946 29922 136998 29931
rect 136946 29629 136998 29638
rect 136946 29595 136955 29629
rect 136955 29595 136989 29629
rect 136989 29595 136998 29629
rect 136946 29586 136998 29595
rect 136946 29293 136998 29302
rect 136946 29259 136955 29293
rect 136955 29259 136989 29293
rect 136989 29259 136998 29293
rect 136946 29250 136998 29259
rect 136946 28957 136998 28966
rect 136946 28923 136955 28957
rect 136955 28923 136989 28957
rect 136989 28923 136998 28957
rect 136946 28914 136998 28923
rect 136946 28621 136998 28630
rect 136946 28587 136955 28621
rect 136955 28587 136989 28621
rect 136989 28587 136998 28621
rect 136946 28578 136998 28587
rect 136946 28285 136998 28294
rect 136946 28251 136955 28285
rect 136955 28251 136989 28285
rect 136989 28251 136998 28285
rect 136946 28242 136998 28251
rect 136946 27949 136998 27958
rect 136946 27915 136955 27949
rect 136955 27915 136989 27949
rect 136989 27915 136998 27949
rect 136946 27906 136998 27915
rect 136946 27613 136998 27622
rect 136946 27579 136955 27613
rect 136955 27579 136989 27613
rect 136989 27579 136998 27613
rect 136946 27570 136998 27579
rect 136946 27277 136998 27286
rect 136946 27243 136955 27277
rect 136955 27243 136989 27277
rect 136989 27243 136998 27277
rect 136946 27234 136998 27243
rect 136946 26941 136998 26950
rect 136946 26907 136955 26941
rect 136955 26907 136989 26941
rect 136989 26907 136998 26941
rect 136946 26898 136998 26907
rect 136946 26605 136998 26614
rect 136946 26571 136955 26605
rect 136955 26571 136989 26605
rect 136989 26571 136998 26605
rect 136946 26562 136998 26571
rect 136946 26269 136998 26278
rect 136946 26235 136955 26269
rect 136955 26235 136989 26269
rect 136989 26235 136998 26269
rect 136946 26226 136998 26235
rect 136946 25933 136998 25942
rect 136946 25899 136955 25933
rect 136955 25899 136989 25933
rect 136989 25899 136998 25933
rect 136946 25890 136998 25899
rect 136946 25597 136998 25606
rect 136946 25563 136955 25597
rect 136955 25563 136989 25597
rect 136989 25563 136998 25597
rect 136946 25554 136998 25563
rect 136946 25261 136998 25270
rect 136946 25227 136955 25261
rect 136955 25227 136989 25261
rect 136989 25227 136998 25261
rect 136946 25218 136998 25227
rect 136946 24925 136998 24934
rect 136946 24891 136955 24925
rect 136955 24891 136989 24925
rect 136989 24891 136998 24925
rect 136946 24882 136998 24891
rect 1800 24253 1852 24262
rect 1800 24219 1809 24253
rect 1809 24219 1843 24253
rect 1843 24219 1852 24253
rect 1800 24210 1852 24219
rect 1800 23917 1852 23926
rect 1800 23883 1809 23917
rect 1809 23883 1843 23917
rect 1843 23883 1852 23917
rect 1800 23874 1852 23883
rect 1800 23581 1852 23590
rect 1800 23547 1809 23581
rect 1809 23547 1843 23581
rect 1843 23547 1852 23581
rect 1800 23538 1852 23547
rect 1800 23245 1852 23254
rect 1800 23211 1809 23245
rect 1809 23211 1843 23245
rect 1843 23211 1852 23245
rect 1800 23202 1852 23211
rect 1800 22909 1852 22918
rect 1800 22875 1809 22909
rect 1809 22875 1843 22909
rect 1843 22875 1852 22909
rect 1800 22866 1852 22875
rect 1800 22573 1852 22582
rect 1800 22539 1809 22573
rect 1809 22539 1843 22573
rect 1843 22539 1852 22573
rect 1800 22530 1852 22539
rect 1800 22237 1852 22246
rect 1800 22203 1809 22237
rect 1809 22203 1843 22237
rect 1843 22203 1852 22237
rect 1800 22194 1852 22203
rect 1800 21901 1852 21910
rect 1800 21867 1809 21901
rect 1809 21867 1843 21901
rect 1843 21867 1852 21901
rect 1800 21858 1852 21867
rect 1800 21565 1852 21574
rect 1800 21531 1809 21565
rect 1809 21531 1843 21565
rect 1843 21531 1852 21565
rect 1800 21522 1852 21531
rect 1800 21229 1852 21238
rect 1800 21195 1809 21229
rect 1809 21195 1843 21229
rect 1843 21195 1852 21229
rect 1800 21186 1852 21195
rect 1800 20893 1852 20902
rect 1800 20859 1809 20893
rect 1809 20859 1843 20893
rect 1843 20859 1852 20893
rect 1800 20850 1852 20859
rect 1800 20557 1852 20566
rect 1800 20523 1809 20557
rect 1809 20523 1843 20557
rect 1843 20523 1852 20557
rect 1800 20514 1852 20523
rect 1800 20221 1852 20230
rect 1800 20187 1809 20221
rect 1809 20187 1843 20221
rect 1843 20187 1852 20221
rect 1800 20178 1852 20187
rect 1800 19885 1852 19894
rect 1800 19851 1809 19885
rect 1809 19851 1843 19885
rect 1843 19851 1852 19885
rect 1800 19842 1852 19851
rect 1800 19549 1852 19558
rect 1800 19515 1809 19549
rect 1809 19515 1843 19549
rect 1843 19515 1852 19549
rect 1800 19506 1852 19515
rect 1800 19213 1852 19222
rect 1800 19179 1809 19213
rect 1809 19179 1843 19213
rect 1843 19179 1852 19213
rect 1800 19170 1852 19179
rect 1800 18877 1852 18886
rect 1800 18843 1809 18877
rect 1809 18843 1843 18877
rect 1843 18843 1852 18877
rect 1800 18834 1852 18843
rect 1800 18541 1852 18550
rect 1800 18507 1809 18541
rect 1809 18507 1843 18541
rect 1843 18507 1852 18541
rect 1800 18498 1852 18507
rect 1800 18205 1852 18214
rect 1800 18171 1809 18205
rect 1809 18171 1843 18205
rect 1843 18171 1852 18205
rect 1800 18162 1852 18171
rect 1800 17869 1852 17878
rect 1800 17835 1809 17869
rect 1809 17835 1843 17869
rect 1843 17835 1852 17869
rect 1800 17826 1852 17835
rect 1800 17533 1852 17542
rect 1800 17499 1809 17533
rect 1809 17499 1843 17533
rect 1843 17499 1852 17533
rect 1800 17490 1852 17499
rect 1800 17197 1852 17206
rect 1800 17163 1809 17197
rect 1809 17163 1843 17197
rect 1843 17163 1852 17197
rect 1800 17154 1852 17163
rect 1800 16861 1852 16870
rect 1800 16827 1809 16861
rect 1809 16827 1843 16861
rect 1843 16827 1852 16861
rect 1800 16818 1852 16827
rect 1800 16525 1852 16534
rect 1800 16491 1809 16525
rect 1809 16491 1843 16525
rect 1843 16491 1852 16525
rect 1800 16482 1852 16491
rect 1800 16189 1852 16198
rect 1800 16155 1809 16189
rect 1809 16155 1843 16189
rect 1843 16155 1852 16189
rect 1800 16146 1852 16155
rect 1800 15853 1852 15862
rect 1800 15819 1809 15853
rect 1809 15819 1843 15853
rect 1843 15819 1852 15853
rect 1800 15810 1852 15819
rect 1800 15517 1852 15526
rect 1800 15483 1809 15517
rect 1809 15483 1843 15517
rect 1843 15483 1852 15517
rect 1800 15474 1852 15483
rect 1800 15181 1852 15190
rect 1800 15147 1809 15181
rect 1809 15147 1843 15181
rect 1843 15147 1852 15181
rect 1800 15138 1852 15147
rect 1800 14845 1852 14854
rect 1800 14811 1809 14845
rect 1809 14811 1843 14845
rect 1843 14811 1852 14845
rect 1800 14802 1852 14811
rect 1800 14509 1852 14518
rect 1800 14475 1809 14509
rect 1809 14475 1843 14509
rect 1843 14475 1852 14509
rect 1800 14466 1852 14475
rect 1800 14173 1852 14182
rect 1800 14139 1809 14173
rect 1809 14139 1843 14173
rect 1843 14139 1852 14173
rect 1800 14130 1852 14139
rect 1800 13837 1852 13846
rect 1800 13803 1809 13837
rect 1809 13803 1843 13837
rect 1843 13803 1852 13837
rect 1800 13794 1852 13803
rect 1800 13501 1852 13510
rect 1800 13467 1809 13501
rect 1809 13467 1843 13501
rect 1843 13467 1852 13501
rect 1800 13458 1852 13467
rect 29564 13207 29616 13259
rect 32060 13207 32112 13259
rect 34556 13207 34608 13259
rect 37052 13207 37104 13259
rect 39548 13207 39600 13259
rect 42044 13207 42096 13259
rect 44540 13207 44592 13259
rect 47036 13207 47088 13259
rect 49532 13207 49584 13259
rect 52028 13207 52080 13259
rect 54524 13207 54576 13259
rect 57020 13207 57072 13259
rect 59516 13207 59568 13259
rect 62012 13207 62064 13259
rect 64508 13207 64560 13259
rect 67004 13207 67056 13259
rect 69500 13207 69552 13259
rect 71996 13207 72048 13259
rect 74492 13207 74544 13259
rect 76988 13207 77040 13259
rect 79484 13207 79536 13259
rect 81980 13207 82032 13259
rect 84476 13207 84528 13259
rect 86972 13207 87024 13259
rect 89468 13207 89520 13259
rect 91964 13207 92016 13259
rect 94460 13207 94512 13259
rect 96956 13207 97008 13259
rect 99452 13207 99504 13259
rect 101948 13207 102000 13259
rect 104444 13207 104496 13259
rect 106940 13207 106992 13259
rect 1800 13165 1852 13174
rect 1800 13131 1809 13165
rect 1809 13131 1843 13165
rect 1843 13131 1852 13165
rect 1800 13122 1852 13131
rect 1800 12829 1852 12838
rect 1800 12795 1809 12829
rect 1809 12795 1843 12829
rect 1843 12795 1852 12829
rect 1800 12786 1852 12795
rect 1800 12493 1852 12502
rect 1800 12459 1809 12493
rect 1809 12459 1843 12493
rect 1843 12459 1852 12493
rect 1800 12450 1852 12459
rect 1800 12157 1852 12166
rect 1800 12123 1809 12157
rect 1809 12123 1843 12157
rect 1843 12123 1852 12157
rect 1800 12114 1852 12123
rect 1800 11821 1852 11830
rect 1800 11787 1809 11821
rect 1809 11787 1843 11821
rect 1843 11787 1852 11821
rect 1800 11778 1852 11787
rect 1800 11485 1852 11494
rect 1800 11451 1809 11485
rect 1809 11451 1843 11485
rect 1843 11451 1852 11485
rect 1800 11442 1852 11451
rect 1800 11149 1852 11158
rect 1800 11115 1809 11149
rect 1809 11115 1843 11149
rect 1843 11115 1852 11149
rect 1800 11106 1852 11115
rect 1800 10813 1852 10822
rect 1800 10779 1809 10813
rect 1809 10779 1843 10813
rect 1843 10779 1852 10813
rect 1800 10770 1852 10779
rect 1800 10477 1852 10486
rect 1800 10443 1809 10477
rect 1809 10443 1843 10477
rect 1843 10443 1852 10477
rect 1800 10434 1852 10443
rect 1800 10141 1852 10150
rect 1800 10107 1809 10141
rect 1809 10107 1843 10141
rect 1843 10107 1852 10141
rect 1800 10098 1852 10107
rect 1800 9805 1852 9814
rect 1800 9771 1809 9805
rect 1809 9771 1843 9805
rect 1843 9771 1852 9805
rect 1800 9762 1852 9771
rect 1800 9469 1852 9478
rect 1800 9435 1809 9469
rect 1809 9435 1843 9469
rect 1843 9435 1852 9469
rect 1800 9426 1852 9435
rect 136946 24589 136998 24598
rect 136946 24555 136955 24589
rect 136955 24555 136989 24589
rect 136989 24555 136998 24589
rect 136946 24546 136998 24555
rect 136946 24253 136998 24262
rect 136946 24219 136955 24253
rect 136955 24219 136989 24253
rect 136989 24219 136998 24253
rect 136946 24210 136998 24219
rect 136946 23917 136998 23926
rect 136946 23883 136955 23917
rect 136955 23883 136989 23917
rect 136989 23883 136998 23917
rect 136946 23874 136998 23883
rect 136946 23581 136998 23590
rect 136946 23547 136955 23581
rect 136955 23547 136989 23581
rect 136989 23547 136998 23581
rect 136946 23538 136998 23547
rect 136946 23245 136998 23254
rect 136946 23211 136955 23245
rect 136955 23211 136989 23245
rect 136989 23211 136998 23245
rect 136946 23202 136998 23211
rect 136946 22909 136998 22918
rect 136946 22875 136955 22909
rect 136955 22875 136989 22909
rect 136989 22875 136998 22909
rect 136946 22866 136998 22875
rect 136946 22573 136998 22582
rect 136946 22539 136955 22573
rect 136955 22539 136989 22573
rect 136989 22539 136998 22573
rect 136946 22530 136998 22539
rect 136946 22237 136998 22246
rect 136946 22203 136955 22237
rect 136955 22203 136989 22237
rect 136989 22203 136998 22237
rect 136946 22194 136998 22203
rect 136946 21901 136998 21910
rect 136946 21867 136955 21901
rect 136955 21867 136989 21901
rect 136989 21867 136998 21901
rect 136946 21858 136998 21867
rect 136946 21565 136998 21574
rect 136946 21531 136955 21565
rect 136955 21531 136989 21565
rect 136989 21531 136998 21565
rect 136946 21522 136998 21531
rect 136946 21229 136998 21238
rect 136946 21195 136955 21229
rect 136955 21195 136989 21229
rect 136989 21195 136998 21229
rect 136946 21186 136998 21195
rect 136946 20893 136998 20902
rect 136946 20859 136955 20893
rect 136955 20859 136989 20893
rect 136989 20859 136998 20893
rect 136946 20850 136998 20859
rect 136946 20557 136998 20566
rect 136946 20523 136955 20557
rect 136955 20523 136989 20557
rect 136989 20523 136998 20557
rect 136946 20514 136998 20523
rect 136946 20221 136998 20230
rect 136946 20187 136955 20221
rect 136955 20187 136989 20221
rect 136989 20187 136998 20221
rect 136946 20178 136998 20187
rect 136946 19885 136998 19894
rect 136946 19851 136955 19885
rect 136955 19851 136989 19885
rect 136989 19851 136998 19885
rect 136946 19842 136998 19851
rect 136946 19549 136998 19558
rect 136946 19515 136955 19549
rect 136955 19515 136989 19549
rect 136989 19515 136998 19549
rect 136946 19506 136998 19515
rect 123333 19185 123385 19237
rect 136946 19213 136998 19222
rect 136946 19179 136955 19213
rect 136955 19179 136989 19213
rect 136989 19179 136998 19213
rect 136946 19170 136998 19179
rect 136946 18877 136998 18886
rect 136946 18843 136955 18877
rect 136955 18843 136989 18877
rect 136989 18843 136998 18877
rect 136946 18834 136998 18843
rect 136946 18541 136998 18550
rect 136946 18507 136955 18541
rect 136955 18507 136989 18541
rect 136989 18507 136998 18541
rect 136946 18498 136998 18507
rect 136946 18205 136998 18214
rect 136946 18171 136955 18205
rect 136955 18171 136989 18205
rect 136989 18171 136998 18205
rect 136946 18162 136998 18171
rect 136946 17869 136998 17878
rect 136946 17835 136955 17869
rect 136955 17835 136989 17869
rect 136989 17835 136998 17869
rect 136946 17826 136998 17835
rect 123253 17627 123305 17679
rect 136946 17533 136998 17542
rect 136946 17499 136955 17533
rect 136955 17499 136989 17533
rect 136989 17499 136998 17533
rect 136946 17490 136998 17499
rect 136946 17197 136998 17206
rect 136946 17163 136955 17197
rect 136955 17163 136989 17197
rect 136989 17163 136998 17197
rect 136946 17154 136998 17163
rect 136946 16861 136998 16870
rect 136946 16827 136955 16861
rect 136955 16827 136989 16861
rect 136989 16827 136998 16861
rect 136946 16818 136998 16827
rect 136946 16525 136998 16534
rect 136946 16491 136955 16525
rect 136955 16491 136989 16525
rect 136989 16491 136998 16525
rect 136946 16482 136998 16491
rect 123173 16357 123225 16409
rect 136946 16189 136998 16198
rect 136946 16155 136955 16189
rect 136955 16155 136989 16189
rect 136989 16155 136998 16189
rect 136946 16146 136998 16155
rect 136946 15853 136998 15862
rect 136946 15819 136955 15853
rect 136955 15819 136989 15853
rect 136989 15819 136998 15853
rect 136946 15810 136998 15819
rect 136946 15517 136998 15526
rect 136946 15483 136955 15517
rect 136955 15483 136989 15517
rect 136989 15483 136998 15517
rect 136946 15474 136998 15483
rect 136946 15181 136998 15190
rect 136946 15147 136955 15181
rect 136955 15147 136989 15181
rect 136989 15147 136998 15181
rect 136946 15138 136998 15147
rect 123093 14799 123145 14851
rect 136946 14845 136998 14854
rect 136946 14811 136955 14845
rect 136955 14811 136989 14845
rect 136989 14811 136998 14845
rect 136946 14802 136998 14811
rect 136946 14509 136998 14518
rect 136946 14475 136955 14509
rect 136955 14475 136989 14509
rect 136989 14475 136998 14509
rect 136946 14466 136998 14475
rect 136946 14173 136998 14182
rect 136946 14139 136955 14173
rect 136955 14139 136989 14173
rect 136989 14139 136998 14173
rect 136946 14130 136998 14139
rect 136946 13837 136998 13846
rect 136946 13803 136955 13837
rect 136955 13803 136989 13837
rect 136989 13803 136998 13837
rect 136946 13794 136998 13803
rect 123013 13529 123065 13581
rect 136946 13501 136998 13510
rect 136946 13467 136955 13501
rect 136955 13467 136989 13501
rect 136989 13467 136998 13501
rect 136946 13458 136998 13467
rect 136946 13165 136998 13174
rect 136946 13131 136955 13165
rect 136955 13131 136989 13165
rect 136989 13131 136998 13165
rect 136946 13122 136998 13131
rect 136946 12829 136998 12838
rect 136946 12795 136955 12829
rect 136955 12795 136989 12829
rect 136989 12795 136998 12829
rect 136946 12786 136998 12795
rect 136946 12493 136998 12502
rect 136946 12459 136955 12493
rect 136955 12459 136989 12493
rect 136989 12459 136998 12493
rect 136946 12450 136998 12459
rect 136946 12157 136998 12166
rect 136946 12123 136955 12157
rect 136955 12123 136989 12157
rect 136989 12123 136998 12157
rect 136946 12114 136998 12123
rect 122933 11971 122985 12023
rect 136946 11821 136998 11830
rect 136946 11787 136955 11821
rect 136955 11787 136989 11821
rect 136989 11787 136998 11821
rect 136946 11778 136998 11787
rect 136946 11485 136998 11494
rect 136946 11451 136955 11485
rect 136955 11451 136989 11485
rect 136989 11451 136998 11485
rect 136946 11442 136998 11451
rect 136946 11149 136998 11158
rect 136946 11115 136955 11149
rect 136955 11115 136989 11149
rect 136989 11115 136998 11149
rect 136946 11106 136998 11115
rect 136946 10813 136998 10822
rect 136946 10779 136955 10813
rect 136955 10779 136989 10813
rect 136989 10779 136998 10813
rect 136946 10770 136998 10779
rect 122853 10701 122905 10753
rect 136946 10477 136998 10486
rect 136946 10443 136955 10477
rect 136955 10443 136989 10477
rect 136989 10443 136998 10477
rect 136946 10434 136998 10443
rect 136946 10141 136998 10150
rect 136946 10107 136955 10141
rect 136955 10107 136989 10141
rect 136989 10107 136998 10141
rect 136946 10098 136998 10107
rect 136946 9805 136998 9814
rect 136946 9771 136955 9805
rect 136955 9771 136989 9805
rect 136989 9771 136998 9805
rect 136946 9762 136998 9771
rect 136946 9469 136998 9478
rect 136946 9435 136955 9469
rect 136955 9435 136989 9469
rect 136989 9435 136998 9469
rect 136946 9426 136998 9435
rect 122773 9143 122825 9195
rect 1800 9133 1852 9142
rect 1800 9099 1809 9133
rect 1809 9099 1843 9133
rect 1843 9099 1852 9133
rect 1800 9090 1852 9099
rect 136946 9133 136998 9142
rect 136946 9099 136955 9133
rect 136955 9099 136989 9133
rect 136989 9099 136998 9133
rect 136946 9090 136998 9099
rect 1800 8797 1852 8806
rect 1800 8763 1809 8797
rect 1809 8763 1843 8797
rect 1843 8763 1852 8797
rect 1800 8754 1852 8763
rect 136946 8797 136998 8806
rect 136946 8763 136955 8797
rect 136955 8763 136989 8797
rect 136989 8763 136998 8797
rect 136946 8754 136998 8763
rect 1800 8461 1852 8470
rect 1800 8427 1809 8461
rect 1809 8427 1843 8461
rect 1843 8427 1852 8461
rect 1800 8418 1852 8427
rect 136946 8461 136998 8470
rect 136946 8427 136955 8461
rect 136955 8427 136989 8461
rect 136989 8427 136998 8461
rect 136946 8418 136998 8427
rect 1800 8125 1852 8134
rect 1800 8091 1809 8125
rect 1809 8091 1843 8125
rect 1843 8091 1852 8125
rect 1800 8082 1852 8091
rect 136946 8125 136998 8134
rect 136946 8091 136955 8125
rect 136955 8091 136989 8125
rect 136989 8091 136998 8125
rect 136946 8082 136998 8091
rect 1800 7789 1852 7798
rect 1800 7755 1809 7789
rect 1809 7755 1843 7789
rect 1843 7755 1852 7789
rect 1800 7746 1852 7755
rect 136946 7789 136998 7798
rect 136946 7755 136955 7789
rect 136955 7755 136989 7789
rect 136989 7755 136998 7789
rect 136946 7746 136998 7755
rect 1800 7453 1852 7462
rect 1800 7419 1809 7453
rect 1809 7419 1843 7453
rect 1843 7419 1852 7453
rect 1800 7410 1852 7419
rect 136946 7453 136998 7462
rect 136946 7419 136955 7453
rect 136955 7419 136989 7453
rect 136989 7419 136998 7453
rect 136946 7410 136998 7419
rect 1800 7117 1852 7126
rect 1800 7083 1809 7117
rect 1809 7083 1843 7117
rect 1843 7083 1852 7117
rect 1800 7074 1852 7083
rect 136946 7117 136998 7126
rect 136946 7083 136955 7117
rect 136955 7083 136989 7117
rect 136989 7083 136998 7117
rect 136946 7074 136998 7083
rect 1800 6781 1852 6790
rect 1800 6747 1809 6781
rect 1809 6747 1843 6781
rect 1843 6747 1852 6781
rect 1800 6738 1852 6747
rect 136946 6781 136998 6790
rect 136946 6747 136955 6781
rect 136955 6747 136989 6781
rect 136989 6747 136998 6781
rect 136946 6738 136998 6747
rect 1800 6445 1852 6454
rect 1800 6411 1809 6445
rect 1809 6411 1843 6445
rect 1843 6411 1852 6445
rect 1800 6402 1852 6411
rect 136946 6445 136998 6454
rect 136946 6411 136955 6445
rect 136955 6411 136989 6445
rect 136989 6411 136998 6445
rect 136946 6402 136998 6411
rect 1800 6109 1852 6118
rect 1800 6075 1809 6109
rect 1809 6075 1843 6109
rect 1843 6075 1852 6109
rect 1800 6066 1852 6075
rect 136946 6109 136998 6118
rect 136946 6075 136955 6109
rect 136955 6075 136989 6109
rect 136989 6075 136998 6109
rect 136946 6066 136998 6075
rect 1800 5773 1852 5782
rect 1800 5739 1809 5773
rect 1809 5739 1843 5773
rect 1843 5739 1852 5773
rect 1800 5730 1852 5739
rect 136946 5773 136998 5782
rect 136946 5739 136955 5773
rect 136955 5739 136989 5773
rect 136989 5739 136998 5773
rect 136946 5730 136998 5739
rect 1800 5437 1852 5446
rect 1800 5403 1809 5437
rect 1809 5403 1843 5437
rect 1843 5403 1852 5437
rect 1800 5394 1852 5403
rect 136946 5437 136998 5446
rect 136946 5403 136955 5437
rect 136955 5403 136989 5437
rect 136989 5403 136998 5437
rect 136946 5394 136998 5403
rect 1800 5101 1852 5110
rect 1800 5067 1809 5101
rect 1809 5067 1843 5101
rect 1843 5067 1852 5101
rect 1800 5058 1852 5067
rect 136946 5101 136998 5110
rect 136946 5067 136955 5101
rect 136955 5067 136989 5101
rect 136989 5067 136998 5101
rect 136946 5058 136998 5067
rect 1800 4765 1852 4774
rect 1800 4731 1809 4765
rect 1809 4731 1843 4765
rect 1843 4731 1852 4765
rect 1800 4722 1852 4731
rect 136946 4765 136998 4774
rect 136946 4731 136955 4765
rect 136955 4731 136989 4765
rect 136989 4731 136998 4765
rect 136946 4722 136998 4731
rect 1800 4429 1852 4438
rect 1800 4395 1809 4429
rect 1809 4395 1843 4429
rect 1843 4395 1852 4429
rect 1800 4386 1852 4395
rect 136946 4429 136998 4438
rect 136946 4395 136955 4429
rect 136955 4395 136989 4429
rect 136989 4395 136998 4429
rect 136946 4386 136998 4395
rect 1800 4093 1852 4102
rect 1800 4059 1809 4093
rect 1809 4059 1843 4093
rect 1843 4059 1852 4093
rect 1800 4050 1852 4059
rect 136946 4093 136998 4102
rect 136946 4059 136955 4093
rect 136955 4059 136989 4093
rect 136989 4059 136998 4093
rect 136946 4050 136998 4059
rect 1800 3757 1852 3766
rect 1800 3723 1809 3757
rect 1809 3723 1843 3757
rect 1843 3723 1852 3757
rect 1800 3714 1852 3723
rect 136946 3757 136998 3766
rect 136946 3723 136955 3757
rect 136955 3723 136989 3757
rect 136989 3723 136998 3757
rect 136946 3714 136998 3723
rect 1800 3421 1852 3430
rect 1800 3387 1809 3421
rect 1809 3387 1843 3421
rect 1843 3387 1852 3421
rect 1800 3378 1852 3387
rect 136946 3421 136998 3430
rect 136946 3387 136955 3421
rect 136955 3387 136989 3421
rect 136989 3387 136998 3421
rect 136946 3378 136998 3387
rect 1800 3085 1852 3094
rect 1800 3051 1809 3085
rect 1809 3051 1843 3085
rect 1843 3051 1852 3085
rect 1800 3042 1852 3051
rect 136946 3085 136998 3094
rect 136946 3051 136955 3085
rect 136955 3051 136989 3085
rect 136989 3051 136998 3085
rect 136946 3042 136998 3051
rect 1800 2749 1852 2758
rect 1800 2715 1809 2749
rect 1809 2715 1843 2749
rect 1843 2715 1852 2749
rect 1800 2706 1852 2715
rect 136946 2749 136998 2758
rect 136946 2715 136955 2749
rect 136955 2715 136989 2749
rect 136989 2715 136998 2749
rect 136946 2706 136998 2715
rect 1800 2413 1852 2422
rect 1800 2379 1809 2413
rect 1809 2379 1843 2413
rect 1843 2379 1852 2413
rect 1800 2370 1852 2379
rect 136946 2413 136998 2422
rect 136946 2379 136955 2413
rect 136955 2379 136989 2413
rect 136989 2379 136998 2413
rect 136946 2370 136998 2379
rect 1800 2077 1852 2086
rect 1800 2043 1809 2077
rect 1809 2043 1843 2077
rect 1843 2043 1852 2077
rect 1800 2034 1852 2043
rect 136946 2077 136998 2086
rect 136946 2043 136955 2077
rect 136955 2043 136989 2077
rect 136989 2043 136998 2077
rect 136946 2034 136998 2043
rect 2136 1741 2188 1750
rect 3816 1741 3868 1750
rect 5496 1741 5548 1750
rect 7176 1741 7228 1750
rect 8856 1741 8908 1750
rect 10536 1741 10588 1750
rect 12216 1741 12268 1750
rect 13896 1741 13948 1750
rect 15576 1741 15628 1750
rect 17256 1741 17308 1750
rect 18936 1741 18988 1750
rect 20616 1741 20668 1750
rect 22296 1741 22348 1750
rect 23976 1741 24028 1750
rect 25656 1741 25708 1750
rect 27336 1741 27388 1750
rect 29016 1741 29068 1750
rect 30696 1741 30748 1750
rect 32376 1741 32428 1750
rect 34056 1741 34108 1750
rect 35736 1741 35788 1750
rect 37416 1741 37468 1750
rect 39096 1741 39148 1750
rect 40776 1741 40828 1750
rect 42456 1741 42508 1750
rect 44136 1741 44188 1750
rect 45816 1741 45868 1750
rect 47496 1741 47548 1750
rect 49176 1741 49228 1750
rect 50856 1741 50908 1750
rect 52536 1741 52588 1750
rect 54216 1741 54268 1750
rect 55896 1741 55948 1750
rect 57576 1741 57628 1750
rect 59256 1741 59308 1750
rect 60936 1741 60988 1750
rect 62616 1741 62668 1750
rect 64296 1741 64348 1750
rect 65976 1741 66028 1750
rect 67656 1741 67708 1750
rect 69336 1741 69388 1750
rect 71016 1741 71068 1750
rect 72696 1741 72748 1750
rect 74376 1741 74428 1750
rect 76056 1741 76108 1750
rect 77736 1741 77788 1750
rect 79416 1741 79468 1750
rect 81096 1741 81148 1750
rect 82776 1741 82828 1750
rect 84456 1741 84508 1750
rect 86136 1741 86188 1750
rect 87816 1741 87868 1750
rect 89496 1741 89548 1750
rect 91176 1741 91228 1750
rect 92856 1741 92908 1750
rect 94536 1741 94588 1750
rect 96216 1741 96268 1750
rect 97896 1741 97948 1750
rect 99576 1741 99628 1750
rect 101256 1741 101308 1750
rect 102936 1741 102988 1750
rect 104616 1741 104668 1750
rect 106296 1741 106348 1750
rect 107976 1741 108028 1750
rect 109656 1741 109708 1750
rect 111336 1741 111388 1750
rect 113016 1741 113068 1750
rect 114696 1741 114748 1750
rect 116376 1741 116428 1750
rect 118056 1741 118108 1750
rect 119736 1741 119788 1750
rect 121416 1741 121468 1750
rect 123096 1741 123148 1750
rect 124776 1741 124828 1750
rect 126456 1741 126508 1750
rect 128136 1741 128188 1750
rect 129816 1741 129868 1750
rect 131496 1741 131548 1750
rect 133176 1741 133228 1750
rect 134856 1741 134908 1750
rect 136536 1741 136588 1750
rect 2136 1707 2145 1741
rect 2145 1707 2179 1741
rect 2179 1707 2188 1741
rect 3816 1707 3825 1741
rect 3825 1707 3859 1741
rect 3859 1707 3868 1741
rect 5496 1707 5505 1741
rect 5505 1707 5539 1741
rect 5539 1707 5548 1741
rect 7176 1707 7185 1741
rect 7185 1707 7219 1741
rect 7219 1707 7228 1741
rect 8856 1707 8865 1741
rect 8865 1707 8899 1741
rect 8899 1707 8908 1741
rect 10536 1707 10545 1741
rect 10545 1707 10579 1741
rect 10579 1707 10588 1741
rect 12216 1707 12225 1741
rect 12225 1707 12259 1741
rect 12259 1707 12268 1741
rect 13896 1707 13905 1741
rect 13905 1707 13939 1741
rect 13939 1707 13948 1741
rect 15576 1707 15585 1741
rect 15585 1707 15619 1741
rect 15619 1707 15628 1741
rect 17256 1707 17265 1741
rect 17265 1707 17299 1741
rect 17299 1707 17308 1741
rect 18936 1707 18945 1741
rect 18945 1707 18979 1741
rect 18979 1707 18988 1741
rect 20616 1707 20625 1741
rect 20625 1707 20659 1741
rect 20659 1707 20668 1741
rect 22296 1707 22305 1741
rect 22305 1707 22339 1741
rect 22339 1707 22348 1741
rect 23976 1707 23985 1741
rect 23985 1707 24019 1741
rect 24019 1707 24028 1741
rect 25656 1707 25665 1741
rect 25665 1707 25699 1741
rect 25699 1707 25708 1741
rect 27336 1707 27345 1741
rect 27345 1707 27379 1741
rect 27379 1707 27388 1741
rect 29016 1707 29025 1741
rect 29025 1707 29059 1741
rect 29059 1707 29068 1741
rect 30696 1707 30705 1741
rect 30705 1707 30739 1741
rect 30739 1707 30748 1741
rect 32376 1707 32385 1741
rect 32385 1707 32419 1741
rect 32419 1707 32428 1741
rect 34056 1707 34065 1741
rect 34065 1707 34099 1741
rect 34099 1707 34108 1741
rect 35736 1707 35745 1741
rect 35745 1707 35779 1741
rect 35779 1707 35788 1741
rect 37416 1707 37425 1741
rect 37425 1707 37459 1741
rect 37459 1707 37468 1741
rect 39096 1707 39105 1741
rect 39105 1707 39139 1741
rect 39139 1707 39148 1741
rect 40776 1707 40785 1741
rect 40785 1707 40819 1741
rect 40819 1707 40828 1741
rect 42456 1707 42465 1741
rect 42465 1707 42499 1741
rect 42499 1707 42508 1741
rect 44136 1707 44145 1741
rect 44145 1707 44179 1741
rect 44179 1707 44188 1741
rect 45816 1707 45825 1741
rect 45825 1707 45859 1741
rect 45859 1707 45868 1741
rect 47496 1707 47505 1741
rect 47505 1707 47539 1741
rect 47539 1707 47548 1741
rect 49176 1707 49185 1741
rect 49185 1707 49219 1741
rect 49219 1707 49228 1741
rect 50856 1707 50865 1741
rect 50865 1707 50899 1741
rect 50899 1707 50908 1741
rect 52536 1707 52545 1741
rect 52545 1707 52579 1741
rect 52579 1707 52588 1741
rect 54216 1707 54225 1741
rect 54225 1707 54259 1741
rect 54259 1707 54268 1741
rect 55896 1707 55905 1741
rect 55905 1707 55939 1741
rect 55939 1707 55948 1741
rect 57576 1707 57585 1741
rect 57585 1707 57619 1741
rect 57619 1707 57628 1741
rect 59256 1707 59265 1741
rect 59265 1707 59299 1741
rect 59299 1707 59308 1741
rect 60936 1707 60945 1741
rect 60945 1707 60979 1741
rect 60979 1707 60988 1741
rect 62616 1707 62625 1741
rect 62625 1707 62659 1741
rect 62659 1707 62668 1741
rect 64296 1707 64305 1741
rect 64305 1707 64339 1741
rect 64339 1707 64348 1741
rect 65976 1707 65985 1741
rect 65985 1707 66019 1741
rect 66019 1707 66028 1741
rect 67656 1707 67665 1741
rect 67665 1707 67699 1741
rect 67699 1707 67708 1741
rect 69336 1707 69345 1741
rect 69345 1707 69379 1741
rect 69379 1707 69388 1741
rect 71016 1707 71025 1741
rect 71025 1707 71059 1741
rect 71059 1707 71068 1741
rect 72696 1707 72705 1741
rect 72705 1707 72739 1741
rect 72739 1707 72748 1741
rect 74376 1707 74385 1741
rect 74385 1707 74419 1741
rect 74419 1707 74428 1741
rect 76056 1707 76065 1741
rect 76065 1707 76099 1741
rect 76099 1707 76108 1741
rect 77736 1707 77745 1741
rect 77745 1707 77779 1741
rect 77779 1707 77788 1741
rect 79416 1707 79425 1741
rect 79425 1707 79459 1741
rect 79459 1707 79468 1741
rect 81096 1707 81105 1741
rect 81105 1707 81139 1741
rect 81139 1707 81148 1741
rect 82776 1707 82785 1741
rect 82785 1707 82819 1741
rect 82819 1707 82828 1741
rect 84456 1707 84465 1741
rect 84465 1707 84499 1741
rect 84499 1707 84508 1741
rect 86136 1707 86145 1741
rect 86145 1707 86179 1741
rect 86179 1707 86188 1741
rect 87816 1707 87825 1741
rect 87825 1707 87859 1741
rect 87859 1707 87868 1741
rect 89496 1707 89505 1741
rect 89505 1707 89539 1741
rect 89539 1707 89548 1741
rect 91176 1707 91185 1741
rect 91185 1707 91219 1741
rect 91219 1707 91228 1741
rect 92856 1707 92865 1741
rect 92865 1707 92899 1741
rect 92899 1707 92908 1741
rect 94536 1707 94545 1741
rect 94545 1707 94579 1741
rect 94579 1707 94588 1741
rect 96216 1707 96225 1741
rect 96225 1707 96259 1741
rect 96259 1707 96268 1741
rect 97896 1707 97905 1741
rect 97905 1707 97939 1741
rect 97939 1707 97948 1741
rect 99576 1707 99585 1741
rect 99585 1707 99619 1741
rect 99619 1707 99628 1741
rect 101256 1707 101265 1741
rect 101265 1707 101299 1741
rect 101299 1707 101308 1741
rect 102936 1707 102945 1741
rect 102945 1707 102979 1741
rect 102979 1707 102988 1741
rect 104616 1707 104625 1741
rect 104625 1707 104659 1741
rect 104659 1707 104668 1741
rect 106296 1707 106305 1741
rect 106305 1707 106339 1741
rect 106339 1707 106348 1741
rect 107976 1707 107985 1741
rect 107985 1707 108019 1741
rect 108019 1707 108028 1741
rect 109656 1707 109665 1741
rect 109665 1707 109699 1741
rect 109699 1707 109708 1741
rect 111336 1707 111345 1741
rect 111345 1707 111379 1741
rect 111379 1707 111388 1741
rect 113016 1707 113025 1741
rect 113025 1707 113059 1741
rect 113059 1707 113068 1741
rect 114696 1707 114705 1741
rect 114705 1707 114739 1741
rect 114739 1707 114748 1741
rect 116376 1707 116385 1741
rect 116385 1707 116419 1741
rect 116419 1707 116428 1741
rect 118056 1707 118065 1741
rect 118065 1707 118099 1741
rect 118099 1707 118108 1741
rect 119736 1707 119745 1741
rect 119745 1707 119779 1741
rect 119779 1707 119788 1741
rect 121416 1707 121425 1741
rect 121425 1707 121459 1741
rect 121459 1707 121468 1741
rect 123096 1707 123105 1741
rect 123105 1707 123139 1741
rect 123139 1707 123148 1741
rect 124776 1707 124785 1741
rect 124785 1707 124819 1741
rect 124819 1707 124828 1741
rect 126456 1707 126465 1741
rect 126465 1707 126499 1741
rect 126499 1707 126508 1741
rect 128136 1707 128145 1741
rect 128145 1707 128179 1741
rect 128179 1707 128188 1741
rect 129816 1707 129825 1741
rect 129825 1707 129859 1741
rect 129859 1707 129868 1741
rect 131496 1707 131505 1741
rect 131505 1707 131539 1741
rect 131539 1707 131548 1741
rect 133176 1707 133185 1741
rect 133185 1707 133219 1741
rect 133219 1707 133228 1741
rect 134856 1707 134865 1741
rect 134865 1707 134899 1741
rect 134899 1707 134908 1741
rect 136536 1707 136545 1741
rect 136545 1707 136579 1741
rect 136579 1707 136588 1741
rect 2136 1698 2188 1707
rect 3816 1698 3868 1707
rect 5496 1698 5548 1707
rect 7176 1698 7228 1707
rect 8856 1698 8908 1707
rect 10536 1698 10588 1707
rect 12216 1698 12268 1707
rect 13896 1698 13948 1707
rect 15576 1698 15628 1707
rect 17256 1698 17308 1707
rect 18936 1698 18988 1707
rect 20616 1698 20668 1707
rect 22296 1698 22348 1707
rect 23976 1698 24028 1707
rect 25656 1698 25708 1707
rect 27336 1698 27388 1707
rect 29016 1698 29068 1707
rect 30696 1698 30748 1707
rect 32376 1698 32428 1707
rect 34056 1698 34108 1707
rect 35736 1698 35788 1707
rect 37416 1698 37468 1707
rect 39096 1698 39148 1707
rect 40776 1698 40828 1707
rect 42456 1698 42508 1707
rect 44136 1698 44188 1707
rect 45816 1698 45868 1707
rect 47496 1698 47548 1707
rect 49176 1698 49228 1707
rect 50856 1698 50908 1707
rect 52536 1698 52588 1707
rect 54216 1698 54268 1707
rect 55896 1698 55948 1707
rect 57576 1698 57628 1707
rect 59256 1698 59308 1707
rect 60936 1698 60988 1707
rect 62616 1698 62668 1707
rect 64296 1698 64348 1707
rect 65976 1698 66028 1707
rect 67656 1698 67708 1707
rect 69336 1698 69388 1707
rect 71016 1698 71068 1707
rect 72696 1698 72748 1707
rect 74376 1698 74428 1707
rect 76056 1698 76108 1707
rect 77736 1698 77788 1707
rect 79416 1698 79468 1707
rect 81096 1698 81148 1707
rect 82776 1698 82828 1707
rect 84456 1698 84508 1707
rect 86136 1698 86188 1707
rect 87816 1698 87868 1707
rect 89496 1698 89548 1707
rect 91176 1698 91228 1707
rect 92856 1698 92908 1707
rect 94536 1698 94588 1707
rect 96216 1698 96268 1707
rect 97896 1698 97948 1707
rect 99576 1698 99628 1707
rect 101256 1698 101308 1707
rect 102936 1698 102988 1707
rect 104616 1698 104668 1707
rect 106296 1698 106348 1707
rect 107976 1698 108028 1707
rect 109656 1698 109708 1707
rect 111336 1698 111388 1707
rect 113016 1698 113068 1707
rect 114696 1698 114748 1707
rect 116376 1698 116428 1707
rect 118056 1698 118108 1707
rect 119736 1698 119788 1707
rect 121416 1698 121468 1707
rect 123096 1698 123148 1707
rect 124776 1698 124828 1707
rect 126456 1698 126508 1707
rect 128136 1698 128188 1707
rect 129816 1698 129868 1707
rect 131496 1698 131548 1707
rect 133176 1698 133228 1707
rect 134856 1698 134908 1707
rect 136536 1698 136588 1707
<< metal2 >>
rect 1714 131448 1938 132145
rect 2134 132061 2190 132070
rect 2134 131996 2190 132005
rect 3814 132061 3870 132070
rect 3814 131996 3870 132005
rect 5494 132061 5550 132070
rect 5494 131996 5550 132005
rect 7174 132061 7230 132070
rect 7174 131996 7230 132005
rect 8854 132061 8910 132070
rect 8854 131996 8910 132005
rect 10534 132061 10590 132070
rect 10534 131996 10590 132005
rect 12214 132061 12270 132070
rect 12214 131996 12270 132005
rect 13894 132061 13950 132070
rect 13894 131996 13950 132005
rect 15574 132061 15630 132070
rect 15574 131996 15630 132005
rect 17254 132061 17310 132070
rect 17254 131996 17310 132005
rect 18934 132061 18990 132070
rect 18934 131996 18990 132005
rect 20614 132061 20670 132070
rect 20614 131996 20670 132005
rect 22294 132061 22350 132070
rect 22294 131996 22350 132005
rect 23974 132061 24030 132070
rect 23974 131996 24030 132005
rect 25654 132061 25710 132070
rect 25654 131996 25710 132005
rect 27334 132061 27390 132070
rect 27334 131996 27390 132005
rect 29014 132061 29070 132070
rect 29014 131996 29070 132005
rect 30694 132061 30750 132070
rect 30694 131996 30750 132005
rect 32374 132061 32430 132070
rect 32374 131996 32430 132005
rect 34054 132061 34110 132070
rect 34054 131996 34110 132005
rect 35734 132061 35790 132070
rect 35734 131996 35790 132005
rect 37414 132061 37470 132070
rect 37414 131996 37470 132005
rect 39094 132061 39150 132070
rect 39094 131996 39150 132005
rect 40774 132061 40830 132070
rect 40774 131996 40830 132005
rect 42454 132061 42510 132070
rect 42454 131996 42510 132005
rect 44134 132061 44190 132070
rect 44134 131996 44190 132005
rect 45814 132061 45870 132070
rect 45814 131996 45870 132005
rect 47494 132061 47550 132070
rect 47494 131996 47550 132005
rect 49174 132061 49230 132070
rect 49174 131996 49230 132005
rect 50854 132061 50910 132070
rect 50854 131996 50910 132005
rect 52534 132061 52590 132070
rect 52534 131996 52590 132005
rect 54214 132061 54270 132070
rect 54214 131996 54270 132005
rect 55894 132061 55950 132070
rect 55894 131996 55950 132005
rect 57574 132061 57630 132070
rect 57574 131996 57630 132005
rect 59254 132061 59310 132070
rect 59254 131996 59310 132005
rect 60934 132061 60990 132070
rect 60934 131996 60990 132005
rect 62614 132061 62670 132070
rect 62614 131996 62670 132005
rect 64294 132061 64350 132070
rect 64294 131996 64350 132005
rect 65974 132061 66030 132070
rect 65974 131996 66030 132005
rect 67654 132061 67710 132070
rect 67654 131996 67710 132005
rect 69334 132061 69390 132070
rect 69334 131996 69390 132005
rect 71014 132061 71070 132070
rect 71014 131996 71070 132005
rect 72694 132061 72750 132070
rect 72694 131996 72750 132005
rect 74374 132061 74430 132070
rect 74374 131996 74430 132005
rect 76054 132061 76110 132070
rect 76054 131996 76110 132005
rect 77734 132061 77790 132070
rect 77734 131996 77790 132005
rect 79414 132061 79470 132070
rect 79414 131996 79470 132005
rect 81094 132061 81150 132070
rect 81094 131996 81150 132005
rect 82774 132061 82830 132070
rect 82774 131996 82830 132005
rect 84454 132061 84510 132070
rect 84454 131996 84510 132005
rect 86134 132061 86190 132070
rect 86134 131996 86190 132005
rect 87814 132061 87870 132070
rect 87814 131996 87870 132005
rect 89494 132061 89550 132070
rect 89494 131996 89550 132005
rect 91174 132061 91230 132070
rect 91174 131996 91230 132005
rect 92854 132061 92910 132070
rect 92854 131996 92910 132005
rect 94534 132061 94590 132070
rect 94534 131996 94590 132005
rect 96214 132061 96270 132070
rect 96214 131996 96270 132005
rect 97894 132061 97950 132070
rect 97894 131996 97950 132005
rect 99574 132061 99630 132070
rect 99574 131996 99630 132005
rect 101254 132061 101310 132070
rect 101254 131996 101310 132005
rect 102934 132061 102990 132070
rect 102934 131996 102990 132005
rect 104614 132061 104670 132070
rect 104614 131996 104670 132005
rect 106294 132061 106350 132070
rect 106294 131996 106350 132005
rect 107974 132061 108030 132070
rect 107974 131996 108030 132005
rect 109654 132061 109710 132070
rect 109654 131996 109710 132005
rect 111334 132061 111390 132070
rect 111334 131996 111390 132005
rect 113014 132061 113070 132070
rect 113014 131996 113070 132005
rect 114694 132061 114750 132070
rect 114694 131996 114750 132005
rect 116374 132061 116430 132070
rect 116374 131996 116430 132005
rect 118054 132061 118110 132070
rect 118054 131996 118110 132005
rect 119734 132061 119790 132070
rect 119734 131996 119790 132005
rect 121414 132061 121470 132070
rect 121414 131996 121470 132005
rect 123094 132061 123150 132070
rect 123094 131996 123150 132005
rect 124774 132061 124830 132070
rect 124774 131996 124830 132005
rect 126454 132061 126510 132070
rect 126454 131996 126510 132005
rect 128134 132061 128190 132070
rect 128134 131996 128190 132005
rect 129814 132061 129870 132070
rect 129814 131996 129870 132005
rect 131494 132061 131550 132070
rect 131494 131996 131550 132005
rect 133174 132061 133230 132070
rect 133174 131996 133230 132005
rect 134854 132061 134910 132070
rect 134854 131996 134910 132005
rect 136534 132061 136590 132070
rect 136534 131996 136590 132005
rect 1714 131392 1798 131448
rect 1854 131392 1938 131448
rect 1714 131110 1938 131392
rect 1714 131058 1800 131110
rect 1852 131058 1938 131110
rect 136860 131448 137084 132145
rect 136860 131392 136944 131448
rect 137000 131392 137084 131448
rect 136860 131110 137084 131392
rect 1714 130774 1938 131058
rect 123532 131081 123588 131090
rect 123532 131016 123588 131025
rect 136860 131058 136946 131110
rect 136998 131058 137084 131110
rect 1714 130722 1800 130774
rect 1852 130722 1938 130774
rect 119942 130825 119998 130834
rect 119942 130760 119998 130769
rect 121110 130825 121166 130834
rect 121110 130760 121166 130769
rect 1714 130438 1938 130722
rect 1714 130386 1800 130438
rect 1852 130386 1938 130438
rect 1714 130102 1938 130386
rect 1714 130050 1800 130102
rect 1852 130050 1938 130102
rect 1714 129768 1938 130050
rect 1714 129712 1798 129768
rect 1854 129712 1938 129768
rect 1714 129430 1938 129712
rect 1714 129378 1800 129430
rect 1852 129378 1938 129430
rect 1714 129094 1938 129378
rect 1714 129042 1800 129094
rect 1852 129042 1938 129094
rect 1714 128758 1938 129042
rect 1714 128706 1800 128758
rect 1852 128706 1938 128758
rect 1714 128422 1938 128706
rect 1714 128370 1800 128422
rect 1852 128370 1938 128422
rect 1714 128088 1938 128370
rect 1714 128032 1798 128088
rect 1854 128032 1938 128088
rect 1714 127750 1938 128032
rect 1714 127698 1800 127750
rect 1852 127698 1938 127750
rect 1714 127414 1938 127698
rect 123546 129671 123574 131016
rect 136860 130774 137084 131058
rect 136860 130722 136946 130774
rect 136998 130722 137084 130774
rect 136860 130438 137084 130722
rect 136860 130386 136946 130438
rect 136998 130386 137084 130438
rect 136860 130102 137084 130386
rect 136860 130050 136946 130102
rect 136998 130050 137084 130102
rect 135984 129828 136040 129837
rect 135984 129763 136040 129772
rect 136860 129768 137084 130050
rect 132847 129723 132903 129732
rect 123546 129643 123644 129671
rect 132847 129658 132903 129667
rect 136860 129712 136944 129768
rect 137000 129712 137084 129768
rect 29562 127607 29618 127616
rect 29562 127542 29618 127551
rect 32058 127607 32114 127616
rect 32058 127542 32114 127551
rect 34554 127607 34610 127616
rect 34554 127542 34610 127551
rect 37050 127607 37106 127616
rect 37050 127542 37106 127551
rect 39546 127607 39602 127616
rect 39546 127542 39602 127551
rect 42042 127607 42098 127616
rect 42042 127542 42098 127551
rect 44538 127607 44594 127616
rect 44538 127542 44594 127551
rect 47034 127607 47090 127616
rect 47034 127542 47090 127551
rect 49530 127607 49586 127616
rect 49530 127542 49586 127551
rect 52026 127607 52082 127616
rect 52026 127542 52082 127551
rect 54522 127607 54578 127616
rect 54522 127542 54578 127551
rect 57018 127607 57074 127616
rect 57018 127542 57074 127551
rect 59514 127607 59570 127616
rect 59514 127542 59570 127551
rect 62010 127607 62066 127616
rect 62010 127542 62066 127551
rect 64506 127607 64562 127616
rect 64506 127542 64562 127551
rect 67002 127607 67058 127616
rect 67002 127542 67058 127551
rect 69498 127607 69554 127616
rect 69498 127542 69554 127551
rect 71994 127607 72050 127616
rect 71994 127542 72050 127551
rect 74490 127607 74546 127616
rect 74490 127542 74546 127551
rect 76986 127607 77042 127616
rect 76986 127542 77042 127551
rect 79482 127607 79538 127616
rect 79482 127542 79538 127551
rect 81978 127607 82034 127616
rect 81978 127542 82034 127551
rect 84474 127607 84530 127616
rect 84474 127542 84530 127551
rect 86970 127607 87026 127616
rect 86970 127542 87026 127551
rect 89466 127607 89522 127616
rect 89466 127542 89522 127551
rect 91962 127607 92018 127616
rect 91962 127542 92018 127551
rect 94458 127607 94514 127616
rect 94458 127542 94514 127551
rect 96954 127607 97010 127616
rect 96954 127542 97010 127551
rect 99450 127607 99506 127616
rect 99450 127542 99506 127551
rect 101946 127607 102002 127616
rect 101946 127542 102002 127551
rect 104442 127607 104498 127616
rect 104442 127542 104498 127551
rect 106938 127607 106994 127616
rect 106938 127542 106994 127551
rect 1714 127362 1800 127414
rect 1852 127362 1938 127414
rect 1714 127078 1938 127362
rect 1714 127026 1800 127078
rect 1852 127026 1938 127078
rect 1714 126742 1938 127026
rect 1714 126690 1800 126742
rect 1852 126690 1938 126742
rect 1714 126408 1938 126690
rect 1714 126352 1798 126408
rect 1854 126352 1938 126408
rect 1714 126070 1938 126352
rect 1714 126018 1800 126070
rect 1852 126018 1938 126070
rect 1714 125734 1938 126018
rect 1714 125682 1800 125734
rect 1852 125682 1938 125734
rect 1714 125398 1938 125682
rect 1714 125346 1800 125398
rect 1852 125346 1938 125398
rect 111005 125443 111061 125452
rect 111005 125378 111061 125387
rect 1714 125062 1938 125346
rect 1714 125010 1800 125062
rect 1852 125010 1938 125062
rect 1714 124728 1938 125010
rect 1714 124672 1798 124728
rect 1854 124672 1938 124728
rect 1714 124390 1938 124672
rect 1714 124338 1800 124390
rect 1852 124338 1938 124390
rect 1714 124054 1938 124338
rect 1714 124002 1800 124054
rect 1852 124002 1938 124054
rect 1714 123718 1938 124002
rect 1714 123666 1800 123718
rect 1852 123666 1938 123718
rect 1714 123382 1938 123666
rect 1714 123330 1800 123382
rect 1852 123330 1938 123382
rect 1714 123048 1938 123330
rect 1714 122992 1798 123048
rect 1854 122992 1938 123048
rect 1714 122710 1938 122992
rect 1714 122658 1800 122710
rect 1852 122658 1938 122710
rect 1714 122374 1938 122658
rect 1714 122322 1800 122374
rect 1852 122322 1938 122374
rect 1714 122038 1938 122322
rect 1714 121986 1800 122038
rect 1852 121986 1938 122038
rect 1714 121702 1938 121986
rect 111019 121742 111047 125378
rect 111129 124029 111185 124038
rect 111129 123964 111185 123973
rect 111143 121742 111171 123964
rect 114990 122615 115046 122624
rect 114990 122550 115046 122559
rect 1714 121650 1800 121702
rect 1852 121650 1938 121702
rect 1714 121368 1938 121650
rect 1714 121312 1798 121368
rect 1854 121312 1938 121368
rect 1714 121030 1938 121312
rect 115004 121265 115032 122550
rect 1714 120978 1800 121030
rect 1852 120978 1938 121030
rect 1714 120694 1938 120978
rect 1714 120642 1800 120694
rect 1852 120642 1938 120694
rect 1714 120358 1938 120642
rect 1714 120306 1800 120358
rect 1852 120306 1938 120358
rect 1714 120022 1938 120306
rect 1714 119970 1800 120022
rect 1852 119970 1938 120022
rect 1714 119688 1938 119970
rect 1714 119632 1798 119688
rect 1854 119632 1938 119688
rect 1714 119350 1938 119632
rect 1714 119298 1800 119350
rect 1852 119298 1938 119350
rect 1714 119014 1938 119298
rect 1714 118962 1800 119014
rect 1852 118962 1938 119014
rect 1714 118678 1938 118962
rect 1714 118626 1800 118678
rect 1852 118626 1938 118678
rect 1714 118342 1938 118626
rect 1714 118290 1800 118342
rect 1852 118290 1938 118342
rect 1714 118008 1938 118290
rect 1714 117952 1798 118008
rect 1854 117952 1938 118008
rect 1714 117670 1938 117952
rect 1714 117618 1800 117670
rect 1852 117618 1938 117670
rect 1714 117334 1938 117618
rect 1714 117282 1800 117334
rect 1852 117282 1938 117334
rect 1714 116998 1938 117282
rect 1714 116946 1800 116998
rect 1852 116946 1938 116998
rect 1714 116662 1938 116946
rect 1714 116610 1800 116662
rect 1852 116610 1938 116662
rect 1714 116328 1938 116610
rect 1714 116272 1798 116328
rect 1854 116272 1938 116328
rect 1714 115990 1938 116272
rect 1714 115938 1800 115990
rect 1852 115938 1938 115990
rect 1714 115654 1938 115938
rect 1714 115602 1800 115654
rect 1852 115602 1938 115654
rect 1714 115318 1938 115602
rect 1714 115266 1800 115318
rect 1852 115266 1938 115318
rect 1714 114982 1938 115266
rect 1714 114930 1800 114982
rect 1852 114930 1938 114982
rect 1714 114648 1938 114930
rect 1714 114592 1798 114648
rect 1854 114592 1938 114648
rect 1714 114310 1938 114592
rect 1714 114258 1800 114310
rect 1852 114258 1938 114310
rect 1714 113974 1938 114258
rect 1714 113922 1800 113974
rect 1852 113922 1938 113974
rect 1714 113638 1938 113922
rect 1714 113586 1800 113638
rect 1852 113586 1938 113638
rect 1714 113302 1938 113586
rect 1714 113250 1800 113302
rect 1852 113250 1938 113302
rect 1714 112968 1938 113250
rect 1714 112912 1798 112968
rect 1854 112912 1938 112968
rect 1714 112630 1938 112912
rect 1714 112578 1800 112630
rect 1852 112578 1938 112630
rect 1714 112294 1938 112578
rect 1714 112242 1800 112294
rect 1852 112242 1938 112294
rect 1714 111958 1938 112242
rect 1714 111906 1800 111958
rect 1852 111906 1938 111958
rect 1714 111622 1938 111906
rect 1714 111570 1800 111622
rect 1852 111570 1938 111622
rect 1714 111288 1938 111570
rect 1714 111232 1798 111288
rect 1854 111232 1938 111288
rect 1714 110950 1938 111232
rect 1714 110898 1800 110950
rect 1852 110898 1938 110950
rect 1714 110614 1938 110898
rect 1714 110562 1800 110614
rect 1852 110562 1938 110614
rect 1714 110278 1938 110562
rect 1714 110226 1800 110278
rect 1852 110226 1938 110278
rect 1714 109942 1938 110226
rect 1714 109890 1800 109942
rect 1852 109890 1938 109942
rect 1714 109608 1938 109890
rect 1714 109552 1798 109608
rect 1854 109552 1938 109608
rect 1714 109270 1938 109552
rect 1714 109218 1800 109270
rect 1852 109218 1938 109270
rect 1714 108934 1938 109218
rect 1714 108882 1800 108934
rect 1852 108882 1938 108934
rect 1714 108598 1938 108882
rect 1714 108546 1800 108598
rect 1852 108546 1938 108598
rect 1714 108262 1938 108546
rect 1714 108210 1800 108262
rect 1852 108210 1938 108262
rect 1714 107928 1938 108210
rect 1714 107872 1798 107928
rect 1854 107872 1938 107928
rect 1714 107590 1938 107872
rect 1714 107538 1800 107590
rect 1852 107538 1938 107590
rect 1714 107254 1938 107538
rect 1714 107202 1800 107254
rect 1852 107202 1938 107254
rect 1714 106918 1938 107202
rect 1714 106866 1800 106918
rect 1852 106866 1938 106918
rect 1714 106582 1938 106866
rect 1714 106530 1800 106582
rect 1852 106530 1938 106582
rect 1714 106248 1938 106530
rect 1714 106192 1798 106248
rect 1854 106192 1938 106248
rect 1714 105910 1938 106192
rect 1714 105858 1800 105910
rect 1852 105858 1938 105910
rect 1714 105574 1938 105858
rect 1714 105522 1800 105574
rect 1852 105522 1938 105574
rect 1714 105238 1938 105522
rect 1714 105186 1800 105238
rect 1852 105186 1938 105238
rect 1714 104902 1938 105186
rect 1714 104850 1800 104902
rect 1852 104850 1938 104902
rect 1714 104568 1938 104850
rect 1714 104512 1798 104568
rect 1854 104512 1938 104568
rect 1714 104230 1938 104512
rect 1714 104178 1800 104230
rect 1852 104178 1938 104230
rect 1714 103894 1938 104178
rect 1714 103842 1800 103894
rect 1852 103842 1938 103894
rect 1714 103558 1938 103842
rect 1714 103506 1800 103558
rect 1852 103506 1938 103558
rect 1714 103222 1938 103506
rect 1714 103170 1800 103222
rect 1852 103170 1938 103222
rect 1714 102888 1938 103170
rect 1714 102832 1798 102888
rect 1854 102832 1938 102888
rect 1714 102550 1938 102832
rect 1714 102498 1800 102550
rect 1852 102498 1938 102550
rect 1714 102214 1938 102498
rect 1714 102162 1800 102214
rect 1852 102162 1938 102214
rect 1714 101878 1938 102162
rect 1714 101826 1800 101878
rect 1852 101826 1938 101878
rect 1714 101542 1938 101826
rect 1714 101490 1800 101542
rect 1852 101490 1938 101542
rect 1714 101208 1938 101490
rect 1714 101152 1798 101208
rect 1854 101152 1938 101208
rect 1714 100870 1938 101152
rect 1714 100818 1800 100870
rect 1852 100818 1938 100870
rect 1714 100534 1938 100818
rect 1714 100482 1800 100534
rect 1852 100482 1938 100534
rect 1714 100198 1938 100482
rect 1714 100146 1800 100198
rect 1852 100146 1938 100198
rect 1714 99862 1938 100146
rect 1714 99810 1800 99862
rect 1852 99810 1938 99862
rect 1714 99528 1938 99810
rect 1714 99472 1798 99528
rect 1854 99472 1938 99528
rect 1714 99190 1938 99472
rect 1714 99138 1800 99190
rect 1852 99138 1938 99190
rect 1714 98854 1938 99138
rect 1714 98802 1800 98854
rect 1852 98802 1938 98854
rect 1714 98518 1938 98802
rect 1714 98466 1800 98518
rect 1852 98466 1938 98518
rect 1714 98182 1938 98466
rect 1714 98130 1800 98182
rect 1852 98130 1938 98182
rect 1714 97848 1938 98130
rect 1714 97792 1798 97848
rect 1854 97792 1938 97848
rect 1714 97510 1938 97792
rect 1714 97458 1800 97510
rect 1852 97458 1938 97510
rect 1714 97174 1938 97458
rect 1714 97122 1800 97174
rect 1852 97122 1938 97174
rect 1714 96838 1938 97122
rect 1714 96786 1800 96838
rect 1852 96786 1938 96838
rect 1714 96502 1938 96786
rect 1714 96450 1800 96502
rect 1852 96450 1938 96502
rect 1714 96168 1938 96450
rect 1714 96112 1798 96168
rect 1854 96112 1938 96168
rect 1714 95830 1938 96112
rect 1714 95778 1800 95830
rect 1852 95778 1938 95830
rect 1714 95494 1938 95778
rect 1714 95442 1800 95494
rect 1852 95442 1938 95494
rect 1714 95158 1938 95442
rect 1714 95106 1800 95158
rect 1852 95106 1938 95158
rect 1714 94822 1938 95106
rect 1714 94770 1800 94822
rect 1852 94770 1938 94822
rect 1714 94488 1938 94770
rect 1714 94432 1798 94488
rect 1854 94432 1938 94488
rect 1714 94150 1938 94432
rect 1714 94098 1800 94150
rect 1852 94098 1938 94150
rect 1714 93814 1938 94098
rect 1714 93762 1800 93814
rect 1852 93762 1938 93814
rect 1714 93478 1938 93762
rect 1714 93426 1800 93478
rect 1852 93426 1938 93478
rect 1714 93142 1938 93426
rect 1714 93090 1800 93142
rect 1852 93090 1938 93142
rect 1714 92808 1938 93090
rect 1714 92752 1798 92808
rect 1854 92752 1938 92808
rect 1714 92470 1938 92752
rect 1714 92418 1800 92470
rect 1852 92418 1938 92470
rect 1714 92134 1938 92418
rect 1714 92082 1800 92134
rect 1852 92082 1938 92134
rect 1714 91798 1938 92082
rect 1714 91746 1800 91798
rect 1852 91746 1938 91798
rect 1714 91462 1938 91746
rect 1714 91410 1800 91462
rect 1852 91410 1938 91462
rect 1714 91128 1938 91410
rect 1714 91072 1798 91128
rect 1854 91072 1938 91128
rect 1714 90790 1938 91072
rect 1714 90738 1800 90790
rect 1852 90738 1938 90790
rect 1714 90454 1938 90738
rect 1714 90402 1800 90454
rect 1852 90402 1938 90454
rect 1714 90118 1938 90402
rect 1714 90066 1800 90118
rect 1852 90066 1938 90118
rect 1714 89782 1938 90066
rect 1714 89730 1800 89782
rect 1852 89730 1938 89782
rect 1714 89448 1938 89730
rect 1714 89392 1798 89448
rect 1854 89392 1938 89448
rect 1714 89110 1938 89392
rect 1714 89058 1800 89110
rect 1852 89058 1938 89110
rect 1714 88774 1938 89058
rect 1714 88722 1800 88774
rect 1852 88722 1938 88774
rect 1714 88438 1938 88722
rect 1714 88386 1800 88438
rect 1852 88386 1938 88438
rect 1714 88102 1938 88386
rect 1714 88050 1800 88102
rect 1852 88050 1938 88102
rect 1714 87768 1938 88050
rect 1714 87712 1798 87768
rect 1854 87712 1938 87768
rect 1714 87430 1938 87712
rect 1714 87378 1800 87430
rect 1852 87378 1938 87430
rect 1714 87094 1938 87378
rect 1714 87042 1800 87094
rect 1852 87042 1938 87094
rect 1714 86758 1938 87042
rect 1714 86706 1800 86758
rect 1852 86706 1938 86758
rect 1714 86422 1938 86706
rect 1714 86370 1800 86422
rect 1852 86370 1938 86422
rect 1714 86088 1938 86370
rect 1714 86032 1798 86088
rect 1854 86032 1938 86088
rect 1714 85750 1938 86032
rect 1714 85698 1800 85750
rect 1852 85698 1938 85750
rect 1714 85414 1938 85698
rect 1714 85362 1800 85414
rect 1852 85362 1938 85414
rect 1714 85078 1938 85362
rect 1714 85026 1800 85078
rect 1852 85026 1938 85078
rect 1714 84742 1938 85026
rect 1714 84690 1800 84742
rect 1852 84690 1938 84742
rect 1714 84408 1938 84690
rect 1714 84352 1798 84408
rect 1854 84352 1938 84408
rect 1714 84070 1938 84352
rect 1714 84018 1800 84070
rect 1852 84018 1938 84070
rect 1714 83734 1938 84018
rect 1714 83682 1800 83734
rect 1852 83682 1938 83734
rect 1714 83398 1938 83682
rect 1714 83346 1800 83398
rect 1852 83346 1938 83398
rect 1714 83062 1938 83346
rect 1714 83010 1800 83062
rect 1852 83010 1938 83062
rect 1714 82728 1938 83010
rect 1714 82672 1798 82728
rect 1854 82672 1938 82728
rect 1714 82390 1938 82672
rect 1714 82338 1800 82390
rect 1852 82338 1938 82390
rect 1714 82054 1938 82338
rect 1714 82002 1800 82054
rect 1852 82002 1938 82054
rect 1714 81718 1938 82002
rect 1714 81666 1800 81718
rect 1852 81666 1938 81718
rect 1714 81382 1938 81666
rect 1714 81330 1800 81382
rect 1852 81330 1938 81382
rect 1714 81048 1938 81330
rect 1714 80992 1798 81048
rect 1854 80992 1938 81048
rect 1714 80710 1938 80992
rect 1714 80658 1800 80710
rect 1852 80658 1938 80710
rect 1714 80374 1938 80658
rect 1714 80322 1800 80374
rect 1852 80322 1938 80374
rect 1714 80038 1938 80322
rect 1714 79986 1800 80038
rect 1852 79986 1938 80038
rect 1714 79702 1938 79986
rect 1714 79650 1800 79702
rect 1852 79650 1938 79702
rect 1714 79368 1938 79650
rect 1714 79312 1798 79368
rect 1854 79312 1938 79368
rect 1714 79030 1938 79312
rect 1714 78978 1800 79030
rect 1852 78978 1938 79030
rect 1714 78694 1938 78978
rect 1714 78642 1800 78694
rect 1852 78642 1938 78694
rect 1714 78358 1938 78642
rect 1714 78306 1800 78358
rect 1852 78306 1938 78358
rect 1714 78022 1938 78306
rect 1714 77970 1800 78022
rect 1852 77970 1938 78022
rect 1714 77688 1938 77970
rect 1714 77632 1798 77688
rect 1854 77632 1938 77688
rect 1714 77350 1938 77632
rect 1714 77298 1800 77350
rect 1852 77298 1938 77350
rect 1714 77014 1938 77298
rect 1714 76962 1800 77014
rect 1852 76962 1938 77014
rect 1714 76678 1938 76962
rect 1714 76626 1800 76678
rect 1852 76626 1938 76678
rect 1714 76342 1938 76626
rect 1714 76290 1800 76342
rect 1852 76290 1938 76342
rect 1714 76008 1938 76290
rect 1714 75952 1798 76008
rect 1854 75952 1938 76008
rect 1714 75670 1938 75952
rect 1714 75618 1800 75670
rect 1852 75618 1938 75670
rect 1714 75334 1938 75618
rect 1714 75282 1800 75334
rect 1852 75282 1938 75334
rect 1714 74998 1938 75282
rect 1714 74946 1800 74998
rect 1852 74946 1938 74998
rect 1714 74662 1938 74946
rect 1714 74610 1800 74662
rect 1852 74610 1938 74662
rect 1714 74328 1938 74610
rect 1714 74272 1798 74328
rect 1854 74272 1938 74328
rect 1714 73990 1938 74272
rect 1714 73938 1800 73990
rect 1852 73938 1938 73990
rect 1714 73654 1938 73938
rect 1714 73602 1800 73654
rect 1852 73602 1938 73654
rect 1714 73318 1938 73602
rect 1714 73266 1800 73318
rect 1852 73266 1938 73318
rect 1714 72982 1938 73266
rect 1714 72930 1800 72982
rect 1852 72930 1938 72982
rect 1714 72648 1938 72930
rect 1714 72592 1798 72648
rect 1854 72592 1938 72648
rect 1714 72310 1938 72592
rect 1714 72258 1800 72310
rect 1852 72258 1938 72310
rect 1714 71974 1938 72258
rect 1714 71922 1800 71974
rect 1852 71922 1938 71974
rect 1714 71638 1938 71922
rect 1714 71586 1800 71638
rect 1852 71586 1938 71638
rect 1714 71302 1938 71586
rect 1714 71250 1800 71302
rect 1852 71250 1938 71302
rect 1714 70968 1938 71250
rect 1714 70912 1798 70968
rect 1854 70912 1938 70968
rect 1714 70630 1938 70912
rect 1714 70578 1800 70630
rect 1852 70578 1938 70630
rect 1714 70294 1938 70578
rect 1714 70242 1800 70294
rect 1852 70242 1938 70294
rect 1714 69958 1938 70242
rect 1714 69906 1800 69958
rect 1852 69906 1938 69958
rect 1714 69622 1938 69906
rect 1714 69570 1800 69622
rect 1852 69570 1938 69622
rect 1714 69288 1938 69570
rect 1714 69232 1798 69288
rect 1854 69232 1938 69288
rect 1714 68950 1938 69232
rect 1714 68898 1800 68950
rect 1852 68898 1938 68950
rect 1714 68614 1938 68898
rect 1714 68562 1800 68614
rect 1852 68562 1938 68614
rect 1714 68278 1938 68562
rect 1714 68226 1800 68278
rect 1852 68226 1938 68278
rect 1714 67942 1938 68226
rect 1714 67890 1800 67942
rect 1852 67890 1938 67942
rect 1714 67608 1938 67890
rect 1714 67552 1798 67608
rect 1854 67552 1938 67608
rect 1714 67270 1938 67552
rect 1714 67218 1800 67270
rect 1852 67218 1938 67270
rect 1714 66934 1938 67218
rect 1714 66882 1800 66934
rect 1852 66882 1938 66934
rect 1714 66598 1938 66882
rect 1714 66546 1800 66598
rect 1852 66546 1938 66598
rect 1714 66262 1938 66546
rect 1714 66210 1800 66262
rect 1852 66210 1938 66262
rect 1714 65928 1938 66210
rect 1714 65872 1798 65928
rect 1854 65872 1938 65928
rect 1714 65590 1938 65872
rect 1714 65538 1800 65590
rect 1852 65538 1938 65590
rect 1714 65254 1938 65538
rect 1714 65202 1800 65254
rect 1852 65202 1938 65254
rect 1714 64918 1938 65202
rect 1714 64866 1800 64918
rect 1852 64866 1938 64918
rect 1714 64582 1938 64866
rect 1714 64530 1800 64582
rect 1852 64530 1938 64582
rect 1714 64248 1938 64530
rect 1714 64192 1798 64248
rect 1854 64192 1938 64248
rect 1714 63910 1938 64192
rect 1714 63858 1800 63910
rect 1852 63858 1938 63910
rect 1714 63574 1938 63858
rect 1714 63522 1800 63574
rect 1852 63522 1938 63574
rect 1714 63238 1938 63522
rect 1714 63186 1800 63238
rect 1852 63186 1938 63238
rect 1714 62902 1938 63186
rect 1714 62850 1800 62902
rect 1852 62850 1938 62902
rect 1714 62568 1938 62850
rect 1714 62512 1798 62568
rect 1854 62512 1938 62568
rect 1714 62230 1938 62512
rect 1714 62178 1800 62230
rect 1852 62178 1938 62230
rect 1714 61894 1938 62178
rect 1714 61842 1800 61894
rect 1852 61842 1938 61894
rect 1714 61558 1938 61842
rect 1714 61506 1800 61558
rect 1852 61506 1938 61558
rect 1714 61222 1938 61506
rect 1714 61170 1800 61222
rect 1852 61170 1938 61222
rect 1714 60888 1938 61170
rect 1714 60832 1798 60888
rect 1854 60832 1938 60888
rect 1714 60550 1938 60832
rect 1714 60498 1800 60550
rect 1852 60498 1938 60550
rect 1714 60214 1938 60498
rect 1714 60162 1800 60214
rect 1852 60162 1938 60214
rect 1714 59878 1938 60162
rect 1714 59826 1800 59878
rect 1852 59826 1938 59878
rect 1714 59542 1938 59826
rect 1714 59490 1800 59542
rect 1852 59490 1938 59542
rect 1714 59208 1938 59490
rect 1714 59152 1798 59208
rect 1854 59152 1938 59208
rect 1714 58870 1938 59152
rect 1714 58818 1800 58870
rect 1852 58818 1938 58870
rect 1714 58534 1938 58818
rect 1714 58482 1800 58534
rect 1852 58482 1938 58534
rect 1714 58198 1938 58482
rect 1714 58146 1800 58198
rect 1852 58146 1938 58198
rect 1714 57862 1938 58146
rect 1714 57810 1800 57862
rect 1852 57810 1938 57862
rect 1714 57528 1938 57810
rect 1714 57472 1798 57528
rect 1854 57472 1938 57528
rect 1714 57190 1938 57472
rect 1714 57138 1800 57190
rect 1852 57138 1938 57190
rect 1714 56854 1938 57138
rect 1714 56802 1800 56854
rect 1852 56802 1938 56854
rect 1714 56518 1938 56802
rect 1714 56466 1800 56518
rect 1852 56466 1938 56518
rect 1714 56182 1938 56466
rect 1714 56130 1800 56182
rect 1852 56130 1938 56182
rect 1714 55848 1938 56130
rect 1714 55792 1798 55848
rect 1854 55792 1938 55848
rect 1714 55510 1938 55792
rect 1714 55458 1800 55510
rect 1852 55458 1938 55510
rect 1714 55174 1938 55458
rect 1714 55122 1800 55174
rect 1852 55122 1938 55174
rect 1714 54838 1938 55122
rect 1714 54786 1800 54838
rect 1852 54786 1938 54838
rect 1714 54502 1938 54786
rect 1714 54450 1800 54502
rect 1852 54450 1938 54502
rect 1714 54168 1938 54450
rect 1714 54112 1798 54168
rect 1854 54112 1938 54168
rect 1714 53830 1938 54112
rect 1714 53778 1800 53830
rect 1852 53778 1938 53830
rect 1714 53494 1938 53778
rect 1714 53442 1800 53494
rect 1852 53442 1938 53494
rect 1714 53158 1938 53442
rect 1714 53106 1800 53158
rect 1852 53106 1938 53158
rect 1714 52822 1938 53106
rect 1714 52770 1800 52822
rect 1852 52770 1938 52822
rect 1714 52488 1938 52770
rect 1714 52432 1798 52488
rect 1854 52432 1938 52488
rect 1714 52150 1938 52432
rect 1714 52098 1800 52150
rect 1852 52098 1938 52150
rect 1714 51814 1938 52098
rect 1714 51762 1800 51814
rect 1852 51762 1938 51814
rect 1714 51478 1938 51762
rect 1714 51426 1800 51478
rect 1852 51426 1938 51478
rect 1714 51142 1938 51426
rect 1714 51090 1800 51142
rect 1852 51090 1938 51142
rect 1714 50808 1938 51090
rect 1714 50752 1798 50808
rect 1854 50752 1938 50808
rect 1714 50470 1938 50752
rect 1714 50418 1800 50470
rect 1852 50418 1938 50470
rect 1714 50134 1938 50418
rect 1714 50082 1800 50134
rect 1852 50082 1938 50134
rect 1714 49798 1938 50082
rect 1714 49746 1800 49798
rect 1852 49746 1938 49798
rect 1714 49462 1938 49746
rect 1714 49410 1800 49462
rect 1852 49410 1938 49462
rect 1714 49128 1938 49410
rect 1714 49072 1798 49128
rect 1854 49072 1938 49128
rect 1714 48790 1938 49072
rect 1714 48738 1800 48790
rect 1852 48738 1938 48790
rect 1714 48454 1938 48738
rect 1714 48402 1800 48454
rect 1852 48402 1938 48454
rect 1714 48118 1938 48402
rect 1714 48066 1800 48118
rect 1852 48066 1938 48118
rect 1714 47782 1938 48066
rect 1714 47730 1800 47782
rect 1852 47730 1938 47782
rect 1714 47448 1938 47730
rect 1714 47392 1798 47448
rect 1854 47392 1938 47448
rect 1714 47110 1938 47392
rect 1714 47058 1800 47110
rect 1852 47058 1938 47110
rect 1714 46774 1938 47058
rect 1714 46722 1800 46774
rect 1852 46722 1938 46774
rect 1714 46438 1938 46722
rect 1714 46386 1800 46438
rect 1852 46386 1938 46438
rect 1714 46102 1938 46386
rect 1714 46050 1800 46102
rect 1852 46050 1938 46102
rect 1714 45768 1938 46050
rect 1714 45712 1798 45768
rect 1854 45712 1938 45768
rect 1714 45430 1938 45712
rect 1714 45378 1800 45430
rect 1852 45378 1938 45430
rect 1714 45094 1938 45378
rect 1714 45042 1800 45094
rect 1852 45042 1938 45094
rect 1714 44758 1938 45042
rect 1714 44706 1800 44758
rect 1852 44706 1938 44758
rect 1714 44422 1938 44706
rect 1714 44370 1800 44422
rect 1852 44370 1938 44422
rect 1714 44088 1938 44370
rect 1714 44032 1798 44088
rect 1854 44032 1938 44088
rect 1714 43750 1938 44032
rect 1714 43698 1800 43750
rect 1852 43698 1938 43750
rect 1714 43414 1938 43698
rect 1714 43362 1800 43414
rect 1852 43362 1938 43414
rect 1714 43078 1938 43362
rect 1714 43026 1800 43078
rect 1852 43026 1938 43078
rect 1714 42742 1938 43026
rect 1714 42690 1800 42742
rect 1852 42690 1938 42742
rect 1714 42408 1938 42690
rect 1714 42352 1798 42408
rect 1854 42352 1938 42408
rect 1714 42070 1938 42352
rect 1714 42018 1800 42070
rect 1852 42018 1938 42070
rect 1714 41734 1938 42018
rect 1714 41682 1800 41734
rect 1852 41682 1938 41734
rect 1714 41398 1938 41682
rect 1714 41346 1800 41398
rect 1852 41346 1938 41398
rect 1714 41062 1938 41346
rect 1714 41010 1800 41062
rect 1852 41010 1938 41062
rect 1714 40728 1938 41010
rect 1714 40672 1798 40728
rect 1854 40672 1938 40728
rect 1714 40390 1938 40672
rect 1714 40338 1800 40390
rect 1852 40338 1938 40390
rect 1714 40054 1938 40338
rect 1714 40002 1800 40054
rect 1852 40002 1938 40054
rect 14212 40102 14268 40111
rect 14212 40037 14268 40046
rect 1714 39718 1938 40002
rect 15157 40031 15213 40040
rect 15157 39966 15213 39975
rect 15971 40031 16027 40040
rect 15971 39966 16027 39975
rect 1714 39666 1800 39718
rect 1852 39666 1938 39718
rect 1714 39382 1938 39666
rect 1714 39330 1800 39382
rect 1852 39330 1938 39382
rect 1714 39048 1938 39330
rect 1714 38992 1798 39048
rect 1854 38992 1938 39048
rect 1714 38710 1938 38992
rect 1714 38658 1800 38710
rect 1852 38658 1938 38710
rect 1714 38374 1938 38658
rect 15157 38473 15213 38482
rect 1714 38322 1800 38374
rect 1852 38322 1938 38374
rect 14212 38402 14268 38411
rect 15157 38408 15213 38417
rect 15891 38473 15947 38482
rect 15891 38408 15947 38417
rect 14212 38337 14268 38346
rect 1714 38038 1938 38322
rect 1714 37986 1800 38038
rect 1852 37986 1938 38038
rect 1714 37702 1938 37986
rect 1714 37650 1800 37702
rect 1852 37650 1938 37702
rect 1714 37368 1938 37650
rect 1714 37312 1798 37368
rect 1854 37312 1938 37368
rect 1714 37030 1938 37312
rect 14212 37274 14268 37283
rect 14212 37209 14268 37218
rect 15157 37203 15213 37212
rect 15157 37138 15213 37147
rect 15811 37203 15867 37212
rect 15811 37138 15867 37147
rect 1714 36978 1800 37030
rect 1852 36978 1938 37030
rect 1714 36694 1938 36978
rect 1714 36642 1800 36694
rect 1852 36642 1938 36694
rect 1714 36358 1938 36642
rect 1714 36306 1800 36358
rect 1852 36306 1938 36358
rect 1714 36022 1938 36306
rect 1714 35970 1800 36022
rect 1852 35970 1938 36022
rect 1714 35688 1938 35970
rect 1714 35632 1798 35688
rect 1854 35632 1938 35688
rect 1714 35350 1938 35632
rect 15157 35645 15213 35654
rect 14212 35574 14268 35583
rect 15157 35580 15213 35589
rect 15731 35645 15787 35654
rect 15731 35580 15787 35589
rect 14212 35509 14268 35518
rect 1714 35298 1800 35350
rect 1852 35298 1938 35350
rect 1714 35014 1938 35298
rect 1714 34962 1800 35014
rect 1852 34962 1938 35014
rect 1714 34678 1938 34962
rect 1714 34626 1800 34678
rect 1852 34626 1938 34678
rect 1714 34342 1938 34626
rect 14212 34446 14268 34455
rect 14212 34381 14268 34390
rect 1714 34290 1800 34342
rect 1852 34290 1938 34342
rect 15157 34375 15213 34384
rect 15157 34310 15213 34319
rect 15651 34375 15707 34384
rect 15651 34310 15707 34319
rect 1714 34008 1938 34290
rect 1714 33952 1798 34008
rect 1854 33952 1938 34008
rect 1714 33670 1938 33952
rect 1714 33618 1800 33670
rect 1852 33618 1938 33670
rect 1714 33334 1938 33618
rect 1714 33282 1800 33334
rect 1852 33282 1938 33334
rect 1714 32998 1938 33282
rect 1714 32946 1800 32998
rect 1852 32946 1938 32998
rect 1714 32662 1938 32946
rect 15157 32817 15213 32826
rect 14212 32746 14268 32755
rect 15157 32752 15213 32761
rect 15571 32817 15627 32826
rect 15571 32752 15627 32761
rect 14212 32681 14268 32690
rect 1714 32610 1800 32662
rect 1852 32610 1938 32662
rect 1714 32328 1938 32610
rect 1714 32272 1798 32328
rect 1854 32272 1938 32328
rect 1714 31990 1938 32272
rect 1714 31938 1800 31990
rect 1852 31938 1938 31990
rect 1714 31654 1938 31938
rect 1714 31602 1800 31654
rect 1852 31602 1938 31654
rect 1714 31318 1938 31602
rect 14212 31618 14268 31627
rect 14212 31553 14268 31562
rect 15157 31547 15213 31556
rect 15157 31482 15213 31491
rect 15491 31547 15547 31556
rect 15491 31482 15547 31491
rect 1714 31266 1800 31318
rect 1852 31266 1938 31318
rect 1714 30982 1938 31266
rect 1714 30930 1800 30982
rect 1852 30930 1938 30982
rect 1714 30648 1938 30930
rect 1714 30592 1798 30648
rect 1854 30592 1938 30648
rect 1714 30310 1938 30592
rect 1714 30258 1800 30310
rect 1852 30258 1938 30310
rect 1714 29974 1938 30258
rect 1714 29922 1800 29974
rect 1852 29922 1938 29974
rect 15157 29989 15213 29998
rect 1714 29638 1938 29922
rect 14212 29918 14268 29927
rect 15157 29924 15213 29933
rect 15411 29989 15467 29998
rect 15411 29924 15467 29933
rect 14212 29853 14268 29862
rect 1714 29586 1800 29638
rect 1852 29586 1938 29638
rect 15294 29662 15350 29671
rect 15294 29597 15350 29606
rect 1714 29302 1938 29586
rect 1714 29250 1800 29302
rect 1852 29250 1938 29302
rect 1714 28968 1938 29250
rect 1714 28912 1798 28968
rect 1854 28912 1938 28968
rect 1714 28630 1938 28912
rect 1714 28578 1800 28630
rect 1852 28578 1938 28630
rect 1714 28294 1938 28578
rect 1714 28242 1800 28294
rect 1852 28242 1938 28294
rect 1714 27958 1938 28242
rect 1714 27906 1800 27958
rect 1852 27906 1938 27958
rect 1714 27622 1938 27906
rect 1714 27570 1800 27622
rect 1852 27570 1938 27622
rect 1714 27288 1938 27570
rect 1714 27232 1798 27288
rect 1854 27232 1938 27288
rect 1714 26950 1938 27232
rect 1714 26898 1800 26950
rect 1852 26898 1938 26950
rect 1714 26614 1938 26898
rect 1714 26562 1800 26614
rect 1852 26562 1938 26614
rect 1714 26278 1938 26562
rect 1714 26226 1800 26278
rect 1852 26226 1938 26278
rect 1714 25942 1938 26226
rect 1714 25890 1800 25942
rect 1852 25890 1938 25942
rect 1714 25608 1938 25890
rect 1714 25552 1798 25608
rect 1854 25552 1938 25608
rect 1714 25270 1938 25552
rect 2545 25361 2601 25370
rect 2545 25296 2601 25305
rect 1714 25218 1800 25270
rect 1852 25218 1938 25270
rect 1714 24934 1938 25218
rect 1714 24882 1800 24934
rect 1852 24882 1938 24934
rect 1714 24598 1938 24882
rect 1714 24546 1800 24598
rect 1852 24546 1938 24598
rect 1714 24262 1938 24546
rect 1714 24210 1800 24262
rect 1852 24210 1938 24262
rect 1714 23928 1938 24210
rect 1714 23872 1798 23928
rect 1854 23872 1938 23928
rect 1714 23590 1938 23872
rect 1714 23538 1800 23590
rect 1852 23538 1938 23590
rect 1714 23254 1938 23538
rect 1714 23202 1800 23254
rect 1852 23202 1938 23254
rect 1714 22918 1938 23202
rect 1714 22866 1800 22918
rect 1852 22866 1938 22918
rect 1714 22582 1938 22866
rect 1714 22530 1800 22582
rect 1852 22530 1938 22582
rect 1714 22248 1938 22530
rect 1714 22192 1798 22248
rect 1854 22192 1938 22248
rect 1714 21910 1938 22192
rect 1714 21858 1800 21910
rect 1852 21858 1938 21910
rect 1714 21574 1938 21858
rect 1714 21522 1800 21574
rect 1852 21522 1938 21574
rect 1714 21238 1938 21522
rect 1714 21186 1800 21238
rect 1852 21186 1938 21238
rect 1714 20902 1938 21186
rect 1714 20850 1800 20902
rect 1852 20850 1938 20902
rect 1714 20568 1938 20850
rect 1714 20512 1798 20568
rect 1854 20512 1938 20568
rect 1714 20230 1938 20512
rect 1714 20178 1800 20230
rect 1852 20178 1938 20230
rect 1714 19894 1938 20178
rect 1714 19842 1800 19894
rect 1852 19842 1938 19894
rect 1714 19558 1938 19842
rect 1714 19506 1800 19558
rect 1852 19506 1938 19558
rect 1714 19222 1938 19506
rect 1714 19170 1800 19222
rect 1852 19170 1938 19222
rect 1714 18888 1938 19170
rect 1714 18832 1798 18888
rect 1854 18832 1938 18888
rect 1714 18550 1938 18832
rect 1714 18498 1800 18550
rect 1852 18498 1938 18550
rect 1714 18214 1938 18498
rect 1714 18162 1800 18214
rect 1852 18162 1938 18214
rect 15210 18253 15266 18262
rect 15210 18188 15266 18197
rect 1714 17878 1938 18162
rect 1714 17826 1800 17878
rect 1852 17826 1938 17878
rect 1714 17542 1938 17826
rect 1714 17490 1800 17542
rect 1852 17490 1938 17542
rect 1714 17208 1938 17490
rect 1714 17152 1798 17208
rect 1854 17152 1938 17208
rect 1714 16870 1938 17152
rect 1714 16818 1800 16870
rect 1852 16818 1938 16870
rect 1714 16534 1938 16818
rect 1714 16482 1800 16534
rect 1852 16482 1938 16534
rect 1714 16198 1938 16482
rect 1714 16146 1800 16198
rect 1852 16146 1938 16198
rect 1714 15862 1938 16146
rect 1714 15810 1800 15862
rect 1852 15810 1938 15862
rect 1714 15528 1938 15810
rect 1714 15472 1798 15528
rect 1854 15472 1938 15528
rect 1714 15190 1938 15472
rect 15210 15425 15266 15434
rect 15210 15360 15266 15369
rect 1714 15138 1800 15190
rect 1852 15138 1938 15190
rect 1714 14854 1938 15138
rect 1714 14802 1800 14854
rect 1852 14802 1938 14854
rect 1714 14518 1938 14802
rect 1714 14466 1800 14518
rect 1852 14466 1938 14518
rect 1714 14182 1938 14466
rect 1714 14130 1800 14182
rect 1852 14130 1938 14182
rect 1714 13848 1938 14130
rect 15210 14011 15266 14020
rect 15210 13946 15266 13955
rect 1714 13792 1798 13848
rect 1854 13792 1938 13848
rect 1714 13510 1938 13792
rect 1714 13458 1800 13510
rect 1852 13458 1938 13510
rect 1714 13174 1938 13458
rect 1714 13122 1800 13174
rect 1852 13122 1938 13174
rect 1714 12838 1938 13122
rect 1714 12786 1800 12838
rect 1852 12786 1938 12838
rect 1714 12502 1938 12786
rect 15210 12597 15266 12606
rect 15210 12532 15266 12541
rect 1714 12450 1800 12502
rect 1852 12450 1938 12502
rect 1714 12168 1938 12450
rect 1714 12112 1798 12168
rect 1854 12112 1938 12168
rect 1714 11830 1938 12112
rect 1714 11778 1800 11830
rect 1852 11778 1938 11830
rect 1714 11494 1938 11778
rect 1714 11442 1800 11494
rect 1852 11442 1938 11494
rect 1714 11158 1938 11442
rect 1714 11106 1800 11158
rect 1852 11106 1938 11158
rect 1714 10822 1938 11106
rect 1714 10770 1800 10822
rect 1852 10770 1938 10822
rect 1714 10488 1938 10770
rect 1714 10432 1798 10488
rect 1854 10432 1938 10488
rect 1714 10150 1938 10432
rect 1714 10098 1800 10150
rect 1852 10098 1938 10150
rect 1714 9814 1938 10098
rect 2758 9912 2814 9921
rect 2758 9847 2814 9856
rect 1714 9762 1800 9814
rect 1852 9762 1938 9814
rect 1714 9478 1938 9762
rect 1714 9426 1800 9478
rect 1852 9426 1938 9478
rect 1714 9142 1938 9426
rect 1714 9090 1800 9142
rect 1852 9090 1938 9142
rect 1714 8808 1938 9090
rect 1714 8752 1798 8808
rect 1854 8752 1938 8808
rect 1714 8470 1938 8752
rect 1714 8418 1800 8470
rect 1852 8418 1938 8470
rect 1714 8134 1938 8418
rect 15308 8341 15336 29597
rect 123546 19575 123574 129643
rect 136860 129430 137084 129712
rect 136860 129378 136946 129430
rect 136998 129378 137084 129430
rect 136860 129094 137084 129378
rect 136860 129042 136946 129094
rect 136998 129042 137084 129094
rect 136860 128758 137084 129042
rect 136860 128706 136946 128758
rect 136998 128706 137084 128758
rect 136860 128422 137084 128706
rect 136860 128370 136946 128422
rect 136998 128370 137084 128422
rect 136860 128088 137084 128370
rect 136860 128032 136944 128088
rect 137000 128032 137084 128088
rect 136860 127750 137084 128032
rect 136860 127698 136946 127750
rect 136998 127698 137084 127750
rect 136860 127414 137084 127698
rect 136860 127362 136946 127414
rect 136998 127362 137084 127414
rect 136860 127078 137084 127362
rect 136860 127026 136946 127078
rect 136998 127026 137084 127078
rect 136860 126742 137084 127026
rect 136860 126690 136946 126742
rect 136998 126690 137084 126742
rect 136860 126408 137084 126690
rect 136860 126352 136944 126408
rect 137000 126352 137084 126408
rect 136860 126070 137084 126352
rect 136860 126018 136946 126070
rect 136998 126018 137084 126070
rect 136860 125734 137084 126018
rect 136860 125682 136946 125734
rect 136998 125682 137084 125734
rect 123616 125443 123672 125452
rect 123616 125378 123672 125387
rect 136860 125398 137084 125682
rect 136860 125346 136946 125398
rect 136998 125346 137084 125398
rect 136860 125062 137084 125346
rect 136860 125010 136946 125062
rect 136998 125010 137084 125062
rect 136860 124728 137084 125010
rect 136860 124672 136944 124728
rect 137000 124672 137084 124728
rect 136860 124390 137084 124672
rect 136860 124338 136946 124390
rect 136998 124338 137084 124390
rect 136860 124054 137084 124338
rect 123616 124029 123672 124038
rect 123616 123964 123672 123973
rect 136860 124002 136946 124054
rect 136998 124002 137084 124054
rect 136860 123718 137084 124002
rect 136860 123666 136946 123718
rect 136998 123666 137084 123718
rect 136860 123382 137084 123666
rect 136860 123330 136946 123382
rect 136998 123330 137084 123382
rect 136860 123048 137084 123330
rect 136860 122992 136944 123048
rect 137000 122992 137084 123048
rect 136860 122710 137084 122992
rect 136860 122658 136946 122710
rect 136998 122658 137084 122710
rect 123616 122615 123672 122624
rect 123616 122550 123672 122559
rect 136860 122374 137084 122658
rect 136860 122322 136946 122374
rect 136998 122322 137084 122374
rect 136860 122038 137084 122322
rect 136860 121986 136946 122038
rect 136998 121986 137084 122038
rect 136860 121702 137084 121986
rect 136860 121650 136946 121702
rect 136998 121650 137084 121702
rect 136860 121368 137084 121650
rect 136860 121312 136944 121368
rect 137000 121312 137084 121368
rect 136860 121030 137084 121312
rect 136860 120978 136946 121030
rect 136998 120978 137084 121030
rect 136860 120694 137084 120978
rect 136860 120642 136946 120694
rect 136998 120642 137084 120694
rect 136860 120358 137084 120642
rect 136860 120306 136946 120358
rect 136998 120306 137084 120358
rect 136860 120022 137084 120306
rect 136860 119970 136946 120022
rect 136998 119970 137084 120022
rect 136860 119688 137084 119970
rect 136860 119632 136944 119688
rect 137000 119632 137084 119688
rect 136860 119350 137084 119632
rect 136860 119298 136946 119350
rect 136998 119298 137084 119350
rect 136860 119014 137084 119298
rect 136860 118962 136946 119014
rect 136998 118962 137084 119014
rect 136860 118678 137084 118962
rect 136860 118626 136946 118678
rect 136998 118626 137084 118678
rect 136860 118342 137084 118626
rect 136860 118290 136946 118342
rect 136998 118290 137084 118342
rect 136860 118008 137084 118290
rect 136860 117952 136944 118008
rect 137000 117952 137084 118008
rect 136860 117670 137084 117952
rect 136860 117618 136946 117670
rect 136998 117618 137084 117670
rect 136860 117334 137084 117618
rect 136860 117282 136946 117334
rect 136998 117282 137084 117334
rect 136860 116998 137084 117282
rect 136860 116946 136946 116998
rect 136998 116946 137084 116998
rect 136860 116662 137084 116946
rect 136860 116610 136946 116662
rect 136998 116610 137084 116662
rect 136860 116328 137084 116610
rect 136860 116272 136944 116328
rect 137000 116272 137084 116328
rect 136860 115990 137084 116272
rect 136860 115938 136946 115990
rect 136998 115938 137084 115990
rect 136860 115654 137084 115938
rect 136860 115602 136946 115654
rect 136998 115602 137084 115654
rect 136860 115318 137084 115602
rect 136860 115266 136946 115318
rect 136998 115266 137084 115318
rect 136860 114982 137084 115266
rect 136860 114930 136946 114982
rect 136998 114930 137084 114982
rect 136860 114648 137084 114930
rect 136860 114592 136944 114648
rect 137000 114592 137084 114648
rect 136860 114310 137084 114592
rect 136860 114258 136946 114310
rect 136998 114258 137084 114310
rect 136860 113974 137084 114258
rect 136860 113922 136946 113974
rect 136998 113922 137084 113974
rect 136860 113638 137084 113922
rect 136860 113586 136946 113638
rect 136998 113586 137084 113638
rect 136860 113302 137084 113586
rect 136860 113250 136946 113302
rect 136998 113250 137084 113302
rect 136860 112968 137084 113250
rect 136860 112912 136944 112968
rect 137000 112912 137084 112968
rect 136197 112679 136253 112688
rect 136197 112614 136253 112623
rect 136860 112630 137084 112912
rect 136860 112578 136946 112630
rect 136998 112578 137084 112630
rect 136860 112294 137084 112578
rect 136860 112242 136946 112294
rect 136998 112242 137084 112294
rect 136860 111958 137084 112242
rect 136860 111906 136946 111958
rect 136998 111906 137084 111958
rect 136860 111622 137084 111906
rect 136860 111570 136946 111622
rect 136998 111570 137084 111622
rect 136860 111288 137084 111570
rect 136860 111232 136944 111288
rect 137000 111232 137084 111288
rect 136860 110950 137084 111232
rect 136860 110898 136946 110950
rect 136998 110898 137084 110950
rect 136860 110614 137084 110898
rect 136860 110562 136946 110614
rect 136998 110562 137084 110614
rect 136860 110278 137084 110562
rect 136860 110226 136946 110278
rect 136998 110226 137084 110278
rect 136860 109942 137084 110226
rect 136860 109890 136946 109942
rect 136998 109890 137084 109942
rect 136860 109608 137084 109890
rect 136860 109552 136944 109608
rect 137000 109552 137084 109608
rect 136860 109270 137084 109552
rect 136860 109218 136946 109270
rect 136998 109218 137084 109270
rect 136860 108934 137084 109218
rect 136860 108882 136946 108934
rect 136998 108882 137084 108934
rect 136860 108598 137084 108882
rect 136860 108546 136946 108598
rect 136998 108546 137084 108598
rect 136860 108262 137084 108546
rect 136860 108210 136946 108262
rect 136998 108210 137084 108262
rect 136860 107928 137084 108210
rect 136860 107872 136944 107928
rect 137000 107872 137084 107928
rect 136860 107590 137084 107872
rect 136860 107538 136946 107590
rect 136998 107538 137084 107590
rect 136860 107254 137084 107538
rect 136860 107202 136946 107254
rect 136998 107202 137084 107254
rect 136860 106918 137084 107202
rect 136860 106866 136946 106918
rect 136998 106866 137084 106918
rect 136860 106582 137084 106866
rect 136860 106530 136946 106582
rect 136998 106530 137084 106582
rect 136860 106248 137084 106530
rect 136860 106192 136944 106248
rect 137000 106192 137084 106248
rect 136860 105910 137084 106192
rect 136860 105858 136946 105910
rect 136998 105858 137084 105910
rect 136860 105574 137084 105858
rect 136860 105522 136946 105574
rect 136998 105522 137084 105574
rect 136860 105238 137084 105522
rect 136860 105186 136946 105238
rect 136998 105186 137084 105238
rect 136860 104902 137084 105186
rect 136860 104850 136946 104902
rect 136998 104850 137084 104902
rect 136860 104568 137084 104850
rect 136860 104512 136944 104568
rect 137000 104512 137084 104568
rect 136860 104230 137084 104512
rect 136860 104178 136946 104230
rect 136998 104178 137084 104230
rect 136860 103894 137084 104178
rect 136860 103842 136946 103894
rect 136998 103842 137084 103894
rect 136860 103558 137084 103842
rect 136860 103506 136946 103558
rect 136998 103506 137084 103558
rect 136860 103222 137084 103506
rect 136860 103170 136946 103222
rect 136998 103170 137084 103222
rect 136860 102888 137084 103170
rect 136860 102832 136944 102888
rect 137000 102832 137084 102888
rect 136860 102550 137084 102832
rect 136860 102498 136946 102550
rect 136998 102498 137084 102550
rect 136860 102214 137084 102498
rect 136860 102162 136946 102214
rect 136998 102162 137084 102214
rect 136860 101878 137084 102162
rect 136860 101826 136946 101878
rect 136998 101826 137084 101878
rect 136860 101542 137084 101826
rect 136860 101490 136946 101542
rect 136998 101490 137084 101542
rect 136860 101208 137084 101490
rect 136860 101152 136944 101208
rect 137000 101152 137084 101208
rect 136860 100870 137084 101152
rect 136860 100818 136946 100870
rect 136998 100818 137084 100870
rect 136860 100534 137084 100818
rect 136860 100482 136946 100534
rect 136998 100482 137084 100534
rect 136860 100198 137084 100482
rect 136860 100146 136946 100198
rect 136998 100146 137084 100198
rect 136860 99862 137084 100146
rect 136860 99810 136946 99862
rect 136998 99810 137084 99862
rect 136860 99528 137084 99810
rect 136860 99472 136944 99528
rect 137000 99472 137084 99528
rect 136860 99190 137084 99472
rect 136860 99138 136946 99190
rect 136998 99138 137084 99190
rect 136860 98854 137084 99138
rect 136860 98802 136946 98854
rect 136998 98802 137084 98854
rect 136860 98518 137084 98802
rect 136860 98466 136946 98518
rect 136998 98466 137084 98518
rect 136860 98182 137084 98466
rect 136860 98130 136946 98182
rect 136998 98130 137084 98182
rect 136860 97848 137084 98130
rect 136860 97792 136944 97848
rect 137000 97792 137084 97848
rect 136860 97510 137084 97792
rect 136860 97458 136946 97510
rect 136998 97458 137084 97510
rect 136860 97174 137084 97458
rect 136860 97122 136946 97174
rect 136998 97122 137084 97174
rect 136860 96838 137084 97122
rect 136860 96786 136946 96838
rect 136998 96786 137084 96838
rect 136860 96502 137084 96786
rect 136860 96450 136946 96502
rect 136998 96450 137084 96502
rect 136860 96168 137084 96450
rect 136860 96112 136944 96168
rect 137000 96112 137084 96168
rect 136860 95830 137084 96112
rect 136860 95778 136946 95830
rect 136998 95778 137084 95830
rect 136860 95494 137084 95778
rect 136860 95442 136946 95494
rect 136998 95442 137084 95494
rect 136860 95158 137084 95442
rect 136860 95106 136946 95158
rect 136998 95106 137084 95158
rect 136860 94822 137084 95106
rect 136860 94770 136946 94822
rect 136998 94770 137084 94822
rect 136860 94488 137084 94770
rect 136860 94432 136944 94488
rect 137000 94432 137084 94488
rect 136860 94150 137084 94432
rect 136860 94098 136946 94150
rect 136998 94098 137084 94150
rect 136860 93814 137084 94098
rect 136860 93762 136946 93814
rect 136998 93762 137084 93814
rect 136860 93478 137084 93762
rect 136860 93426 136946 93478
rect 136998 93426 137084 93478
rect 136860 93142 137084 93426
rect 136860 93090 136946 93142
rect 136998 93090 137084 93142
rect 136860 92808 137084 93090
rect 136860 92752 136944 92808
rect 137000 92752 137084 92808
rect 136860 92470 137084 92752
rect 136860 92418 136946 92470
rect 136998 92418 137084 92470
rect 136860 92134 137084 92418
rect 136860 92082 136946 92134
rect 136998 92082 137084 92134
rect 136860 91798 137084 92082
rect 136860 91746 136946 91798
rect 136998 91746 137084 91798
rect 136860 91462 137084 91746
rect 136860 91410 136946 91462
rect 136998 91410 137084 91462
rect 136860 91128 137084 91410
rect 136860 91072 136944 91128
rect 137000 91072 137084 91128
rect 136860 90790 137084 91072
rect 136860 90738 136946 90790
rect 136998 90738 137084 90790
rect 136860 90454 137084 90738
rect 136860 90402 136946 90454
rect 136998 90402 137084 90454
rect 136860 90118 137084 90402
rect 136860 90066 136946 90118
rect 136998 90066 137084 90118
rect 136860 89782 137084 90066
rect 136860 89730 136946 89782
rect 136998 89730 137084 89782
rect 136860 89448 137084 89730
rect 136860 89392 136944 89448
rect 137000 89392 137084 89448
rect 136860 89110 137084 89392
rect 136860 89058 136946 89110
rect 136998 89058 137084 89110
rect 136860 88774 137084 89058
rect 136860 88722 136946 88774
rect 136998 88722 137084 88774
rect 136860 88438 137084 88722
rect 136860 88386 136946 88438
rect 136998 88386 137084 88438
rect 136860 88102 137084 88386
rect 136860 88050 136946 88102
rect 136998 88050 137084 88102
rect 136860 87768 137084 88050
rect 136860 87712 136944 87768
rect 137000 87712 137084 87768
rect 136860 87430 137084 87712
rect 136860 87378 136946 87430
rect 136998 87378 137084 87430
rect 136860 87094 137084 87378
rect 136860 87042 136946 87094
rect 136998 87042 137084 87094
rect 136860 86758 137084 87042
rect 136860 86706 136946 86758
rect 136998 86706 137084 86758
rect 136860 86422 137084 86706
rect 136860 86370 136946 86422
rect 136998 86370 137084 86422
rect 136860 86088 137084 86370
rect 136860 86032 136944 86088
rect 137000 86032 137084 86088
rect 136860 85750 137084 86032
rect 136860 85698 136946 85750
rect 136998 85698 137084 85750
rect 136860 85414 137084 85698
rect 136860 85362 136946 85414
rect 136998 85362 137084 85414
rect 136860 85078 137084 85362
rect 136860 85026 136946 85078
rect 136998 85026 137084 85078
rect 136860 84742 137084 85026
rect 136860 84690 136946 84742
rect 136998 84690 137084 84742
rect 136860 84408 137084 84690
rect 136860 84352 136944 84408
rect 137000 84352 137084 84408
rect 136860 84070 137084 84352
rect 136860 84018 136946 84070
rect 136998 84018 137084 84070
rect 136860 83734 137084 84018
rect 136860 83682 136946 83734
rect 136998 83682 137084 83734
rect 136860 83398 137084 83682
rect 136860 83346 136946 83398
rect 136998 83346 137084 83398
rect 136860 83062 137084 83346
rect 136860 83010 136946 83062
rect 136998 83010 137084 83062
rect 136860 82728 137084 83010
rect 136860 82672 136944 82728
rect 137000 82672 137084 82728
rect 136860 82390 137084 82672
rect 136860 82338 136946 82390
rect 136998 82338 137084 82390
rect 136860 82054 137084 82338
rect 136860 82002 136946 82054
rect 136998 82002 137084 82054
rect 136860 81718 137084 82002
rect 136860 81666 136946 81718
rect 136998 81666 137084 81718
rect 136860 81382 137084 81666
rect 136860 81330 136946 81382
rect 136998 81330 137084 81382
rect 136860 81048 137084 81330
rect 136860 80992 136944 81048
rect 137000 80992 137084 81048
rect 136860 80710 137084 80992
rect 136860 80658 136946 80710
rect 136998 80658 137084 80710
rect 136860 80374 137084 80658
rect 136860 80322 136946 80374
rect 136998 80322 137084 80374
rect 136860 80038 137084 80322
rect 136860 79986 136946 80038
rect 136998 79986 137084 80038
rect 136860 79702 137084 79986
rect 136860 79650 136946 79702
rect 136998 79650 137084 79702
rect 136860 79368 137084 79650
rect 136860 79312 136944 79368
rect 137000 79312 137084 79368
rect 136860 79030 137084 79312
rect 136860 78978 136946 79030
rect 136998 78978 137084 79030
rect 136860 78694 137084 78978
rect 136860 78642 136946 78694
rect 136998 78642 137084 78694
rect 136860 78358 137084 78642
rect 136860 78306 136946 78358
rect 136998 78306 137084 78358
rect 136860 78022 137084 78306
rect 136860 77970 136946 78022
rect 136998 77970 137084 78022
rect 136860 77688 137084 77970
rect 136860 77632 136944 77688
rect 137000 77632 137084 77688
rect 136860 77350 137084 77632
rect 136860 77298 136946 77350
rect 136998 77298 137084 77350
rect 136860 77014 137084 77298
rect 136860 76962 136946 77014
rect 136998 76962 137084 77014
rect 136860 76678 137084 76962
rect 136860 76626 136946 76678
rect 136998 76626 137084 76678
rect 136860 76342 137084 76626
rect 136860 76290 136946 76342
rect 136998 76290 137084 76342
rect 136860 76008 137084 76290
rect 136860 75952 136944 76008
rect 137000 75952 137084 76008
rect 136860 75670 137084 75952
rect 136860 75618 136946 75670
rect 136998 75618 137084 75670
rect 136860 75334 137084 75618
rect 136860 75282 136946 75334
rect 136998 75282 137084 75334
rect 136860 74998 137084 75282
rect 136860 74946 136946 74998
rect 136998 74946 137084 74998
rect 136860 74662 137084 74946
rect 136860 74610 136946 74662
rect 136998 74610 137084 74662
rect 136860 74328 137084 74610
rect 136860 74272 136944 74328
rect 137000 74272 137084 74328
rect 136860 73990 137084 74272
rect 136860 73938 136946 73990
rect 136998 73938 137084 73990
rect 136860 73654 137084 73938
rect 136860 73602 136946 73654
rect 136998 73602 137084 73654
rect 136860 73318 137084 73602
rect 136860 73266 136946 73318
rect 136998 73266 137084 73318
rect 136860 72982 137084 73266
rect 136860 72930 136946 72982
rect 136998 72930 137084 72982
rect 136860 72648 137084 72930
rect 136860 72592 136944 72648
rect 137000 72592 137084 72648
rect 136860 72310 137084 72592
rect 136860 72258 136946 72310
rect 136998 72258 137084 72310
rect 136860 71974 137084 72258
rect 136860 71922 136946 71974
rect 136998 71922 137084 71974
rect 136860 71638 137084 71922
rect 136860 71586 136946 71638
rect 136998 71586 137084 71638
rect 136860 71302 137084 71586
rect 136860 71250 136946 71302
rect 136998 71250 137084 71302
rect 136860 70968 137084 71250
rect 136860 70912 136944 70968
rect 137000 70912 137084 70968
rect 136860 70630 137084 70912
rect 136860 70578 136946 70630
rect 136998 70578 137084 70630
rect 136860 70294 137084 70578
rect 136860 70242 136946 70294
rect 136998 70242 137084 70294
rect 136860 69958 137084 70242
rect 136860 69906 136946 69958
rect 136998 69906 137084 69958
rect 136860 69622 137084 69906
rect 136860 69570 136946 69622
rect 136998 69570 137084 69622
rect 136860 69288 137084 69570
rect 136860 69232 136944 69288
rect 137000 69232 137084 69288
rect 136860 68950 137084 69232
rect 136860 68898 136946 68950
rect 136998 68898 137084 68950
rect 136860 68614 137084 68898
rect 136860 68562 136946 68614
rect 136998 68562 137084 68614
rect 136860 68278 137084 68562
rect 136860 68226 136946 68278
rect 136998 68226 137084 68278
rect 136860 67942 137084 68226
rect 136860 67890 136946 67942
rect 136998 67890 137084 67942
rect 136860 67608 137084 67890
rect 136860 67552 136944 67608
rect 137000 67552 137084 67608
rect 136860 67270 137084 67552
rect 136860 67218 136946 67270
rect 136998 67218 137084 67270
rect 136860 66934 137084 67218
rect 136860 66882 136946 66934
rect 136998 66882 137084 66934
rect 136860 66598 137084 66882
rect 136860 66546 136946 66598
rect 136998 66546 137084 66598
rect 136860 66262 137084 66546
rect 136860 66210 136946 66262
rect 136998 66210 137084 66262
rect 136860 65928 137084 66210
rect 136860 65872 136944 65928
rect 137000 65872 137084 65928
rect 136860 65590 137084 65872
rect 136860 65538 136946 65590
rect 136998 65538 137084 65590
rect 136860 65254 137084 65538
rect 136860 65202 136946 65254
rect 136998 65202 137084 65254
rect 136860 64918 137084 65202
rect 136860 64866 136946 64918
rect 136998 64866 137084 64918
rect 136860 64582 137084 64866
rect 136860 64530 136946 64582
rect 136998 64530 137084 64582
rect 136860 64248 137084 64530
rect 136860 64192 136944 64248
rect 137000 64192 137084 64248
rect 136860 63910 137084 64192
rect 136860 63858 136946 63910
rect 136998 63858 137084 63910
rect 136860 63574 137084 63858
rect 136860 63522 136946 63574
rect 136998 63522 137084 63574
rect 136860 63238 137084 63522
rect 136860 63186 136946 63238
rect 136998 63186 137084 63238
rect 136860 62902 137084 63186
rect 136860 62850 136946 62902
rect 136998 62850 137084 62902
rect 136860 62568 137084 62850
rect 136860 62512 136944 62568
rect 137000 62512 137084 62568
rect 136860 62230 137084 62512
rect 136860 62178 136946 62230
rect 136998 62178 137084 62230
rect 136860 61894 137084 62178
rect 136860 61842 136946 61894
rect 136998 61842 137084 61894
rect 136860 61558 137084 61842
rect 136860 61506 136946 61558
rect 136998 61506 137084 61558
rect 136860 61222 137084 61506
rect 136860 61170 136946 61222
rect 136998 61170 137084 61222
rect 136860 60888 137084 61170
rect 136860 60832 136944 60888
rect 137000 60832 137084 60888
rect 136860 60550 137084 60832
rect 136860 60498 136946 60550
rect 136998 60498 137084 60550
rect 136860 60214 137084 60498
rect 136860 60162 136946 60214
rect 136998 60162 137084 60214
rect 136860 59878 137084 60162
rect 136860 59826 136946 59878
rect 136998 59826 137084 59878
rect 136860 59542 137084 59826
rect 136860 59490 136946 59542
rect 136998 59490 137084 59542
rect 136860 59208 137084 59490
rect 136860 59152 136944 59208
rect 137000 59152 137084 59208
rect 136860 58870 137084 59152
rect 136860 58818 136946 58870
rect 136998 58818 137084 58870
rect 136860 58534 137084 58818
rect 136860 58482 136946 58534
rect 136998 58482 137084 58534
rect 136860 58198 137084 58482
rect 136860 58146 136946 58198
rect 136998 58146 137084 58198
rect 136860 57862 137084 58146
rect 136860 57810 136946 57862
rect 136998 57810 137084 57862
rect 136860 57528 137084 57810
rect 136860 57472 136944 57528
rect 137000 57472 137084 57528
rect 136860 57190 137084 57472
rect 136860 57138 136946 57190
rect 136998 57138 137084 57190
rect 136860 56854 137084 57138
rect 136860 56802 136946 56854
rect 136998 56802 137084 56854
rect 136860 56518 137084 56802
rect 136860 56466 136946 56518
rect 136998 56466 137084 56518
rect 136860 56182 137084 56466
rect 136860 56130 136946 56182
rect 136998 56130 137084 56182
rect 136860 55848 137084 56130
rect 136860 55792 136944 55848
rect 137000 55792 137084 55848
rect 136860 55510 137084 55792
rect 136860 55458 136946 55510
rect 136998 55458 137084 55510
rect 136860 55174 137084 55458
rect 136860 55122 136946 55174
rect 136998 55122 137084 55174
rect 136860 54838 137084 55122
rect 136860 54786 136946 54838
rect 136998 54786 137084 54838
rect 136860 54502 137084 54786
rect 136860 54450 136946 54502
rect 136998 54450 137084 54502
rect 136860 54168 137084 54450
rect 136860 54112 136944 54168
rect 137000 54112 137084 54168
rect 136860 53830 137084 54112
rect 136860 53778 136946 53830
rect 136998 53778 137084 53830
rect 136860 53494 137084 53778
rect 136860 53442 136946 53494
rect 136998 53442 137084 53494
rect 136860 53158 137084 53442
rect 136860 53106 136946 53158
rect 136998 53106 137084 53158
rect 136860 52822 137084 53106
rect 136860 52770 136946 52822
rect 136998 52770 137084 52822
rect 136860 52488 137084 52770
rect 136860 52432 136944 52488
rect 137000 52432 137084 52488
rect 136860 52150 137084 52432
rect 136860 52098 136946 52150
rect 136998 52098 137084 52150
rect 136860 51814 137084 52098
rect 136860 51762 136946 51814
rect 136998 51762 137084 51814
rect 136860 51478 137084 51762
rect 136860 51426 136946 51478
rect 136998 51426 137084 51478
rect 136860 51142 137084 51426
rect 136860 51090 136946 51142
rect 136998 51090 137084 51142
rect 136860 50808 137084 51090
rect 136860 50752 136944 50808
rect 137000 50752 137084 50808
rect 136860 50470 137084 50752
rect 136860 50418 136946 50470
rect 136998 50418 137084 50470
rect 136860 50134 137084 50418
rect 136860 50082 136946 50134
rect 136998 50082 137084 50134
rect 136860 49798 137084 50082
rect 136860 49746 136946 49798
rect 136998 49746 137084 49798
rect 136860 49462 137084 49746
rect 136860 49410 136946 49462
rect 136998 49410 137084 49462
rect 136860 49128 137084 49410
rect 136860 49072 136944 49128
rect 137000 49072 137084 49128
rect 136860 48790 137084 49072
rect 136860 48738 136946 48790
rect 136998 48738 137084 48790
rect 136860 48454 137084 48738
rect 136860 48402 136946 48454
rect 136998 48402 137084 48454
rect 136860 48118 137084 48402
rect 136860 48066 136946 48118
rect 136998 48066 137084 48118
rect 136860 47782 137084 48066
rect 136860 47730 136946 47782
rect 136998 47730 137084 47782
rect 136860 47448 137084 47730
rect 136860 47392 136944 47448
rect 137000 47392 137084 47448
rect 136860 47110 137084 47392
rect 136860 47058 136946 47110
rect 136998 47058 137084 47110
rect 136860 46774 137084 47058
rect 136860 46722 136946 46774
rect 136998 46722 137084 46774
rect 136860 46438 137084 46722
rect 136860 46386 136946 46438
rect 136998 46386 137084 46438
rect 136860 46102 137084 46386
rect 136860 46050 136946 46102
rect 136998 46050 137084 46102
rect 136860 45768 137084 46050
rect 136860 45712 136944 45768
rect 137000 45712 137084 45768
rect 136860 45430 137084 45712
rect 136860 45378 136946 45430
rect 136998 45378 137084 45430
rect 136860 45094 137084 45378
rect 136860 45042 136946 45094
rect 136998 45042 137084 45094
rect 136860 44758 137084 45042
rect 136860 44706 136946 44758
rect 136998 44706 137084 44758
rect 136860 44422 137084 44706
rect 136860 44370 136946 44422
rect 136998 44370 137084 44422
rect 136860 44088 137084 44370
rect 136860 44032 136944 44088
rect 137000 44032 137084 44088
rect 136860 43750 137084 44032
rect 136860 43698 136946 43750
rect 136998 43698 137084 43750
rect 136860 43414 137084 43698
rect 136860 43362 136946 43414
rect 136998 43362 137084 43414
rect 136860 43078 137084 43362
rect 136860 43026 136946 43078
rect 136998 43026 137084 43078
rect 136860 42742 137084 43026
rect 136860 42690 136946 42742
rect 136998 42690 137084 42742
rect 136860 42408 137084 42690
rect 136860 42352 136944 42408
rect 137000 42352 137084 42408
rect 136860 42070 137084 42352
rect 136860 42018 136946 42070
rect 136998 42018 137084 42070
rect 136860 41734 137084 42018
rect 136860 41682 136946 41734
rect 136998 41682 137084 41734
rect 136860 41398 137084 41682
rect 136860 41346 136946 41398
rect 136998 41346 137084 41398
rect 136860 41062 137084 41346
rect 136860 41010 136946 41062
rect 136998 41010 137084 41062
rect 136860 40728 137084 41010
rect 136860 40672 136944 40728
rect 137000 40672 137084 40728
rect 136860 40390 137084 40672
rect 136860 40338 136946 40390
rect 136998 40338 137084 40390
rect 136860 40054 137084 40338
rect 136860 40002 136946 40054
rect 136998 40002 137084 40054
rect 136860 39718 137084 40002
rect 136860 39666 136946 39718
rect 136998 39666 137084 39718
rect 136860 39382 137084 39666
rect 136860 39330 136946 39382
rect 136998 39330 137084 39382
rect 136860 39048 137084 39330
rect 136860 38992 136944 39048
rect 137000 38992 137084 39048
rect 136860 38710 137084 38992
rect 136860 38658 136946 38710
rect 136998 38658 137084 38710
rect 136860 38374 137084 38658
rect 136860 38322 136946 38374
rect 136998 38322 137084 38374
rect 136860 38038 137084 38322
rect 136860 37986 136946 38038
rect 136998 37986 137084 38038
rect 136860 37702 137084 37986
rect 136860 37650 136946 37702
rect 136998 37650 137084 37702
rect 136860 37368 137084 37650
rect 136860 37312 136944 37368
rect 137000 37312 137084 37368
rect 136860 37030 137084 37312
rect 136860 36978 136946 37030
rect 136998 36978 137084 37030
rect 136860 36694 137084 36978
rect 136860 36642 136946 36694
rect 136998 36642 137084 36694
rect 136860 36358 137084 36642
rect 136860 36306 136946 36358
rect 136998 36306 137084 36358
rect 136860 36022 137084 36306
rect 136860 35970 136946 36022
rect 136998 35970 137084 36022
rect 136860 35688 137084 35970
rect 136860 35632 136944 35688
rect 137000 35632 137084 35688
rect 136860 35350 137084 35632
rect 136860 35298 136946 35350
rect 136998 35298 137084 35350
rect 136860 35014 137084 35298
rect 136860 34962 136946 35014
rect 136998 34962 137084 35014
rect 136860 34678 137084 34962
rect 136860 34626 136946 34678
rect 136998 34626 137084 34678
rect 136860 34342 137084 34626
rect 136860 34290 136946 34342
rect 136998 34290 137084 34342
rect 136860 34008 137084 34290
rect 136860 33952 136944 34008
rect 137000 33952 137084 34008
rect 136860 33670 137084 33952
rect 136860 33618 136946 33670
rect 136998 33618 137084 33670
rect 136860 33334 137084 33618
rect 136860 33282 136946 33334
rect 136998 33282 137084 33334
rect 136860 32998 137084 33282
rect 136860 32946 136946 32998
rect 136998 32946 137084 32998
rect 136860 32662 137084 32946
rect 136860 32610 136946 32662
rect 136998 32610 137084 32662
rect 136860 32328 137084 32610
rect 136860 32272 136944 32328
rect 137000 32272 137084 32328
rect 136860 31990 137084 32272
rect 136860 31938 136946 31990
rect 136998 31938 137084 31990
rect 136860 31654 137084 31938
rect 136860 31602 136946 31654
rect 136998 31602 137084 31654
rect 136860 31318 137084 31602
rect 136860 31266 136946 31318
rect 136998 31266 137084 31318
rect 136860 30982 137084 31266
rect 136860 30930 136946 30982
rect 136998 30930 137084 30982
rect 136860 30648 137084 30930
rect 136860 30592 136944 30648
rect 137000 30592 137084 30648
rect 136860 30310 137084 30592
rect 136860 30258 136946 30310
rect 136998 30258 137084 30310
rect 136860 29974 137084 30258
rect 136860 29922 136946 29974
rect 136998 29922 137084 29974
rect 136860 29638 137084 29922
rect 136860 29586 136946 29638
rect 136998 29586 137084 29638
rect 136860 29302 137084 29586
rect 136860 29250 136946 29302
rect 136998 29250 137084 29302
rect 136860 28968 137084 29250
rect 136860 28912 136944 28968
rect 137000 28912 137084 28968
rect 136860 28630 137084 28912
rect 136860 28578 136946 28630
rect 136998 28578 137084 28630
rect 136860 28294 137084 28578
rect 136860 28242 136946 28294
rect 136998 28242 137084 28294
rect 136860 27958 137084 28242
rect 136860 27906 136946 27958
rect 136998 27906 137084 27958
rect 136860 27622 137084 27906
rect 136860 27570 136946 27622
rect 136998 27570 137084 27622
rect 136860 27288 137084 27570
rect 136860 27232 136944 27288
rect 137000 27232 137084 27288
rect 136860 26950 137084 27232
rect 136860 26898 136946 26950
rect 136998 26898 137084 26950
rect 136860 26614 137084 26898
rect 136860 26562 136946 26614
rect 136998 26562 137084 26614
rect 136860 26278 137084 26562
rect 136860 26226 136946 26278
rect 136998 26226 137084 26278
rect 136860 25942 137084 26226
rect 136860 25890 136946 25942
rect 136998 25890 137084 25942
rect 136860 25608 137084 25890
rect 136860 25552 136944 25608
rect 137000 25552 137084 25608
rect 136860 25270 137084 25552
rect 136860 25218 136946 25270
rect 136998 25218 137084 25270
rect 136860 24934 137084 25218
rect 136860 24882 136946 24934
rect 136998 24882 137084 24934
rect 136860 24598 137084 24882
rect 136860 24546 136946 24598
rect 136998 24546 137084 24598
rect 136860 24262 137084 24546
rect 136860 24210 136946 24262
rect 136998 24210 137084 24262
rect 136860 23928 137084 24210
rect 136860 23872 136944 23928
rect 137000 23872 137084 23928
rect 136860 23590 137084 23872
rect 136860 23538 136946 23590
rect 136998 23538 137084 23590
rect 136860 23254 137084 23538
rect 136860 23202 136946 23254
rect 136998 23202 137084 23254
rect 136860 22918 137084 23202
rect 136860 22866 136946 22918
rect 136998 22866 137084 22918
rect 136860 22582 137084 22866
rect 136860 22530 136946 22582
rect 136998 22530 137084 22582
rect 136860 22248 137084 22530
rect 136860 22192 136944 22248
rect 137000 22192 137084 22248
rect 136860 21910 137084 22192
rect 136860 21858 136946 21910
rect 136998 21858 137084 21910
rect 136860 21574 137084 21858
rect 136860 21522 136946 21574
rect 136998 21522 137084 21574
rect 136860 21238 137084 21522
rect 136860 21186 136946 21238
rect 136998 21186 137084 21238
rect 136860 20902 137084 21186
rect 136860 20850 136946 20902
rect 136998 20850 137084 20902
rect 136860 20568 137084 20850
rect 136860 20512 136944 20568
rect 137000 20512 137084 20568
rect 136860 20230 137084 20512
rect 136860 20178 136946 20230
rect 136998 20178 137084 20230
rect 136860 19894 137084 20178
rect 136860 19842 136946 19894
rect 136998 19842 137084 19894
rect 123532 19566 123588 19575
rect 23766 18262 23794 19547
rect 123532 19501 123588 19510
rect 136860 19558 137084 19842
rect 136860 19506 136946 19558
rect 136998 19506 137084 19558
rect 124614 19310 124670 19319
rect 123331 19239 123387 19248
rect 123331 19174 123387 19183
rect 123669 19239 123725 19248
rect 124614 19245 124670 19254
rect 123669 19174 123725 19183
rect 136860 19222 137084 19506
rect 136860 19170 136946 19222
rect 136998 19170 137084 19222
rect 23752 18253 23808 18262
rect 23752 18188 23808 18197
rect 27469 15434 27497 19070
rect 136860 18888 137084 19170
rect 136860 18832 136944 18888
rect 137000 18832 137084 18888
rect 136860 18550 137084 18832
rect 136860 18498 136946 18550
rect 136998 18498 137084 18550
rect 136860 18214 137084 18498
rect 136860 18162 136946 18214
rect 136998 18162 137084 18214
rect 136860 17878 137084 18162
rect 136860 17826 136946 17878
rect 136998 17826 137084 17878
rect 123251 17681 123307 17690
rect 123251 17616 123307 17625
rect 123669 17681 123725 17690
rect 123669 17616 123725 17625
rect 124614 17610 124670 17619
rect 124614 17545 124670 17554
rect 136860 17542 137084 17826
rect 136860 17490 136946 17542
rect 136998 17490 137084 17542
rect 136860 17208 137084 17490
rect 136860 17152 136944 17208
rect 137000 17152 137084 17208
rect 136860 16870 137084 17152
rect 136860 16818 136946 16870
rect 136998 16818 137084 16870
rect 136860 16534 137084 16818
rect 124614 16482 124670 16491
rect 123171 16411 123227 16420
rect 123171 16346 123227 16355
rect 123669 16411 123725 16420
rect 124614 16417 124670 16426
rect 136860 16482 136946 16534
rect 136998 16482 137084 16534
rect 123669 16346 123725 16355
rect 136860 16198 137084 16482
rect 136860 16146 136946 16198
rect 136998 16146 137084 16198
rect 136860 15862 137084 16146
rect 136860 15810 136946 15862
rect 136998 15810 137084 15862
rect 136860 15528 137084 15810
rect 136860 15472 136944 15528
rect 137000 15472 137084 15528
rect 27455 15425 27511 15434
rect 27455 15360 27511 15369
rect 136860 15190 137084 15472
rect 136860 15138 136946 15190
rect 136998 15138 137084 15190
rect 123091 14853 123147 14862
rect 123091 14788 123147 14797
rect 123669 14853 123725 14862
rect 123669 14788 123725 14797
rect 136860 14854 137084 15138
rect 136860 14802 136946 14854
rect 136998 14802 137084 14854
rect 124614 14782 124670 14791
rect 124614 14717 124670 14726
rect 136860 14518 137084 14802
rect 136860 14466 136946 14518
rect 136998 14466 137084 14518
rect 136860 14182 137084 14466
rect 136860 14130 136946 14182
rect 136998 14130 137084 14182
rect 27703 14011 27759 14020
rect 27703 13946 27759 13955
rect 27579 12597 27635 12606
rect 27579 12532 27635 12541
rect 27593 9457 27621 12532
rect 27717 9457 27745 13946
rect 136860 13848 137084 14130
rect 136860 13792 136944 13848
rect 137000 13792 137084 13848
rect 124614 13654 124670 13663
rect 123011 13583 123067 13592
rect 123011 13518 123067 13527
rect 123669 13583 123725 13592
rect 124614 13589 124670 13598
rect 123669 13518 123725 13527
rect 136860 13510 137084 13792
rect 136860 13458 136946 13510
rect 136998 13458 137084 13510
rect 29562 13261 29618 13270
rect 29562 13196 29618 13205
rect 32058 13261 32114 13270
rect 32058 13196 32114 13205
rect 34554 13261 34610 13270
rect 34554 13196 34610 13205
rect 37050 13261 37106 13270
rect 37050 13196 37106 13205
rect 39546 13261 39602 13270
rect 39546 13196 39602 13205
rect 42042 13261 42098 13270
rect 42042 13196 42098 13205
rect 44538 13261 44594 13270
rect 44538 13196 44594 13205
rect 47034 13261 47090 13270
rect 47034 13196 47090 13205
rect 49530 13261 49586 13270
rect 49530 13196 49586 13205
rect 52026 13261 52082 13270
rect 52026 13196 52082 13205
rect 54522 13261 54578 13270
rect 54522 13196 54578 13205
rect 57018 13261 57074 13270
rect 57018 13196 57074 13205
rect 59514 13261 59570 13270
rect 59514 13196 59570 13205
rect 62010 13261 62066 13270
rect 62010 13196 62066 13205
rect 64506 13261 64562 13270
rect 64506 13196 64562 13205
rect 67002 13261 67058 13270
rect 67002 13196 67058 13205
rect 69498 13261 69554 13270
rect 69498 13196 69554 13205
rect 71994 13261 72050 13270
rect 71994 13196 72050 13205
rect 74490 13261 74546 13270
rect 74490 13196 74546 13205
rect 76986 13261 77042 13270
rect 76986 13196 77042 13205
rect 79482 13261 79538 13270
rect 79482 13196 79538 13205
rect 81978 13261 82034 13270
rect 81978 13196 82034 13205
rect 84474 13261 84530 13270
rect 84474 13196 84530 13205
rect 86970 13261 87026 13270
rect 86970 13196 87026 13205
rect 89466 13261 89522 13270
rect 89466 13196 89522 13205
rect 91962 13261 92018 13270
rect 91962 13196 92018 13205
rect 94458 13261 94514 13270
rect 94458 13196 94514 13205
rect 96954 13261 97010 13270
rect 96954 13196 97010 13205
rect 99450 13261 99506 13270
rect 99450 13196 99506 13205
rect 101946 13261 102002 13270
rect 101946 13196 102002 13205
rect 104442 13261 104498 13270
rect 104442 13196 104498 13205
rect 106938 13261 106994 13270
rect 106938 13196 106994 13205
rect 136860 13174 137084 13458
rect 136860 13122 136946 13174
rect 136998 13122 137084 13174
rect 136860 12838 137084 13122
rect 136860 12786 136946 12838
rect 136998 12786 137084 12838
rect 136860 12502 137084 12786
rect 136860 12450 136946 12502
rect 136998 12450 137084 12502
rect 136860 12168 137084 12450
rect 136860 12112 136944 12168
rect 137000 12112 137084 12168
rect 122931 12025 122987 12034
rect 122931 11960 122987 11969
rect 123669 12025 123725 12034
rect 123669 11960 123725 11969
rect 124614 11954 124670 11963
rect 124614 11889 124670 11898
rect 136860 11830 137084 12112
rect 136860 11778 136946 11830
rect 136998 11778 137084 11830
rect 136860 11494 137084 11778
rect 136860 11442 136946 11494
rect 136998 11442 137084 11494
rect 136860 11158 137084 11442
rect 136860 11106 136946 11158
rect 136998 11106 137084 11158
rect 124614 10826 124670 10835
rect 122851 10755 122907 10764
rect 122851 10690 122907 10699
rect 123669 10755 123725 10764
rect 124614 10761 124670 10770
rect 136860 10822 137084 11106
rect 136860 10770 136946 10822
rect 136998 10770 137084 10822
rect 123669 10690 123725 10699
rect 136860 10488 137084 10770
rect 136860 10432 136944 10488
rect 137000 10432 137084 10488
rect 136860 10150 137084 10432
rect 136860 10098 136946 10150
rect 136998 10098 137084 10150
rect 136860 9814 137084 10098
rect 136860 9762 136946 9814
rect 136998 9762 137084 9814
rect 136860 9478 137084 9762
rect 136860 9426 136946 9478
rect 136998 9426 137084 9478
rect 122771 9197 122827 9206
rect 122771 9132 122827 9141
rect 123669 9197 123725 9206
rect 123669 9132 123725 9141
rect 136860 9142 137084 9426
rect 124614 9126 124670 9135
rect 124614 9061 124670 9070
rect 136860 9090 136946 9142
rect 136998 9090 137084 9142
rect 5979 8317 6035 8326
rect 15238 8313 15336 8341
rect 5979 8252 6035 8261
rect 2758 8212 2814 8221
rect 2758 8147 2814 8156
rect 1714 8082 1800 8134
rect 1852 8082 1938 8134
rect 1714 7798 1938 8082
rect 1714 7746 1800 7798
rect 1852 7746 1938 7798
rect 1714 7462 1938 7746
rect 1714 7410 1800 7462
rect 1852 7410 1938 7462
rect 1714 7128 1938 7410
rect 1714 7072 1798 7128
rect 1854 7072 1938 7128
rect 1714 6790 1938 7072
rect 1714 6738 1800 6790
rect 1852 6738 1938 6790
rect 1714 6454 1938 6738
rect 1714 6402 1800 6454
rect 1852 6402 1938 6454
rect 1714 6118 1938 6402
rect 1714 6066 1800 6118
rect 1852 6066 1938 6118
rect 1714 5782 1938 6066
rect 1714 5730 1800 5782
rect 1852 5730 1938 5782
rect 1714 5448 1938 5730
rect 1714 5392 1798 5448
rect 1854 5392 1938 5448
rect 1714 5110 1938 5392
rect 1714 5058 1800 5110
rect 1852 5058 1938 5110
rect 1714 4774 1938 5058
rect 1714 4722 1800 4774
rect 1852 4722 1938 4774
rect 1714 4438 1938 4722
rect 1714 4386 1800 4438
rect 1852 4386 1938 4438
rect 1714 4102 1938 4386
rect 1714 4050 1800 4102
rect 1852 4050 1938 4102
rect 1714 3768 1938 4050
rect 1714 3712 1798 3768
rect 1854 3712 1938 3768
rect 1714 3430 1938 3712
rect 1714 3378 1800 3430
rect 1852 3378 1938 3430
rect 1714 3094 1938 3378
rect 1714 3042 1800 3094
rect 1852 3042 1938 3094
rect 1714 2758 1938 3042
rect 1714 2706 1800 2758
rect 1852 2706 1938 2758
rect 15308 2741 15336 8313
rect 136860 8808 137084 9090
rect 136860 8752 136944 8808
rect 137000 8752 137084 8808
rect 136860 8470 137084 8752
rect 136860 8418 136946 8470
rect 136998 8418 137084 8470
rect 136860 8134 137084 8418
rect 136860 8082 136946 8134
rect 136998 8082 137084 8134
rect 136860 7798 137084 8082
rect 136860 7746 136946 7798
rect 136998 7746 137084 7798
rect 136860 7462 137084 7746
rect 136860 7410 136946 7462
rect 136998 7410 137084 7462
rect 136860 7128 137084 7410
rect 136860 7072 136944 7128
rect 137000 7072 137084 7128
rect 136860 6790 137084 7072
rect 136860 6738 136946 6790
rect 136998 6738 137084 6790
rect 136860 6454 137084 6738
rect 136860 6402 136946 6454
rect 136998 6402 137084 6454
rect 136860 6118 137084 6402
rect 136860 6066 136946 6118
rect 136998 6066 137084 6118
rect 136860 5782 137084 6066
rect 136860 5730 136946 5782
rect 136998 5730 137084 5782
rect 136860 5448 137084 5730
rect 136860 5392 136944 5448
rect 137000 5392 137084 5448
rect 136860 5110 137084 5392
rect 136860 5058 136946 5110
rect 136998 5058 137084 5110
rect 136860 4774 137084 5058
rect 136860 4722 136946 4774
rect 136998 4722 137084 4774
rect 136860 4438 137084 4722
rect 136860 4386 136946 4438
rect 136998 4386 137084 4438
rect 136860 4102 137084 4386
rect 136860 4050 136946 4102
rect 136998 4050 137084 4102
rect 136860 3768 137084 4050
rect 136860 3712 136944 3768
rect 137000 3712 137084 3768
rect 136860 3430 137084 3712
rect 136860 3378 136946 3430
rect 136998 3378 137084 3430
rect 136860 3094 137084 3378
rect 136860 3042 136946 3094
rect 136998 3042 137084 3094
rect 16548 2988 16604 2997
rect 16548 2923 16604 2932
rect 17716 2988 17772 2997
rect 17716 2923 17772 2932
rect 18884 2988 18940 2997
rect 18884 2923 18940 2932
rect 20052 2988 20108 2997
rect 20052 2923 20108 2932
rect 21220 2988 21276 2997
rect 21220 2923 21276 2932
rect 22388 2988 22444 2997
rect 22388 2923 22444 2932
rect 23556 2988 23612 2997
rect 23556 2923 23612 2932
rect 24724 2988 24780 2997
rect 24724 2923 24780 2932
rect 25892 2988 25948 2997
rect 25892 2923 25948 2932
rect 27060 2988 27116 2997
rect 27060 2923 27116 2932
rect 28228 2988 28284 2997
rect 28228 2923 28284 2932
rect 29396 2988 29452 2997
rect 29396 2923 29452 2932
rect 30564 2988 30620 2997
rect 30564 2923 30620 2932
rect 31732 2988 31788 2997
rect 31732 2923 31788 2932
rect 32900 2988 32956 2997
rect 32900 2923 32956 2932
rect 34068 2988 34124 2997
rect 34068 2923 34124 2932
rect 35236 2988 35292 2997
rect 35236 2923 35292 2932
rect 36404 2988 36460 2997
rect 36404 2923 36460 2932
rect 37572 2988 37628 2997
rect 37572 2923 37628 2932
rect 38740 2988 38796 2997
rect 38740 2923 38796 2932
rect 39908 2988 39964 2997
rect 39908 2923 39964 2932
rect 41076 2988 41132 2997
rect 41076 2923 41132 2932
rect 42244 2988 42300 2997
rect 42244 2923 42300 2932
rect 43412 2988 43468 2997
rect 43412 2923 43468 2932
rect 44580 2988 44636 2997
rect 44580 2923 44636 2932
rect 45748 2988 45804 2997
rect 45748 2923 45804 2932
rect 46916 2988 46972 2997
rect 46916 2923 46972 2932
rect 48084 2988 48140 2997
rect 48084 2923 48140 2932
rect 49252 2988 49308 2997
rect 49252 2923 49308 2932
rect 50420 2988 50476 2997
rect 50420 2923 50476 2932
rect 51588 2988 51644 2997
rect 51588 2923 51644 2932
rect 52756 2988 52812 2997
rect 52756 2923 52812 2932
rect 53924 2988 53980 2997
rect 53924 2923 53980 2932
rect 55092 2988 55148 2997
rect 55092 2923 55148 2932
rect 56260 2988 56316 2997
rect 56260 2923 56316 2932
rect 57428 2988 57484 2997
rect 57428 2923 57484 2932
rect 58596 2988 58652 2997
rect 58596 2923 58652 2932
rect 59764 2988 59820 2997
rect 59764 2923 59820 2932
rect 136860 2758 137084 3042
rect 1714 2422 1938 2706
rect 15294 2732 15350 2741
rect 15294 2667 15350 2676
rect 136860 2706 136946 2758
rect 136998 2706 137084 2758
rect 1714 2370 1800 2422
rect 1852 2370 1938 2422
rect 1714 2088 1938 2370
rect 1714 2032 1798 2088
rect 1854 2032 1938 2088
rect 1714 1612 1938 2032
rect 136860 2422 137084 2706
rect 136860 2370 136946 2422
rect 136998 2370 137084 2422
rect 136860 2088 137084 2370
rect 136860 2032 136944 2088
rect 137000 2032 137084 2088
rect 2134 1752 2190 1761
rect 2134 1687 2190 1696
rect 3814 1752 3870 1761
rect 3814 1687 3870 1696
rect 5494 1752 5550 1761
rect 5494 1687 5550 1696
rect 7174 1752 7230 1761
rect 7174 1687 7230 1696
rect 8854 1752 8910 1761
rect 8854 1687 8910 1696
rect 10534 1752 10590 1761
rect 10534 1687 10590 1696
rect 12214 1752 12270 1761
rect 12214 1687 12270 1696
rect 13894 1752 13950 1761
rect 13894 1687 13950 1696
rect 15574 1752 15630 1761
rect 15574 1687 15630 1696
rect 17254 1752 17310 1761
rect 17254 1687 17310 1696
rect 18934 1752 18990 1761
rect 18934 1687 18990 1696
rect 20614 1752 20670 1761
rect 20614 1687 20670 1696
rect 22294 1752 22350 1761
rect 22294 1687 22350 1696
rect 23974 1752 24030 1761
rect 23974 1687 24030 1696
rect 25654 1752 25710 1761
rect 25654 1687 25710 1696
rect 27334 1752 27390 1761
rect 27334 1687 27390 1696
rect 29014 1752 29070 1761
rect 29014 1687 29070 1696
rect 30694 1752 30750 1761
rect 30694 1687 30750 1696
rect 32374 1752 32430 1761
rect 32374 1687 32430 1696
rect 34054 1752 34110 1761
rect 34054 1687 34110 1696
rect 35734 1752 35790 1761
rect 35734 1687 35790 1696
rect 37414 1752 37470 1761
rect 37414 1687 37470 1696
rect 39094 1752 39150 1761
rect 39094 1687 39150 1696
rect 40774 1752 40830 1761
rect 40774 1687 40830 1696
rect 42454 1752 42510 1761
rect 42454 1687 42510 1696
rect 44134 1752 44190 1761
rect 44134 1687 44190 1696
rect 45814 1752 45870 1761
rect 45814 1687 45870 1696
rect 47494 1752 47550 1761
rect 47494 1687 47550 1696
rect 49174 1752 49230 1761
rect 49174 1687 49230 1696
rect 50854 1752 50910 1761
rect 50854 1687 50910 1696
rect 52534 1752 52590 1761
rect 52534 1687 52590 1696
rect 54214 1752 54270 1761
rect 54214 1687 54270 1696
rect 55894 1752 55950 1761
rect 55894 1687 55950 1696
rect 57574 1752 57630 1761
rect 57574 1687 57630 1696
rect 59254 1752 59310 1761
rect 59254 1687 59310 1696
rect 60934 1752 60990 1761
rect 60934 1687 60990 1696
rect 62614 1752 62670 1761
rect 62614 1687 62670 1696
rect 64294 1752 64350 1761
rect 64294 1687 64350 1696
rect 65974 1752 66030 1761
rect 65974 1687 66030 1696
rect 67654 1752 67710 1761
rect 67654 1687 67710 1696
rect 69334 1752 69390 1761
rect 69334 1687 69390 1696
rect 71014 1752 71070 1761
rect 71014 1687 71070 1696
rect 72694 1752 72750 1761
rect 72694 1687 72750 1696
rect 74374 1752 74430 1761
rect 74374 1687 74430 1696
rect 76054 1752 76110 1761
rect 76054 1687 76110 1696
rect 77734 1752 77790 1761
rect 77734 1687 77790 1696
rect 79414 1752 79470 1761
rect 79414 1687 79470 1696
rect 81094 1752 81150 1761
rect 81094 1687 81150 1696
rect 82774 1752 82830 1761
rect 82774 1687 82830 1696
rect 84454 1752 84510 1761
rect 84454 1687 84510 1696
rect 86134 1752 86190 1761
rect 86134 1687 86190 1696
rect 87814 1752 87870 1761
rect 87814 1687 87870 1696
rect 89494 1752 89550 1761
rect 89494 1687 89550 1696
rect 91174 1752 91230 1761
rect 91174 1687 91230 1696
rect 92854 1752 92910 1761
rect 92854 1687 92910 1696
rect 94534 1752 94590 1761
rect 94534 1687 94590 1696
rect 96214 1752 96270 1761
rect 96214 1687 96270 1696
rect 97894 1752 97950 1761
rect 97894 1687 97950 1696
rect 99574 1752 99630 1761
rect 99574 1687 99630 1696
rect 101254 1752 101310 1761
rect 101254 1687 101310 1696
rect 102934 1752 102990 1761
rect 102934 1687 102990 1696
rect 104614 1752 104670 1761
rect 104614 1687 104670 1696
rect 106294 1752 106350 1761
rect 106294 1687 106350 1696
rect 107974 1752 108030 1761
rect 107974 1687 108030 1696
rect 109654 1752 109710 1761
rect 109654 1687 109710 1696
rect 111334 1752 111390 1761
rect 111334 1687 111390 1696
rect 113014 1752 113070 1761
rect 113014 1687 113070 1696
rect 114694 1752 114750 1761
rect 114694 1687 114750 1696
rect 116374 1752 116430 1761
rect 116374 1687 116430 1696
rect 118054 1752 118110 1761
rect 118054 1687 118110 1696
rect 119734 1752 119790 1761
rect 119734 1687 119790 1696
rect 121414 1752 121470 1761
rect 121414 1687 121470 1696
rect 123094 1752 123150 1761
rect 123094 1687 123150 1696
rect 124774 1752 124830 1761
rect 124774 1687 124830 1696
rect 126454 1752 126510 1761
rect 126454 1687 126510 1696
rect 128134 1752 128190 1761
rect 128134 1687 128190 1696
rect 129814 1752 129870 1761
rect 129814 1687 129870 1696
rect 131494 1752 131550 1761
rect 131494 1687 131550 1696
rect 133174 1752 133230 1761
rect 133174 1687 133230 1696
rect 134854 1752 134910 1761
rect 134854 1687 134910 1696
rect 136534 1752 136590 1761
rect 136534 1687 136590 1696
rect 136860 1612 137084 2032
<< via2 >>
rect 2134 132059 2190 132061
rect 2134 132007 2136 132059
rect 2136 132007 2188 132059
rect 2188 132007 2190 132059
rect 2134 132005 2190 132007
rect 3814 132059 3870 132061
rect 3814 132007 3816 132059
rect 3816 132007 3868 132059
rect 3868 132007 3870 132059
rect 3814 132005 3870 132007
rect 5494 132059 5550 132061
rect 5494 132007 5496 132059
rect 5496 132007 5548 132059
rect 5548 132007 5550 132059
rect 5494 132005 5550 132007
rect 7174 132059 7230 132061
rect 7174 132007 7176 132059
rect 7176 132007 7228 132059
rect 7228 132007 7230 132059
rect 7174 132005 7230 132007
rect 8854 132059 8910 132061
rect 8854 132007 8856 132059
rect 8856 132007 8908 132059
rect 8908 132007 8910 132059
rect 8854 132005 8910 132007
rect 10534 132059 10590 132061
rect 10534 132007 10536 132059
rect 10536 132007 10588 132059
rect 10588 132007 10590 132059
rect 10534 132005 10590 132007
rect 12214 132059 12270 132061
rect 12214 132007 12216 132059
rect 12216 132007 12268 132059
rect 12268 132007 12270 132059
rect 12214 132005 12270 132007
rect 13894 132059 13950 132061
rect 13894 132007 13896 132059
rect 13896 132007 13948 132059
rect 13948 132007 13950 132059
rect 13894 132005 13950 132007
rect 15574 132059 15630 132061
rect 15574 132007 15576 132059
rect 15576 132007 15628 132059
rect 15628 132007 15630 132059
rect 15574 132005 15630 132007
rect 17254 132059 17310 132061
rect 17254 132007 17256 132059
rect 17256 132007 17308 132059
rect 17308 132007 17310 132059
rect 17254 132005 17310 132007
rect 18934 132059 18990 132061
rect 18934 132007 18936 132059
rect 18936 132007 18988 132059
rect 18988 132007 18990 132059
rect 18934 132005 18990 132007
rect 20614 132059 20670 132061
rect 20614 132007 20616 132059
rect 20616 132007 20668 132059
rect 20668 132007 20670 132059
rect 20614 132005 20670 132007
rect 22294 132059 22350 132061
rect 22294 132007 22296 132059
rect 22296 132007 22348 132059
rect 22348 132007 22350 132059
rect 22294 132005 22350 132007
rect 23974 132059 24030 132061
rect 23974 132007 23976 132059
rect 23976 132007 24028 132059
rect 24028 132007 24030 132059
rect 23974 132005 24030 132007
rect 25654 132059 25710 132061
rect 25654 132007 25656 132059
rect 25656 132007 25708 132059
rect 25708 132007 25710 132059
rect 25654 132005 25710 132007
rect 27334 132059 27390 132061
rect 27334 132007 27336 132059
rect 27336 132007 27388 132059
rect 27388 132007 27390 132059
rect 27334 132005 27390 132007
rect 29014 132059 29070 132061
rect 29014 132007 29016 132059
rect 29016 132007 29068 132059
rect 29068 132007 29070 132059
rect 29014 132005 29070 132007
rect 30694 132059 30750 132061
rect 30694 132007 30696 132059
rect 30696 132007 30748 132059
rect 30748 132007 30750 132059
rect 30694 132005 30750 132007
rect 32374 132059 32430 132061
rect 32374 132007 32376 132059
rect 32376 132007 32428 132059
rect 32428 132007 32430 132059
rect 32374 132005 32430 132007
rect 34054 132059 34110 132061
rect 34054 132007 34056 132059
rect 34056 132007 34108 132059
rect 34108 132007 34110 132059
rect 34054 132005 34110 132007
rect 35734 132059 35790 132061
rect 35734 132007 35736 132059
rect 35736 132007 35788 132059
rect 35788 132007 35790 132059
rect 35734 132005 35790 132007
rect 37414 132059 37470 132061
rect 37414 132007 37416 132059
rect 37416 132007 37468 132059
rect 37468 132007 37470 132059
rect 37414 132005 37470 132007
rect 39094 132059 39150 132061
rect 39094 132007 39096 132059
rect 39096 132007 39148 132059
rect 39148 132007 39150 132059
rect 39094 132005 39150 132007
rect 40774 132059 40830 132061
rect 40774 132007 40776 132059
rect 40776 132007 40828 132059
rect 40828 132007 40830 132059
rect 40774 132005 40830 132007
rect 42454 132059 42510 132061
rect 42454 132007 42456 132059
rect 42456 132007 42508 132059
rect 42508 132007 42510 132059
rect 42454 132005 42510 132007
rect 44134 132059 44190 132061
rect 44134 132007 44136 132059
rect 44136 132007 44188 132059
rect 44188 132007 44190 132059
rect 44134 132005 44190 132007
rect 45814 132059 45870 132061
rect 45814 132007 45816 132059
rect 45816 132007 45868 132059
rect 45868 132007 45870 132059
rect 45814 132005 45870 132007
rect 47494 132059 47550 132061
rect 47494 132007 47496 132059
rect 47496 132007 47548 132059
rect 47548 132007 47550 132059
rect 47494 132005 47550 132007
rect 49174 132059 49230 132061
rect 49174 132007 49176 132059
rect 49176 132007 49228 132059
rect 49228 132007 49230 132059
rect 49174 132005 49230 132007
rect 50854 132059 50910 132061
rect 50854 132007 50856 132059
rect 50856 132007 50908 132059
rect 50908 132007 50910 132059
rect 50854 132005 50910 132007
rect 52534 132059 52590 132061
rect 52534 132007 52536 132059
rect 52536 132007 52588 132059
rect 52588 132007 52590 132059
rect 52534 132005 52590 132007
rect 54214 132059 54270 132061
rect 54214 132007 54216 132059
rect 54216 132007 54268 132059
rect 54268 132007 54270 132059
rect 54214 132005 54270 132007
rect 55894 132059 55950 132061
rect 55894 132007 55896 132059
rect 55896 132007 55948 132059
rect 55948 132007 55950 132059
rect 55894 132005 55950 132007
rect 57574 132059 57630 132061
rect 57574 132007 57576 132059
rect 57576 132007 57628 132059
rect 57628 132007 57630 132059
rect 57574 132005 57630 132007
rect 59254 132059 59310 132061
rect 59254 132007 59256 132059
rect 59256 132007 59308 132059
rect 59308 132007 59310 132059
rect 59254 132005 59310 132007
rect 60934 132059 60990 132061
rect 60934 132007 60936 132059
rect 60936 132007 60988 132059
rect 60988 132007 60990 132059
rect 60934 132005 60990 132007
rect 62614 132059 62670 132061
rect 62614 132007 62616 132059
rect 62616 132007 62668 132059
rect 62668 132007 62670 132059
rect 62614 132005 62670 132007
rect 64294 132059 64350 132061
rect 64294 132007 64296 132059
rect 64296 132007 64348 132059
rect 64348 132007 64350 132059
rect 64294 132005 64350 132007
rect 65974 132059 66030 132061
rect 65974 132007 65976 132059
rect 65976 132007 66028 132059
rect 66028 132007 66030 132059
rect 65974 132005 66030 132007
rect 67654 132059 67710 132061
rect 67654 132007 67656 132059
rect 67656 132007 67708 132059
rect 67708 132007 67710 132059
rect 67654 132005 67710 132007
rect 69334 132059 69390 132061
rect 69334 132007 69336 132059
rect 69336 132007 69388 132059
rect 69388 132007 69390 132059
rect 69334 132005 69390 132007
rect 71014 132059 71070 132061
rect 71014 132007 71016 132059
rect 71016 132007 71068 132059
rect 71068 132007 71070 132059
rect 71014 132005 71070 132007
rect 72694 132059 72750 132061
rect 72694 132007 72696 132059
rect 72696 132007 72748 132059
rect 72748 132007 72750 132059
rect 72694 132005 72750 132007
rect 74374 132059 74430 132061
rect 74374 132007 74376 132059
rect 74376 132007 74428 132059
rect 74428 132007 74430 132059
rect 74374 132005 74430 132007
rect 76054 132059 76110 132061
rect 76054 132007 76056 132059
rect 76056 132007 76108 132059
rect 76108 132007 76110 132059
rect 76054 132005 76110 132007
rect 77734 132059 77790 132061
rect 77734 132007 77736 132059
rect 77736 132007 77788 132059
rect 77788 132007 77790 132059
rect 77734 132005 77790 132007
rect 79414 132059 79470 132061
rect 79414 132007 79416 132059
rect 79416 132007 79468 132059
rect 79468 132007 79470 132059
rect 79414 132005 79470 132007
rect 81094 132059 81150 132061
rect 81094 132007 81096 132059
rect 81096 132007 81148 132059
rect 81148 132007 81150 132059
rect 81094 132005 81150 132007
rect 82774 132059 82830 132061
rect 82774 132007 82776 132059
rect 82776 132007 82828 132059
rect 82828 132007 82830 132059
rect 82774 132005 82830 132007
rect 84454 132059 84510 132061
rect 84454 132007 84456 132059
rect 84456 132007 84508 132059
rect 84508 132007 84510 132059
rect 84454 132005 84510 132007
rect 86134 132059 86190 132061
rect 86134 132007 86136 132059
rect 86136 132007 86188 132059
rect 86188 132007 86190 132059
rect 86134 132005 86190 132007
rect 87814 132059 87870 132061
rect 87814 132007 87816 132059
rect 87816 132007 87868 132059
rect 87868 132007 87870 132059
rect 87814 132005 87870 132007
rect 89494 132059 89550 132061
rect 89494 132007 89496 132059
rect 89496 132007 89548 132059
rect 89548 132007 89550 132059
rect 89494 132005 89550 132007
rect 91174 132059 91230 132061
rect 91174 132007 91176 132059
rect 91176 132007 91228 132059
rect 91228 132007 91230 132059
rect 91174 132005 91230 132007
rect 92854 132059 92910 132061
rect 92854 132007 92856 132059
rect 92856 132007 92908 132059
rect 92908 132007 92910 132059
rect 92854 132005 92910 132007
rect 94534 132059 94590 132061
rect 94534 132007 94536 132059
rect 94536 132007 94588 132059
rect 94588 132007 94590 132059
rect 94534 132005 94590 132007
rect 96214 132059 96270 132061
rect 96214 132007 96216 132059
rect 96216 132007 96268 132059
rect 96268 132007 96270 132059
rect 96214 132005 96270 132007
rect 97894 132059 97950 132061
rect 97894 132007 97896 132059
rect 97896 132007 97948 132059
rect 97948 132007 97950 132059
rect 97894 132005 97950 132007
rect 99574 132059 99630 132061
rect 99574 132007 99576 132059
rect 99576 132007 99628 132059
rect 99628 132007 99630 132059
rect 99574 132005 99630 132007
rect 101254 132059 101310 132061
rect 101254 132007 101256 132059
rect 101256 132007 101308 132059
rect 101308 132007 101310 132059
rect 101254 132005 101310 132007
rect 102934 132059 102990 132061
rect 102934 132007 102936 132059
rect 102936 132007 102988 132059
rect 102988 132007 102990 132059
rect 102934 132005 102990 132007
rect 104614 132059 104670 132061
rect 104614 132007 104616 132059
rect 104616 132007 104668 132059
rect 104668 132007 104670 132059
rect 104614 132005 104670 132007
rect 106294 132059 106350 132061
rect 106294 132007 106296 132059
rect 106296 132007 106348 132059
rect 106348 132007 106350 132059
rect 106294 132005 106350 132007
rect 107974 132059 108030 132061
rect 107974 132007 107976 132059
rect 107976 132007 108028 132059
rect 108028 132007 108030 132059
rect 107974 132005 108030 132007
rect 109654 132059 109710 132061
rect 109654 132007 109656 132059
rect 109656 132007 109708 132059
rect 109708 132007 109710 132059
rect 109654 132005 109710 132007
rect 111334 132059 111390 132061
rect 111334 132007 111336 132059
rect 111336 132007 111388 132059
rect 111388 132007 111390 132059
rect 111334 132005 111390 132007
rect 113014 132059 113070 132061
rect 113014 132007 113016 132059
rect 113016 132007 113068 132059
rect 113068 132007 113070 132059
rect 113014 132005 113070 132007
rect 114694 132059 114750 132061
rect 114694 132007 114696 132059
rect 114696 132007 114748 132059
rect 114748 132007 114750 132059
rect 114694 132005 114750 132007
rect 116374 132059 116430 132061
rect 116374 132007 116376 132059
rect 116376 132007 116428 132059
rect 116428 132007 116430 132059
rect 116374 132005 116430 132007
rect 118054 132059 118110 132061
rect 118054 132007 118056 132059
rect 118056 132007 118108 132059
rect 118108 132007 118110 132059
rect 118054 132005 118110 132007
rect 119734 132059 119790 132061
rect 119734 132007 119736 132059
rect 119736 132007 119788 132059
rect 119788 132007 119790 132059
rect 119734 132005 119790 132007
rect 121414 132059 121470 132061
rect 121414 132007 121416 132059
rect 121416 132007 121468 132059
rect 121468 132007 121470 132059
rect 121414 132005 121470 132007
rect 123094 132059 123150 132061
rect 123094 132007 123096 132059
rect 123096 132007 123148 132059
rect 123148 132007 123150 132059
rect 123094 132005 123150 132007
rect 124774 132059 124830 132061
rect 124774 132007 124776 132059
rect 124776 132007 124828 132059
rect 124828 132007 124830 132059
rect 124774 132005 124830 132007
rect 126454 132059 126510 132061
rect 126454 132007 126456 132059
rect 126456 132007 126508 132059
rect 126508 132007 126510 132059
rect 126454 132005 126510 132007
rect 128134 132059 128190 132061
rect 128134 132007 128136 132059
rect 128136 132007 128188 132059
rect 128188 132007 128190 132059
rect 128134 132005 128190 132007
rect 129814 132059 129870 132061
rect 129814 132007 129816 132059
rect 129816 132007 129868 132059
rect 129868 132007 129870 132059
rect 129814 132005 129870 132007
rect 131494 132059 131550 132061
rect 131494 132007 131496 132059
rect 131496 132007 131548 132059
rect 131548 132007 131550 132059
rect 131494 132005 131550 132007
rect 133174 132059 133230 132061
rect 133174 132007 133176 132059
rect 133176 132007 133228 132059
rect 133228 132007 133230 132059
rect 133174 132005 133230 132007
rect 134854 132059 134910 132061
rect 134854 132007 134856 132059
rect 134856 132007 134908 132059
rect 134908 132007 134910 132059
rect 134854 132005 134910 132007
rect 136534 132059 136590 132061
rect 136534 132007 136536 132059
rect 136536 132007 136588 132059
rect 136588 132007 136590 132059
rect 136534 132005 136590 132007
rect 1798 131446 1854 131448
rect 1798 131394 1800 131446
rect 1800 131394 1852 131446
rect 1852 131394 1854 131446
rect 1798 131392 1854 131394
rect 136944 131446 137000 131448
rect 136944 131394 136946 131446
rect 136946 131394 136998 131446
rect 136998 131394 137000 131446
rect 136944 131392 137000 131394
rect 123532 131025 123588 131081
rect 119942 130769 119998 130825
rect 121110 130769 121166 130825
rect 1798 129766 1854 129768
rect 1798 129714 1800 129766
rect 1800 129714 1852 129766
rect 1852 129714 1854 129766
rect 1798 129712 1854 129714
rect 1798 128086 1854 128088
rect 1798 128034 1800 128086
rect 1800 128034 1852 128086
rect 1852 128034 1854 128086
rect 1798 128032 1854 128034
rect 135984 129772 136040 129828
rect 132847 129667 132903 129723
rect 136944 129766 137000 129768
rect 136944 129714 136946 129766
rect 136946 129714 136998 129766
rect 136998 129714 137000 129766
rect 136944 129712 137000 129714
rect 29562 127605 29618 127607
rect 29562 127553 29564 127605
rect 29564 127553 29616 127605
rect 29616 127553 29618 127605
rect 29562 127551 29618 127553
rect 32058 127605 32114 127607
rect 32058 127553 32060 127605
rect 32060 127553 32112 127605
rect 32112 127553 32114 127605
rect 32058 127551 32114 127553
rect 34554 127605 34610 127607
rect 34554 127553 34556 127605
rect 34556 127553 34608 127605
rect 34608 127553 34610 127605
rect 34554 127551 34610 127553
rect 37050 127605 37106 127607
rect 37050 127553 37052 127605
rect 37052 127553 37104 127605
rect 37104 127553 37106 127605
rect 37050 127551 37106 127553
rect 39546 127605 39602 127607
rect 39546 127553 39548 127605
rect 39548 127553 39600 127605
rect 39600 127553 39602 127605
rect 39546 127551 39602 127553
rect 42042 127605 42098 127607
rect 42042 127553 42044 127605
rect 42044 127553 42096 127605
rect 42096 127553 42098 127605
rect 42042 127551 42098 127553
rect 44538 127605 44594 127607
rect 44538 127553 44540 127605
rect 44540 127553 44592 127605
rect 44592 127553 44594 127605
rect 44538 127551 44594 127553
rect 47034 127605 47090 127607
rect 47034 127553 47036 127605
rect 47036 127553 47088 127605
rect 47088 127553 47090 127605
rect 47034 127551 47090 127553
rect 49530 127605 49586 127607
rect 49530 127553 49532 127605
rect 49532 127553 49584 127605
rect 49584 127553 49586 127605
rect 49530 127551 49586 127553
rect 52026 127605 52082 127607
rect 52026 127553 52028 127605
rect 52028 127553 52080 127605
rect 52080 127553 52082 127605
rect 52026 127551 52082 127553
rect 54522 127605 54578 127607
rect 54522 127553 54524 127605
rect 54524 127553 54576 127605
rect 54576 127553 54578 127605
rect 54522 127551 54578 127553
rect 57018 127605 57074 127607
rect 57018 127553 57020 127605
rect 57020 127553 57072 127605
rect 57072 127553 57074 127605
rect 57018 127551 57074 127553
rect 59514 127605 59570 127607
rect 59514 127553 59516 127605
rect 59516 127553 59568 127605
rect 59568 127553 59570 127605
rect 59514 127551 59570 127553
rect 62010 127605 62066 127607
rect 62010 127553 62012 127605
rect 62012 127553 62064 127605
rect 62064 127553 62066 127605
rect 62010 127551 62066 127553
rect 64506 127605 64562 127607
rect 64506 127553 64508 127605
rect 64508 127553 64560 127605
rect 64560 127553 64562 127605
rect 64506 127551 64562 127553
rect 67002 127605 67058 127607
rect 67002 127553 67004 127605
rect 67004 127553 67056 127605
rect 67056 127553 67058 127605
rect 67002 127551 67058 127553
rect 69498 127605 69554 127607
rect 69498 127553 69500 127605
rect 69500 127553 69552 127605
rect 69552 127553 69554 127605
rect 69498 127551 69554 127553
rect 71994 127605 72050 127607
rect 71994 127553 71996 127605
rect 71996 127553 72048 127605
rect 72048 127553 72050 127605
rect 71994 127551 72050 127553
rect 74490 127605 74546 127607
rect 74490 127553 74492 127605
rect 74492 127553 74544 127605
rect 74544 127553 74546 127605
rect 74490 127551 74546 127553
rect 76986 127605 77042 127607
rect 76986 127553 76988 127605
rect 76988 127553 77040 127605
rect 77040 127553 77042 127605
rect 76986 127551 77042 127553
rect 79482 127605 79538 127607
rect 79482 127553 79484 127605
rect 79484 127553 79536 127605
rect 79536 127553 79538 127605
rect 79482 127551 79538 127553
rect 81978 127605 82034 127607
rect 81978 127553 81980 127605
rect 81980 127553 82032 127605
rect 82032 127553 82034 127605
rect 81978 127551 82034 127553
rect 84474 127605 84530 127607
rect 84474 127553 84476 127605
rect 84476 127553 84528 127605
rect 84528 127553 84530 127605
rect 84474 127551 84530 127553
rect 86970 127605 87026 127607
rect 86970 127553 86972 127605
rect 86972 127553 87024 127605
rect 87024 127553 87026 127605
rect 86970 127551 87026 127553
rect 89466 127605 89522 127607
rect 89466 127553 89468 127605
rect 89468 127553 89520 127605
rect 89520 127553 89522 127605
rect 89466 127551 89522 127553
rect 91962 127605 92018 127607
rect 91962 127553 91964 127605
rect 91964 127553 92016 127605
rect 92016 127553 92018 127605
rect 91962 127551 92018 127553
rect 94458 127605 94514 127607
rect 94458 127553 94460 127605
rect 94460 127553 94512 127605
rect 94512 127553 94514 127605
rect 94458 127551 94514 127553
rect 96954 127605 97010 127607
rect 96954 127553 96956 127605
rect 96956 127553 97008 127605
rect 97008 127553 97010 127605
rect 96954 127551 97010 127553
rect 99450 127605 99506 127607
rect 99450 127553 99452 127605
rect 99452 127553 99504 127605
rect 99504 127553 99506 127605
rect 99450 127551 99506 127553
rect 101946 127605 102002 127607
rect 101946 127553 101948 127605
rect 101948 127553 102000 127605
rect 102000 127553 102002 127605
rect 101946 127551 102002 127553
rect 104442 127605 104498 127607
rect 104442 127553 104444 127605
rect 104444 127553 104496 127605
rect 104496 127553 104498 127605
rect 104442 127551 104498 127553
rect 106938 127605 106994 127607
rect 106938 127553 106940 127605
rect 106940 127553 106992 127605
rect 106992 127553 106994 127605
rect 106938 127551 106994 127553
rect 1798 126406 1854 126408
rect 1798 126354 1800 126406
rect 1800 126354 1852 126406
rect 1852 126354 1854 126406
rect 1798 126352 1854 126354
rect 111005 125387 111061 125443
rect 1798 124726 1854 124728
rect 1798 124674 1800 124726
rect 1800 124674 1852 124726
rect 1852 124674 1854 124726
rect 1798 124672 1854 124674
rect 1798 123046 1854 123048
rect 1798 122994 1800 123046
rect 1800 122994 1852 123046
rect 1852 122994 1854 123046
rect 1798 122992 1854 122994
rect 111129 123973 111185 124029
rect 114990 122559 115046 122615
rect 1798 121366 1854 121368
rect 1798 121314 1800 121366
rect 1800 121314 1852 121366
rect 1852 121314 1854 121366
rect 1798 121312 1854 121314
rect 1798 119686 1854 119688
rect 1798 119634 1800 119686
rect 1800 119634 1852 119686
rect 1852 119634 1854 119686
rect 1798 119632 1854 119634
rect 1798 118006 1854 118008
rect 1798 117954 1800 118006
rect 1800 117954 1852 118006
rect 1852 117954 1854 118006
rect 1798 117952 1854 117954
rect 1798 116326 1854 116328
rect 1798 116274 1800 116326
rect 1800 116274 1852 116326
rect 1852 116274 1854 116326
rect 1798 116272 1854 116274
rect 1798 114646 1854 114648
rect 1798 114594 1800 114646
rect 1800 114594 1852 114646
rect 1852 114594 1854 114646
rect 1798 114592 1854 114594
rect 1798 112966 1854 112968
rect 1798 112914 1800 112966
rect 1800 112914 1852 112966
rect 1852 112914 1854 112966
rect 1798 112912 1854 112914
rect 1798 111286 1854 111288
rect 1798 111234 1800 111286
rect 1800 111234 1852 111286
rect 1852 111234 1854 111286
rect 1798 111232 1854 111234
rect 1798 109606 1854 109608
rect 1798 109554 1800 109606
rect 1800 109554 1852 109606
rect 1852 109554 1854 109606
rect 1798 109552 1854 109554
rect 1798 107926 1854 107928
rect 1798 107874 1800 107926
rect 1800 107874 1852 107926
rect 1852 107874 1854 107926
rect 1798 107872 1854 107874
rect 1798 106246 1854 106248
rect 1798 106194 1800 106246
rect 1800 106194 1852 106246
rect 1852 106194 1854 106246
rect 1798 106192 1854 106194
rect 1798 104566 1854 104568
rect 1798 104514 1800 104566
rect 1800 104514 1852 104566
rect 1852 104514 1854 104566
rect 1798 104512 1854 104514
rect 1798 102886 1854 102888
rect 1798 102834 1800 102886
rect 1800 102834 1852 102886
rect 1852 102834 1854 102886
rect 1798 102832 1854 102834
rect 1798 101206 1854 101208
rect 1798 101154 1800 101206
rect 1800 101154 1852 101206
rect 1852 101154 1854 101206
rect 1798 101152 1854 101154
rect 1798 99526 1854 99528
rect 1798 99474 1800 99526
rect 1800 99474 1852 99526
rect 1852 99474 1854 99526
rect 1798 99472 1854 99474
rect 1798 97846 1854 97848
rect 1798 97794 1800 97846
rect 1800 97794 1852 97846
rect 1852 97794 1854 97846
rect 1798 97792 1854 97794
rect 1798 96166 1854 96168
rect 1798 96114 1800 96166
rect 1800 96114 1852 96166
rect 1852 96114 1854 96166
rect 1798 96112 1854 96114
rect 1798 94486 1854 94488
rect 1798 94434 1800 94486
rect 1800 94434 1852 94486
rect 1852 94434 1854 94486
rect 1798 94432 1854 94434
rect 1798 92806 1854 92808
rect 1798 92754 1800 92806
rect 1800 92754 1852 92806
rect 1852 92754 1854 92806
rect 1798 92752 1854 92754
rect 1798 91126 1854 91128
rect 1798 91074 1800 91126
rect 1800 91074 1852 91126
rect 1852 91074 1854 91126
rect 1798 91072 1854 91074
rect 1798 89446 1854 89448
rect 1798 89394 1800 89446
rect 1800 89394 1852 89446
rect 1852 89394 1854 89446
rect 1798 89392 1854 89394
rect 1798 87766 1854 87768
rect 1798 87714 1800 87766
rect 1800 87714 1852 87766
rect 1852 87714 1854 87766
rect 1798 87712 1854 87714
rect 1798 86086 1854 86088
rect 1798 86034 1800 86086
rect 1800 86034 1852 86086
rect 1852 86034 1854 86086
rect 1798 86032 1854 86034
rect 1798 84406 1854 84408
rect 1798 84354 1800 84406
rect 1800 84354 1852 84406
rect 1852 84354 1854 84406
rect 1798 84352 1854 84354
rect 1798 82726 1854 82728
rect 1798 82674 1800 82726
rect 1800 82674 1852 82726
rect 1852 82674 1854 82726
rect 1798 82672 1854 82674
rect 1798 81046 1854 81048
rect 1798 80994 1800 81046
rect 1800 80994 1852 81046
rect 1852 80994 1854 81046
rect 1798 80992 1854 80994
rect 1798 79366 1854 79368
rect 1798 79314 1800 79366
rect 1800 79314 1852 79366
rect 1852 79314 1854 79366
rect 1798 79312 1854 79314
rect 1798 77686 1854 77688
rect 1798 77634 1800 77686
rect 1800 77634 1852 77686
rect 1852 77634 1854 77686
rect 1798 77632 1854 77634
rect 1798 76006 1854 76008
rect 1798 75954 1800 76006
rect 1800 75954 1852 76006
rect 1852 75954 1854 76006
rect 1798 75952 1854 75954
rect 1798 74326 1854 74328
rect 1798 74274 1800 74326
rect 1800 74274 1852 74326
rect 1852 74274 1854 74326
rect 1798 74272 1854 74274
rect 1798 72646 1854 72648
rect 1798 72594 1800 72646
rect 1800 72594 1852 72646
rect 1852 72594 1854 72646
rect 1798 72592 1854 72594
rect 1798 70966 1854 70968
rect 1798 70914 1800 70966
rect 1800 70914 1852 70966
rect 1852 70914 1854 70966
rect 1798 70912 1854 70914
rect 1798 69286 1854 69288
rect 1798 69234 1800 69286
rect 1800 69234 1852 69286
rect 1852 69234 1854 69286
rect 1798 69232 1854 69234
rect 1798 67606 1854 67608
rect 1798 67554 1800 67606
rect 1800 67554 1852 67606
rect 1852 67554 1854 67606
rect 1798 67552 1854 67554
rect 1798 65926 1854 65928
rect 1798 65874 1800 65926
rect 1800 65874 1852 65926
rect 1852 65874 1854 65926
rect 1798 65872 1854 65874
rect 1798 64246 1854 64248
rect 1798 64194 1800 64246
rect 1800 64194 1852 64246
rect 1852 64194 1854 64246
rect 1798 64192 1854 64194
rect 1798 62566 1854 62568
rect 1798 62514 1800 62566
rect 1800 62514 1852 62566
rect 1852 62514 1854 62566
rect 1798 62512 1854 62514
rect 1798 60886 1854 60888
rect 1798 60834 1800 60886
rect 1800 60834 1852 60886
rect 1852 60834 1854 60886
rect 1798 60832 1854 60834
rect 1798 59206 1854 59208
rect 1798 59154 1800 59206
rect 1800 59154 1852 59206
rect 1852 59154 1854 59206
rect 1798 59152 1854 59154
rect 1798 57526 1854 57528
rect 1798 57474 1800 57526
rect 1800 57474 1852 57526
rect 1852 57474 1854 57526
rect 1798 57472 1854 57474
rect 1798 55846 1854 55848
rect 1798 55794 1800 55846
rect 1800 55794 1852 55846
rect 1852 55794 1854 55846
rect 1798 55792 1854 55794
rect 1798 54166 1854 54168
rect 1798 54114 1800 54166
rect 1800 54114 1852 54166
rect 1852 54114 1854 54166
rect 1798 54112 1854 54114
rect 1798 52486 1854 52488
rect 1798 52434 1800 52486
rect 1800 52434 1852 52486
rect 1852 52434 1854 52486
rect 1798 52432 1854 52434
rect 1798 50806 1854 50808
rect 1798 50754 1800 50806
rect 1800 50754 1852 50806
rect 1852 50754 1854 50806
rect 1798 50752 1854 50754
rect 1798 49126 1854 49128
rect 1798 49074 1800 49126
rect 1800 49074 1852 49126
rect 1852 49074 1854 49126
rect 1798 49072 1854 49074
rect 1798 47446 1854 47448
rect 1798 47394 1800 47446
rect 1800 47394 1852 47446
rect 1852 47394 1854 47446
rect 1798 47392 1854 47394
rect 1798 45766 1854 45768
rect 1798 45714 1800 45766
rect 1800 45714 1852 45766
rect 1852 45714 1854 45766
rect 1798 45712 1854 45714
rect 1798 44086 1854 44088
rect 1798 44034 1800 44086
rect 1800 44034 1852 44086
rect 1852 44034 1854 44086
rect 1798 44032 1854 44034
rect 1798 42406 1854 42408
rect 1798 42354 1800 42406
rect 1800 42354 1852 42406
rect 1852 42354 1854 42406
rect 1798 42352 1854 42354
rect 1798 40726 1854 40728
rect 1798 40674 1800 40726
rect 1800 40674 1852 40726
rect 1852 40674 1854 40726
rect 1798 40672 1854 40674
rect 14212 40046 14268 40102
rect 15157 39975 15213 40031
rect 15971 40029 16027 40031
rect 15971 39977 15973 40029
rect 15973 39977 16025 40029
rect 16025 39977 16027 40029
rect 15971 39975 16027 39977
rect 1798 39046 1854 39048
rect 1798 38994 1800 39046
rect 1800 38994 1852 39046
rect 1852 38994 1854 39046
rect 1798 38992 1854 38994
rect 15157 38417 15213 38473
rect 15891 38471 15947 38473
rect 15891 38419 15893 38471
rect 15893 38419 15945 38471
rect 15945 38419 15947 38471
rect 15891 38417 15947 38419
rect 14212 38346 14268 38402
rect 1798 37366 1854 37368
rect 1798 37314 1800 37366
rect 1800 37314 1852 37366
rect 1852 37314 1854 37366
rect 1798 37312 1854 37314
rect 14212 37218 14268 37274
rect 15157 37147 15213 37203
rect 15811 37201 15867 37203
rect 15811 37149 15813 37201
rect 15813 37149 15865 37201
rect 15865 37149 15867 37201
rect 15811 37147 15867 37149
rect 1798 35686 1854 35688
rect 1798 35634 1800 35686
rect 1800 35634 1852 35686
rect 1852 35634 1854 35686
rect 1798 35632 1854 35634
rect 15157 35589 15213 35645
rect 15731 35643 15787 35645
rect 15731 35591 15733 35643
rect 15733 35591 15785 35643
rect 15785 35591 15787 35643
rect 15731 35589 15787 35591
rect 14212 35518 14268 35574
rect 14212 34390 14268 34446
rect 15157 34319 15213 34375
rect 15651 34373 15707 34375
rect 15651 34321 15653 34373
rect 15653 34321 15705 34373
rect 15705 34321 15707 34373
rect 15651 34319 15707 34321
rect 1798 34006 1854 34008
rect 1798 33954 1800 34006
rect 1800 33954 1852 34006
rect 1852 33954 1854 34006
rect 1798 33952 1854 33954
rect 15157 32761 15213 32817
rect 15571 32815 15627 32817
rect 15571 32763 15573 32815
rect 15573 32763 15625 32815
rect 15625 32763 15627 32815
rect 15571 32761 15627 32763
rect 14212 32690 14268 32746
rect 1798 32326 1854 32328
rect 1798 32274 1800 32326
rect 1800 32274 1852 32326
rect 1852 32274 1854 32326
rect 1798 32272 1854 32274
rect 14212 31562 14268 31618
rect 15157 31491 15213 31547
rect 15491 31545 15547 31547
rect 15491 31493 15493 31545
rect 15493 31493 15545 31545
rect 15545 31493 15547 31545
rect 15491 31491 15547 31493
rect 1798 30646 1854 30648
rect 1798 30594 1800 30646
rect 1800 30594 1852 30646
rect 1852 30594 1854 30646
rect 1798 30592 1854 30594
rect 15157 29933 15213 29989
rect 15411 29987 15467 29989
rect 15411 29935 15413 29987
rect 15413 29935 15465 29987
rect 15465 29935 15467 29987
rect 15411 29933 15467 29935
rect 14212 29862 14268 29918
rect 15294 29606 15350 29662
rect 1798 28966 1854 28968
rect 1798 28914 1800 28966
rect 1800 28914 1852 28966
rect 1852 28914 1854 28966
rect 1798 28912 1854 28914
rect 1798 27286 1854 27288
rect 1798 27234 1800 27286
rect 1800 27234 1852 27286
rect 1852 27234 1854 27286
rect 1798 27232 1854 27234
rect 1798 25606 1854 25608
rect 1798 25554 1800 25606
rect 1800 25554 1852 25606
rect 1852 25554 1854 25606
rect 1798 25552 1854 25554
rect 2545 25305 2601 25361
rect 1798 23926 1854 23928
rect 1798 23874 1800 23926
rect 1800 23874 1852 23926
rect 1852 23874 1854 23926
rect 1798 23872 1854 23874
rect 1798 22246 1854 22248
rect 1798 22194 1800 22246
rect 1800 22194 1852 22246
rect 1852 22194 1854 22246
rect 1798 22192 1854 22194
rect 1798 20566 1854 20568
rect 1798 20514 1800 20566
rect 1800 20514 1852 20566
rect 1852 20514 1854 20566
rect 1798 20512 1854 20514
rect 1798 18886 1854 18888
rect 1798 18834 1800 18886
rect 1800 18834 1852 18886
rect 1852 18834 1854 18886
rect 1798 18832 1854 18834
rect 15210 18197 15266 18253
rect 1798 17206 1854 17208
rect 1798 17154 1800 17206
rect 1800 17154 1852 17206
rect 1852 17154 1854 17206
rect 1798 17152 1854 17154
rect 1798 15526 1854 15528
rect 1798 15474 1800 15526
rect 1800 15474 1852 15526
rect 1852 15474 1854 15526
rect 1798 15472 1854 15474
rect 15210 15369 15266 15425
rect 15210 13955 15266 14011
rect 1798 13846 1854 13848
rect 1798 13794 1800 13846
rect 1800 13794 1852 13846
rect 1852 13794 1854 13846
rect 1798 13792 1854 13794
rect 15210 12541 15266 12597
rect 1798 12166 1854 12168
rect 1798 12114 1800 12166
rect 1800 12114 1852 12166
rect 1852 12114 1854 12166
rect 1798 12112 1854 12114
rect 1798 10486 1854 10488
rect 1798 10434 1800 10486
rect 1800 10434 1852 10486
rect 1852 10434 1854 10486
rect 1798 10432 1854 10434
rect 2758 9856 2814 9912
rect 1798 8806 1854 8808
rect 1798 8754 1800 8806
rect 1800 8754 1852 8806
rect 1852 8754 1854 8806
rect 1798 8752 1854 8754
rect 136944 128086 137000 128088
rect 136944 128034 136946 128086
rect 136946 128034 136998 128086
rect 136998 128034 137000 128086
rect 136944 128032 137000 128034
rect 136944 126406 137000 126408
rect 136944 126354 136946 126406
rect 136946 126354 136998 126406
rect 136998 126354 137000 126406
rect 136944 126352 137000 126354
rect 123616 125387 123672 125443
rect 136944 124726 137000 124728
rect 136944 124674 136946 124726
rect 136946 124674 136998 124726
rect 136998 124674 137000 124726
rect 136944 124672 137000 124674
rect 123616 123973 123672 124029
rect 136944 123046 137000 123048
rect 136944 122994 136946 123046
rect 136946 122994 136998 123046
rect 136998 122994 137000 123046
rect 136944 122992 137000 122994
rect 123616 122559 123672 122615
rect 136944 121366 137000 121368
rect 136944 121314 136946 121366
rect 136946 121314 136998 121366
rect 136998 121314 137000 121366
rect 136944 121312 137000 121314
rect 136944 119686 137000 119688
rect 136944 119634 136946 119686
rect 136946 119634 136998 119686
rect 136998 119634 137000 119686
rect 136944 119632 137000 119634
rect 136944 118006 137000 118008
rect 136944 117954 136946 118006
rect 136946 117954 136998 118006
rect 136998 117954 137000 118006
rect 136944 117952 137000 117954
rect 136944 116326 137000 116328
rect 136944 116274 136946 116326
rect 136946 116274 136998 116326
rect 136998 116274 137000 116326
rect 136944 116272 137000 116274
rect 136944 114646 137000 114648
rect 136944 114594 136946 114646
rect 136946 114594 136998 114646
rect 136998 114594 137000 114646
rect 136944 114592 137000 114594
rect 136944 112966 137000 112968
rect 136944 112914 136946 112966
rect 136946 112914 136998 112966
rect 136998 112914 137000 112966
rect 136944 112912 137000 112914
rect 136197 112623 136253 112679
rect 136944 111286 137000 111288
rect 136944 111234 136946 111286
rect 136946 111234 136998 111286
rect 136998 111234 137000 111286
rect 136944 111232 137000 111234
rect 136944 109606 137000 109608
rect 136944 109554 136946 109606
rect 136946 109554 136998 109606
rect 136998 109554 137000 109606
rect 136944 109552 137000 109554
rect 136944 107926 137000 107928
rect 136944 107874 136946 107926
rect 136946 107874 136998 107926
rect 136998 107874 137000 107926
rect 136944 107872 137000 107874
rect 136944 106246 137000 106248
rect 136944 106194 136946 106246
rect 136946 106194 136998 106246
rect 136998 106194 137000 106246
rect 136944 106192 137000 106194
rect 136944 104566 137000 104568
rect 136944 104514 136946 104566
rect 136946 104514 136998 104566
rect 136998 104514 137000 104566
rect 136944 104512 137000 104514
rect 136944 102886 137000 102888
rect 136944 102834 136946 102886
rect 136946 102834 136998 102886
rect 136998 102834 137000 102886
rect 136944 102832 137000 102834
rect 136944 101206 137000 101208
rect 136944 101154 136946 101206
rect 136946 101154 136998 101206
rect 136998 101154 137000 101206
rect 136944 101152 137000 101154
rect 136944 99526 137000 99528
rect 136944 99474 136946 99526
rect 136946 99474 136998 99526
rect 136998 99474 137000 99526
rect 136944 99472 137000 99474
rect 136944 97846 137000 97848
rect 136944 97794 136946 97846
rect 136946 97794 136998 97846
rect 136998 97794 137000 97846
rect 136944 97792 137000 97794
rect 136944 96166 137000 96168
rect 136944 96114 136946 96166
rect 136946 96114 136998 96166
rect 136998 96114 137000 96166
rect 136944 96112 137000 96114
rect 136944 94486 137000 94488
rect 136944 94434 136946 94486
rect 136946 94434 136998 94486
rect 136998 94434 137000 94486
rect 136944 94432 137000 94434
rect 136944 92806 137000 92808
rect 136944 92754 136946 92806
rect 136946 92754 136998 92806
rect 136998 92754 137000 92806
rect 136944 92752 137000 92754
rect 136944 91126 137000 91128
rect 136944 91074 136946 91126
rect 136946 91074 136998 91126
rect 136998 91074 137000 91126
rect 136944 91072 137000 91074
rect 136944 89446 137000 89448
rect 136944 89394 136946 89446
rect 136946 89394 136998 89446
rect 136998 89394 137000 89446
rect 136944 89392 137000 89394
rect 136944 87766 137000 87768
rect 136944 87714 136946 87766
rect 136946 87714 136998 87766
rect 136998 87714 137000 87766
rect 136944 87712 137000 87714
rect 136944 86086 137000 86088
rect 136944 86034 136946 86086
rect 136946 86034 136998 86086
rect 136998 86034 137000 86086
rect 136944 86032 137000 86034
rect 136944 84406 137000 84408
rect 136944 84354 136946 84406
rect 136946 84354 136998 84406
rect 136998 84354 137000 84406
rect 136944 84352 137000 84354
rect 136944 82726 137000 82728
rect 136944 82674 136946 82726
rect 136946 82674 136998 82726
rect 136998 82674 137000 82726
rect 136944 82672 137000 82674
rect 136944 81046 137000 81048
rect 136944 80994 136946 81046
rect 136946 80994 136998 81046
rect 136998 80994 137000 81046
rect 136944 80992 137000 80994
rect 136944 79366 137000 79368
rect 136944 79314 136946 79366
rect 136946 79314 136998 79366
rect 136998 79314 137000 79366
rect 136944 79312 137000 79314
rect 136944 77686 137000 77688
rect 136944 77634 136946 77686
rect 136946 77634 136998 77686
rect 136998 77634 137000 77686
rect 136944 77632 137000 77634
rect 136944 76006 137000 76008
rect 136944 75954 136946 76006
rect 136946 75954 136998 76006
rect 136998 75954 137000 76006
rect 136944 75952 137000 75954
rect 136944 74326 137000 74328
rect 136944 74274 136946 74326
rect 136946 74274 136998 74326
rect 136998 74274 137000 74326
rect 136944 74272 137000 74274
rect 136944 72646 137000 72648
rect 136944 72594 136946 72646
rect 136946 72594 136998 72646
rect 136998 72594 137000 72646
rect 136944 72592 137000 72594
rect 136944 70966 137000 70968
rect 136944 70914 136946 70966
rect 136946 70914 136998 70966
rect 136998 70914 137000 70966
rect 136944 70912 137000 70914
rect 136944 69286 137000 69288
rect 136944 69234 136946 69286
rect 136946 69234 136998 69286
rect 136998 69234 137000 69286
rect 136944 69232 137000 69234
rect 136944 67606 137000 67608
rect 136944 67554 136946 67606
rect 136946 67554 136998 67606
rect 136998 67554 137000 67606
rect 136944 67552 137000 67554
rect 136944 65926 137000 65928
rect 136944 65874 136946 65926
rect 136946 65874 136998 65926
rect 136998 65874 137000 65926
rect 136944 65872 137000 65874
rect 136944 64246 137000 64248
rect 136944 64194 136946 64246
rect 136946 64194 136998 64246
rect 136998 64194 137000 64246
rect 136944 64192 137000 64194
rect 136944 62566 137000 62568
rect 136944 62514 136946 62566
rect 136946 62514 136998 62566
rect 136998 62514 137000 62566
rect 136944 62512 137000 62514
rect 136944 60886 137000 60888
rect 136944 60834 136946 60886
rect 136946 60834 136998 60886
rect 136998 60834 137000 60886
rect 136944 60832 137000 60834
rect 136944 59206 137000 59208
rect 136944 59154 136946 59206
rect 136946 59154 136998 59206
rect 136998 59154 137000 59206
rect 136944 59152 137000 59154
rect 136944 57526 137000 57528
rect 136944 57474 136946 57526
rect 136946 57474 136998 57526
rect 136998 57474 137000 57526
rect 136944 57472 137000 57474
rect 136944 55846 137000 55848
rect 136944 55794 136946 55846
rect 136946 55794 136998 55846
rect 136998 55794 137000 55846
rect 136944 55792 137000 55794
rect 136944 54166 137000 54168
rect 136944 54114 136946 54166
rect 136946 54114 136998 54166
rect 136998 54114 137000 54166
rect 136944 54112 137000 54114
rect 136944 52486 137000 52488
rect 136944 52434 136946 52486
rect 136946 52434 136998 52486
rect 136998 52434 137000 52486
rect 136944 52432 137000 52434
rect 136944 50806 137000 50808
rect 136944 50754 136946 50806
rect 136946 50754 136998 50806
rect 136998 50754 137000 50806
rect 136944 50752 137000 50754
rect 136944 49126 137000 49128
rect 136944 49074 136946 49126
rect 136946 49074 136998 49126
rect 136998 49074 137000 49126
rect 136944 49072 137000 49074
rect 136944 47446 137000 47448
rect 136944 47394 136946 47446
rect 136946 47394 136998 47446
rect 136998 47394 137000 47446
rect 136944 47392 137000 47394
rect 136944 45766 137000 45768
rect 136944 45714 136946 45766
rect 136946 45714 136998 45766
rect 136998 45714 137000 45766
rect 136944 45712 137000 45714
rect 136944 44086 137000 44088
rect 136944 44034 136946 44086
rect 136946 44034 136998 44086
rect 136998 44034 137000 44086
rect 136944 44032 137000 44034
rect 136944 42406 137000 42408
rect 136944 42354 136946 42406
rect 136946 42354 136998 42406
rect 136998 42354 137000 42406
rect 136944 42352 137000 42354
rect 136944 40726 137000 40728
rect 136944 40674 136946 40726
rect 136946 40674 136998 40726
rect 136998 40674 137000 40726
rect 136944 40672 137000 40674
rect 136944 39046 137000 39048
rect 136944 38994 136946 39046
rect 136946 38994 136998 39046
rect 136998 38994 137000 39046
rect 136944 38992 137000 38994
rect 136944 37366 137000 37368
rect 136944 37314 136946 37366
rect 136946 37314 136998 37366
rect 136998 37314 137000 37366
rect 136944 37312 137000 37314
rect 136944 35686 137000 35688
rect 136944 35634 136946 35686
rect 136946 35634 136998 35686
rect 136998 35634 137000 35686
rect 136944 35632 137000 35634
rect 136944 34006 137000 34008
rect 136944 33954 136946 34006
rect 136946 33954 136998 34006
rect 136998 33954 137000 34006
rect 136944 33952 137000 33954
rect 136944 32326 137000 32328
rect 136944 32274 136946 32326
rect 136946 32274 136998 32326
rect 136998 32274 137000 32326
rect 136944 32272 137000 32274
rect 136944 30646 137000 30648
rect 136944 30594 136946 30646
rect 136946 30594 136998 30646
rect 136998 30594 137000 30646
rect 136944 30592 137000 30594
rect 136944 28966 137000 28968
rect 136944 28914 136946 28966
rect 136946 28914 136998 28966
rect 136998 28914 137000 28966
rect 136944 28912 137000 28914
rect 136944 27286 137000 27288
rect 136944 27234 136946 27286
rect 136946 27234 136998 27286
rect 136998 27234 137000 27286
rect 136944 27232 137000 27234
rect 136944 25606 137000 25608
rect 136944 25554 136946 25606
rect 136946 25554 136998 25606
rect 136998 25554 137000 25606
rect 136944 25552 137000 25554
rect 136944 23926 137000 23928
rect 136944 23874 136946 23926
rect 136946 23874 136998 23926
rect 136998 23874 137000 23926
rect 136944 23872 137000 23874
rect 136944 22246 137000 22248
rect 136944 22194 136946 22246
rect 136946 22194 136998 22246
rect 136998 22194 137000 22246
rect 136944 22192 137000 22194
rect 136944 20566 137000 20568
rect 136944 20514 136946 20566
rect 136946 20514 136998 20566
rect 136998 20514 137000 20566
rect 136944 20512 137000 20514
rect 123532 19510 123588 19566
rect 124614 19254 124670 19310
rect 123331 19237 123387 19239
rect 123331 19185 123333 19237
rect 123333 19185 123385 19237
rect 123385 19185 123387 19237
rect 123331 19183 123387 19185
rect 123669 19183 123725 19239
rect 23752 18197 23808 18253
rect 136944 18886 137000 18888
rect 136944 18834 136946 18886
rect 136946 18834 136998 18886
rect 136998 18834 137000 18886
rect 136944 18832 137000 18834
rect 123251 17679 123307 17681
rect 123251 17627 123253 17679
rect 123253 17627 123305 17679
rect 123305 17627 123307 17679
rect 123251 17625 123307 17627
rect 123669 17625 123725 17681
rect 124614 17554 124670 17610
rect 136944 17206 137000 17208
rect 136944 17154 136946 17206
rect 136946 17154 136998 17206
rect 136998 17154 137000 17206
rect 136944 17152 137000 17154
rect 124614 16426 124670 16482
rect 123171 16409 123227 16411
rect 123171 16357 123173 16409
rect 123173 16357 123225 16409
rect 123225 16357 123227 16409
rect 123171 16355 123227 16357
rect 123669 16355 123725 16411
rect 136944 15526 137000 15528
rect 136944 15474 136946 15526
rect 136946 15474 136998 15526
rect 136998 15474 137000 15526
rect 136944 15472 137000 15474
rect 27455 15369 27511 15425
rect 123091 14851 123147 14853
rect 123091 14799 123093 14851
rect 123093 14799 123145 14851
rect 123145 14799 123147 14851
rect 123091 14797 123147 14799
rect 123669 14797 123725 14853
rect 124614 14726 124670 14782
rect 27703 13955 27759 14011
rect 27579 12541 27635 12597
rect 136944 13846 137000 13848
rect 136944 13794 136946 13846
rect 136946 13794 136998 13846
rect 136998 13794 137000 13846
rect 136944 13792 137000 13794
rect 124614 13598 124670 13654
rect 123011 13581 123067 13583
rect 123011 13529 123013 13581
rect 123013 13529 123065 13581
rect 123065 13529 123067 13581
rect 123011 13527 123067 13529
rect 123669 13527 123725 13583
rect 29562 13259 29618 13261
rect 29562 13207 29564 13259
rect 29564 13207 29616 13259
rect 29616 13207 29618 13259
rect 29562 13205 29618 13207
rect 32058 13259 32114 13261
rect 32058 13207 32060 13259
rect 32060 13207 32112 13259
rect 32112 13207 32114 13259
rect 32058 13205 32114 13207
rect 34554 13259 34610 13261
rect 34554 13207 34556 13259
rect 34556 13207 34608 13259
rect 34608 13207 34610 13259
rect 34554 13205 34610 13207
rect 37050 13259 37106 13261
rect 37050 13207 37052 13259
rect 37052 13207 37104 13259
rect 37104 13207 37106 13259
rect 37050 13205 37106 13207
rect 39546 13259 39602 13261
rect 39546 13207 39548 13259
rect 39548 13207 39600 13259
rect 39600 13207 39602 13259
rect 39546 13205 39602 13207
rect 42042 13259 42098 13261
rect 42042 13207 42044 13259
rect 42044 13207 42096 13259
rect 42096 13207 42098 13259
rect 42042 13205 42098 13207
rect 44538 13259 44594 13261
rect 44538 13207 44540 13259
rect 44540 13207 44592 13259
rect 44592 13207 44594 13259
rect 44538 13205 44594 13207
rect 47034 13259 47090 13261
rect 47034 13207 47036 13259
rect 47036 13207 47088 13259
rect 47088 13207 47090 13259
rect 47034 13205 47090 13207
rect 49530 13259 49586 13261
rect 49530 13207 49532 13259
rect 49532 13207 49584 13259
rect 49584 13207 49586 13259
rect 49530 13205 49586 13207
rect 52026 13259 52082 13261
rect 52026 13207 52028 13259
rect 52028 13207 52080 13259
rect 52080 13207 52082 13259
rect 52026 13205 52082 13207
rect 54522 13259 54578 13261
rect 54522 13207 54524 13259
rect 54524 13207 54576 13259
rect 54576 13207 54578 13259
rect 54522 13205 54578 13207
rect 57018 13259 57074 13261
rect 57018 13207 57020 13259
rect 57020 13207 57072 13259
rect 57072 13207 57074 13259
rect 57018 13205 57074 13207
rect 59514 13259 59570 13261
rect 59514 13207 59516 13259
rect 59516 13207 59568 13259
rect 59568 13207 59570 13259
rect 59514 13205 59570 13207
rect 62010 13259 62066 13261
rect 62010 13207 62012 13259
rect 62012 13207 62064 13259
rect 62064 13207 62066 13259
rect 62010 13205 62066 13207
rect 64506 13259 64562 13261
rect 64506 13207 64508 13259
rect 64508 13207 64560 13259
rect 64560 13207 64562 13259
rect 64506 13205 64562 13207
rect 67002 13259 67058 13261
rect 67002 13207 67004 13259
rect 67004 13207 67056 13259
rect 67056 13207 67058 13259
rect 67002 13205 67058 13207
rect 69498 13259 69554 13261
rect 69498 13207 69500 13259
rect 69500 13207 69552 13259
rect 69552 13207 69554 13259
rect 69498 13205 69554 13207
rect 71994 13259 72050 13261
rect 71994 13207 71996 13259
rect 71996 13207 72048 13259
rect 72048 13207 72050 13259
rect 71994 13205 72050 13207
rect 74490 13259 74546 13261
rect 74490 13207 74492 13259
rect 74492 13207 74544 13259
rect 74544 13207 74546 13259
rect 74490 13205 74546 13207
rect 76986 13259 77042 13261
rect 76986 13207 76988 13259
rect 76988 13207 77040 13259
rect 77040 13207 77042 13259
rect 76986 13205 77042 13207
rect 79482 13259 79538 13261
rect 79482 13207 79484 13259
rect 79484 13207 79536 13259
rect 79536 13207 79538 13259
rect 79482 13205 79538 13207
rect 81978 13259 82034 13261
rect 81978 13207 81980 13259
rect 81980 13207 82032 13259
rect 82032 13207 82034 13259
rect 81978 13205 82034 13207
rect 84474 13259 84530 13261
rect 84474 13207 84476 13259
rect 84476 13207 84528 13259
rect 84528 13207 84530 13259
rect 84474 13205 84530 13207
rect 86970 13259 87026 13261
rect 86970 13207 86972 13259
rect 86972 13207 87024 13259
rect 87024 13207 87026 13259
rect 86970 13205 87026 13207
rect 89466 13259 89522 13261
rect 89466 13207 89468 13259
rect 89468 13207 89520 13259
rect 89520 13207 89522 13259
rect 89466 13205 89522 13207
rect 91962 13259 92018 13261
rect 91962 13207 91964 13259
rect 91964 13207 92016 13259
rect 92016 13207 92018 13259
rect 91962 13205 92018 13207
rect 94458 13259 94514 13261
rect 94458 13207 94460 13259
rect 94460 13207 94512 13259
rect 94512 13207 94514 13259
rect 94458 13205 94514 13207
rect 96954 13259 97010 13261
rect 96954 13207 96956 13259
rect 96956 13207 97008 13259
rect 97008 13207 97010 13259
rect 96954 13205 97010 13207
rect 99450 13259 99506 13261
rect 99450 13207 99452 13259
rect 99452 13207 99504 13259
rect 99504 13207 99506 13259
rect 99450 13205 99506 13207
rect 101946 13259 102002 13261
rect 101946 13207 101948 13259
rect 101948 13207 102000 13259
rect 102000 13207 102002 13259
rect 101946 13205 102002 13207
rect 104442 13259 104498 13261
rect 104442 13207 104444 13259
rect 104444 13207 104496 13259
rect 104496 13207 104498 13259
rect 104442 13205 104498 13207
rect 106938 13259 106994 13261
rect 106938 13207 106940 13259
rect 106940 13207 106992 13259
rect 106992 13207 106994 13259
rect 106938 13205 106994 13207
rect 136944 12166 137000 12168
rect 136944 12114 136946 12166
rect 136946 12114 136998 12166
rect 136998 12114 137000 12166
rect 136944 12112 137000 12114
rect 122931 12023 122987 12025
rect 122931 11971 122933 12023
rect 122933 11971 122985 12023
rect 122985 11971 122987 12023
rect 122931 11969 122987 11971
rect 123669 11969 123725 12025
rect 124614 11898 124670 11954
rect 124614 10770 124670 10826
rect 122851 10753 122907 10755
rect 122851 10701 122853 10753
rect 122853 10701 122905 10753
rect 122905 10701 122907 10753
rect 122851 10699 122907 10701
rect 123669 10699 123725 10755
rect 136944 10486 137000 10488
rect 136944 10434 136946 10486
rect 136946 10434 136998 10486
rect 136998 10434 137000 10486
rect 136944 10432 137000 10434
rect 122771 9195 122827 9197
rect 122771 9143 122773 9195
rect 122773 9143 122825 9195
rect 122825 9143 122827 9195
rect 122771 9141 122827 9143
rect 123669 9141 123725 9197
rect 124614 9070 124670 9126
rect 5979 8261 6035 8317
rect 2758 8156 2814 8212
rect 1798 7126 1854 7128
rect 1798 7074 1800 7126
rect 1800 7074 1852 7126
rect 1852 7074 1854 7126
rect 1798 7072 1854 7074
rect 1798 5446 1854 5448
rect 1798 5394 1800 5446
rect 1800 5394 1852 5446
rect 1852 5394 1854 5446
rect 1798 5392 1854 5394
rect 1798 3766 1854 3768
rect 1798 3714 1800 3766
rect 1800 3714 1852 3766
rect 1852 3714 1854 3766
rect 1798 3712 1854 3714
rect 136944 8806 137000 8808
rect 136944 8754 136946 8806
rect 136946 8754 136998 8806
rect 136998 8754 137000 8806
rect 136944 8752 137000 8754
rect 136944 7126 137000 7128
rect 136944 7074 136946 7126
rect 136946 7074 136998 7126
rect 136998 7074 137000 7126
rect 136944 7072 137000 7074
rect 136944 5446 137000 5448
rect 136944 5394 136946 5446
rect 136946 5394 136998 5446
rect 136998 5394 137000 5446
rect 136944 5392 137000 5394
rect 136944 3766 137000 3768
rect 136944 3714 136946 3766
rect 136946 3714 136998 3766
rect 136998 3714 137000 3766
rect 136944 3712 137000 3714
rect 16548 2932 16604 2988
rect 17716 2932 17772 2988
rect 18884 2932 18940 2988
rect 20052 2932 20108 2988
rect 21220 2932 21276 2988
rect 22388 2932 22444 2988
rect 23556 2932 23612 2988
rect 24724 2932 24780 2988
rect 25892 2932 25948 2988
rect 27060 2932 27116 2988
rect 28228 2932 28284 2988
rect 29396 2932 29452 2988
rect 30564 2932 30620 2988
rect 31732 2932 31788 2988
rect 32900 2932 32956 2988
rect 34068 2932 34124 2988
rect 35236 2932 35292 2988
rect 36404 2932 36460 2988
rect 37572 2932 37628 2988
rect 38740 2932 38796 2988
rect 39908 2932 39964 2988
rect 41076 2932 41132 2988
rect 42244 2932 42300 2988
rect 43412 2932 43468 2988
rect 44580 2932 44636 2988
rect 45748 2932 45804 2988
rect 46916 2932 46972 2988
rect 48084 2932 48140 2988
rect 49252 2932 49308 2988
rect 50420 2932 50476 2988
rect 51588 2932 51644 2988
rect 52756 2932 52812 2988
rect 53924 2932 53980 2988
rect 55092 2932 55148 2988
rect 56260 2932 56316 2988
rect 57428 2932 57484 2988
rect 58596 2932 58652 2988
rect 59764 2932 59820 2988
rect 15294 2676 15350 2732
rect 1798 2086 1854 2088
rect 1798 2034 1800 2086
rect 1800 2034 1852 2086
rect 1852 2034 1854 2086
rect 1798 2032 1854 2034
rect 136944 2086 137000 2088
rect 136944 2034 136946 2086
rect 136946 2034 136998 2086
rect 136998 2034 137000 2086
rect 136944 2032 137000 2034
rect 2134 1750 2190 1752
rect 2134 1698 2136 1750
rect 2136 1698 2188 1750
rect 2188 1698 2190 1750
rect 2134 1696 2190 1698
rect 3814 1750 3870 1752
rect 3814 1698 3816 1750
rect 3816 1698 3868 1750
rect 3868 1698 3870 1750
rect 3814 1696 3870 1698
rect 5494 1750 5550 1752
rect 5494 1698 5496 1750
rect 5496 1698 5548 1750
rect 5548 1698 5550 1750
rect 5494 1696 5550 1698
rect 7174 1750 7230 1752
rect 7174 1698 7176 1750
rect 7176 1698 7228 1750
rect 7228 1698 7230 1750
rect 7174 1696 7230 1698
rect 8854 1750 8910 1752
rect 8854 1698 8856 1750
rect 8856 1698 8908 1750
rect 8908 1698 8910 1750
rect 8854 1696 8910 1698
rect 10534 1750 10590 1752
rect 10534 1698 10536 1750
rect 10536 1698 10588 1750
rect 10588 1698 10590 1750
rect 10534 1696 10590 1698
rect 12214 1750 12270 1752
rect 12214 1698 12216 1750
rect 12216 1698 12268 1750
rect 12268 1698 12270 1750
rect 12214 1696 12270 1698
rect 13894 1750 13950 1752
rect 13894 1698 13896 1750
rect 13896 1698 13948 1750
rect 13948 1698 13950 1750
rect 13894 1696 13950 1698
rect 15574 1750 15630 1752
rect 15574 1698 15576 1750
rect 15576 1698 15628 1750
rect 15628 1698 15630 1750
rect 15574 1696 15630 1698
rect 17254 1750 17310 1752
rect 17254 1698 17256 1750
rect 17256 1698 17308 1750
rect 17308 1698 17310 1750
rect 17254 1696 17310 1698
rect 18934 1750 18990 1752
rect 18934 1698 18936 1750
rect 18936 1698 18988 1750
rect 18988 1698 18990 1750
rect 18934 1696 18990 1698
rect 20614 1750 20670 1752
rect 20614 1698 20616 1750
rect 20616 1698 20668 1750
rect 20668 1698 20670 1750
rect 20614 1696 20670 1698
rect 22294 1750 22350 1752
rect 22294 1698 22296 1750
rect 22296 1698 22348 1750
rect 22348 1698 22350 1750
rect 22294 1696 22350 1698
rect 23974 1750 24030 1752
rect 23974 1698 23976 1750
rect 23976 1698 24028 1750
rect 24028 1698 24030 1750
rect 23974 1696 24030 1698
rect 25654 1750 25710 1752
rect 25654 1698 25656 1750
rect 25656 1698 25708 1750
rect 25708 1698 25710 1750
rect 25654 1696 25710 1698
rect 27334 1750 27390 1752
rect 27334 1698 27336 1750
rect 27336 1698 27388 1750
rect 27388 1698 27390 1750
rect 27334 1696 27390 1698
rect 29014 1750 29070 1752
rect 29014 1698 29016 1750
rect 29016 1698 29068 1750
rect 29068 1698 29070 1750
rect 29014 1696 29070 1698
rect 30694 1750 30750 1752
rect 30694 1698 30696 1750
rect 30696 1698 30748 1750
rect 30748 1698 30750 1750
rect 30694 1696 30750 1698
rect 32374 1750 32430 1752
rect 32374 1698 32376 1750
rect 32376 1698 32428 1750
rect 32428 1698 32430 1750
rect 32374 1696 32430 1698
rect 34054 1750 34110 1752
rect 34054 1698 34056 1750
rect 34056 1698 34108 1750
rect 34108 1698 34110 1750
rect 34054 1696 34110 1698
rect 35734 1750 35790 1752
rect 35734 1698 35736 1750
rect 35736 1698 35788 1750
rect 35788 1698 35790 1750
rect 35734 1696 35790 1698
rect 37414 1750 37470 1752
rect 37414 1698 37416 1750
rect 37416 1698 37468 1750
rect 37468 1698 37470 1750
rect 37414 1696 37470 1698
rect 39094 1750 39150 1752
rect 39094 1698 39096 1750
rect 39096 1698 39148 1750
rect 39148 1698 39150 1750
rect 39094 1696 39150 1698
rect 40774 1750 40830 1752
rect 40774 1698 40776 1750
rect 40776 1698 40828 1750
rect 40828 1698 40830 1750
rect 40774 1696 40830 1698
rect 42454 1750 42510 1752
rect 42454 1698 42456 1750
rect 42456 1698 42508 1750
rect 42508 1698 42510 1750
rect 42454 1696 42510 1698
rect 44134 1750 44190 1752
rect 44134 1698 44136 1750
rect 44136 1698 44188 1750
rect 44188 1698 44190 1750
rect 44134 1696 44190 1698
rect 45814 1750 45870 1752
rect 45814 1698 45816 1750
rect 45816 1698 45868 1750
rect 45868 1698 45870 1750
rect 45814 1696 45870 1698
rect 47494 1750 47550 1752
rect 47494 1698 47496 1750
rect 47496 1698 47548 1750
rect 47548 1698 47550 1750
rect 47494 1696 47550 1698
rect 49174 1750 49230 1752
rect 49174 1698 49176 1750
rect 49176 1698 49228 1750
rect 49228 1698 49230 1750
rect 49174 1696 49230 1698
rect 50854 1750 50910 1752
rect 50854 1698 50856 1750
rect 50856 1698 50908 1750
rect 50908 1698 50910 1750
rect 50854 1696 50910 1698
rect 52534 1750 52590 1752
rect 52534 1698 52536 1750
rect 52536 1698 52588 1750
rect 52588 1698 52590 1750
rect 52534 1696 52590 1698
rect 54214 1750 54270 1752
rect 54214 1698 54216 1750
rect 54216 1698 54268 1750
rect 54268 1698 54270 1750
rect 54214 1696 54270 1698
rect 55894 1750 55950 1752
rect 55894 1698 55896 1750
rect 55896 1698 55948 1750
rect 55948 1698 55950 1750
rect 55894 1696 55950 1698
rect 57574 1750 57630 1752
rect 57574 1698 57576 1750
rect 57576 1698 57628 1750
rect 57628 1698 57630 1750
rect 57574 1696 57630 1698
rect 59254 1750 59310 1752
rect 59254 1698 59256 1750
rect 59256 1698 59308 1750
rect 59308 1698 59310 1750
rect 59254 1696 59310 1698
rect 60934 1750 60990 1752
rect 60934 1698 60936 1750
rect 60936 1698 60988 1750
rect 60988 1698 60990 1750
rect 60934 1696 60990 1698
rect 62614 1750 62670 1752
rect 62614 1698 62616 1750
rect 62616 1698 62668 1750
rect 62668 1698 62670 1750
rect 62614 1696 62670 1698
rect 64294 1750 64350 1752
rect 64294 1698 64296 1750
rect 64296 1698 64348 1750
rect 64348 1698 64350 1750
rect 64294 1696 64350 1698
rect 65974 1750 66030 1752
rect 65974 1698 65976 1750
rect 65976 1698 66028 1750
rect 66028 1698 66030 1750
rect 65974 1696 66030 1698
rect 67654 1750 67710 1752
rect 67654 1698 67656 1750
rect 67656 1698 67708 1750
rect 67708 1698 67710 1750
rect 67654 1696 67710 1698
rect 69334 1750 69390 1752
rect 69334 1698 69336 1750
rect 69336 1698 69388 1750
rect 69388 1698 69390 1750
rect 69334 1696 69390 1698
rect 71014 1750 71070 1752
rect 71014 1698 71016 1750
rect 71016 1698 71068 1750
rect 71068 1698 71070 1750
rect 71014 1696 71070 1698
rect 72694 1750 72750 1752
rect 72694 1698 72696 1750
rect 72696 1698 72748 1750
rect 72748 1698 72750 1750
rect 72694 1696 72750 1698
rect 74374 1750 74430 1752
rect 74374 1698 74376 1750
rect 74376 1698 74428 1750
rect 74428 1698 74430 1750
rect 74374 1696 74430 1698
rect 76054 1750 76110 1752
rect 76054 1698 76056 1750
rect 76056 1698 76108 1750
rect 76108 1698 76110 1750
rect 76054 1696 76110 1698
rect 77734 1750 77790 1752
rect 77734 1698 77736 1750
rect 77736 1698 77788 1750
rect 77788 1698 77790 1750
rect 77734 1696 77790 1698
rect 79414 1750 79470 1752
rect 79414 1698 79416 1750
rect 79416 1698 79468 1750
rect 79468 1698 79470 1750
rect 79414 1696 79470 1698
rect 81094 1750 81150 1752
rect 81094 1698 81096 1750
rect 81096 1698 81148 1750
rect 81148 1698 81150 1750
rect 81094 1696 81150 1698
rect 82774 1750 82830 1752
rect 82774 1698 82776 1750
rect 82776 1698 82828 1750
rect 82828 1698 82830 1750
rect 82774 1696 82830 1698
rect 84454 1750 84510 1752
rect 84454 1698 84456 1750
rect 84456 1698 84508 1750
rect 84508 1698 84510 1750
rect 84454 1696 84510 1698
rect 86134 1750 86190 1752
rect 86134 1698 86136 1750
rect 86136 1698 86188 1750
rect 86188 1698 86190 1750
rect 86134 1696 86190 1698
rect 87814 1750 87870 1752
rect 87814 1698 87816 1750
rect 87816 1698 87868 1750
rect 87868 1698 87870 1750
rect 87814 1696 87870 1698
rect 89494 1750 89550 1752
rect 89494 1698 89496 1750
rect 89496 1698 89548 1750
rect 89548 1698 89550 1750
rect 89494 1696 89550 1698
rect 91174 1750 91230 1752
rect 91174 1698 91176 1750
rect 91176 1698 91228 1750
rect 91228 1698 91230 1750
rect 91174 1696 91230 1698
rect 92854 1750 92910 1752
rect 92854 1698 92856 1750
rect 92856 1698 92908 1750
rect 92908 1698 92910 1750
rect 92854 1696 92910 1698
rect 94534 1750 94590 1752
rect 94534 1698 94536 1750
rect 94536 1698 94588 1750
rect 94588 1698 94590 1750
rect 94534 1696 94590 1698
rect 96214 1750 96270 1752
rect 96214 1698 96216 1750
rect 96216 1698 96268 1750
rect 96268 1698 96270 1750
rect 96214 1696 96270 1698
rect 97894 1750 97950 1752
rect 97894 1698 97896 1750
rect 97896 1698 97948 1750
rect 97948 1698 97950 1750
rect 97894 1696 97950 1698
rect 99574 1750 99630 1752
rect 99574 1698 99576 1750
rect 99576 1698 99628 1750
rect 99628 1698 99630 1750
rect 99574 1696 99630 1698
rect 101254 1750 101310 1752
rect 101254 1698 101256 1750
rect 101256 1698 101308 1750
rect 101308 1698 101310 1750
rect 101254 1696 101310 1698
rect 102934 1750 102990 1752
rect 102934 1698 102936 1750
rect 102936 1698 102988 1750
rect 102988 1698 102990 1750
rect 102934 1696 102990 1698
rect 104614 1750 104670 1752
rect 104614 1698 104616 1750
rect 104616 1698 104668 1750
rect 104668 1698 104670 1750
rect 104614 1696 104670 1698
rect 106294 1750 106350 1752
rect 106294 1698 106296 1750
rect 106296 1698 106348 1750
rect 106348 1698 106350 1750
rect 106294 1696 106350 1698
rect 107974 1750 108030 1752
rect 107974 1698 107976 1750
rect 107976 1698 108028 1750
rect 108028 1698 108030 1750
rect 107974 1696 108030 1698
rect 109654 1750 109710 1752
rect 109654 1698 109656 1750
rect 109656 1698 109708 1750
rect 109708 1698 109710 1750
rect 109654 1696 109710 1698
rect 111334 1750 111390 1752
rect 111334 1698 111336 1750
rect 111336 1698 111388 1750
rect 111388 1698 111390 1750
rect 111334 1696 111390 1698
rect 113014 1750 113070 1752
rect 113014 1698 113016 1750
rect 113016 1698 113068 1750
rect 113068 1698 113070 1750
rect 113014 1696 113070 1698
rect 114694 1750 114750 1752
rect 114694 1698 114696 1750
rect 114696 1698 114748 1750
rect 114748 1698 114750 1750
rect 114694 1696 114750 1698
rect 116374 1750 116430 1752
rect 116374 1698 116376 1750
rect 116376 1698 116428 1750
rect 116428 1698 116430 1750
rect 116374 1696 116430 1698
rect 118054 1750 118110 1752
rect 118054 1698 118056 1750
rect 118056 1698 118108 1750
rect 118108 1698 118110 1750
rect 118054 1696 118110 1698
rect 119734 1750 119790 1752
rect 119734 1698 119736 1750
rect 119736 1698 119788 1750
rect 119788 1698 119790 1750
rect 119734 1696 119790 1698
rect 121414 1750 121470 1752
rect 121414 1698 121416 1750
rect 121416 1698 121468 1750
rect 121468 1698 121470 1750
rect 121414 1696 121470 1698
rect 123094 1750 123150 1752
rect 123094 1698 123096 1750
rect 123096 1698 123148 1750
rect 123148 1698 123150 1750
rect 123094 1696 123150 1698
rect 124774 1750 124830 1752
rect 124774 1698 124776 1750
rect 124776 1698 124828 1750
rect 124828 1698 124830 1750
rect 124774 1696 124830 1698
rect 126454 1750 126510 1752
rect 126454 1698 126456 1750
rect 126456 1698 126508 1750
rect 126508 1698 126510 1750
rect 126454 1696 126510 1698
rect 128134 1750 128190 1752
rect 128134 1698 128136 1750
rect 128136 1698 128188 1750
rect 128188 1698 128190 1750
rect 128134 1696 128190 1698
rect 129814 1750 129870 1752
rect 129814 1698 129816 1750
rect 129816 1698 129868 1750
rect 129868 1698 129870 1750
rect 129814 1696 129870 1698
rect 131494 1750 131550 1752
rect 131494 1698 131496 1750
rect 131496 1698 131548 1750
rect 131548 1698 131550 1750
rect 131494 1696 131550 1698
rect 133174 1750 133230 1752
rect 133174 1698 133176 1750
rect 133176 1698 133228 1750
rect 133228 1698 133230 1750
rect 133174 1696 133230 1698
rect 134854 1750 134910 1752
rect 134854 1698 134856 1750
rect 134856 1698 134908 1750
rect 134908 1698 134910 1750
rect 134854 1696 134910 1698
rect 136534 1750 136590 1752
rect 136534 1698 136536 1750
rect 136536 1698 136588 1750
rect 136588 1698 136590 1750
rect 136534 1696 136590 1698
<< metal3 >>
rect 272 133486 138524 133492
rect 272 133422 278 133486
rect 342 133422 414 133486
rect 478 133422 550 133486
rect 614 133422 138182 133486
rect 138246 133422 138318 133486
rect 138382 133422 138454 133486
rect 138518 133422 138524 133486
rect 272 133350 138524 133422
rect 272 133286 278 133350
rect 342 133286 414 133350
rect 478 133286 550 133350
rect 614 133286 138182 133350
rect 138246 133286 138318 133350
rect 138382 133286 138454 133350
rect 138518 133286 138524 133350
rect 272 133214 138524 133286
rect 272 133150 278 133214
rect 342 133150 414 133214
rect 478 133150 550 133214
rect 614 133150 120638 133214
rect 120702 133150 123630 133214
rect 123694 133150 138182 133214
rect 138246 133150 138318 133214
rect 138382 133150 138454 133214
rect 138518 133150 138524 133214
rect 272 133144 138524 133150
rect 952 132806 137844 132812
rect 952 132742 958 132806
rect 1022 132742 1094 132806
rect 1158 132742 1230 132806
rect 1294 132742 137502 132806
rect 137566 132742 137638 132806
rect 137702 132742 137774 132806
rect 137838 132742 137844 132806
rect 952 132670 137844 132742
rect 952 132606 958 132670
rect 1022 132606 1094 132670
rect 1158 132606 1230 132670
rect 1294 132606 137502 132670
rect 137566 132606 137638 132670
rect 137702 132606 137774 132670
rect 137838 132606 137844 132670
rect 952 132534 137844 132606
rect 952 132470 958 132534
rect 1022 132470 1094 132534
rect 1158 132470 1230 132534
rect 1294 132470 2182 132534
rect 2246 132470 3678 132534
rect 3742 132470 5446 132534
rect 5510 132470 7214 132534
rect 7278 132470 8982 132534
rect 9046 132470 10478 132534
rect 10542 132470 12110 132534
rect 12174 132470 13878 132534
rect 13942 132470 15646 132534
rect 15710 132470 17142 132534
rect 17206 132470 18910 132534
rect 18974 132470 20678 132534
rect 20742 132470 22174 132534
rect 22238 132470 23942 132534
rect 24006 132470 25710 132534
rect 25774 132470 27206 132534
rect 27270 132470 28974 132534
rect 29038 132470 30742 132534
rect 30806 132470 32238 132534
rect 32302 132470 34142 132534
rect 34206 132470 35638 132534
rect 35702 132470 37406 132534
rect 37470 132470 39174 132534
rect 39238 132470 40670 132534
rect 40734 132470 42438 132534
rect 42502 132470 44206 132534
rect 44270 132470 45702 132534
rect 45766 132470 47470 132534
rect 47534 132470 49102 132534
rect 49166 132470 50734 132534
rect 50798 132470 52638 132534
rect 52702 132470 54134 132534
rect 54198 132470 55902 132534
rect 55966 132470 57670 132534
rect 57734 132470 59166 132534
rect 59230 132470 61070 132534
rect 61134 132470 62702 132534
rect 62766 132470 64198 132534
rect 64262 132470 66102 132534
rect 66166 132470 67734 132534
rect 67798 132470 69230 132534
rect 69294 132470 71134 132534
rect 71198 132470 72630 132534
rect 72694 132470 74262 132534
rect 74326 132470 76166 132534
rect 76230 132470 77662 132534
rect 77726 132470 79294 132534
rect 79358 132470 81198 132534
rect 81262 132470 82694 132534
rect 82758 132470 84326 132534
rect 84390 132470 86094 132534
rect 86158 132470 87726 132534
rect 87790 132470 89766 132534
rect 89830 132470 91126 132534
rect 91190 132470 92894 132534
rect 92958 132470 94662 132534
rect 94726 132470 96158 132534
rect 96222 132470 97926 132534
rect 97990 132470 99694 132534
rect 99758 132470 101190 132534
rect 101254 132470 102958 132534
rect 103022 132470 104726 132534
rect 104790 132470 106222 132534
rect 106286 132470 107854 132534
rect 107918 132470 109622 132534
rect 109686 132470 111390 132534
rect 111454 132470 112886 132534
rect 112950 132470 114654 132534
rect 114718 132470 116422 132534
rect 116486 132470 117918 132534
rect 117982 132470 119686 132534
rect 119750 132470 121454 132534
rect 121518 132470 123086 132534
rect 123150 132470 124718 132534
rect 124782 132470 126350 132534
rect 126414 132470 128118 132534
rect 128182 132470 129886 132534
rect 129950 132470 131382 132534
rect 131446 132470 133150 132534
rect 133214 132470 134918 132534
rect 134982 132470 136414 132534
rect 136478 132470 137502 132534
rect 137566 132470 137638 132534
rect 137702 132470 137774 132534
rect 137838 132470 137844 132534
rect 952 132464 137844 132470
rect 2040 132126 2252 132132
rect 2040 132062 2182 132126
rect 2246 132062 2252 132126
rect 2040 132061 2252 132062
rect 2040 132005 2134 132061
rect 2190 132005 2252 132061
rect 2040 131990 2252 132005
rect 2040 131926 2046 131990
rect 2110 131926 2252 131990
rect 2040 131920 2252 131926
rect 3672 132126 4020 132132
rect 3672 132062 3678 132126
rect 3742 132062 4020 132126
rect 3672 132061 4020 132062
rect 3672 132005 3814 132061
rect 3870 132005 4020 132061
rect 3672 131920 4020 132005
rect 5440 132126 5652 132132
rect 5440 132062 5446 132126
rect 5510 132062 5652 132126
rect 5440 132061 5652 132062
rect 5440 132005 5494 132061
rect 5550 132005 5652 132061
rect 5440 131920 5652 132005
rect 7072 132126 7284 132132
rect 7072 132062 7214 132126
rect 7278 132062 7284 132126
rect 7072 132061 7284 132062
rect 7072 132005 7174 132061
rect 7230 132005 7284 132061
rect 7072 131920 7284 132005
rect 8704 132126 9052 132132
rect 8704 132062 8982 132126
rect 9046 132062 9052 132126
rect 8704 132061 9052 132062
rect 8704 132005 8854 132061
rect 8910 132005 9052 132061
rect 8704 131920 9052 132005
rect 10472 132126 10684 132132
rect 10472 132062 10478 132126
rect 10542 132062 10684 132126
rect 10472 132061 10684 132062
rect 10472 132005 10534 132061
rect 10590 132005 10684 132061
rect 10472 131920 10684 132005
rect 12104 132126 12316 132132
rect 12104 132062 12110 132126
rect 12174 132062 12316 132126
rect 12104 132061 12316 132062
rect 12104 132005 12214 132061
rect 12270 132005 12316 132061
rect 12104 131920 12316 132005
rect 13872 132126 14084 132132
rect 13872 132062 13878 132126
rect 13942 132062 14084 132126
rect 13872 132061 14084 132062
rect 13872 132005 13894 132061
rect 13950 132005 14084 132061
rect 13872 131920 14084 132005
rect 15504 132126 15716 132132
rect 15504 132062 15646 132126
rect 15710 132062 15716 132126
rect 15504 132061 15716 132062
rect 15504 132005 15574 132061
rect 15630 132005 15716 132061
rect 15504 131920 15716 132005
rect 17136 132126 17348 132132
rect 17136 132062 17142 132126
rect 17206 132062 17348 132126
rect 17136 132061 17348 132062
rect 17136 132005 17254 132061
rect 17310 132005 17348 132061
rect 17136 131920 17348 132005
rect 18904 132126 19116 132132
rect 18904 132062 18910 132126
rect 18974 132062 19116 132126
rect 18904 132061 19116 132062
rect 18904 132005 18934 132061
rect 18990 132005 19116 132061
rect 18904 131920 19116 132005
rect 20536 132126 20748 132132
rect 20536 132062 20678 132126
rect 20742 132062 20748 132126
rect 20536 132061 20748 132062
rect 20536 132005 20614 132061
rect 20670 132005 20748 132061
rect 20536 131920 20748 132005
rect 22168 132126 22380 132132
rect 22168 132062 22174 132126
rect 22238 132062 22380 132126
rect 22168 132061 22380 132062
rect 22168 132005 22294 132061
rect 22350 132005 22380 132061
rect 22168 131920 22380 132005
rect 23936 132126 24148 132132
rect 23936 132062 23942 132126
rect 24006 132062 24148 132126
rect 23936 132061 24148 132062
rect 23936 132005 23974 132061
rect 24030 132005 24148 132061
rect 23936 131920 24148 132005
rect 25568 132126 25780 132132
rect 25568 132062 25710 132126
rect 25774 132062 25780 132126
rect 25568 132061 25780 132062
rect 25568 132005 25654 132061
rect 25710 132005 25780 132061
rect 25568 131920 25780 132005
rect 27200 132126 27412 132132
rect 27200 132062 27206 132126
rect 27270 132062 27412 132126
rect 27200 132061 27412 132062
rect 27200 132005 27334 132061
rect 27390 132005 27412 132061
rect 27200 131920 27412 132005
rect 28968 132126 29180 132132
rect 28968 132062 28974 132126
rect 29038 132062 29180 132126
rect 28968 132061 29180 132062
rect 28968 132005 29014 132061
rect 29070 132005 29180 132061
rect 28968 131920 29180 132005
rect 30600 132126 30812 132132
rect 30600 132062 30742 132126
rect 30806 132062 30812 132126
rect 30600 132061 30812 132062
rect 30600 132005 30694 132061
rect 30750 132005 30812 132061
rect 30600 131920 30812 132005
rect 32232 132126 32580 132132
rect 32232 132062 32238 132126
rect 32302 132062 32580 132126
rect 32232 132061 32580 132062
rect 32232 132005 32374 132061
rect 32430 132005 32580 132061
rect 32232 131920 32580 132005
rect 34000 132126 34212 132132
rect 34000 132062 34142 132126
rect 34206 132062 34212 132126
rect 34000 132061 34212 132062
rect 34000 132005 34054 132061
rect 34110 132005 34212 132061
rect 34000 131920 34212 132005
rect 35632 132126 35844 132132
rect 35632 132062 35638 132126
rect 35702 132062 35844 132126
rect 35632 132061 35844 132062
rect 35632 132005 35734 132061
rect 35790 132005 35844 132061
rect 35632 131920 35844 132005
rect 37264 132126 37612 132132
rect 37264 132062 37406 132126
rect 37470 132062 37612 132126
rect 37264 132061 37612 132062
rect 37264 132005 37414 132061
rect 37470 132005 37612 132061
rect 37264 131920 37612 132005
rect 39032 132126 39244 132132
rect 39032 132062 39174 132126
rect 39238 132062 39244 132126
rect 39032 132061 39244 132062
rect 39032 132005 39094 132061
rect 39150 132005 39244 132061
rect 39032 131920 39244 132005
rect 40664 132126 40876 132132
rect 40664 132062 40670 132126
rect 40734 132062 40876 132126
rect 40664 132061 40876 132062
rect 40664 132005 40774 132061
rect 40830 132005 40876 132061
rect 40664 131920 40876 132005
rect 42432 132126 42644 132132
rect 42432 132062 42438 132126
rect 42502 132062 42644 132126
rect 42432 132061 42644 132062
rect 42432 132005 42454 132061
rect 42510 132005 42644 132061
rect 42432 131920 42644 132005
rect 44064 132126 44276 132132
rect 44064 132062 44206 132126
rect 44270 132062 44276 132126
rect 44064 132061 44276 132062
rect 44064 132005 44134 132061
rect 44190 132005 44276 132061
rect 44064 131920 44276 132005
rect 45696 132126 45908 132132
rect 45696 132062 45702 132126
rect 45766 132062 45908 132126
rect 45696 132061 45908 132062
rect 45696 132005 45814 132061
rect 45870 132005 45908 132061
rect 45696 131920 45908 132005
rect 47464 132126 47676 132132
rect 47464 132062 47470 132126
rect 47534 132062 47676 132126
rect 47464 132061 47676 132062
rect 47464 132005 47494 132061
rect 47550 132005 47676 132061
rect 47464 131920 47676 132005
rect 49096 132126 49308 132132
rect 49096 132062 49102 132126
rect 49166 132062 49308 132126
rect 49096 132061 49308 132062
rect 49096 132005 49174 132061
rect 49230 132005 49308 132061
rect 49096 131920 49308 132005
rect 50728 132126 50940 132132
rect 50728 132062 50734 132126
rect 50798 132062 50940 132126
rect 50728 132061 50940 132062
rect 50728 132005 50854 132061
rect 50910 132005 50940 132061
rect 50728 131920 50940 132005
rect 52496 132126 52708 132132
rect 52496 132062 52638 132126
rect 52702 132062 52708 132126
rect 52496 132061 52708 132062
rect 52496 132005 52534 132061
rect 52590 132005 52708 132061
rect 52496 131920 52708 132005
rect 54128 132126 54340 132132
rect 54128 132062 54134 132126
rect 54198 132062 54340 132126
rect 54128 132061 54340 132062
rect 54128 132005 54214 132061
rect 54270 132005 54340 132061
rect 54128 131920 54340 132005
rect 55760 132126 55972 132132
rect 55760 132062 55902 132126
rect 55966 132062 55972 132126
rect 55760 132061 55972 132062
rect 55760 132005 55894 132061
rect 55950 132005 55972 132061
rect 55760 131920 55972 132005
rect 57528 132126 57740 132132
rect 57528 132062 57670 132126
rect 57734 132062 57740 132126
rect 57528 132061 57740 132062
rect 57528 132005 57574 132061
rect 57630 132005 57740 132061
rect 57528 131920 57740 132005
rect 59160 132126 59372 132132
rect 59160 132062 59166 132126
rect 59230 132062 59372 132126
rect 59160 132061 59372 132062
rect 59160 132005 59254 132061
rect 59310 132005 59372 132061
rect 59160 131920 59372 132005
rect 60792 132126 61140 132132
rect 60792 132062 61070 132126
rect 61134 132062 61140 132126
rect 60792 132061 61140 132062
rect 60792 132005 60934 132061
rect 60990 132005 61140 132061
rect 60792 131920 61140 132005
rect 62560 132126 62772 132132
rect 62560 132062 62702 132126
rect 62766 132062 62772 132126
rect 62560 132061 62772 132062
rect 62560 132005 62614 132061
rect 62670 132005 62772 132061
rect 62560 131920 62772 132005
rect 64192 132126 64404 132132
rect 64192 132062 64198 132126
rect 64262 132062 64404 132126
rect 64192 132061 64404 132062
rect 64192 132005 64294 132061
rect 64350 132005 64404 132061
rect 64192 131920 64404 132005
rect 65824 132126 66172 132132
rect 65824 132062 66102 132126
rect 66166 132062 66172 132126
rect 65824 132061 66172 132062
rect 65824 132005 65974 132061
rect 66030 132005 66172 132061
rect 65824 131920 66172 132005
rect 67592 132126 67804 132132
rect 67592 132062 67734 132126
rect 67798 132062 67804 132126
rect 67592 132061 67804 132062
rect 67592 132005 67654 132061
rect 67710 132005 67804 132061
rect 67592 131920 67804 132005
rect 69224 132126 69436 132132
rect 69224 132062 69230 132126
rect 69294 132062 69436 132126
rect 69224 132061 69436 132062
rect 69224 132005 69334 132061
rect 69390 132005 69436 132061
rect 69224 131920 69436 132005
rect 70992 132126 71204 132132
rect 70992 132062 71134 132126
rect 71198 132062 71204 132126
rect 70992 132061 71204 132062
rect 70992 132005 71014 132061
rect 71070 132005 71204 132061
rect 70992 131920 71204 132005
rect 72624 132126 72836 132132
rect 72624 132062 72630 132126
rect 72694 132062 72836 132126
rect 72624 132061 72836 132062
rect 72624 132005 72694 132061
rect 72750 132005 72836 132061
rect 72624 131920 72836 132005
rect 74256 132126 74468 132132
rect 74256 132062 74262 132126
rect 74326 132062 74468 132126
rect 74256 132061 74468 132062
rect 74256 132005 74374 132061
rect 74430 132005 74468 132061
rect 74256 131920 74468 132005
rect 76024 132126 76236 132132
rect 76024 132062 76166 132126
rect 76230 132062 76236 132126
rect 76024 132061 76236 132062
rect 76024 132005 76054 132061
rect 76110 132005 76236 132061
rect 76024 131920 76236 132005
rect 77656 132126 77868 132132
rect 77656 132062 77662 132126
rect 77726 132062 77868 132126
rect 77656 132061 77868 132062
rect 77656 132005 77734 132061
rect 77790 132005 77868 132061
rect 77656 131920 77868 132005
rect 79288 132126 79500 132132
rect 79288 132062 79294 132126
rect 79358 132062 79500 132126
rect 79288 132061 79500 132062
rect 79288 132005 79414 132061
rect 79470 132005 79500 132061
rect 79288 131920 79500 132005
rect 81056 132126 81268 132132
rect 81056 132062 81198 132126
rect 81262 132062 81268 132126
rect 81056 132061 81268 132062
rect 81056 132005 81094 132061
rect 81150 132005 81268 132061
rect 81056 131920 81268 132005
rect 82688 132126 82900 132132
rect 82688 132062 82694 132126
rect 82758 132062 82900 132126
rect 82688 132061 82900 132062
rect 82688 132005 82774 132061
rect 82830 132005 82900 132061
rect 82688 131920 82900 132005
rect 84320 132126 84532 132132
rect 84320 132062 84326 132126
rect 84390 132062 84532 132126
rect 84320 132061 84532 132062
rect 84320 132005 84454 132061
rect 84510 132005 84532 132061
rect 84320 131920 84532 132005
rect 86088 132126 86300 132132
rect 86088 132062 86094 132126
rect 86158 132062 86300 132126
rect 86088 132061 86300 132062
rect 86088 132005 86134 132061
rect 86190 132005 86300 132061
rect 86088 131920 86300 132005
rect 87720 132126 87932 132132
rect 87720 132062 87726 132126
rect 87790 132062 87932 132126
rect 87720 132061 87932 132062
rect 87720 132005 87814 132061
rect 87870 132005 87932 132061
rect 87720 131920 87932 132005
rect 89352 132126 89836 132132
rect 89352 132062 89766 132126
rect 89830 132062 89836 132126
rect 89352 132061 89836 132062
rect 89352 132005 89494 132061
rect 89550 132056 89836 132061
rect 91120 132126 91332 132132
rect 91120 132062 91126 132126
rect 91190 132062 91332 132126
rect 91120 132061 91332 132062
rect 89550 132005 89700 132056
rect 89352 131920 89700 132005
rect 91120 132005 91174 132061
rect 91230 132005 91332 132061
rect 91120 131920 91332 132005
rect 92752 132126 92964 132132
rect 92752 132062 92894 132126
rect 92958 132062 92964 132126
rect 92752 132061 92964 132062
rect 92752 132005 92854 132061
rect 92910 132005 92964 132061
rect 92752 131920 92964 132005
rect 94384 132126 94732 132132
rect 94384 132062 94662 132126
rect 94726 132062 94732 132126
rect 94384 132061 94732 132062
rect 94384 132005 94534 132061
rect 94590 132005 94732 132061
rect 94384 131920 94732 132005
rect 96152 132126 96364 132132
rect 96152 132062 96158 132126
rect 96222 132062 96364 132126
rect 96152 132061 96364 132062
rect 96152 132005 96214 132061
rect 96270 132005 96364 132061
rect 96152 131920 96364 132005
rect 97784 132126 97996 132132
rect 97784 132062 97926 132126
rect 97990 132062 97996 132126
rect 97784 132061 97996 132062
rect 97784 132005 97894 132061
rect 97950 132005 97996 132061
rect 97784 131920 97996 132005
rect 99552 132126 99764 132132
rect 99552 132062 99694 132126
rect 99758 132062 99764 132126
rect 99552 132061 99764 132062
rect 99552 132005 99574 132061
rect 99630 132005 99764 132061
rect 99552 131920 99764 132005
rect 101184 132126 101396 132132
rect 101184 132062 101190 132126
rect 101254 132062 101396 132126
rect 101184 132061 101396 132062
rect 101184 132005 101254 132061
rect 101310 132005 101396 132061
rect 101184 131920 101396 132005
rect 102816 132126 103028 132132
rect 102816 132062 102958 132126
rect 103022 132062 103028 132126
rect 102816 132061 103028 132062
rect 102816 132005 102934 132061
rect 102990 132005 103028 132061
rect 102816 131920 103028 132005
rect 104584 132126 104796 132132
rect 104584 132062 104726 132126
rect 104790 132062 104796 132126
rect 104584 132061 104796 132062
rect 104584 132005 104614 132061
rect 104670 132005 104796 132061
rect 104584 131920 104796 132005
rect 106216 132126 106428 132132
rect 106216 132062 106222 132126
rect 106286 132062 106428 132126
rect 106216 132061 106428 132062
rect 106216 132005 106294 132061
rect 106350 132005 106428 132061
rect 106216 131920 106428 132005
rect 107848 132126 108060 132132
rect 107848 132062 107854 132126
rect 107918 132062 108060 132126
rect 107848 132061 108060 132062
rect 107848 132005 107974 132061
rect 108030 132005 108060 132061
rect 107848 131920 108060 132005
rect 109616 132126 109828 132132
rect 109616 132062 109622 132126
rect 109686 132062 109828 132126
rect 109616 132061 109828 132062
rect 109616 132005 109654 132061
rect 109710 132005 109828 132061
rect 109616 131920 109828 132005
rect 111248 132126 111460 132132
rect 111248 132062 111390 132126
rect 111454 132062 111460 132126
rect 111248 132061 111460 132062
rect 111248 132005 111334 132061
rect 111390 132005 111460 132061
rect 111248 131920 111460 132005
rect 112880 132126 113092 132132
rect 112880 132062 112886 132126
rect 112950 132062 113092 132126
rect 112880 132061 113092 132062
rect 112880 132005 113014 132061
rect 113070 132005 113092 132061
rect 112880 131920 113092 132005
rect 114648 132126 114860 132132
rect 114648 132062 114654 132126
rect 114718 132062 114860 132126
rect 114648 132061 114860 132062
rect 114648 132005 114694 132061
rect 114750 132005 114860 132061
rect 114648 131920 114860 132005
rect 116280 132126 116492 132132
rect 116280 132062 116422 132126
rect 116486 132062 116492 132126
rect 116280 132061 116492 132062
rect 116280 132005 116374 132061
rect 116430 132005 116492 132061
rect 116280 131920 116492 132005
rect 117912 132126 118260 132132
rect 117912 132062 117918 132126
rect 117982 132062 118260 132126
rect 117912 132061 118260 132062
rect 117912 132005 118054 132061
rect 118110 132005 118260 132061
rect 117912 131920 118260 132005
rect 119680 132126 119892 132132
rect 119680 132062 119686 132126
rect 119750 132062 119892 132126
rect 119680 132061 119892 132062
rect 119680 132005 119734 132061
rect 119790 132005 119892 132061
rect 119680 131990 119892 132005
rect 119680 131926 119686 131990
rect 119750 131926 119892 131990
rect 119680 131920 119892 131926
rect 121312 132126 121524 132132
rect 121312 132062 121454 132126
rect 121518 132062 121524 132126
rect 121312 132061 121524 132062
rect 121312 132005 121414 132061
rect 121470 132005 121524 132061
rect 121312 131920 121524 132005
rect 122944 132126 123292 132132
rect 122944 132062 123086 132126
rect 123150 132062 123292 132126
rect 122944 132061 123292 132062
rect 122944 132005 123094 132061
rect 123150 132005 123292 132061
rect 122944 131920 123292 132005
rect 124712 132126 124924 132132
rect 124712 132062 124718 132126
rect 124782 132062 124924 132126
rect 124712 132061 124924 132062
rect 124712 132005 124774 132061
rect 124830 132005 124924 132061
rect 124712 131920 124924 132005
rect 126344 132126 126556 132132
rect 126344 132062 126350 132126
rect 126414 132062 126556 132126
rect 126344 132061 126556 132062
rect 126344 132005 126454 132061
rect 126510 132005 126556 132061
rect 126344 131920 126556 132005
rect 128112 132126 128324 132132
rect 128112 132062 128118 132126
rect 128182 132062 128324 132126
rect 128112 132061 128324 132062
rect 128112 132005 128134 132061
rect 128190 132005 128324 132061
rect 128112 131920 128324 132005
rect 129744 132126 129956 132132
rect 129744 132062 129886 132126
rect 129950 132062 129956 132126
rect 129744 132061 129956 132062
rect 129744 132005 129814 132061
rect 129870 132005 129956 132061
rect 129744 131920 129956 132005
rect 131376 132126 131588 132132
rect 131376 132062 131382 132126
rect 131446 132062 131588 132126
rect 131376 132061 131588 132062
rect 131376 132005 131494 132061
rect 131550 132005 131588 132061
rect 131376 131920 131588 132005
rect 133144 132126 133356 132132
rect 133144 132062 133150 132126
rect 133214 132062 133356 132126
rect 133144 132061 133356 132062
rect 133144 132005 133174 132061
rect 133230 132005 133356 132061
rect 133144 131920 133356 132005
rect 134776 132126 134988 132132
rect 134776 132062 134918 132126
rect 134982 132062 134988 132126
rect 134776 132061 134988 132062
rect 134776 132005 134854 132061
rect 134910 132005 134988 132061
rect 134776 131920 134988 132005
rect 136408 132126 136620 132132
rect 136408 132062 136414 132126
rect 136478 132062 136620 132126
rect 136408 132061 136620 132062
rect 136408 132005 136534 132061
rect 136590 132005 136620 132061
rect 136408 131996 136620 132005
rect 136408 131990 136892 131996
rect 136408 131926 136822 131990
rect 136886 131926 136892 131990
rect 136408 131920 136892 131926
rect 1768 131582 2116 131588
rect 1768 131518 2046 131582
rect 2110 131518 2116 131582
rect 1768 131512 2116 131518
rect 136816 131582 137028 131588
rect 136816 131518 136822 131582
rect 136886 131518 137028 131582
rect 1768 131448 1980 131512
rect 1768 131392 1798 131448
rect 1854 131392 1980 131448
rect 1768 131240 1980 131392
rect 119408 131446 120844 131452
rect 119408 131382 120638 131446
rect 120702 131382 120844 131446
rect 119408 131376 120844 131382
rect 119408 131310 119620 131376
rect 119408 131246 119550 131310
rect 119614 131246 119620 131310
rect 119408 131240 119620 131246
rect 120632 131240 120844 131376
rect 136816 131448 137028 131518
rect 136816 131392 136944 131448
rect 137000 131392 137028 131448
rect 136816 131240 137028 131392
rect 123527 131083 123593 131086
rect 120140 131081 123593 131083
rect 120140 131025 123532 131081
rect 123588 131025 123593 131081
rect 120140 131023 123593 131025
rect 123527 131020 123593 131023
rect 119816 130902 120028 130908
rect 119816 130838 119958 130902
rect 120022 130838 120028 130902
rect 119816 130825 120028 130838
rect 119816 130769 119942 130825
rect 119998 130769 120028 130825
rect 119816 130696 120028 130769
rect 121040 130902 121252 130908
rect 121040 130838 121182 130902
rect 121246 130838 121252 130902
rect 121040 130825 121252 130838
rect 121040 130769 121110 130825
rect 121166 130769 121252 130825
rect 121040 130696 121252 130769
rect 123624 130494 123836 130500
rect 123624 130430 123630 130494
rect 123694 130430 123836 130494
rect 123624 130358 123836 130430
rect 123624 130294 123766 130358
rect 123830 130294 123836 130358
rect 123624 130288 123836 130294
rect 136000 130494 138252 130500
rect 136000 130430 138182 130494
rect 138246 130430 138252 130494
rect 136000 130424 138252 130430
rect 136000 130288 136348 130424
rect 119408 130086 119756 130092
rect 119408 130022 119686 130086
rect 119750 130022 119756 130086
rect 119408 130016 119756 130022
rect 119408 129956 119620 130016
rect 120632 129956 120844 130092
rect 119408 129950 123700 129956
rect 119408 129886 119414 129950
rect 119478 129886 123630 129950
rect 123694 129886 123700 129950
rect 119408 129880 123700 129886
rect 135864 129880 138796 129956
rect 135864 129828 136076 129880
rect 1224 129814 1980 129820
rect 1224 129750 1230 129814
rect 1294 129768 1980 129814
rect 1294 129750 1798 129768
rect 1224 129744 1798 129750
rect 1768 129712 1798 129744
rect 1854 129712 1980 129768
rect 1768 129608 1980 129712
rect 132736 129814 132948 129820
rect 132736 129750 132742 129814
rect 132806 129750 132948 129814
rect 132736 129723 132948 129750
rect 135864 129772 135984 129828
rect 136040 129772 136076 129828
rect 135864 129744 136076 129772
rect 136816 129814 137572 129820
rect 136816 129768 137502 129814
rect 132736 129667 132847 129723
rect 132903 129667 132948 129723
rect 132736 129608 132948 129667
rect 136816 129712 136944 129768
rect 137000 129750 137502 129768
rect 137566 129750 137572 129814
rect 137000 129744 137572 129750
rect 137000 129712 137028 129744
rect 136816 129608 137028 129712
rect 116280 129140 116492 129276
rect 117368 129270 119620 129276
rect 117368 129206 119550 129270
rect 119614 129206 119620 129270
rect 117368 129200 119620 129206
rect 117368 129140 117580 129200
rect 116280 129134 117580 129140
rect 116280 129070 117510 129134
rect 117574 129070 117580 129134
rect 116280 129064 117580 129070
rect 123624 128998 123836 129004
rect 123624 128934 123630 128998
rect 123694 128934 123836 128998
rect 123624 128862 123836 128934
rect 123624 128798 123630 128862
rect 123694 128798 123836 128862
rect 123624 128792 123836 128798
rect 136000 128868 136348 129004
rect 136000 128862 136892 128868
rect 136000 128798 136822 128862
rect 136886 128798 136892 128862
rect 136000 128792 136892 128798
rect 1224 128182 1980 128188
rect 1224 128118 1230 128182
rect 1294 128118 1980 128182
rect 1224 128112 1980 128118
rect 1768 128088 1980 128112
rect 1768 128032 1798 128088
rect 1854 128032 1980 128088
rect 1768 127976 1980 128032
rect 136816 128182 137572 128188
rect 136816 128118 136822 128182
rect 136886 128118 137502 128182
rect 137566 128118 137572 128182
rect 136816 128112 137572 128118
rect 136816 128088 137028 128112
rect 136816 128032 136944 128088
rect 137000 128032 137028 128088
rect 136816 127976 137028 128032
rect 116280 127780 116492 127916
rect 117368 127910 119484 127916
rect 117368 127846 119414 127910
rect 119478 127846 119484 127910
rect 117368 127840 119484 127846
rect 117368 127780 117580 127840
rect 29920 127647 29996 127780
rect 32368 127647 32444 127780
rect 34816 127647 34892 127780
rect 29512 127638 29724 127644
rect 29512 127607 29654 127638
rect 29512 127551 29562 127607
rect 29618 127574 29654 127607
rect 29718 127574 29724 127638
rect 29618 127551 29724 127574
rect 29512 127432 29724 127551
rect 29795 127549 29996 127647
rect 29920 127502 29996 127549
rect 29920 127438 29926 127502
rect 29990 127438 29996 127502
rect 29920 127432 29996 127438
rect 31960 127638 32172 127644
rect 31960 127574 31966 127638
rect 32030 127607 32172 127638
rect 32030 127574 32058 127607
rect 31960 127551 32058 127574
rect 32114 127551 32172 127607
rect 31960 127432 32172 127551
rect 32291 127549 32444 127647
rect 32368 127508 32444 127549
rect 34408 127638 34620 127644
rect 34408 127574 34550 127638
rect 34614 127628 34620 127638
rect 34614 127574 34631 127628
rect 34408 127551 34554 127574
rect 34610 127551 34631 127574
rect 34408 127530 34631 127551
rect 34787 127549 34892 127647
rect 32368 127502 32580 127508
rect 32368 127438 32510 127502
rect 32574 127438 32580 127502
rect 32368 127432 32580 127438
rect 34408 127432 34620 127530
rect 34816 127508 34892 127549
rect 36992 127638 37204 127644
rect 36992 127574 36998 127638
rect 37062 127607 37204 127638
rect 36992 127551 37050 127574
rect 37106 127551 37204 127607
rect 34816 127502 35028 127508
rect 34816 127438 34958 127502
rect 35022 127438 35028 127502
rect 34816 127432 35028 127438
rect 36992 127432 37204 127551
rect 37264 127502 37476 127780
rect 37264 127438 37270 127502
rect 37334 127438 37476 127502
rect 37264 127432 37476 127438
rect 39440 127638 39652 127644
rect 39440 127607 39582 127638
rect 39440 127551 39546 127607
rect 39646 127574 39652 127638
rect 39602 127551 39652 127574
rect 39440 127432 39652 127551
rect 39712 127508 39924 127780
rect 42296 127647 42508 127780
rect 44880 127647 44956 127780
rect 47328 127647 47404 127780
rect 49776 127647 49988 127780
rect 41888 127638 42100 127644
rect 41888 127574 42030 127638
rect 42094 127628 42100 127638
rect 42094 127607 42119 127628
rect 41888 127551 42042 127574
rect 42098 127551 42119 127607
rect 41888 127530 42119 127551
rect 42275 127549 42508 127647
rect 39712 127502 40060 127508
rect 39712 127438 39990 127502
rect 40054 127438 40060 127502
rect 39712 127432 40060 127438
rect 41888 127432 42100 127530
rect 42296 127502 42508 127549
rect 42296 127438 42438 127502
rect 42502 127438 42508 127502
rect 42296 127432 42508 127438
rect 44472 127638 44684 127644
rect 44472 127607 44614 127638
rect 44472 127551 44538 127607
rect 44594 127574 44614 127607
rect 44678 127574 44684 127638
rect 44594 127551 44684 127574
rect 44472 127432 44684 127551
rect 44771 127549 44956 127647
rect 44880 127502 44956 127549
rect 44880 127438 44886 127502
rect 44950 127438 44956 127502
rect 44880 127432 44956 127438
rect 46920 127638 47132 127644
rect 46920 127607 47062 127638
rect 46920 127551 47034 127607
rect 47126 127574 47132 127638
rect 47090 127551 47132 127574
rect 46920 127432 47132 127551
rect 47267 127549 47404 127647
rect 47328 127502 47404 127549
rect 47328 127438 47334 127502
rect 47398 127438 47404 127502
rect 47328 127432 47404 127438
rect 49504 127638 49580 127644
rect 49504 127574 49510 127638
rect 49574 127628 49580 127638
rect 49574 127607 49607 127628
rect 49504 127551 49530 127574
rect 49586 127551 49607 127607
rect 49504 127530 49607 127551
rect 49763 127549 49988 127647
rect 49504 127432 49580 127530
rect 49776 127502 49988 127549
rect 49776 127438 49918 127502
rect 49982 127438 49988 127502
rect 49776 127432 49988 127438
rect 51952 127638 52164 127644
rect 51952 127574 51958 127638
rect 52022 127607 52164 127638
rect 52022 127574 52026 127607
rect 51952 127551 52026 127574
rect 52082 127551 52164 127607
rect 51952 127432 52164 127551
rect 52224 127502 52436 127780
rect 54808 127647 54884 127780
rect 57256 127647 57468 127780
rect 59840 127647 59916 127780
rect 62288 127647 62364 127780
rect 52224 127438 52366 127502
rect 52430 127438 52436 127502
rect 52224 127432 52436 127438
rect 54400 127638 54612 127644
rect 54400 127574 54406 127638
rect 54470 127607 54612 127638
rect 54470 127574 54522 127607
rect 54400 127551 54522 127574
rect 54578 127551 54612 127607
rect 54400 127432 54612 127551
rect 54755 127549 54884 127647
rect 54808 127508 54884 127549
rect 56984 127638 57060 127644
rect 56984 127574 56990 127638
rect 57054 127628 57060 127638
rect 57054 127607 57095 127628
rect 56984 127551 57018 127574
rect 57074 127551 57095 127607
rect 56984 127530 57095 127551
rect 57251 127549 57468 127647
rect 54808 127502 55020 127508
rect 54808 127438 54950 127502
rect 55014 127438 55020 127502
rect 54808 127432 55020 127438
rect 56984 127432 57060 127530
rect 57256 127502 57468 127549
rect 57256 127438 57398 127502
rect 57462 127438 57468 127502
rect 57256 127432 57468 127438
rect 59432 127638 59644 127644
rect 59432 127607 59574 127638
rect 59432 127551 59514 127607
rect 59570 127574 59574 127607
rect 59638 127574 59644 127638
rect 59570 127551 59644 127574
rect 59432 127432 59644 127551
rect 59747 127549 59916 127647
rect 59840 127502 59916 127549
rect 59840 127438 59846 127502
rect 59910 127438 59916 127502
rect 59840 127432 59916 127438
rect 61880 127638 62092 127644
rect 61880 127607 62022 127638
rect 61880 127551 62010 127607
rect 62086 127574 62092 127638
rect 62066 127551 62092 127574
rect 61880 127432 62092 127551
rect 62243 127549 62364 127647
rect 62288 127508 62364 127549
rect 64464 127638 64676 127644
rect 64464 127607 64606 127638
rect 64464 127551 64506 127607
rect 64562 127574 64606 127607
rect 64670 127574 64676 127638
rect 64562 127551 64676 127574
rect 62288 127502 62500 127508
rect 62288 127438 62430 127502
rect 62494 127438 62500 127502
rect 62288 127432 62500 127438
rect 64464 127432 64676 127551
rect 64736 127502 64948 127780
rect 67320 127647 67396 127780
rect 69768 127647 69844 127780
rect 72352 127647 72428 127780
rect 74800 127647 74876 127780
rect 77248 127647 77324 127780
rect 79832 127647 79908 127780
rect 82280 127647 82356 127780
rect 84728 127647 84940 127780
rect 87312 127647 87388 127780
rect 89760 127647 89836 127780
rect 92208 127647 92420 127780
rect 94792 127647 94868 127780
rect 97240 127647 97316 127780
rect 99552 127704 99900 127780
rect 64736 127438 64742 127502
rect 64806 127438 64948 127502
rect 64736 127432 64948 127438
rect 66912 127638 67124 127644
rect 66912 127607 67054 127638
rect 66912 127551 67002 127607
rect 67118 127574 67124 127638
rect 67058 127551 67124 127574
rect 66912 127432 67124 127551
rect 67235 127549 67396 127647
rect 67320 127502 67396 127549
rect 67320 127438 67326 127502
rect 67390 127438 67396 127502
rect 67320 127432 67396 127438
rect 69360 127638 69572 127644
rect 69360 127574 69366 127638
rect 69430 127628 69572 127638
rect 69430 127607 69575 127628
rect 69430 127574 69498 127607
rect 69360 127551 69498 127574
rect 69554 127551 69575 127607
rect 69360 127530 69575 127551
rect 69731 127549 69844 127647
rect 69360 127432 69572 127530
rect 69768 127502 69844 127549
rect 69768 127438 69774 127502
rect 69838 127438 69844 127502
rect 69768 127432 69844 127438
rect 71944 127638 72156 127644
rect 71944 127607 72086 127638
rect 71944 127551 71994 127607
rect 72050 127574 72086 127607
rect 72150 127574 72156 127638
rect 72050 127551 72156 127574
rect 71944 127432 72156 127551
rect 72227 127549 72428 127647
rect 72352 127502 72428 127549
rect 72352 127438 72358 127502
rect 72422 127438 72428 127502
rect 72352 127432 72428 127438
rect 74392 127638 74604 127644
rect 74392 127574 74398 127638
rect 74462 127607 74604 127638
rect 74462 127574 74490 127607
rect 74392 127551 74490 127574
rect 74546 127551 74604 127607
rect 74392 127432 74604 127551
rect 74723 127549 74876 127647
rect 74800 127508 74876 127549
rect 76840 127638 77052 127644
rect 76840 127574 76982 127638
rect 77046 127628 77052 127638
rect 77046 127574 77063 127628
rect 76840 127551 76986 127574
rect 77042 127551 77063 127574
rect 76840 127530 77063 127551
rect 77219 127549 77324 127647
rect 74800 127502 75012 127508
rect 74800 127438 74942 127502
rect 75006 127438 75012 127502
rect 74800 127432 75012 127438
rect 76840 127432 77052 127530
rect 77248 127508 77324 127549
rect 79424 127638 79636 127644
rect 79424 127574 79430 127638
rect 79494 127607 79636 127638
rect 79424 127551 79482 127574
rect 79538 127551 79636 127607
rect 77248 127502 77460 127508
rect 77248 127438 77390 127502
rect 77454 127438 77460 127502
rect 77248 127432 77460 127438
rect 79424 127432 79636 127551
rect 79715 127549 79908 127647
rect 79832 127502 79908 127549
rect 79832 127438 79838 127502
rect 79902 127438 79908 127502
rect 79832 127432 79908 127438
rect 81872 127638 82084 127644
rect 81872 127607 82014 127638
rect 81872 127551 81978 127607
rect 82078 127574 82084 127638
rect 82034 127551 82084 127574
rect 81872 127432 82084 127551
rect 82211 127549 82356 127647
rect 82280 127508 82356 127549
rect 84320 127638 84532 127644
rect 84320 127574 84462 127638
rect 84526 127628 84532 127638
rect 84526 127607 84551 127628
rect 84320 127551 84474 127574
rect 84530 127551 84551 127607
rect 84320 127530 84551 127551
rect 84707 127549 84940 127647
rect 82280 127502 82492 127508
rect 82280 127438 82422 127502
rect 82486 127438 82492 127502
rect 82280 127432 82492 127438
rect 84320 127432 84532 127530
rect 84728 127502 84940 127549
rect 84728 127438 84870 127502
rect 84934 127438 84940 127502
rect 84728 127432 84940 127438
rect 86904 127638 87116 127644
rect 86904 127607 87046 127638
rect 86904 127551 86970 127607
rect 87026 127574 87046 127607
rect 87110 127574 87116 127638
rect 87026 127551 87116 127574
rect 86904 127432 87116 127551
rect 87203 127549 87388 127647
rect 87312 127502 87388 127549
rect 87312 127438 87318 127502
rect 87382 127438 87388 127502
rect 87312 127432 87388 127438
rect 89352 127638 89564 127644
rect 89352 127607 89494 127638
rect 89352 127551 89466 127607
rect 89558 127574 89564 127638
rect 89522 127551 89564 127574
rect 89352 127432 89564 127551
rect 89699 127549 89836 127647
rect 89760 127502 89836 127549
rect 89760 127438 89766 127502
rect 89830 127438 89836 127502
rect 89760 127432 89836 127438
rect 91936 127638 92012 127644
rect 91936 127574 91942 127638
rect 92006 127628 92012 127638
rect 92006 127607 92039 127628
rect 91936 127551 91962 127574
rect 92018 127551 92039 127607
rect 91936 127530 92039 127551
rect 92195 127549 92420 127647
rect 91936 127432 92012 127530
rect 92208 127502 92420 127549
rect 92208 127438 92350 127502
rect 92414 127438 92420 127502
rect 92208 127432 92420 127438
rect 94384 127638 94596 127644
rect 94384 127574 94390 127638
rect 94454 127607 94596 127638
rect 94454 127574 94458 127607
rect 94384 127551 94458 127574
rect 94514 127551 94596 127607
rect 94384 127432 94596 127551
rect 94691 127549 94868 127647
rect 94792 127502 94868 127549
rect 94792 127438 94798 127502
rect 94862 127438 94868 127502
rect 94792 127432 94868 127438
rect 96832 127638 97044 127644
rect 96832 127574 96838 127638
rect 96902 127607 97044 127638
rect 96902 127574 96954 127607
rect 96832 127551 96954 127574
rect 97010 127551 97044 127607
rect 96832 127432 97044 127551
rect 97187 127549 97316 127647
rect 97240 127508 97316 127549
rect 99416 127638 99492 127644
rect 99416 127574 99422 127638
rect 99486 127628 99492 127638
rect 99486 127607 99527 127628
rect 99416 127551 99450 127574
rect 99506 127551 99527 127607
rect 99416 127530 99527 127551
rect 99683 127549 99900 127704
rect 102272 127647 102348 127780
rect 104720 127647 104796 127780
rect 107304 127647 107380 127780
rect 116280 127774 117580 127780
rect 116280 127710 117374 127774
rect 117438 127710 117580 127774
rect 116280 127704 117580 127710
rect 97240 127502 97452 127508
rect 97240 127438 97382 127502
rect 97446 127438 97452 127502
rect 97240 127432 97452 127438
rect 99416 127432 99492 127530
rect 99688 127502 99900 127549
rect 99688 127438 99830 127502
rect 99894 127438 99900 127502
rect 99688 127432 99900 127438
rect 101864 127638 102076 127644
rect 101864 127607 102006 127638
rect 101864 127551 101946 127607
rect 102002 127574 102006 127607
rect 102070 127574 102076 127638
rect 102002 127551 102076 127574
rect 101864 127432 102076 127551
rect 102179 127549 102348 127647
rect 102272 127502 102348 127549
rect 102272 127438 102278 127502
rect 102342 127438 102348 127502
rect 102272 127432 102348 127438
rect 104312 127638 104524 127644
rect 104312 127607 104454 127638
rect 104312 127551 104442 127607
rect 104518 127574 104524 127638
rect 104498 127551 104524 127574
rect 104312 127432 104524 127551
rect 104675 127549 104796 127647
rect 104720 127508 104796 127549
rect 106896 127638 107108 127644
rect 106896 127607 107038 127638
rect 106896 127551 106938 127607
rect 106994 127574 107038 127607
rect 107102 127574 107108 127638
rect 106994 127551 107108 127574
rect 104720 127502 104932 127508
rect 104720 127438 104862 127502
rect 104926 127438 104932 127502
rect 104720 127432 104932 127438
rect 106896 127432 107108 127551
rect 107171 127549 107380 127647
rect 107304 127502 107380 127549
rect 107304 127438 107310 127502
rect 107374 127438 107380 127502
rect 107304 127432 107380 127438
rect 123624 127638 123836 127644
rect 123624 127574 123766 127638
rect 123830 127574 123836 127638
rect 123624 127508 123836 127574
rect 123624 127502 123934 127508
rect 123624 127438 123902 127502
rect 123966 127438 123972 127502
rect 123624 127432 123934 127438
rect 29784 127236 29996 127372
rect 29784 127230 32172 127236
rect 29784 127166 29790 127230
rect 29854 127166 32102 127230
rect 32166 127166 32172 127230
rect 29784 127160 32172 127166
rect 32232 127230 32444 127372
rect 32232 127166 32374 127230
rect 32438 127166 32444 127230
rect 32232 127160 32444 127166
rect 34680 127230 34892 127372
rect 37264 127236 37476 127372
rect 37166 127230 37476 127236
rect 34680 127166 34822 127230
rect 34886 127166 34892 127230
rect 37128 127166 37134 127230
rect 37198 127166 37406 127230
rect 37470 127166 37476 127230
rect 34680 127160 34892 127166
rect 37166 127160 37476 127166
rect 39712 127230 39924 127372
rect 39712 127166 39854 127230
rect 39918 127166 39924 127230
rect 39712 127160 39924 127166
rect 42160 127296 44956 127372
rect 42160 127230 42508 127296
rect 42160 127166 42166 127230
rect 42230 127166 42508 127230
rect 42160 127160 42508 127166
rect 44744 127230 44956 127296
rect 44744 127166 44886 127230
rect 44950 127166 44956 127230
rect 44744 127160 44956 127166
rect 47192 127236 47404 127372
rect 49640 127236 49988 127372
rect 52224 127296 54884 127372
rect 52224 127236 52436 127296
rect 47192 127230 49580 127236
rect 47192 127166 47198 127230
rect 47262 127166 49510 127230
rect 49574 127166 49580 127230
rect 47192 127160 49580 127166
rect 49640 127230 52436 127236
rect 49640 127166 49782 127230
rect 49846 127166 52230 127230
rect 52294 127166 52436 127230
rect 49640 127160 52436 127166
rect 54672 127230 54884 127296
rect 57120 127236 57468 127372
rect 59704 127236 59916 127372
rect 57022 127230 57468 127236
rect 59606 127230 59916 127236
rect 54672 127166 54814 127230
rect 54878 127166 54884 127230
rect 56984 127166 56990 127230
rect 57054 127166 57262 127230
rect 57326 127166 57468 127230
rect 59568 127166 59574 127230
rect 59638 127166 59846 127230
rect 59910 127166 59916 127230
rect 54672 127160 54884 127166
rect 57022 127160 57468 127166
rect 59606 127160 59916 127166
rect 62152 127230 62364 127372
rect 62152 127166 62294 127230
rect 62358 127166 62364 127230
rect 62152 127160 62364 127166
rect 64736 127236 64948 127372
rect 67184 127296 72428 127372
rect 64736 127230 67124 127236
rect 64736 127166 64878 127230
rect 64942 127166 67054 127230
rect 67118 127166 67124 127230
rect 64736 127160 67124 127166
rect 67184 127230 67396 127296
rect 67184 127166 67190 127230
rect 67254 127166 67396 127230
rect 67184 127160 67396 127166
rect 69632 127230 69844 127296
rect 69632 127166 69638 127230
rect 69702 127166 69844 127230
rect 69632 127160 69844 127166
rect 72216 127236 72428 127296
rect 72216 127230 74604 127236
rect 72216 127166 72222 127230
rect 72286 127166 74534 127230
rect 74598 127166 74604 127230
rect 72216 127160 74604 127166
rect 74664 127230 74876 127372
rect 74664 127166 74806 127230
rect 74870 127166 74876 127230
rect 74664 127160 74876 127166
rect 77112 127230 77324 127372
rect 79696 127236 79908 127372
rect 82144 127236 82356 127372
rect 84592 127296 87388 127372
rect 84592 127236 84940 127296
rect 79598 127230 79908 127236
rect 82046 127230 82356 127236
rect 84494 127230 84940 127236
rect 77112 127166 77254 127230
rect 77318 127166 77324 127230
rect 79560 127166 79566 127230
rect 79630 127166 79838 127230
rect 79902 127166 79908 127230
rect 82008 127166 82014 127230
rect 82078 127166 82286 127230
rect 82350 127166 82356 127230
rect 84456 127166 84462 127230
rect 84526 127166 84598 127230
rect 84662 127166 84940 127230
rect 77112 127160 77324 127166
rect 79598 127160 79908 127166
rect 82046 127160 82356 127166
rect 84494 127160 84940 127166
rect 87176 127230 87388 127296
rect 87176 127166 87318 127230
rect 87382 127166 87388 127230
rect 87176 127160 87388 127166
rect 89624 127236 89836 127372
rect 92072 127236 92420 127372
rect 94656 127296 97316 127372
rect 94656 127236 94868 127296
rect 89624 127230 94868 127236
rect 89624 127166 89630 127230
rect 89694 127166 92214 127230
rect 92278 127166 94662 127230
rect 94726 127166 94868 127230
rect 89624 127160 94868 127166
rect 97104 127230 97316 127296
rect 99552 127236 99900 127372
rect 99454 127230 99900 127236
rect 97104 127166 97246 127230
rect 97310 127166 97316 127230
rect 99416 127166 99422 127230
rect 99486 127166 99694 127230
rect 99758 127166 99900 127230
rect 97104 127160 97316 127166
rect 99454 127160 99900 127166
rect 102136 127230 102348 127372
rect 102136 127166 102278 127230
rect 102342 127166 102348 127230
rect 102136 127160 102348 127166
rect 104584 127230 104796 127372
rect 104584 127166 104726 127230
rect 104790 127166 104796 127230
rect 104584 127160 104796 127166
rect 107168 127230 107380 127372
rect 107168 127166 107174 127230
rect 107238 127166 107380 127230
rect 107168 127160 107380 127166
rect 1768 126420 1980 126556
rect 1224 126414 1980 126420
rect 1224 126350 1230 126414
rect 1294 126408 1980 126414
rect 1294 126352 1798 126408
rect 1854 126352 1980 126408
rect 1294 126350 1980 126352
rect 1224 126344 1980 126350
rect 29648 126550 29996 126556
rect 32134 126550 32444 126556
rect 29648 126486 29790 126550
rect 29854 126486 29996 126550
rect 32096 126486 32102 126550
rect 32166 126486 32374 126550
rect 32438 126486 32444 126550
rect 29648 126344 29996 126486
rect 32134 126480 32444 126486
rect 32232 126420 32444 126480
rect 34680 126550 37204 126556
rect 34680 126486 34822 126550
rect 34886 126486 37134 126550
rect 37198 126486 37204 126550
rect 34680 126480 37204 126486
rect 37264 126550 42372 126556
rect 37264 126486 37406 126550
rect 37470 126486 39854 126550
rect 39918 126486 42166 126550
rect 42230 126486 42372 126550
rect 37264 126480 42372 126486
rect 34680 126420 34892 126480
rect 32232 126344 34892 126420
rect 37264 126344 37476 126480
rect 39712 126344 39924 126480
rect 42160 126344 42372 126480
rect 44744 126550 44956 126556
rect 44744 126486 44886 126550
rect 44950 126486 44956 126550
rect 44744 126420 44956 126486
rect 47192 126550 47404 126556
rect 49542 126550 49852 126556
rect 47192 126486 47198 126550
rect 47262 126486 47404 126550
rect 49504 126486 49510 126550
rect 49574 126486 49782 126550
rect 49846 126486 49852 126550
rect 47192 126420 47404 126486
rect 49542 126480 49852 126486
rect 44744 126344 47404 126420
rect 49640 126344 49852 126480
rect 52224 126550 52436 126556
rect 52224 126486 52230 126550
rect 52294 126486 52436 126550
rect 52224 126344 52436 126486
rect 54672 126550 57060 126556
rect 54672 126486 54814 126550
rect 54878 126486 56990 126550
rect 57054 126486 57060 126550
rect 54672 126480 57060 126486
rect 57120 126550 59644 126556
rect 57120 126486 57262 126550
rect 57326 126486 59574 126550
rect 59638 126486 59644 126550
rect 57120 126480 59644 126486
rect 59704 126550 59916 126556
rect 59704 126486 59846 126550
rect 59910 126486 59916 126550
rect 54672 126344 54884 126480
rect 57120 126344 57468 126480
rect 59704 126420 59916 126486
rect 62152 126550 62364 126556
rect 62152 126486 62294 126550
rect 62358 126486 62364 126550
rect 62152 126420 62364 126486
rect 64600 126550 64948 126556
rect 67086 126550 67396 126556
rect 64600 126486 64878 126550
rect 64942 126486 64948 126550
rect 67048 126486 67054 126550
rect 67118 126486 67190 126550
rect 67254 126486 67396 126550
rect 64600 126420 64948 126486
rect 67086 126480 67396 126486
rect 59704 126344 64948 126420
rect 67184 126344 67396 126480
rect 69632 126550 69844 126556
rect 69632 126486 69638 126550
rect 69702 126486 69844 126550
rect 69632 126344 69844 126486
rect 72080 126550 72428 126556
rect 74566 126550 74876 126556
rect 72080 126486 72222 126550
rect 72286 126486 72428 126550
rect 74528 126486 74534 126550
rect 74598 126486 74806 126550
rect 74870 126486 74876 126550
rect 72080 126344 72428 126486
rect 74566 126480 74876 126486
rect 74664 126420 74876 126480
rect 77112 126550 79636 126556
rect 77112 126486 77254 126550
rect 77318 126486 79566 126550
rect 79630 126486 79636 126550
rect 77112 126480 79636 126486
rect 79696 126550 82084 126556
rect 79696 126486 79838 126550
rect 79902 126486 82014 126550
rect 82078 126486 82084 126550
rect 79696 126480 82084 126486
rect 82144 126550 84532 126556
rect 82144 126486 82286 126550
rect 82350 126486 84462 126550
rect 84526 126486 84532 126550
rect 82144 126480 84532 126486
rect 84592 126550 84804 126556
rect 84592 126486 84598 126550
rect 84662 126486 84804 126550
rect 77112 126420 77324 126480
rect 74664 126344 77324 126420
rect 79696 126344 79908 126480
rect 82144 126344 82356 126480
rect 84592 126344 84804 126486
rect 87176 126550 89836 126556
rect 87176 126486 87318 126550
rect 87382 126486 89630 126550
rect 89694 126486 89836 126550
rect 87176 126480 89836 126486
rect 87176 126420 87388 126480
rect 87176 126414 87932 126420
rect 87176 126350 87862 126414
rect 87926 126350 87932 126414
rect 87176 126344 87932 126350
rect 89624 126344 89836 126480
rect 92072 126550 92284 126556
rect 92072 126486 92214 126550
rect 92278 126486 92284 126550
rect 92072 126344 92284 126486
rect 94656 126550 94868 126556
rect 94656 126486 94662 126550
rect 94726 126486 94868 126550
rect 94656 126344 94868 126486
rect 97104 126550 99492 126556
rect 97104 126486 97246 126550
rect 97310 126486 99422 126550
rect 99486 126486 99492 126550
rect 97104 126480 99492 126486
rect 99552 126550 102348 126556
rect 99552 126486 99694 126550
rect 99758 126486 102278 126550
rect 102342 126486 102348 126550
rect 99552 126480 102348 126486
rect 97104 126344 97316 126480
rect 99552 126344 99900 126480
rect 102136 126420 102348 126480
rect 104584 126550 104796 126556
rect 104584 126486 104726 126550
rect 104790 126486 104796 126550
rect 104584 126420 104796 126486
rect 107032 126550 107380 126556
rect 107032 126486 107174 126550
rect 107238 126486 107380 126550
rect 107032 126420 107380 126486
rect 136816 126550 137572 126556
rect 136816 126486 137502 126550
rect 137566 126486 137572 126550
rect 136816 126480 137572 126486
rect 102136 126344 107380 126420
rect 116280 126414 117580 126420
rect 116280 126350 117510 126414
rect 117574 126350 117580 126414
rect 116280 126344 117580 126350
rect 1768 126208 1980 126344
rect 116280 126284 116492 126344
rect 116280 126278 117308 126284
rect 116280 126214 117238 126278
rect 117302 126214 117308 126278
rect 116280 126208 117308 126214
rect 117368 126208 117580 126344
rect 136816 126408 137028 126480
rect 136816 126352 136944 126408
rect 137000 126352 137028 126408
rect 123624 126278 123836 126284
rect 123624 126214 123630 126278
rect 123694 126214 123836 126278
rect 123624 126142 123836 126214
rect 136816 126208 137028 126352
rect 123624 126078 123766 126142
rect 123830 126078 123836 126142
rect 123624 126072 123836 126078
rect 29784 125734 30132 125740
rect 29784 125670 29926 125734
rect 29990 125670 30062 125734
rect 30126 125670 30132 125734
rect 29784 125664 30132 125670
rect 32232 125734 32716 125740
rect 32232 125670 32510 125734
rect 32574 125670 32646 125734
rect 32710 125670 32716 125734
rect 32232 125664 32716 125670
rect 34816 125734 35164 125740
rect 34816 125670 34958 125734
rect 35022 125670 35094 125734
rect 35158 125670 35164 125734
rect 34816 125664 35164 125670
rect 37264 125734 37476 125740
rect 37264 125670 37270 125734
rect 37334 125670 37406 125734
rect 37470 125670 37476 125734
rect 37264 125664 37476 125670
rect 39848 125734 40196 125740
rect 39848 125670 39990 125734
rect 40054 125670 40126 125734
rect 40190 125670 40196 125734
rect 39848 125664 40196 125670
rect 42296 125734 42644 125740
rect 42296 125670 42438 125734
rect 42502 125670 42574 125734
rect 42638 125670 42644 125734
rect 42296 125664 42644 125670
rect 44744 125734 44956 125740
rect 44744 125670 44750 125734
rect 44814 125670 44886 125734
rect 44950 125670 44956 125734
rect 44744 125664 44956 125670
rect 47328 125734 47540 125740
rect 47328 125670 47334 125734
rect 47398 125670 47470 125734
rect 47534 125670 47540 125734
rect 47328 125664 47540 125670
rect 49776 125734 50124 125740
rect 49776 125670 49918 125734
rect 49982 125670 50054 125734
rect 50118 125670 50124 125734
rect 49776 125664 50124 125670
rect 52224 125734 52572 125740
rect 52224 125670 52366 125734
rect 52430 125670 52502 125734
rect 52566 125670 52572 125734
rect 52224 125664 52572 125670
rect 54808 125734 55156 125740
rect 54808 125670 54950 125734
rect 55014 125670 55086 125734
rect 55150 125670 55156 125734
rect 54808 125664 55156 125670
rect 57256 125734 57604 125740
rect 57256 125670 57398 125734
rect 57462 125670 57534 125734
rect 57598 125670 57604 125734
rect 57256 125664 57604 125670
rect 59704 125734 60052 125740
rect 59704 125670 59710 125734
rect 59774 125670 59982 125734
rect 60046 125670 60052 125734
rect 59704 125664 60052 125670
rect 62288 125734 62636 125740
rect 62288 125670 62430 125734
rect 62494 125670 62566 125734
rect 62630 125670 62636 125734
rect 62288 125664 62636 125670
rect 64736 125734 64948 125740
rect 64736 125670 64742 125734
rect 64806 125670 64878 125734
rect 64942 125670 64948 125734
rect 64736 125664 64948 125670
rect 67184 125734 67532 125740
rect 67184 125670 67326 125734
rect 67390 125670 67462 125734
rect 67526 125670 67532 125734
rect 67184 125664 67532 125670
rect 69768 125734 69980 125740
rect 69768 125670 69774 125734
rect 69838 125670 69910 125734
rect 69974 125670 69980 125734
rect 69768 125664 69980 125670
rect 72216 125734 72564 125740
rect 72216 125670 72358 125734
rect 72422 125670 72494 125734
rect 72558 125670 72564 125734
rect 72216 125664 72564 125670
rect 74664 125734 75148 125740
rect 74664 125670 74942 125734
rect 75006 125670 75078 125734
rect 75142 125670 75148 125734
rect 74664 125664 75148 125670
rect 77248 125734 77596 125740
rect 77248 125670 77390 125734
rect 77454 125670 77526 125734
rect 77590 125670 77596 125734
rect 77248 125664 77596 125670
rect 79696 125734 79908 125740
rect 79696 125670 79702 125734
rect 79766 125670 79838 125734
rect 79902 125670 79908 125734
rect 79696 125664 79908 125670
rect 82280 125734 82628 125740
rect 82280 125670 82422 125734
rect 82486 125670 82558 125734
rect 82622 125670 82628 125734
rect 82280 125664 82628 125670
rect 84728 125734 85076 125740
rect 84728 125670 84870 125734
rect 84934 125670 85006 125734
rect 85070 125670 85076 125734
rect 84728 125664 85076 125670
rect 87176 125734 87388 125740
rect 87176 125670 87182 125734
rect 87246 125670 87318 125734
rect 87382 125670 87388 125734
rect 87176 125664 87388 125670
rect 89760 125734 89972 125740
rect 89760 125670 89766 125734
rect 89830 125670 89902 125734
rect 89966 125670 89972 125734
rect 89760 125664 89972 125670
rect 92208 125734 92556 125740
rect 92208 125670 92350 125734
rect 92414 125670 92486 125734
rect 92550 125670 92556 125734
rect 92208 125664 92556 125670
rect 94656 125734 95004 125740
rect 94656 125670 94798 125734
rect 94862 125670 94934 125734
rect 94998 125670 95004 125734
rect 94656 125664 95004 125670
rect 97240 125734 97588 125740
rect 97240 125670 97382 125734
rect 97446 125670 97518 125734
rect 97582 125670 97588 125734
rect 97240 125664 97588 125670
rect 99688 125734 100036 125740
rect 99688 125670 99830 125734
rect 99894 125670 99966 125734
rect 100030 125670 100036 125734
rect 99688 125664 100036 125670
rect 102136 125734 102484 125740
rect 102136 125670 102142 125734
rect 102206 125670 102414 125734
rect 102478 125670 102484 125734
rect 102136 125664 102484 125670
rect 104720 125734 105068 125740
rect 104720 125670 104862 125734
rect 104926 125670 104998 125734
rect 105062 125670 105068 125734
rect 104720 125664 105068 125670
rect 107168 125734 107516 125740
rect 107168 125670 107310 125734
rect 107374 125670 107446 125734
rect 107510 125670 107516 125734
rect 107168 125664 107516 125670
rect 29865 125615 29963 125664
rect 32361 125615 32459 125664
rect 34857 125615 34955 125664
rect 37353 125615 37451 125664
rect 39849 125615 39947 125664
rect 42345 125615 42443 125664
rect 44841 125615 44939 125664
rect 47337 125615 47435 125664
rect 49833 125615 49931 125664
rect 52329 125615 52427 125664
rect 54825 125615 54923 125664
rect 57321 125615 57419 125664
rect 59817 125615 59915 125664
rect 62313 125615 62411 125664
rect 64809 125615 64907 125664
rect 67305 125615 67403 125664
rect 69801 125615 69899 125664
rect 72297 125615 72395 125664
rect 74793 125615 74891 125664
rect 77289 125615 77387 125664
rect 79785 125615 79883 125664
rect 82281 125615 82379 125664
rect 84777 125615 84875 125664
rect 87273 125615 87371 125664
rect 89769 125615 89867 125664
rect 92265 125615 92363 125664
rect 94761 125615 94859 125664
rect 97257 125615 97355 125664
rect 99753 125615 99851 125664
rect 102249 125615 102347 125664
rect 104745 125615 104843 125664
rect 107241 125615 107339 125664
rect 111000 125445 111066 125448
rect 123611 125445 123677 125448
rect 111000 125443 123677 125445
rect 111000 125387 111005 125443
rect 111061 125387 123616 125443
rect 123672 125387 123677 125443
rect 111000 125385 123677 125387
rect 111000 125382 111066 125385
rect 123611 125382 123677 125385
rect 116280 125054 117580 125060
rect 116280 124990 117374 125054
rect 117438 124990 117580 125054
rect 116280 124984 117580 124990
rect 116280 124918 116492 124984
rect 116280 124854 116286 124918
rect 116350 124854 116492 124918
rect 116280 124848 116492 124854
rect 117368 124848 117580 124984
rect 1768 124728 1980 124788
rect 1768 124672 1798 124728
rect 1854 124672 1980 124728
rect 1768 124652 1980 124672
rect 1224 124646 1980 124652
rect 1224 124582 1230 124646
rect 1294 124582 1980 124646
rect 1224 124576 1980 124582
rect 123624 124782 123972 124788
rect 123624 124718 123902 124782
rect 123966 124718 123972 124782
rect 123624 124712 123972 124718
rect 134640 124712 135668 124788
rect 123624 124646 123836 124712
rect 123624 124582 123630 124646
rect 123694 124582 123836 124646
rect 123624 124576 123836 124582
rect 134640 124576 134852 124712
rect 135456 124652 135668 124712
rect 136816 124782 137572 124788
rect 136816 124728 137502 124782
rect 136816 124672 136944 124728
rect 137000 124718 137502 124728
rect 137566 124718 137572 124782
rect 137000 124712 137572 124718
rect 137000 124672 137028 124712
rect 136816 124652 137028 124672
rect 135456 124576 137028 124652
rect 111124 124031 111190 124034
rect 123611 124031 123677 124034
rect 111124 124029 123677 124031
rect 111124 123973 111129 124029
rect 111185 123973 123616 124029
rect 123672 123973 123677 124029
rect 111124 123971 123677 123973
rect 111124 123968 111190 123971
rect 123611 123968 123677 123971
rect 29920 123830 30268 123836
rect 29920 123766 30062 123830
rect 30126 123766 30268 123830
rect 29920 123564 30268 123766
rect 31280 123700 31492 123836
rect 32504 123830 32716 123836
rect 32504 123766 32646 123830
rect 32710 123766 32716 123830
rect 32504 123700 32716 123766
rect 33728 123700 33940 123836
rect 34952 123830 35164 123836
rect 34952 123766 35094 123830
rect 35158 123766 35164 123830
rect 34952 123700 35164 123766
rect 36176 123700 36388 123836
rect 31280 123624 36388 123700
rect 31280 123564 31492 123624
rect 29920 123558 31492 123564
rect 29920 123494 29926 123558
rect 29990 123494 31492 123558
rect 29920 123488 31492 123494
rect 32504 123488 32716 123624
rect 33728 123488 33940 123624
rect 34952 123488 35164 123624
rect 36176 123564 36388 123624
rect 37400 123830 37748 123836
rect 37400 123766 37406 123830
rect 37470 123766 37748 123830
rect 37400 123564 37748 123766
rect 38760 123564 38972 123836
rect 39984 123830 40196 123836
rect 39984 123766 40126 123830
rect 40190 123766 40196 123830
rect 39984 123700 40196 123766
rect 41208 123700 41420 123836
rect 42432 123830 42644 123836
rect 42432 123766 42574 123830
rect 42638 123766 42644 123830
rect 42432 123700 42644 123766
rect 43656 123700 43868 123836
rect 44880 123830 45228 123836
rect 44880 123766 44886 123830
rect 44950 123766 45228 123830
rect 44880 123700 45228 123766
rect 46240 123700 46452 123836
rect 39984 123624 46452 123700
rect 39984 123564 40196 123624
rect 36176 123488 40196 123564
rect 41208 123488 41420 123624
rect 42432 123488 42644 123624
rect 43656 123488 43868 123624
rect 44880 123488 45228 123624
rect 46240 123564 46452 123624
rect 47464 123830 47676 123836
rect 47464 123766 47470 123830
rect 47534 123766 47676 123830
rect 47464 123564 47676 123766
rect 48688 123700 48900 123836
rect 49912 123830 50124 123836
rect 49912 123766 50054 123830
rect 50118 123766 50124 123830
rect 49912 123700 50124 123766
rect 51136 123700 51484 123836
rect 48688 123624 51484 123700
rect 48688 123564 48900 123624
rect 46240 123488 48900 123564
rect 49912 123488 50124 123624
rect 51136 123564 51484 123624
rect 52496 123830 52708 123836
rect 52496 123766 52502 123830
rect 52566 123766 52708 123830
rect 52496 123564 52708 123766
rect 53720 123700 53932 123836
rect 54944 123830 55156 123836
rect 54944 123766 55086 123830
rect 55150 123766 55156 123830
rect 54944 123700 55156 123766
rect 53720 123624 55156 123700
rect 53720 123564 53932 123624
rect 51136 123488 53932 123564
rect 54944 123564 55156 123624
rect 56168 123564 56380 123836
rect 57392 123830 57604 123836
rect 57392 123766 57534 123830
rect 57598 123766 57604 123830
rect 57392 123700 57604 123766
rect 58616 123830 60188 123836
rect 58616 123766 59982 123830
rect 60046 123766 60188 123830
rect 58616 123760 60188 123766
rect 58616 123700 58964 123760
rect 57392 123624 58964 123700
rect 57392 123564 57604 123624
rect 54944 123488 57604 123564
rect 58616 123488 58964 123624
rect 59976 123564 60188 123760
rect 61200 123564 61412 123836
rect 62424 123830 62636 123836
rect 62424 123766 62566 123830
rect 62630 123766 62636 123830
rect 62424 123700 62636 123766
rect 63648 123700 63860 123836
rect 62424 123624 63860 123700
rect 62424 123564 62636 123624
rect 59976 123488 62636 123564
rect 63648 123564 63860 123624
rect 64872 123830 65084 123836
rect 64872 123766 64878 123830
rect 64942 123766 65084 123830
rect 64872 123564 65084 123766
rect 66096 123564 66444 123836
rect 67456 123830 68892 123836
rect 67456 123766 67462 123830
rect 67526 123766 68892 123830
rect 67456 123760 68892 123766
rect 67456 123564 67668 123760
rect 63648 123488 67668 123564
rect 68680 123564 68892 123760
rect 69904 123830 70116 123836
rect 69904 123766 69910 123830
rect 69974 123766 70116 123830
rect 69904 123564 70116 123766
rect 71128 123700 71340 123836
rect 72352 123830 72700 123836
rect 72352 123766 72494 123830
rect 72558 123766 72700 123830
rect 72352 123700 72700 123766
rect 71128 123624 72700 123700
rect 71128 123564 71340 123624
rect 68680 123488 71340 123564
rect 72352 123564 72700 123624
rect 73712 123700 73924 123836
rect 74936 123830 75148 123836
rect 74936 123766 75078 123830
rect 75142 123766 75148 123830
rect 74936 123700 75148 123766
rect 73712 123624 75148 123700
rect 73712 123564 73924 123624
rect 72352 123488 73924 123564
rect 74936 123564 75148 123624
rect 76160 123830 77596 123836
rect 76160 123766 77526 123830
rect 77590 123766 77596 123830
rect 76160 123760 77596 123766
rect 76160 123564 76372 123760
rect 74936 123488 76372 123564
rect 77384 123564 77596 123760
rect 78608 123564 78820 123836
rect 79832 123830 80180 123836
rect 79832 123766 79838 123830
rect 79902 123766 80180 123830
rect 79832 123564 80180 123766
rect 81192 123564 81404 123836
rect 82416 123830 82628 123836
rect 82416 123766 82558 123830
rect 82622 123766 82628 123830
rect 82416 123700 82628 123766
rect 83640 123700 83852 123836
rect 82416 123624 83852 123700
rect 82416 123564 82628 123624
rect 77384 123488 82628 123564
rect 83640 123564 83852 123624
rect 84864 123830 86300 123836
rect 84864 123766 85006 123830
rect 85070 123766 86300 123830
rect 84864 123760 86300 123766
rect 84864 123564 85076 123760
rect 83640 123488 85076 123564
rect 86088 123564 86300 123760
rect 87312 123830 87660 123836
rect 87312 123766 87318 123830
rect 87382 123766 87660 123830
rect 87312 123564 87660 123766
rect 88672 123564 88884 123836
rect 89896 123830 90108 123836
rect 89896 123766 89902 123830
rect 89966 123766 90108 123830
rect 89896 123564 90108 123766
rect 91120 123700 91332 123836
rect 92344 123830 92556 123836
rect 92344 123766 92486 123830
rect 92550 123766 92556 123830
rect 92344 123700 92556 123766
rect 91120 123624 92556 123700
rect 91120 123564 91332 123624
rect 86088 123488 91332 123564
rect 92344 123564 92556 123624
rect 93568 123830 95140 123836
rect 93568 123766 94934 123830
rect 94998 123766 95140 123830
rect 93568 123760 95140 123766
rect 93568 123564 93916 123760
rect 92344 123488 93916 123564
rect 94928 123700 95140 123760
rect 96152 123700 96364 123836
rect 94928 123624 96364 123700
rect 94928 123488 95140 123624
rect 96152 123564 96364 123624
rect 97376 123830 97588 123836
rect 97376 123766 97518 123830
rect 97582 123766 97588 123830
rect 97376 123564 97588 123766
rect 98600 123564 98812 123836
rect 99824 123830 100036 123836
rect 99824 123766 99966 123830
rect 100030 123766 100036 123830
rect 99824 123700 100036 123766
rect 101048 123700 101396 123836
rect 99824 123624 101396 123700
rect 99824 123564 100036 123624
rect 96152 123488 100036 123564
rect 101048 123564 101396 123624
rect 102408 123830 103844 123836
rect 102408 123766 102414 123830
rect 102478 123766 103844 123830
rect 102408 123760 103844 123766
rect 102408 123564 102620 123760
rect 101048 123488 102620 123564
rect 103632 123700 103844 123760
rect 104856 123830 105068 123836
rect 104856 123766 104998 123830
rect 105062 123766 105068 123830
rect 104856 123700 105068 123766
rect 103632 123624 105068 123700
rect 103632 123488 103844 123624
rect 104856 123564 105068 123624
rect 106080 123564 106292 123836
rect 107304 123830 107516 123836
rect 107304 123766 107446 123830
rect 107510 123766 107516 123830
rect 107304 123564 107516 123766
rect 108528 123564 108876 123836
rect 116280 123694 117580 123700
rect 116280 123630 117374 123694
rect 117438 123630 117580 123694
rect 116280 123624 117580 123630
rect 104856 123558 110236 123564
rect 104856 123494 110166 123558
rect 110230 123494 110236 123558
rect 104856 123488 110236 123494
rect 116280 123352 116492 123624
rect 117368 123422 117580 123624
rect 117368 123358 117374 123422
rect 117438 123358 117580 123422
rect 117368 123352 117580 123358
rect 123624 123422 123836 123428
rect 123624 123358 123766 123422
rect 123830 123358 123836 123422
rect 123624 123216 123836 123358
rect 134640 123292 134852 123428
rect 135456 123422 138252 123428
rect 135456 123358 138182 123422
rect 138246 123358 138252 123422
rect 135456 123352 138252 123358
rect 135456 123292 135668 123352
rect 134640 123286 135668 123292
rect 134640 123222 134646 123286
rect 134710 123222 135668 123286
rect 134640 123216 135668 123222
rect 1224 123150 1980 123156
rect 1224 123086 1230 123150
rect 1294 123086 1980 123150
rect 1224 123080 1980 123086
rect 1768 123048 1980 123080
rect 1768 122992 1798 123048
rect 1854 122992 1980 123048
rect 1768 122944 1980 122992
rect 136816 123048 137028 123156
rect 136816 122992 136944 123048
rect 137000 123020 137028 123048
rect 137000 123014 137572 123020
rect 137000 122992 137502 123014
rect 136816 122950 137502 122992
rect 137566 122950 137572 123014
rect 136816 122944 137572 122950
rect 136187 122916 136193 122918
rect 116416 122856 116476 122916
rect 123476 122856 136193 122916
rect 136187 122854 136193 122856
rect 136257 122854 136263 122918
rect 114985 122617 115051 122620
rect 123611 122617 123677 122620
rect 114985 122615 123677 122617
rect 114985 122559 114990 122615
rect 115046 122559 123616 122615
rect 123672 122559 123677 122615
rect 114985 122557 123677 122559
rect 114985 122554 115051 122557
rect 123611 122554 123677 122557
rect 29512 122068 29724 122204
rect 30464 122128 31084 122204
rect 29512 122062 30404 122068
rect 29512 121998 29654 122062
rect 29718 121998 30334 122062
rect 30398 121998 30404 122062
rect 29512 121992 30404 121998
rect 30464 122062 30676 122128
rect 30464 121998 30470 122062
rect 30534 121998 30676 122062
rect 30464 121992 30676 121998
rect 30736 121992 31084 122128
rect 31688 122068 31900 122204
rect 32096 122068 32308 122204
rect 32912 122128 33532 122204
rect 31688 122062 32852 122068
rect 31688 121998 31694 122062
rect 31758 121998 32782 122062
rect 32846 121998 32852 122062
rect 31688 121992 32852 121998
rect 32912 121992 33124 122128
rect 33320 122062 33532 122128
rect 33320 121998 33462 122062
rect 33526 121998 33532 122062
rect 33320 121992 33532 121998
rect 34136 122068 34348 122204
rect 34544 122068 34756 122204
rect 34136 122062 34756 122068
rect 34136 121998 34142 122062
rect 34206 121998 34686 122062
rect 34750 121998 34756 122062
rect 34136 121992 34756 121998
rect 35360 122128 35980 122204
rect 35360 122062 35572 122128
rect 35360 121998 35366 122062
rect 35430 121998 35572 122062
rect 35360 121992 35572 121998
rect 35768 122062 35980 122128
rect 35768 121998 35910 122062
rect 35974 121998 35980 122062
rect 35768 121992 35980 121998
rect 36584 122128 37204 122204
rect 36584 121992 36932 122128
rect 36992 122062 37204 122128
rect 36992 121998 37134 122062
rect 37198 121998 37204 122062
rect 36992 121992 37204 121998
rect 37944 122068 38156 122204
rect 38216 122068 38564 122204
rect 37944 122062 38564 122068
rect 37944 121998 38494 122062
rect 38558 121998 38564 122062
rect 37944 121992 38564 121998
rect 39168 122128 39788 122204
rect 39168 122062 39380 122128
rect 39168 121998 39174 122062
rect 39238 121998 39380 122062
rect 39168 121992 39380 121998
rect 39576 122062 39788 122128
rect 39576 121998 39582 122062
rect 39646 121998 39788 122062
rect 39576 121992 39788 121998
rect 40392 122068 40604 122204
rect 40800 122068 41012 122204
rect 40392 122062 41012 122068
rect 40392 121998 40398 122062
rect 40462 121998 40942 122062
rect 41006 121998 41012 122062
rect 40392 121992 41012 121998
rect 41616 122128 42236 122204
rect 41616 121992 41828 122128
rect 42024 122062 42236 122128
rect 42024 121998 42166 122062
rect 42230 121998 42236 122062
rect 42024 121992 42236 121998
rect 42840 122068 43052 122204
rect 43248 122068 43460 122204
rect 44064 122128 44684 122204
rect 44064 122068 44412 122128
rect 42840 122062 43460 122068
rect 43966 122062 44412 122068
rect 42840 121998 42846 122062
rect 42910 121998 43390 122062
rect 43454 121998 43460 122062
rect 43928 121998 43934 122062
rect 43998 121998 44070 122062
rect 44134 121998 44412 122062
rect 42840 121992 43460 121998
rect 43966 121992 44412 121998
rect 44472 122062 44684 122128
rect 44472 121998 44614 122062
rect 44678 121998 44684 122062
rect 44472 121992 44684 121998
rect 45424 122128 46044 122204
rect 45424 121992 45636 122128
rect 45696 122062 46044 122128
rect 45696 121998 45702 122062
rect 45766 121998 46044 122062
rect 45696 121992 46044 121998
rect 46648 122068 46860 122204
rect 47056 122068 47268 122204
rect 46648 122062 47268 122068
rect 46648 121998 46654 122062
rect 46718 121998 47268 122062
rect 46648 121992 47268 121998
rect 47872 122128 48492 122204
rect 47872 122062 48084 122128
rect 47872 121998 47878 122062
rect 47942 121998 48084 122062
rect 47872 121992 48084 121998
rect 48280 122062 48492 122128
rect 48280 121998 48422 122062
rect 48486 121998 48492 122062
rect 48280 121992 48492 121998
rect 49096 122068 49308 122204
rect 49504 122068 49716 122204
rect 49096 122062 49716 122068
rect 49096 121998 49102 122062
rect 49166 121998 49238 122062
rect 49302 121998 49716 122062
rect 49096 121992 49716 121998
rect 50320 122128 50940 122204
rect 50320 122062 50668 122128
rect 50320 121998 50326 122062
rect 50390 121998 50668 122062
rect 50320 121992 50668 121998
rect 50728 122062 50940 122128
rect 50728 121998 50870 122062
rect 50934 121998 50940 122062
rect 50728 121992 50940 121998
rect 51680 122128 52300 122204
rect 51680 121992 51892 122128
rect 51952 122062 52300 122128
rect 51952 121998 52230 122062
rect 52294 121998 52300 122062
rect 51952 121992 52300 121998
rect 52904 122068 53116 122204
rect 53312 122068 53524 122204
rect 52904 122062 53524 122068
rect 52904 121998 52910 122062
rect 52974 121998 53318 122062
rect 53382 121998 53524 122062
rect 52904 121992 53524 121998
rect 54128 122128 54748 122204
rect 54128 122062 54340 122128
rect 54128 121998 54134 122062
rect 54198 121998 54340 122062
rect 54128 121992 54340 121998
rect 54536 122062 54748 122128
rect 54536 121998 54678 122062
rect 54742 121998 54748 122062
rect 54536 121992 54748 121998
rect 55352 122068 55564 122204
rect 55760 122068 55972 122204
rect 55352 122062 55972 122068
rect 55352 121998 55358 122062
rect 55422 121998 55972 122062
rect 55352 121992 55972 121998
rect 56576 122128 57196 122204
rect 56576 122062 56788 122128
rect 56576 121998 56718 122062
rect 56782 121998 56788 122062
rect 56576 121992 56788 121998
rect 56984 122062 57196 122128
rect 56984 121998 57126 122062
rect 57190 121998 57196 122062
rect 56984 121992 57196 121998
rect 57800 122068 58148 122204
rect 58208 122068 58420 122204
rect 57800 122062 58420 122068
rect 57800 121998 58078 122062
rect 58142 121998 58420 122062
rect 57800 121992 58420 121998
rect 59160 122068 59372 122204
rect 59432 122068 59780 122204
rect 59160 122062 59780 122068
rect 59160 121998 59166 122062
rect 59230 121998 59780 122062
rect 59160 121992 59780 121998
rect 60384 122128 61004 122204
rect 60384 121992 60596 122128
rect 60792 122062 61004 122128
rect 60792 121998 60934 122062
rect 60998 121998 61004 122062
rect 60792 121992 61004 121998
rect 61608 122068 61820 122204
rect 62016 122068 62228 122204
rect 61608 122062 62228 122068
rect 61608 121998 61614 122062
rect 61678 121998 62158 122062
rect 62222 121998 62228 122062
rect 61608 121992 62228 121998
rect 62832 122128 63452 122204
rect 62832 122062 63044 122128
rect 62832 121998 62838 122062
rect 62902 121998 63044 122062
rect 62832 121992 63044 121998
rect 63240 122062 63452 122128
rect 63240 121998 63382 122062
rect 63446 121998 63452 122062
rect 63240 121992 63452 121998
rect 64056 122068 64268 122204
rect 64464 122068 64676 122204
rect 64056 122062 64676 122068
rect 64056 121998 64062 122062
rect 64126 121998 64606 122062
rect 64670 121998 64676 122062
rect 64056 121992 64676 121998
rect 65280 122128 65900 122204
rect 65280 121992 65628 122128
rect 65688 122062 65900 122128
rect 65688 121998 65694 122062
rect 65758 121998 65900 122062
rect 65688 121992 65900 121998
rect 66640 122128 67260 122204
rect 66640 121992 66852 122128
rect 66912 122062 67260 122128
rect 66912 121998 67190 122062
rect 67254 121998 67260 122062
rect 66912 121992 67260 121998
rect 67864 122068 68076 122204
rect 68272 122068 68484 122204
rect 67864 122062 68484 122068
rect 67864 121998 67870 122062
rect 67934 121998 68414 122062
rect 68478 121998 68484 122062
rect 67864 121992 68484 121998
rect 69088 122128 69708 122204
rect 69088 122062 69300 122128
rect 69088 121998 69094 122062
rect 69158 121998 69300 122062
rect 69088 121992 69300 121998
rect 69496 122062 69708 122128
rect 69496 121998 69638 122062
rect 69702 121998 69708 122062
rect 69496 121992 69708 121998
rect 70312 122068 70524 122204
rect 70720 122068 70932 122204
rect 70312 122062 70932 122068
rect 70312 121998 70318 122062
rect 70382 121998 70862 122062
rect 70926 121998 70932 122062
rect 70312 121992 70932 121998
rect 71536 122128 72156 122204
rect 71536 121992 71884 122128
rect 71944 122068 72156 122128
rect 72896 122128 73516 122204
rect 71944 122062 72836 122068
rect 71944 121998 72086 122062
rect 72150 121998 72766 122062
rect 72830 121998 72836 122062
rect 71944 121992 72836 121998
rect 72896 122062 73108 122128
rect 72896 121998 72902 122062
rect 72966 121998 73108 122062
rect 72896 121992 73108 121998
rect 73168 122062 73516 122128
rect 73168 121998 73310 122062
rect 73374 121998 73516 122062
rect 73168 121992 73516 121998
rect 74120 122068 74332 122204
rect 74528 122068 74740 122204
rect 75344 122128 75964 122204
rect 74120 122062 75284 122068
rect 74120 121998 74126 122062
rect 74190 121998 75214 122062
rect 75278 121998 75284 122062
rect 74120 121992 75284 121998
rect 75344 122062 75556 122128
rect 75344 121998 75350 122062
rect 75414 121998 75556 122062
rect 75344 121992 75556 121998
rect 75752 122062 75964 122128
rect 75752 121998 75894 122062
rect 75958 121998 75964 122062
rect 75752 121992 75964 121998
rect 76568 122068 76780 122204
rect 76976 122068 77188 122204
rect 76568 122062 77188 122068
rect 76568 121998 76574 122062
rect 76638 121998 77118 122062
rect 77182 121998 77188 122062
rect 76568 121992 77188 121998
rect 77792 122128 78412 122204
rect 77792 122062 78004 122128
rect 77792 121998 77798 122062
rect 77862 121998 78004 122062
rect 77792 121992 78004 121998
rect 78200 122062 78412 122128
rect 78200 121998 78342 122062
rect 78406 121998 78412 122062
rect 78200 121992 78412 121998
rect 79016 122068 79364 122204
rect 79424 122068 79636 122204
rect 79016 122062 79636 122068
rect 79016 121998 79566 122062
rect 79630 121998 79636 122062
rect 79016 121992 79636 121998
rect 80376 122068 80588 122204
rect 80648 122068 80996 122204
rect 81600 122128 82220 122204
rect 80376 122062 81540 122068
rect 80376 121998 80518 122062
rect 80582 121998 81470 122062
rect 81534 121998 81540 122062
rect 80376 121992 81540 121998
rect 81600 122062 81812 122128
rect 81600 121998 81606 122062
rect 81670 121998 81812 122062
rect 81600 121992 81812 121998
rect 82008 121992 82220 122128
rect 82824 122068 83036 122204
rect 83232 122068 83444 122204
rect 82824 122062 83444 122068
rect 82824 121998 82830 122062
rect 82894 121998 83374 122062
rect 83438 121998 83444 122062
rect 82824 121992 83444 121998
rect 84048 122128 84668 122204
rect 84048 122062 84260 122128
rect 84048 121998 84054 122062
rect 84118 121998 84260 122062
rect 84048 121992 84260 121998
rect 84456 122062 84668 122128
rect 84456 121998 84598 122062
rect 84662 121998 84668 122062
rect 84456 121992 84668 121998
rect 85272 122068 85484 122204
rect 85680 122068 85892 122204
rect 85272 122062 85892 122068
rect 85272 121998 85414 122062
rect 85478 121998 85822 122062
rect 85886 121998 85892 122062
rect 85272 121992 85892 121998
rect 86496 122128 87116 122204
rect 86496 122062 86844 122128
rect 86496 121998 86502 122062
rect 86566 121998 86844 122062
rect 86496 121992 86844 121998
rect 86904 122062 87116 122128
rect 86904 121998 87046 122062
rect 87110 121998 87116 122062
rect 86904 121992 87116 121998
rect 87856 122198 88476 122204
rect 87856 122134 87862 122198
rect 87926 122134 88476 122198
rect 87856 122128 88476 122134
rect 87856 121992 88068 122128
rect 88128 122062 88476 122128
rect 88128 121998 88406 122062
rect 88470 121998 88476 122062
rect 88128 121992 88476 121998
rect 89080 122068 89292 122204
rect 89488 122068 89700 122204
rect 89080 122062 89700 122068
rect 89080 121998 89086 122062
rect 89150 121998 89222 122062
rect 89286 121998 89700 122062
rect 89080 121992 89700 121998
rect 90304 122128 90924 122204
rect 90304 122062 90516 122128
rect 90304 121998 90310 122062
rect 90374 121998 90516 122062
rect 90304 121992 90516 121998
rect 90712 122062 90924 122128
rect 90712 121998 90854 122062
rect 90918 121998 90924 122062
rect 90712 121992 90924 121998
rect 91528 122068 91740 122204
rect 91936 122068 92148 122204
rect 91528 122062 92148 122068
rect 91528 121998 91534 122062
rect 91598 121998 92148 122062
rect 91528 121992 92148 121998
rect 92752 122128 93372 122204
rect 92752 122062 93100 122128
rect 92752 121998 92758 122062
rect 92822 121998 93100 122062
rect 92752 121992 93100 121998
rect 93160 122062 93372 122128
rect 93160 121998 93302 122062
rect 93366 121998 93372 122062
rect 93160 121992 93372 121998
rect 94112 122128 94732 122204
rect 94112 122062 94324 122128
rect 94112 121998 94254 122062
rect 94318 121998 94324 122062
rect 94112 121992 94324 121998
rect 94384 121992 94732 122128
rect 95336 122068 95548 122204
rect 95744 122068 95956 122204
rect 95336 122062 95956 122068
rect 95336 121998 95478 122062
rect 95542 121998 95956 122062
rect 95336 121992 95956 121998
rect 96560 122128 97180 122204
rect 96560 121992 96772 122128
rect 96968 122062 97180 122128
rect 96968 121998 97110 122062
rect 97174 121998 97180 122062
rect 96968 121992 97180 121998
rect 97784 122068 97996 122204
rect 98192 122068 98404 122204
rect 97784 122062 98404 122068
rect 97784 121998 97790 122062
rect 97854 121998 98334 122062
rect 98398 121998 98404 122062
rect 97784 121992 98404 121998
rect 99008 122128 99628 122204
rect 99008 122062 99220 122128
rect 99008 121998 99014 122062
rect 99078 121998 99220 122062
rect 99008 121992 99220 121998
rect 99416 122062 99628 122128
rect 99416 121998 99558 122062
rect 99622 121998 99628 122062
rect 99416 121992 99628 121998
rect 100232 122068 100580 122204
rect 100640 122068 100852 122204
rect 100232 122062 100852 122068
rect 100232 121998 100782 122062
rect 100846 121998 100852 122062
rect 100232 121992 100852 121998
rect 101592 122068 101804 122204
rect 101864 122068 102212 122204
rect 101592 122062 102212 122068
rect 101592 121998 101598 122062
rect 101662 121998 102006 122062
rect 102070 121998 102212 122062
rect 101592 121992 102212 121998
rect 102816 122128 103436 122204
rect 102816 121992 103028 122128
rect 103224 122068 103436 122128
rect 104040 122068 104252 122204
rect 104448 122068 104660 122204
rect 103224 122062 103980 122068
rect 103224 121998 103366 122062
rect 103430 121998 103910 122062
rect 103974 121998 103980 122062
rect 103224 121992 103980 121998
rect 104040 122062 104660 122068
rect 104040 121998 104046 122062
rect 104110 121998 104590 122062
rect 104654 121998 104660 122062
rect 104040 121992 104660 121998
rect 105264 122128 105884 122204
rect 105264 121992 105476 122128
rect 105672 122062 105884 122128
rect 105672 121998 105814 122062
rect 105878 121998 105884 122062
rect 105672 121992 105884 121998
rect 106488 122068 106700 122204
rect 106896 122068 107108 122204
rect 106488 122062 107108 122068
rect 106488 121998 107038 122062
rect 107102 121998 107108 122062
rect 106488 121992 107108 121998
rect 107712 122068 108060 122204
rect 108120 122068 108332 122204
rect 107712 122062 108332 122068
rect 107712 121998 108126 122062
rect 108190 121998 108332 122062
rect 107712 121992 108332 121998
rect 109072 122128 109692 122204
rect 109072 121992 109284 122128
rect 109344 122062 109692 122128
rect 109344 121998 109486 122062
rect 109550 121998 109692 122062
rect 109344 121992 109692 121998
rect 123624 121926 123836 121932
rect 123624 121862 123630 121926
rect 123694 121862 123836 121926
rect 123624 121720 123836 121862
rect 134640 121856 135668 121932
rect 134640 121720 134852 121856
rect 135456 121796 135668 121856
rect 135456 121790 136892 121796
rect 135456 121726 136822 121790
rect 136886 121726 136892 121790
rect 135456 121720 136892 121726
rect 28968 121524 29316 121660
rect 29648 121654 29860 121660
rect 29648 121590 29654 121654
rect 29718 121590 29860 121654
rect 29648 121524 29860 121590
rect 1224 121518 1980 121524
rect 1224 121454 1230 121518
rect 1294 121454 1980 121518
rect 1224 121448 1980 121454
rect 28968 121448 29860 121524
rect 30328 121654 30540 121660
rect 30328 121590 30334 121654
rect 30398 121590 30470 121654
rect 30534 121590 30540 121654
rect 30328 121524 30540 121590
rect 30872 121524 31084 121660
rect 31552 121654 32444 121660
rect 31552 121590 31694 121654
rect 31758 121590 32444 121654
rect 31552 121584 32444 121590
rect 31552 121524 31764 121584
rect 30328 121448 31764 121524
rect 32096 121448 32444 121584
rect 32776 121654 32988 121660
rect 32776 121590 32782 121654
rect 32846 121590 32988 121654
rect 32776 121524 32988 121590
rect 33456 121654 34212 121660
rect 33456 121590 33462 121654
rect 33526 121590 34142 121654
rect 34206 121590 34212 121654
rect 33456 121584 34212 121590
rect 33456 121524 33668 121584
rect 32776 121448 33668 121524
rect 34000 121448 34212 121584
rect 34680 121654 34892 121660
rect 34680 121590 34686 121654
rect 34750 121590 34892 121654
rect 34680 121524 34892 121590
rect 35224 121654 35572 121660
rect 35224 121590 35366 121654
rect 35430 121590 35572 121654
rect 35224 121524 35572 121590
rect 34680 121448 35572 121524
rect 35904 121654 36796 121660
rect 35904 121590 35910 121654
rect 35974 121590 36796 121654
rect 35904 121584 36796 121590
rect 35904 121448 36116 121584
rect 36584 121524 36796 121584
rect 37128 121654 37340 121660
rect 37128 121590 37134 121654
rect 37198 121590 37340 121654
rect 37128 121524 37340 121590
rect 37808 121654 39244 121660
rect 37808 121590 38494 121654
rect 38558 121590 39174 121654
rect 39238 121590 39244 121654
rect 37808 121584 39244 121590
rect 37808 121524 38020 121584
rect 36584 121448 38020 121524
rect 38352 121448 38564 121584
rect 39032 121448 39244 121584
rect 39576 121654 40468 121660
rect 39576 121590 39582 121654
rect 39646 121590 40398 121654
rect 40462 121590 40468 121654
rect 39576 121584 40468 121590
rect 39576 121448 39924 121584
rect 40256 121448 40468 121584
rect 40936 121654 41148 121660
rect 40936 121590 40942 121654
rect 41006 121590 41148 121654
rect 40936 121524 41148 121590
rect 41480 121524 41692 121660
rect 42160 121654 43052 121660
rect 42160 121590 42166 121654
rect 42230 121590 42846 121654
rect 42910 121590 43052 121654
rect 42160 121584 43052 121590
rect 42160 121524 42372 121584
rect 40936 121448 42372 121524
rect 42704 121448 43052 121584
rect 43384 121654 44004 121660
rect 43384 121590 43390 121654
rect 43454 121590 43934 121654
rect 43998 121590 44004 121654
rect 43384 121584 44004 121590
rect 44064 121654 44276 121660
rect 44064 121590 44070 121654
rect 44134 121590 44276 121654
rect 43384 121448 43596 121584
rect 44064 121448 44276 121590
rect 44608 121654 45772 121660
rect 44608 121590 44614 121654
rect 44678 121590 45702 121654
rect 45766 121590 45772 121654
rect 44608 121584 45772 121590
rect 44608 121448 44820 121584
rect 45288 121524 45500 121584
rect 45832 121524 46180 121660
rect 46512 121654 47404 121660
rect 46512 121590 46654 121654
rect 46718 121590 47404 121654
rect 46512 121584 47404 121590
rect 46512 121524 46724 121584
rect 45288 121448 46724 121524
rect 47192 121524 47404 121584
rect 47736 121654 47948 121660
rect 47736 121590 47878 121654
rect 47942 121590 47948 121654
rect 47736 121524 47948 121590
rect 47192 121448 47948 121524
rect 48416 121654 49172 121660
rect 49270 121654 49852 121660
rect 48416 121590 48422 121654
rect 48486 121590 49102 121654
rect 49166 121590 49172 121654
rect 49232 121590 49238 121654
rect 49302 121590 49852 121654
rect 48416 121584 49172 121590
rect 49270 121584 49852 121590
rect 48416 121448 48628 121584
rect 48960 121448 49172 121584
rect 49640 121524 49852 121584
rect 50184 121654 50532 121660
rect 50184 121590 50326 121654
rect 50390 121590 50532 121654
rect 50184 121524 50532 121590
rect 49640 121448 50532 121524
rect 50864 121654 51756 121660
rect 50864 121590 50870 121654
rect 50934 121590 51756 121654
rect 50864 121584 51756 121590
rect 50864 121448 51076 121584
rect 51544 121524 51756 121584
rect 52088 121654 52300 121660
rect 52088 121590 52230 121654
rect 52294 121590 52300 121654
rect 52088 121524 52300 121590
rect 52768 121654 52980 121660
rect 52768 121590 52910 121654
rect 52974 121590 52980 121654
rect 52768 121524 52980 121590
rect 51544 121448 52980 121524
rect 53312 121654 54204 121660
rect 53312 121590 53318 121654
rect 53382 121590 54134 121654
rect 54198 121590 54204 121654
rect 53312 121584 54204 121590
rect 53312 121448 53660 121584
rect 53992 121448 54204 121584
rect 54672 121654 56108 121660
rect 54672 121590 54678 121654
rect 54742 121590 55358 121654
rect 55422 121590 56108 121654
rect 54672 121584 56108 121590
rect 54672 121448 54884 121584
rect 55216 121448 55428 121584
rect 55896 121524 56108 121584
rect 56440 121654 56788 121660
rect 56440 121590 56718 121654
rect 56782 121590 56788 121654
rect 56440 121524 56788 121590
rect 55896 121448 56788 121524
rect 57120 121654 58012 121660
rect 58110 121654 58556 121660
rect 57120 121590 57126 121654
rect 57190 121590 58012 121654
rect 58072 121590 58078 121654
rect 58142 121590 58556 121654
rect 57120 121584 58012 121590
rect 58110 121584 58556 121590
rect 57120 121448 57332 121584
rect 57800 121524 58012 121584
rect 58344 121524 58556 121584
rect 59024 121654 60460 121660
rect 59024 121590 59166 121654
rect 59230 121590 60460 121654
rect 59024 121584 60460 121590
rect 59024 121524 59236 121584
rect 57800 121448 59236 121524
rect 59568 121448 59780 121584
rect 60248 121524 60460 121584
rect 60792 121654 61684 121660
rect 60792 121590 60934 121654
rect 60998 121590 61614 121654
rect 61678 121590 61684 121654
rect 60792 121584 61684 121590
rect 60792 121524 61140 121584
rect 60248 121448 61140 121524
rect 61472 121448 61684 121584
rect 62152 121654 62364 121660
rect 62152 121590 62158 121654
rect 62222 121590 62364 121654
rect 62152 121524 62364 121590
rect 62696 121654 62908 121660
rect 62696 121590 62838 121654
rect 62902 121590 62908 121654
rect 62696 121524 62908 121590
rect 62152 121448 62908 121524
rect 63376 121654 64268 121660
rect 63376 121590 63382 121654
rect 63446 121590 64062 121654
rect 64126 121590 64268 121654
rect 63376 121584 64268 121590
rect 63376 121448 63588 121584
rect 63920 121448 64268 121584
rect 64600 121654 64812 121660
rect 64600 121590 64606 121654
rect 64670 121590 64812 121654
rect 64600 121524 64812 121590
rect 65280 121654 65764 121660
rect 65280 121590 65694 121654
rect 65758 121590 65764 121654
rect 65280 121584 65764 121590
rect 65824 121584 66716 121660
rect 65280 121524 65492 121584
rect 65824 121524 66036 121584
rect 64600 121448 66036 121524
rect 66504 121524 66716 121584
rect 67048 121654 67396 121660
rect 67048 121590 67190 121654
rect 67254 121590 67396 121654
rect 67048 121524 67396 121590
rect 67728 121654 67940 121660
rect 67728 121590 67870 121654
rect 67934 121590 67940 121654
rect 67728 121524 67940 121590
rect 66504 121448 67940 121524
rect 68408 121654 68620 121660
rect 68408 121590 68414 121654
rect 68478 121590 68620 121654
rect 68408 121524 68620 121590
rect 68952 121654 69164 121660
rect 68952 121590 69094 121654
rect 69158 121590 69164 121654
rect 68952 121524 69164 121590
rect 68408 121448 69164 121524
rect 69632 121654 70388 121660
rect 69632 121590 69638 121654
rect 69702 121590 70318 121654
rect 70382 121590 70388 121654
rect 69632 121584 70388 121590
rect 69632 121448 69844 121584
rect 70176 121448 70388 121584
rect 70856 121654 71068 121660
rect 70856 121590 70862 121654
rect 70926 121590 71068 121654
rect 70856 121524 71068 121590
rect 71400 121524 71748 121660
rect 72080 121654 72292 121660
rect 72080 121590 72086 121654
rect 72150 121590 72292 121654
rect 72080 121524 72292 121590
rect 70856 121448 72292 121524
rect 72760 121654 72972 121660
rect 72760 121590 72766 121654
rect 72830 121590 72902 121654
rect 72966 121590 72972 121654
rect 72760 121448 72972 121590
rect 73304 121654 73516 121660
rect 73304 121590 73310 121654
rect 73374 121590 73516 121654
rect 73304 121524 73516 121590
rect 73984 121654 74876 121660
rect 73984 121590 74126 121654
rect 74190 121590 74876 121654
rect 73984 121584 74876 121590
rect 73984 121524 74196 121584
rect 73304 121448 74196 121524
rect 74528 121448 74876 121584
rect 75208 121654 75420 121660
rect 75208 121590 75214 121654
rect 75278 121590 75350 121654
rect 75414 121590 75420 121654
rect 75208 121448 75420 121590
rect 75888 121654 76644 121660
rect 75888 121590 75894 121654
rect 75958 121590 76574 121654
rect 76638 121590 76644 121654
rect 75888 121584 76644 121590
rect 75888 121448 76100 121584
rect 76432 121448 76644 121584
rect 77112 121654 77324 121660
rect 77112 121590 77118 121654
rect 77182 121590 77324 121654
rect 77112 121524 77324 121590
rect 77656 121654 78004 121660
rect 77656 121590 77798 121654
rect 77862 121590 78004 121654
rect 77656 121524 78004 121590
rect 77112 121448 78004 121524
rect 78336 121654 79228 121660
rect 78336 121590 78342 121654
rect 78406 121590 79228 121654
rect 78336 121584 79228 121590
rect 78336 121448 78548 121584
rect 79016 121524 79228 121584
rect 79560 121654 79772 121660
rect 79560 121590 79566 121654
rect 79630 121590 79772 121654
rect 79560 121524 79772 121590
rect 80240 121584 80996 121660
rect 80240 121524 80452 121584
rect 80784 121524 80996 121584
rect 79016 121448 80452 121524
rect 80550 121518 80996 121524
rect 80512 121454 80518 121518
rect 80582 121454 80996 121518
rect 80550 121448 80996 121454
rect 81464 121654 81676 121660
rect 81464 121590 81470 121654
rect 81534 121590 81606 121654
rect 81670 121590 81676 121654
rect 81464 121524 81676 121590
rect 82008 121524 82356 121660
rect 82688 121654 82900 121660
rect 82688 121590 82830 121654
rect 82894 121590 82900 121654
rect 82688 121524 82900 121590
rect 81464 121448 82900 121524
rect 83368 121654 83580 121660
rect 83368 121590 83374 121654
rect 83438 121590 83580 121654
rect 83368 121524 83580 121590
rect 83912 121654 84124 121660
rect 83912 121590 84054 121654
rect 84118 121590 84124 121654
rect 83912 121524 84124 121590
rect 83368 121448 84124 121524
rect 84592 121654 85484 121660
rect 84592 121590 84598 121654
rect 84662 121590 85414 121654
rect 85478 121590 85484 121654
rect 84592 121584 85484 121590
rect 84592 121448 84804 121584
rect 85136 121448 85484 121584
rect 85816 121654 86028 121660
rect 85816 121590 85822 121654
rect 85886 121590 86028 121654
rect 85816 121524 86028 121590
rect 86496 121654 86708 121660
rect 86496 121590 86502 121654
rect 86566 121590 86708 121654
rect 86496 121524 86708 121590
rect 85816 121448 86708 121524
rect 87040 121654 87932 121660
rect 87040 121590 87046 121654
rect 87110 121590 87932 121654
rect 87040 121584 87932 121590
rect 87040 121448 87252 121584
rect 87720 121524 87932 121584
rect 88264 121654 88612 121660
rect 88264 121590 88406 121654
rect 88470 121590 88612 121654
rect 88264 121524 88612 121590
rect 88944 121654 89156 121660
rect 89254 121654 89836 121660
rect 88944 121590 89086 121654
rect 89150 121590 89156 121654
rect 89216 121590 89222 121654
rect 89286 121590 89836 121654
rect 88944 121524 89156 121590
rect 89254 121584 89836 121590
rect 87720 121448 89156 121524
rect 89624 121524 89836 121584
rect 90168 121654 90380 121660
rect 90168 121590 90310 121654
rect 90374 121590 90380 121654
rect 90168 121524 90380 121590
rect 89624 121448 90380 121524
rect 90848 121654 92284 121660
rect 90848 121590 90854 121654
rect 90918 121590 91534 121654
rect 91598 121590 92284 121654
rect 90848 121584 92284 121590
rect 90848 121448 91060 121584
rect 91392 121448 91604 121584
rect 92072 121524 92284 121584
rect 92616 121654 92964 121660
rect 92616 121590 92758 121654
rect 92822 121590 92964 121654
rect 92616 121524 92964 121590
rect 92072 121448 92964 121524
rect 93296 121654 94188 121660
rect 94286 121654 94732 121660
rect 93296 121590 93302 121654
rect 93366 121590 94188 121654
rect 94248 121590 94254 121654
rect 94318 121590 94732 121654
rect 93296 121584 94188 121590
rect 94286 121584 94732 121590
rect 93296 121448 93508 121584
rect 93976 121524 94188 121584
rect 94520 121524 94732 121584
rect 95200 121584 96636 121660
rect 95200 121524 95412 121584
rect 95744 121524 96092 121584
rect 93976 121448 95412 121524
rect 95510 121518 96092 121524
rect 95472 121454 95478 121518
rect 95542 121454 96092 121518
rect 95510 121448 96092 121454
rect 96424 121524 96636 121584
rect 97104 121654 97860 121660
rect 97104 121590 97110 121654
rect 97174 121590 97790 121654
rect 97854 121590 97860 121654
rect 97104 121584 97860 121590
rect 97104 121524 97316 121584
rect 96424 121448 97316 121524
rect 97648 121448 97860 121584
rect 98328 121654 98540 121660
rect 98328 121590 98334 121654
rect 98398 121590 98540 121654
rect 98328 121524 98540 121590
rect 98872 121654 99220 121660
rect 98872 121590 99014 121654
rect 99078 121590 99220 121654
rect 98872 121524 99220 121590
rect 98328 121448 99220 121524
rect 99552 121654 100444 121660
rect 99552 121590 99558 121654
rect 99622 121590 100444 121654
rect 99552 121584 100444 121590
rect 99552 121448 99764 121584
rect 100232 121524 100444 121584
rect 100776 121654 100988 121660
rect 100776 121590 100782 121654
rect 100846 121590 100988 121654
rect 100776 121524 100988 121590
rect 101456 121654 101668 121660
rect 101456 121590 101598 121654
rect 101662 121590 101668 121654
rect 101456 121524 101668 121590
rect 100232 121448 101668 121524
rect 102000 121654 102892 121660
rect 102000 121590 102006 121654
rect 102070 121590 102892 121654
rect 102000 121584 102892 121590
rect 102000 121448 102212 121584
rect 102680 121524 102892 121584
rect 103224 121654 103572 121660
rect 103224 121590 103366 121654
rect 103430 121590 103572 121654
rect 103224 121524 103572 121590
rect 102680 121448 103572 121524
rect 103904 121654 104116 121660
rect 103904 121590 103910 121654
rect 103974 121590 104046 121654
rect 104110 121590 104116 121654
rect 103904 121448 104116 121590
rect 104584 121654 104796 121660
rect 104584 121590 104590 121654
rect 104654 121590 104796 121654
rect 104584 121524 104796 121590
rect 105128 121524 105340 121660
rect 105808 121654 107244 121660
rect 105808 121590 105814 121654
rect 105878 121590 107038 121654
rect 107102 121590 107244 121654
rect 105808 121584 107244 121590
rect 105808 121524 106020 121584
rect 104584 121448 106020 121524
rect 106352 121448 106700 121584
rect 107032 121524 107244 121584
rect 107712 121654 108196 121660
rect 107712 121590 108126 121654
rect 108190 121590 108196 121654
rect 107712 121584 108196 121590
rect 108256 121584 109148 121660
rect 107712 121524 107924 121584
rect 108256 121524 108468 121584
rect 107032 121448 108468 121524
rect 108936 121524 109148 121584
rect 109480 121654 109828 121660
rect 109480 121590 109486 121654
rect 109550 121590 109828 121654
rect 109480 121524 109828 121590
rect 108936 121518 111732 121524
rect 108936 121454 111662 121518
rect 111726 121454 111732 121518
rect 108936 121448 111732 121454
rect 136816 121518 137572 121524
rect 136816 121454 136822 121518
rect 136886 121454 137502 121518
rect 137566 121454 137572 121518
rect 136816 121448 137572 121454
rect 1768 121368 1980 121448
rect 1768 121312 1798 121368
rect 1854 121312 1980 121368
rect 1768 121176 1980 121312
rect 28016 121252 28228 121388
rect 28016 121176 28364 121252
rect 28288 121116 28364 121176
rect 110568 121176 110780 121388
rect 136816 121368 137028 121448
rect 136816 121312 136944 121368
rect 137000 121312 137028 121368
rect 111656 121246 111868 121252
rect 111656 121182 111662 121246
rect 111726 121182 111868 121246
rect 110568 121116 110644 121176
rect 28288 121110 29996 121116
rect 28288 121046 29926 121110
rect 29990 121046 29996 121110
rect 28288 121040 29996 121046
rect 110160 121110 110644 121116
rect 110160 121046 110166 121110
rect 110230 121046 110644 121110
rect 110160 121040 110644 121046
rect 111656 121116 111868 121182
rect 114376 121116 114588 121252
rect 115192 121246 116356 121252
rect 115192 121182 116286 121246
rect 116350 121182 116356 121246
rect 115192 121176 116356 121182
rect 136816 121176 137028 121312
rect 115192 121116 115404 121176
rect 111656 121110 115404 121116
rect 111656 121046 115334 121110
rect 115398 121046 115404 121110
rect 111656 121040 115404 121046
rect 28288 120904 28636 121040
rect 110160 120904 110508 121040
rect 28288 120844 28364 120904
rect 110160 120844 110236 120904
rect 22032 120768 23060 120844
rect 22032 120708 22108 120768
rect 22984 120708 23060 120768
rect 21760 120632 22108 120708
rect 22168 120632 22788 120708
rect 21760 120566 21972 120632
rect 21760 120502 21766 120566
rect 21830 120502 21972 120566
rect 21760 120496 21972 120502
rect 22168 120566 22380 120632
rect 22168 120502 22310 120566
rect 22374 120502 22380 120566
rect 22168 120496 22380 120502
rect 22576 120566 22788 120632
rect 22576 120502 22582 120566
rect 22646 120502 22788 120566
rect 22576 120496 22788 120502
rect 22984 120566 23196 120708
rect 22984 120502 22990 120566
rect 23054 120502 23196 120566
rect 22984 120496 23196 120502
rect 23392 120566 23604 120708
rect 28288 120632 28636 120844
rect 110160 120632 110508 120844
rect 115192 120702 115404 120708
rect 115192 120638 115334 120702
rect 115398 120638 115404 120702
rect 28560 120572 28636 120632
rect 110296 120572 110372 120632
rect 23392 120502 23398 120566
rect 23462 120502 23604 120566
rect 23392 120496 23604 120502
rect 28288 120360 28636 120572
rect 110160 120360 110508 120572
rect 115192 120566 115404 120638
rect 115192 120502 115198 120566
rect 115262 120502 115404 120566
rect 115192 120496 115404 120502
rect 115600 120566 115812 120708
rect 115600 120502 115742 120566
rect 115806 120502 115812 120566
rect 115600 120496 115812 120502
rect 116008 120572 116220 120708
rect 116416 120572 116628 120708
rect 116008 120566 116628 120572
rect 116008 120502 116014 120566
rect 116078 120502 116628 120566
rect 116008 120496 116628 120502
rect 116824 120702 117444 120708
rect 116824 120638 117374 120702
rect 117438 120638 117444 120702
rect 116824 120632 117444 120638
rect 116824 120566 117036 120632
rect 116824 120502 116966 120566
rect 117030 120502 117036 120566
rect 116824 120496 117036 120502
rect 134640 120566 135668 120572
rect 134640 120502 134646 120566
rect 134710 120502 135668 120566
rect 134640 120496 135668 120502
rect 116144 120436 116220 120496
rect 116144 120360 116492 120436
rect 134640 120430 134852 120496
rect 134640 120366 134646 120430
rect 134710 120366 134852 120430
rect 134640 120360 134852 120366
rect 135456 120360 135668 120496
rect 28424 120300 28500 120360
rect 110160 120300 110236 120360
rect 116416 120300 116492 120360
rect 21760 120294 21972 120300
rect 21760 120230 21766 120294
rect 21830 120230 21972 120294
rect 21760 120158 21972 120230
rect 21760 120094 21766 120158
rect 21830 120094 21972 120158
rect 21760 120088 21972 120094
rect 22168 120294 22380 120300
rect 22168 120230 22310 120294
rect 22374 120230 22380 120294
rect 22168 120088 22380 120230
rect 22576 120294 22788 120300
rect 22576 120230 22582 120294
rect 22646 120230 22788 120294
rect 22576 120158 22788 120230
rect 22576 120094 22582 120158
rect 22646 120094 22788 120158
rect 22576 120088 22788 120094
rect 22984 120294 23196 120300
rect 22984 120230 22990 120294
rect 23054 120230 23196 120294
rect 22984 120158 23196 120230
rect 22984 120094 23126 120158
rect 23190 120094 23196 120158
rect 22984 120088 23196 120094
rect 23392 120294 23604 120300
rect 23392 120230 23398 120294
rect 23462 120230 23604 120294
rect 23392 120158 23604 120230
rect 23392 120094 23534 120158
rect 23598 120094 23604 120158
rect 23392 120088 23604 120094
rect 28288 120088 28636 120300
rect 110160 120088 110508 120300
rect 115192 120294 115404 120300
rect 115192 120230 115198 120294
rect 115262 120230 115404 120294
rect 115192 120158 115404 120230
rect 115192 120094 115334 120158
rect 115398 120094 115404 120158
rect 115192 120088 115404 120094
rect 115600 120294 115812 120300
rect 115600 120230 115742 120294
rect 115806 120230 115812 120294
rect 115600 120158 115812 120230
rect 115600 120094 115742 120158
rect 115806 120094 115812 120158
rect 115600 120088 115812 120094
rect 116008 120294 116220 120300
rect 116008 120230 116014 120294
rect 116078 120230 116220 120294
rect 116008 120088 116220 120230
rect 116416 120088 116628 120300
rect 116824 120294 117036 120300
rect 116824 120230 116966 120294
rect 117030 120230 117036 120294
rect 116824 120158 117036 120230
rect 116824 120094 116830 120158
rect 116894 120094 117036 120158
rect 116824 120088 117036 120094
rect 28424 120028 28500 120088
rect 110296 120028 110372 120088
rect 116416 120028 116492 120088
rect 21760 119886 21972 119892
rect 21760 119822 21766 119886
rect 21830 119822 21972 119886
rect 1224 119750 1980 119756
rect 1224 119686 1230 119750
rect 1294 119688 1980 119750
rect 1294 119686 1798 119688
rect 1224 119680 1798 119686
rect 1768 119632 1798 119680
rect 1854 119632 1980 119688
rect 21760 119750 21972 119822
rect 21760 119686 21902 119750
rect 21966 119686 21972 119750
rect 21760 119680 21972 119686
rect 22168 119886 22788 119892
rect 22168 119822 22582 119886
rect 22646 119822 22788 119886
rect 22168 119816 22788 119822
rect 22168 119756 22380 119816
rect 22168 119680 22516 119756
rect 22576 119680 22788 119816
rect 22984 119886 23196 119892
rect 22984 119822 23126 119886
rect 23190 119822 23196 119886
rect 22984 119750 23196 119822
rect 22984 119686 22990 119750
rect 23054 119686 23196 119750
rect 22984 119680 23196 119686
rect 23392 119886 23604 119892
rect 23392 119822 23534 119886
rect 23598 119822 23604 119886
rect 23392 119750 23604 119822
rect 23392 119686 23398 119750
rect 23462 119686 23604 119750
rect 23392 119680 23604 119686
rect 28288 119816 28636 120028
rect 110160 119816 110508 120028
rect 116144 119952 116492 120028
rect 116144 119892 116220 119952
rect 28288 119756 28364 119816
rect 110432 119756 110508 119816
rect 1768 119544 1980 119632
rect 22440 119620 22516 119680
rect 22440 119544 22652 119620
rect 28288 119544 28636 119756
rect 22576 119484 22652 119544
rect 28560 119484 28636 119544
rect 21760 119478 21972 119484
rect 21760 119414 21902 119478
rect 21966 119414 21972 119478
rect 21760 119342 21972 119414
rect 21760 119278 21766 119342
rect 21830 119278 21972 119342
rect 21760 119272 21972 119278
rect 22168 119408 22788 119484
rect 22168 119348 22380 119408
rect 22168 119342 22516 119348
rect 22168 119278 22310 119342
rect 22374 119278 22446 119342
rect 22510 119278 22516 119342
rect 22168 119272 22516 119278
rect 22576 119272 22788 119408
rect 22984 119478 23196 119484
rect 22984 119414 22990 119478
rect 23054 119414 23196 119478
rect 22984 119342 23196 119414
rect 22984 119278 23126 119342
rect 23190 119278 23196 119342
rect 22984 119272 23196 119278
rect 23392 119478 23604 119484
rect 23392 119414 23398 119478
rect 23462 119414 23604 119478
rect 23392 119342 23604 119414
rect 23392 119278 23398 119342
rect 23462 119278 23604 119342
rect 23392 119272 23604 119278
rect 28288 119272 28636 119484
rect 110160 119544 110508 119756
rect 115192 119886 115404 119892
rect 115192 119822 115334 119886
rect 115398 119822 115404 119886
rect 115192 119750 115404 119822
rect 115192 119686 115198 119750
rect 115262 119686 115404 119750
rect 115192 119680 115404 119686
rect 115600 119886 115812 119892
rect 115600 119822 115742 119886
rect 115806 119822 115812 119886
rect 115600 119750 115812 119822
rect 115600 119686 115606 119750
rect 115670 119686 115812 119750
rect 115600 119680 115812 119686
rect 116008 119816 116628 119892
rect 116008 119680 116220 119816
rect 116416 119750 116628 119816
rect 116416 119686 116558 119750
rect 116622 119686 116628 119750
rect 116416 119680 116628 119686
rect 116824 119886 117036 119892
rect 116824 119822 116830 119886
rect 116894 119822 117036 119886
rect 116824 119750 117036 119822
rect 116824 119686 116966 119750
rect 117030 119686 117036 119750
rect 116824 119680 117036 119686
rect 136816 119750 137572 119756
rect 136816 119688 137502 119750
rect 136816 119632 136944 119688
rect 137000 119686 137502 119688
rect 137566 119686 137572 119750
rect 137000 119680 137572 119686
rect 137000 119632 137028 119680
rect 136816 119614 137028 119632
rect 136816 119550 136822 119614
rect 136886 119550 137028 119614
rect 136816 119544 137028 119550
rect 110160 119484 110236 119544
rect 110160 119272 110508 119484
rect 115192 119478 115404 119484
rect 115192 119414 115198 119478
rect 115262 119414 115404 119478
rect 115192 119342 115404 119414
rect 115192 119278 115334 119342
rect 115398 119278 115404 119342
rect 115192 119272 115404 119278
rect 115600 119478 115812 119484
rect 115600 119414 115606 119478
rect 115670 119414 115812 119478
rect 115600 119342 115812 119414
rect 115600 119278 115742 119342
rect 115806 119278 115812 119342
rect 115600 119272 115812 119278
rect 116008 119478 116628 119484
rect 116008 119414 116558 119478
rect 116622 119414 116628 119478
rect 116008 119408 116628 119414
rect 116008 119348 116220 119408
rect 116008 119342 116356 119348
rect 116008 119278 116014 119342
rect 116078 119278 116286 119342
rect 116350 119278 116356 119342
rect 116008 119272 116356 119278
rect 116416 119272 116628 119408
rect 116824 119478 117036 119484
rect 116824 119414 116966 119478
rect 117030 119414 117036 119478
rect 116824 119342 117036 119414
rect 116824 119278 116966 119342
rect 117030 119278 117036 119342
rect 116824 119272 117036 119278
rect 28288 119212 28364 119272
rect 110432 119212 110508 119272
rect 21760 119070 21972 119076
rect 21760 119006 21766 119070
rect 21830 119006 21972 119070
rect 21760 118864 21972 119006
rect 22168 119070 22380 119076
rect 22478 119070 22788 119076
rect 22168 119006 22310 119070
rect 22374 119006 22380 119070
rect 22440 119006 22446 119070
rect 22510 119006 22788 119070
rect 22168 118864 22380 119006
rect 22478 119000 22788 119006
rect 22576 118934 22788 119000
rect 22576 118870 22582 118934
rect 22646 118870 22788 118934
rect 22576 118864 22788 118870
rect 22984 119070 23196 119076
rect 22984 119006 23126 119070
rect 23190 119006 23196 119070
rect 22984 118934 23196 119006
rect 22984 118870 22990 118934
rect 23054 118870 23196 118934
rect 22984 118864 23196 118870
rect 23392 119070 23604 119076
rect 23392 119006 23398 119070
rect 23462 119006 23604 119070
rect 23392 118934 23604 119006
rect 23392 118870 23398 118934
rect 23462 118870 23604 118934
rect 23392 118864 23604 118870
rect 28288 119000 28636 119212
rect 110160 119000 110508 119212
rect 134640 119206 136892 119212
rect 134640 119142 136822 119206
rect 136886 119142 136892 119206
rect 134640 119136 136892 119142
rect 115192 119070 115404 119076
rect 115192 119006 115334 119070
rect 115398 119006 115404 119070
rect 28288 118940 28364 119000
rect 110160 118940 110236 119000
rect 21760 118804 21836 118864
rect 21760 118456 21972 118804
rect 28288 118798 28636 118940
rect 28288 118734 28566 118798
rect 28630 118734 28636 118798
rect 28288 118728 28636 118734
rect 110160 118798 110508 118940
rect 115192 118934 115404 119006
rect 115192 118870 115198 118934
rect 115262 118870 115404 118934
rect 115192 118864 115404 118870
rect 115600 119070 115812 119076
rect 115600 119006 115742 119070
rect 115806 119006 115812 119070
rect 115600 118934 115812 119006
rect 115600 118870 115606 118934
rect 115670 118870 115812 118934
rect 115600 118864 115812 118870
rect 116008 119070 116220 119076
rect 116318 119070 116628 119076
rect 116008 119006 116014 119070
rect 116078 119006 116220 119070
rect 116280 119006 116286 119070
rect 116350 119006 116628 119070
rect 116008 118864 116220 119006
rect 116318 119000 116628 119006
rect 116416 118940 116628 119000
rect 116318 118934 116628 118940
rect 116280 118870 116286 118934
rect 116350 118870 116628 118934
rect 116318 118864 116628 118870
rect 116824 119070 117036 119076
rect 116824 119006 116966 119070
rect 117030 119006 117036 119070
rect 116824 118864 117036 119006
rect 134640 119000 134852 119136
rect 135456 119000 135668 119136
rect 116960 118804 117036 118864
rect 110160 118734 110302 118798
rect 110366 118734 110508 118798
rect 110160 118728 110508 118734
rect 28560 118668 28636 118728
rect 110296 118668 110372 118728
rect 22168 118532 22380 118668
rect 22576 118662 22788 118668
rect 22576 118598 22582 118662
rect 22646 118598 22788 118662
rect 22168 118456 22516 118532
rect 22576 118456 22788 118598
rect 22984 118662 23196 118668
rect 22984 118598 22990 118662
rect 23054 118598 23196 118662
rect 22984 118526 23196 118598
rect 22984 118462 22990 118526
rect 23054 118462 23196 118526
rect 22984 118456 23196 118462
rect 23392 118662 23604 118668
rect 23392 118598 23398 118662
rect 23462 118598 23604 118662
rect 23392 118526 23604 118598
rect 23392 118462 23398 118526
rect 23462 118462 23604 118526
rect 23392 118456 23604 118462
rect 28288 118526 28636 118668
rect 28288 118462 28430 118526
rect 28494 118462 28566 118526
rect 28630 118462 28636 118526
rect 21760 118396 21836 118456
rect 22304 118396 22380 118456
rect 1224 118118 1980 118124
rect 1224 118054 1230 118118
rect 1294 118054 1980 118118
rect 1224 118048 1980 118054
rect 1768 118008 1980 118048
rect 1768 117952 1798 118008
rect 1854 117952 1980 118008
rect 1768 117912 1980 117952
rect 21760 118048 21972 118396
rect 22168 118118 22380 118396
rect 22440 118396 22516 118456
rect 22712 118396 22788 118456
rect 22440 118320 22788 118396
rect 22168 118054 22174 118118
rect 22238 118054 22380 118118
rect 22168 118048 22380 118054
rect 22576 118048 22788 118320
rect 22984 118254 23196 118260
rect 22984 118190 22990 118254
rect 23054 118190 23196 118254
rect 22984 118048 23196 118190
rect 23392 118254 23604 118260
rect 23392 118190 23398 118254
rect 23462 118190 23604 118254
rect 23392 118048 23604 118190
rect 28288 118184 28636 118462
rect 110160 118526 110508 118668
rect 110160 118462 110302 118526
rect 110366 118462 110508 118526
rect 110160 118254 110508 118462
rect 115192 118662 115404 118668
rect 115192 118598 115198 118662
rect 115262 118598 115404 118662
rect 115192 118526 115404 118598
rect 115192 118462 115198 118526
rect 115262 118462 115404 118526
rect 115192 118456 115404 118462
rect 115600 118662 115812 118668
rect 115600 118598 115606 118662
rect 115670 118598 115812 118662
rect 115600 118526 115812 118598
rect 115600 118462 115606 118526
rect 115670 118462 115812 118526
rect 115600 118456 115812 118462
rect 116008 118662 116356 118668
rect 116008 118598 116286 118662
rect 116350 118598 116356 118662
rect 116008 118592 116356 118598
rect 116008 118456 116220 118592
rect 116416 118456 116628 118668
rect 116008 118396 116084 118456
rect 116552 118396 116628 118456
rect 116008 118320 116628 118396
rect 110160 118190 110302 118254
rect 110366 118190 110508 118254
rect 110160 118184 110508 118190
rect 115192 118254 115404 118260
rect 115192 118190 115198 118254
rect 115262 118190 115404 118254
rect 21760 117988 21836 118048
rect 23120 117988 23196 118048
rect 23528 117988 23604 118048
rect 21760 117846 21972 117988
rect 21760 117782 21766 117846
rect 21830 117782 21972 117846
rect 21760 117776 21972 117782
rect 22168 117846 22380 117852
rect 22168 117782 22174 117846
rect 22238 117782 22380 117846
rect 22168 117640 22380 117782
rect 22304 117580 22380 117640
rect 21760 117574 21972 117580
rect 21760 117510 21766 117574
rect 21830 117510 21972 117574
rect 21760 117438 21972 117510
rect 21760 117374 21902 117438
rect 21966 117374 21972 117438
rect 21760 117368 21972 117374
rect 22168 117444 22380 117580
rect 22576 117640 22788 117852
rect 22984 117640 23196 117988
rect 22576 117580 22652 117640
rect 23120 117580 23196 117640
rect 22168 117438 22516 117444
rect 22168 117374 22446 117438
rect 22510 117374 22516 117438
rect 22168 117368 22516 117374
rect 22576 117368 22788 117580
rect 22576 117308 22652 117368
rect 22304 117232 22652 117308
rect 22984 117232 23196 117580
rect 22304 117172 22380 117232
rect 23120 117172 23196 117232
rect 21760 117166 21972 117172
rect 21760 117102 21902 117166
rect 21966 117102 21972 117166
rect 21760 117030 21972 117102
rect 21760 116966 21766 117030
rect 21830 116966 21972 117030
rect 21760 116960 21972 116966
rect 22168 117036 22380 117172
rect 22478 117166 22788 117172
rect 22440 117102 22446 117166
rect 22510 117102 22788 117166
rect 22478 117096 22788 117102
rect 22576 117036 22788 117096
rect 22168 116960 22788 117036
rect 22984 117030 23196 117172
rect 22984 116966 22990 117030
rect 23054 116966 23196 117030
rect 22984 116960 23196 116966
rect 23392 117640 23604 117988
rect 28288 118118 28636 118124
rect 28288 118054 28430 118118
rect 28494 118054 28636 118118
rect 28288 117982 28636 118054
rect 28288 117918 28430 117982
rect 28494 117918 28636 117982
rect 28288 117710 28636 117918
rect 28288 117646 28430 117710
rect 28494 117646 28636 117710
rect 23392 117580 23468 117640
rect 23392 117232 23604 117580
rect 28288 117574 28636 117646
rect 28288 117510 28566 117574
rect 28630 117510 28636 117574
rect 28288 117504 28636 117510
rect 110160 117982 110508 118124
rect 115192 118048 115404 118190
rect 115600 118254 115812 118260
rect 115600 118190 115606 118254
rect 115670 118190 115812 118254
rect 115600 118048 115812 118190
rect 116008 118124 116220 118320
rect 116008 118118 116356 118124
rect 116008 118054 116286 118118
rect 116350 118054 116356 118118
rect 116008 118048 116356 118054
rect 116416 118048 116628 118320
rect 116824 118456 117036 118804
rect 116824 118396 116900 118456
rect 116824 118048 117036 118396
rect 136816 118118 137572 118124
rect 136816 118054 137502 118118
rect 137566 118054 137572 118118
rect 136816 118048 137572 118054
rect 115328 117988 115404 118048
rect 115736 117988 115812 118048
rect 110160 117918 110302 117982
rect 110366 117918 110438 117982
rect 110502 117918 110508 117982
rect 110160 117710 110508 117918
rect 110160 117646 110438 117710
rect 110502 117646 110508 117710
rect 110160 117574 110508 117646
rect 110160 117510 110166 117574
rect 110230 117510 110508 117574
rect 110160 117504 110508 117510
rect 115192 117640 115404 117988
rect 115600 117640 115812 117988
rect 116824 117988 116900 118048
rect 136816 118008 137028 118048
rect 116008 117716 116220 117852
rect 116318 117846 116628 117852
rect 116280 117782 116286 117846
rect 116350 117782 116628 117846
rect 116318 117776 116628 117782
rect 116824 117846 117036 117988
rect 136816 117952 136944 118008
rect 137000 117952 137028 118008
rect 136816 117912 137028 117952
rect 116824 117782 116830 117846
rect 116894 117782 117036 117846
rect 116824 117776 117036 117782
rect 116416 117716 116628 117776
rect 116008 117640 116628 117716
rect 115192 117580 115268 117640
rect 115736 117580 115812 117640
rect 116144 117580 116220 117640
rect 116552 117580 116628 117640
rect 134640 117710 134852 117716
rect 134640 117646 134646 117710
rect 134710 117646 134852 117710
rect 134640 117580 134852 117646
rect 135456 117580 135668 117716
rect 23392 117172 23468 117232
rect 23392 117030 23604 117172
rect 23392 116966 23534 117030
rect 23598 116966 23604 117030
rect 23392 116960 23604 116966
rect 28288 117166 28636 117308
rect 28288 117102 28430 117166
rect 28494 117102 28566 117166
rect 28630 117102 28636 117166
rect 28288 116960 28636 117102
rect 110160 117302 110508 117308
rect 110160 117238 110166 117302
rect 110230 117238 110508 117302
rect 110160 116960 110508 117238
rect 115192 117232 115404 117580
rect 115600 117232 115812 117580
rect 116008 117368 116220 117580
rect 116416 117438 116628 117580
rect 116416 117374 116558 117438
rect 116622 117374 116628 117438
rect 116416 117368 116628 117374
rect 116824 117574 117036 117580
rect 116824 117510 116830 117574
rect 116894 117510 117036 117574
rect 116824 117438 117036 117510
rect 134640 117504 135668 117580
rect 116824 117374 116966 117438
rect 117030 117374 117036 117438
rect 116824 117368 117036 117374
rect 115192 117172 115268 117232
rect 115600 117172 115676 117232
rect 115192 117030 115404 117172
rect 115192 116966 115334 117030
rect 115398 116966 115404 117030
rect 115192 116960 115404 116966
rect 115600 117030 115812 117172
rect 115600 116966 115742 117030
rect 115806 116966 115812 117030
rect 115600 116960 115812 116966
rect 22168 116824 22380 116960
rect 22576 116824 22788 116960
rect 28288 116900 28364 116960
rect 110160 116900 110236 116960
rect 28288 116894 28636 116900
rect 28288 116830 28430 116894
rect 28494 116830 28636 116894
rect 22168 116764 22244 116824
rect 22576 116764 22652 116824
rect 21760 116758 21972 116764
rect 21760 116694 21766 116758
rect 21830 116694 21972 116758
rect 21760 116622 21972 116694
rect 21760 116558 21902 116622
rect 21966 116558 21972 116622
rect 21760 116552 21972 116558
rect 22168 116552 22380 116764
rect 22576 116552 22788 116764
rect 22984 116758 23196 116764
rect 22984 116694 22990 116758
rect 23054 116694 23196 116758
rect 22984 116622 23196 116694
rect 22984 116558 23126 116622
rect 23190 116558 23196 116622
rect 22984 116552 23196 116558
rect 23392 116758 23604 116764
rect 23392 116694 23534 116758
rect 23598 116694 23604 116758
rect 23392 116622 23604 116694
rect 28288 116758 28636 116830
rect 28288 116694 28566 116758
rect 28630 116694 28636 116758
rect 28288 116688 28636 116694
rect 110160 116688 110508 116900
rect 116008 116824 116220 117172
rect 116416 117166 116628 117172
rect 116416 117102 116558 117166
rect 116622 117102 116628 117166
rect 116416 116900 116628 117102
rect 116824 117166 117036 117172
rect 116824 117102 116966 117166
rect 117030 117102 117036 117166
rect 116824 117030 117036 117102
rect 116824 116966 116830 117030
rect 116894 116966 117036 117030
rect 116824 116960 117036 116966
rect 116144 116764 116220 116824
rect 116280 116824 116628 116900
rect 116280 116764 116356 116824
rect 28424 116628 28500 116688
rect 110432 116628 110508 116688
rect 23392 116558 23398 116622
rect 23462 116558 23604 116622
rect 23392 116552 23604 116558
rect 22576 116492 22652 116552
rect 22304 116416 22652 116492
rect 22304 116356 22380 116416
rect 1224 116350 1980 116356
rect 1224 116286 1230 116350
rect 1294 116328 1980 116350
rect 1294 116286 1798 116328
rect 1224 116280 1798 116286
rect 1768 116272 1798 116280
rect 1854 116272 1980 116328
rect 1768 116144 1980 116272
rect 21760 116350 21972 116356
rect 21760 116286 21902 116350
rect 21966 116286 21972 116350
rect 21760 116214 21972 116286
rect 21760 116150 21902 116214
rect 21966 116150 21972 116214
rect 21760 116144 21972 116150
rect 22168 116280 22788 116356
rect 22168 116144 22380 116280
rect 22576 116220 22788 116280
rect 22478 116214 22788 116220
rect 22440 116150 22446 116214
rect 22510 116150 22788 116214
rect 22478 116144 22788 116150
rect 22984 116350 23196 116356
rect 22984 116286 23126 116350
rect 23190 116286 23196 116350
rect 22984 116214 23196 116286
rect 22984 116150 22990 116214
rect 23054 116150 23196 116214
rect 22984 116144 23196 116150
rect 23392 116350 23604 116356
rect 23392 116286 23398 116350
rect 23462 116286 23604 116350
rect 23392 116214 23604 116286
rect 23392 116150 23398 116214
rect 23462 116150 23604 116214
rect 23392 116144 23604 116150
rect 28288 116350 28636 116628
rect 28288 116286 28566 116350
rect 28630 116286 28636 116350
rect 28288 116144 28636 116286
rect 110160 116144 110508 116628
rect 115192 116758 115404 116764
rect 115192 116694 115334 116758
rect 115398 116694 115404 116758
rect 115192 116622 115404 116694
rect 115192 116558 115198 116622
rect 115262 116558 115404 116622
rect 115192 116552 115404 116558
rect 115600 116758 115812 116764
rect 115600 116694 115742 116758
rect 115806 116694 115812 116758
rect 115600 116622 115812 116694
rect 115600 116558 115742 116622
rect 115806 116558 115812 116622
rect 115600 116552 115812 116558
rect 116008 116688 116356 116764
rect 116008 116628 116220 116688
rect 116416 116628 116628 116764
rect 116008 116622 116628 116628
rect 116008 116558 116558 116622
rect 116622 116558 116628 116622
rect 116008 116552 116628 116558
rect 116824 116758 117036 116764
rect 116824 116694 116830 116758
rect 116894 116694 117036 116758
rect 116824 116622 117036 116694
rect 116824 116558 116966 116622
rect 117030 116558 117036 116622
rect 116824 116552 117036 116558
rect 115192 116350 115404 116356
rect 115192 116286 115198 116350
rect 115262 116286 115404 116350
rect 115192 116214 115404 116286
rect 115192 116150 115198 116214
rect 115262 116150 115404 116214
rect 115192 116144 115404 116150
rect 115600 116350 115812 116356
rect 115600 116286 115742 116350
rect 115806 116286 115812 116350
rect 115600 116214 115812 116286
rect 115600 116150 115742 116214
rect 115806 116150 115812 116214
rect 115600 116144 115812 116150
rect 116008 116350 116628 116356
rect 116008 116286 116558 116350
rect 116622 116286 116628 116350
rect 116008 116280 116628 116286
rect 116008 116220 116220 116280
rect 116008 116214 116356 116220
rect 116008 116150 116014 116214
rect 116078 116150 116286 116214
rect 116350 116150 116356 116214
rect 116008 116144 116356 116150
rect 116416 116144 116628 116280
rect 116824 116350 117036 116356
rect 116824 116286 116966 116350
rect 117030 116286 117036 116350
rect 116824 116214 117036 116286
rect 116824 116150 116966 116214
rect 117030 116150 117036 116214
rect 116824 116144 117036 116150
rect 134640 116220 134852 116356
rect 135456 116328 137028 116356
rect 135456 116280 136944 116328
rect 135456 116220 135668 116280
rect 134640 116144 135668 116220
rect 136816 116272 136944 116280
rect 137000 116272 137028 116328
rect 136816 116220 137028 116272
rect 136816 116214 137572 116220
rect 136816 116150 137502 116214
rect 137566 116150 137572 116214
rect 136816 116144 137572 116150
rect 28424 116084 28500 116144
rect 110160 116084 110236 116144
rect 21760 115942 21972 115948
rect 21760 115878 21902 115942
rect 21966 115878 21972 115942
rect 21760 115806 21972 115878
rect 21760 115742 21766 115806
rect 21830 115742 21972 115806
rect 21760 115736 21972 115742
rect 22168 115942 22516 115948
rect 22168 115878 22446 115942
rect 22510 115878 22516 115942
rect 22168 115872 22516 115878
rect 22168 115812 22380 115872
rect 22576 115812 22788 115948
rect 22168 115806 22788 115812
rect 22168 115742 22174 115806
rect 22238 115742 22582 115806
rect 22646 115742 22788 115806
rect 22168 115736 22788 115742
rect 22984 115942 23196 115948
rect 22984 115878 22990 115942
rect 23054 115878 23196 115942
rect 22984 115806 23196 115878
rect 22984 115742 23126 115806
rect 23190 115742 23196 115806
rect 22984 115736 23196 115742
rect 23392 115942 23604 115948
rect 23392 115878 23398 115942
rect 23462 115878 23604 115942
rect 23392 115806 23604 115878
rect 28288 115872 28636 116084
rect 110160 115872 110508 116084
rect 28424 115812 28500 115872
rect 110432 115812 110508 115872
rect 23392 115742 23534 115806
rect 23598 115742 23604 115806
rect 23392 115736 23604 115742
rect 28288 115600 28636 115812
rect 110160 115600 110508 115812
rect 115192 115942 115404 115948
rect 115192 115878 115198 115942
rect 115262 115878 115404 115942
rect 115192 115806 115404 115878
rect 115192 115742 115334 115806
rect 115398 115742 115404 115806
rect 115192 115736 115404 115742
rect 115600 115942 115812 115948
rect 115600 115878 115742 115942
rect 115806 115878 115812 115942
rect 115600 115806 115812 115878
rect 115600 115742 115742 115806
rect 115806 115742 115812 115806
rect 115600 115736 115812 115742
rect 116008 115942 116220 115948
rect 116318 115942 116628 115948
rect 116008 115878 116014 115942
rect 116078 115878 116220 115942
rect 116280 115878 116286 115942
rect 116350 115878 116628 115942
rect 116008 115736 116220 115878
rect 116318 115872 116628 115878
rect 116416 115736 116628 115872
rect 116824 115942 117036 115948
rect 116824 115878 116966 115942
rect 117030 115878 117036 115942
rect 116824 115806 117036 115878
rect 116824 115742 116830 115806
rect 116894 115742 117036 115806
rect 116824 115736 117036 115742
rect 116416 115676 116492 115736
rect 116144 115600 116492 115676
rect 28288 115540 28364 115600
rect 110296 115540 110372 115600
rect 116144 115540 116220 115600
rect 21760 115534 21972 115540
rect 21760 115470 21766 115534
rect 21830 115470 21972 115534
rect 21760 115398 21972 115470
rect 21760 115334 21902 115398
rect 21966 115334 21972 115398
rect 21760 115328 21972 115334
rect 22168 115534 22380 115540
rect 22168 115470 22174 115534
rect 22238 115470 22380 115534
rect 22168 115328 22380 115470
rect 22576 115534 22788 115540
rect 22576 115470 22582 115534
rect 22646 115470 22788 115534
rect 22576 115398 22788 115470
rect 22576 115334 22718 115398
rect 22782 115334 22788 115398
rect 22576 115328 22788 115334
rect 22984 115534 23196 115540
rect 22984 115470 23126 115534
rect 23190 115470 23196 115534
rect 22984 115398 23196 115470
rect 22984 115334 23126 115398
rect 23190 115334 23196 115398
rect 22984 115328 23196 115334
rect 23392 115534 23604 115540
rect 23392 115470 23534 115534
rect 23598 115470 23604 115534
rect 23392 115398 23604 115470
rect 23392 115334 23398 115398
rect 23462 115334 23604 115398
rect 23392 115328 23604 115334
rect 28288 115328 28636 115540
rect 110160 115328 110508 115540
rect 115192 115534 115404 115540
rect 115192 115470 115334 115534
rect 115398 115470 115404 115534
rect 115192 115398 115404 115470
rect 115192 115334 115334 115398
rect 115398 115334 115404 115398
rect 115192 115328 115404 115334
rect 115600 115534 115812 115540
rect 115600 115470 115742 115534
rect 115806 115470 115812 115534
rect 115600 115398 115812 115470
rect 115600 115334 115606 115398
rect 115670 115334 115812 115398
rect 115600 115328 115812 115334
rect 116008 115464 116628 115540
rect 116008 115328 116220 115464
rect 116416 115398 116628 115464
rect 116416 115334 116558 115398
rect 116622 115334 116628 115398
rect 116416 115328 116628 115334
rect 116824 115534 117036 115540
rect 116824 115470 116830 115534
rect 116894 115470 117036 115534
rect 116824 115398 117036 115470
rect 116824 115334 116966 115398
rect 117030 115334 117036 115398
rect 116824 115328 117036 115334
rect 28560 115268 28636 115328
rect 110432 115268 110508 115328
rect 21760 115126 21972 115132
rect 21760 115062 21902 115126
rect 21966 115062 21972 115126
rect 21760 114920 21972 115062
rect 22168 114996 22380 115132
rect 22576 115126 22788 115132
rect 22576 115062 22718 115126
rect 22782 115062 22788 115126
rect 22576 114996 22788 115062
rect 22168 114920 22788 114996
rect 22984 115126 23196 115132
rect 22984 115062 23126 115126
rect 23190 115062 23196 115126
rect 22984 114990 23196 115062
rect 22984 114926 23126 114990
rect 23190 114926 23196 114990
rect 22984 114920 23196 114926
rect 23392 115126 23604 115132
rect 23392 115062 23398 115126
rect 23462 115062 23604 115126
rect 23392 114990 23604 115062
rect 28288 115056 28636 115268
rect 110160 115056 110508 115268
rect 28424 114996 28500 115056
rect 110432 114996 110508 115056
rect 23392 114926 23534 114990
rect 23598 114926 23604 114990
rect 23392 114920 23604 114926
rect 21896 114860 21972 114920
rect 1224 114718 1980 114724
rect 1224 114654 1230 114718
rect 1294 114654 1980 114718
rect 1224 114648 1980 114654
rect 1768 114592 1798 114648
rect 1854 114592 1980 114648
rect 1768 114512 1980 114592
rect 21760 114512 21972 114860
rect 22304 114860 22380 114920
rect 22304 114784 22652 114860
rect 28288 114784 28636 114996
rect 110160 114854 110508 114996
rect 115192 115126 115404 115132
rect 115192 115062 115334 115126
rect 115398 115062 115404 115126
rect 115192 114990 115404 115062
rect 115192 114926 115334 114990
rect 115398 114926 115404 114990
rect 115192 114920 115404 114926
rect 115600 115126 115812 115132
rect 115600 115062 115606 115126
rect 115670 115062 115812 115126
rect 115600 114990 115812 115062
rect 115600 114926 115742 114990
rect 115806 114926 115812 114990
rect 115600 114920 115812 114926
rect 116008 114996 116220 115132
rect 116416 115126 116628 115132
rect 116416 115062 116558 115126
rect 116622 115062 116628 115126
rect 116416 114996 116628 115062
rect 116008 114990 116628 114996
rect 116008 114926 116150 114990
rect 116214 114926 116628 114990
rect 116008 114920 116628 114926
rect 116824 115126 117036 115132
rect 116824 115062 116966 115126
rect 117030 115062 117036 115126
rect 116824 114920 117036 115062
rect 110160 114790 110302 114854
rect 110366 114790 110508 114854
rect 110160 114784 110508 114790
rect 116144 114860 116220 114920
rect 116960 114860 117036 114920
rect 116144 114784 116492 114860
rect 22576 114724 22652 114784
rect 28424 114724 28500 114784
rect 110432 114724 110508 114784
rect 116416 114724 116492 114784
rect 22168 114512 22380 114724
rect 22576 114512 22788 114724
rect 22984 114718 23196 114724
rect 22984 114654 23126 114718
rect 23190 114654 23196 114718
rect 22984 114582 23196 114654
rect 22984 114518 22990 114582
rect 23054 114518 23196 114582
rect 22984 114512 23196 114518
rect 23392 114718 23604 114724
rect 23392 114654 23534 114718
rect 23598 114654 23604 114718
rect 23392 114582 23604 114654
rect 23392 114518 23398 114582
rect 23462 114518 23604 114582
rect 23392 114512 23604 114518
rect 21760 114452 21836 114512
rect 22168 114452 22244 114512
rect 22576 114452 22652 114512
rect 21760 114104 21972 114452
rect 22168 114316 22380 114452
rect 22576 114316 22788 114452
rect 22168 114240 22788 114316
rect 22168 114180 22380 114240
rect 22168 114174 22516 114180
rect 22168 114110 22446 114174
rect 22510 114110 22516 114174
rect 22168 114104 22516 114110
rect 22576 114104 22788 114240
rect 22984 114310 23196 114316
rect 22984 114246 22990 114310
rect 23054 114246 23196 114310
rect 22984 114174 23196 114246
rect 22984 114110 23126 114174
rect 23190 114110 23196 114174
rect 22984 114104 23196 114110
rect 23392 114310 23604 114316
rect 23392 114246 23398 114310
rect 23462 114246 23604 114310
rect 23392 114174 23604 114246
rect 28288 114240 28636 114724
rect 110160 114582 110508 114724
rect 110160 114518 110302 114582
rect 110366 114518 110508 114582
rect 110160 114240 110508 114518
rect 115192 114718 115404 114724
rect 115192 114654 115334 114718
rect 115398 114654 115404 114718
rect 115192 114582 115404 114654
rect 115192 114518 115198 114582
rect 115262 114518 115404 114582
rect 115192 114512 115404 114518
rect 115600 114718 115812 114724
rect 115600 114654 115742 114718
rect 115806 114654 115812 114718
rect 115600 114582 115812 114654
rect 115600 114518 115742 114582
rect 115806 114518 115812 114582
rect 115600 114512 115812 114518
rect 116008 114718 116220 114724
rect 116008 114654 116150 114718
rect 116214 114654 116220 114718
rect 116008 114512 116220 114654
rect 116416 114512 116628 114724
rect 116144 114452 116220 114512
rect 116552 114452 116628 114512
rect 115192 114310 115404 114316
rect 115192 114246 115198 114310
rect 115262 114246 115404 114310
rect 28424 114180 28500 114240
rect 110160 114180 110236 114240
rect 23392 114110 23398 114174
rect 23462 114110 23604 114174
rect 23392 114104 23604 114110
rect 21760 114044 21836 114104
rect 21760 113902 21972 114044
rect 28288 114038 28636 114180
rect 28288 113974 28566 114038
rect 28630 113974 28636 114038
rect 28288 113968 28636 113974
rect 110160 113968 110508 114180
rect 115192 114174 115404 114246
rect 115192 114110 115198 114174
rect 115262 114110 115404 114174
rect 115192 114104 115404 114110
rect 115600 114310 115812 114316
rect 115600 114246 115742 114310
rect 115806 114246 115812 114310
rect 115600 114174 115812 114246
rect 115600 114110 115606 114174
rect 115670 114110 115812 114174
rect 115600 114104 115812 114110
rect 116008 114104 116220 114452
rect 116416 114174 116628 114452
rect 116416 114110 116422 114174
rect 116486 114110 116628 114174
rect 116416 114104 116628 114110
rect 116824 114512 117036 114860
rect 134640 114854 138252 114860
rect 134640 114790 138182 114854
rect 138246 114790 138252 114854
rect 134640 114784 138252 114790
rect 134640 114648 134852 114784
rect 135456 114724 135668 114784
rect 135358 114718 135668 114724
rect 135320 114654 135326 114718
rect 135390 114654 135668 114718
rect 135358 114648 135668 114654
rect 136816 114648 137028 114724
rect 136816 114592 136944 114648
rect 137000 114592 137028 114648
rect 136816 114588 137028 114592
rect 136816 114582 137572 114588
rect 136816 114518 137502 114582
rect 137566 114518 137572 114582
rect 136816 114512 137572 114518
rect 116824 114452 116900 114512
rect 116824 114104 117036 114452
rect 116824 114044 116900 114104
rect 28560 113908 28636 113968
rect 110296 113908 110372 113968
rect 21760 113838 21766 113902
rect 21830 113838 21972 113902
rect 21760 113832 21972 113838
rect 22168 113696 22380 113908
rect 22478 113902 22788 113908
rect 22440 113838 22446 113902
rect 22510 113838 22788 113902
rect 22478 113832 22788 113838
rect 22576 113696 22788 113832
rect 22984 113902 23196 113908
rect 22984 113838 23126 113902
rect 23190 113838 23196 113902
rect 22984 113696 23196 113838
rect 23392 113902 23604 113908
rect 23392 113838 23398 113902
rect 23462 113838 23604 113902
rect 23392 113696 23604 113838
rect 22168 113636 22244 113696
rect 22576 113636 22652 113696
rect 22984 113636 23060 113696
rect 23528 113636 23604 113696
rect 21760 113630 21972 113636
rect 21760 113566 21766 113630
rect 21830 113566 21972 113630
rect 21760 113494 21972 113566
rect 21760 113430 21902 113494
rect 21966 113430 21972 113494
rect 21760 113424 21972 113430
rect 22168 113494 22380 113636
rect 22576 113500 22788 113636
rect 22478 113494 22788 113500
rect 22168 113430 22174 113494
rect 22238 113430 22380 113494
rect 22440 113430 22446 113494
rect 22510 113430 22788 113494
rect 22168 113424 22380 113430
rect 22478 113424 22788 113430
rect 22984 113288 23196 113636
rect 23392 113288 23604 113636
rect 28288 113766 28636 113908
rect 28288 113702 28294 113766
rect 28358 113702 28566 113766
rect 28630 113702 28636 113766
rect 28288 113560 28636 113702
rect 110160 113630 110508 113908
rect 115192 113902 115404 113908
rect 115192 113838 115198 113902
rect 115262 113838 115404 113902
rect 115192 113696 115404 113838
rect 115600 113902 115812 113908
rect 115600 113838 115606 113902
rect 115670 113838 115812 113902
rect 115600 113696 115812 113838
rect 115328 113636 115404 113696
rect 115736 113636 115812 113696
rect 110160 113566 110438 113630
rect 110502 113566 110508 113630
rect 110160 113560 110508 113566
rect 23120 113228 23196 113288
rect 23528 113228 23604 113288
rect 21760 113222 21972 113228
rect 21760 113158 21902 113222
rect 21966 113158 21972 113222
rect 1224 113086 1980 113092
rect 1224 113022 1230 113086
rect 1294 113022 1980 113086
rect 1224 113016 1980 113022
rect 21760 113086 21972 113158
rect 21760 113022 21902 113086
rect 21966 113022 21972 113086
rect 21760 113016 21972 113022
rect 22168 113222 22516 113228
rect 22168 113158 22174 113222
rect 22238 113158 22446 113222
rect 22510 113158 22516 113222
rect 22168 113152 22516 113158
rect 1768 112968 1980 113016
rect 1768 112912 1798 112968
rect 1854 112912 1980 112968
rect 1768 112880 1980 112912
rect 22168 112956 22380 113152
rect 22576 112956 22788 113228
rect 22984 113086 23196 113228
rect 22984 113022 22990 113086
rect 23054 113022 23196 113086
rect 22984 113016 23196 113022
rect 23392 113086 23604 113228
rect 23392 113022 23398 113086
rect 23462 113022 23604 113086
rect 23392 113016 23604 113022
rect 28288 113358 28636 113364
rect 28288 113294 28294 113358
rect 28358 113294 28636 113358
rect 28288 113222 28636 113294
rect 28288 113158 28294 113222
rect 28358 113158 28636 113222
rect 28288 113016 28636 113158
rect 110160 113358 110508 113364
rect 110160 113294 110438 113358
rect 110502 113294 110508 113358
rect 110160 113016 110508 113294
rect 115192 113288 115404 113636
rect 115600 113288 115812 113636
rect 116008 113696 116220 113908
rect 116416 113902 116628 113908
rect 116416 113838 116422 113902
rect 116486 113838 116628 113902
rect 116416 113696 116628 113838
rect 116824 113902 117036 114044
rect 116824 113838 116830 113902
rect 116894 113838 117036 113902
rect 116824 113832 117036 113838
rect 116008 113636 116084 113696
rect 116416 113636 116492 113696
rect 116008 113560 116628 113636
rect 116008 113424 116220 113560
rect 116416 113424 116628 113560
rect 116824 113630 117036 113636
rect 116824 113566 116830 113630
rect 116894 113566 117036 113630
rect 116824 113494 117036 113566
rect 116824 113430 116830 113494
rect 116894 113430 117036 113494
rect 116824 113424 117036 113430
rect 134640 113424 135668 113500
rect 116416 113364 116492 113424
rect 115192 113228 115268 113288
rect 115736 113228 115812 113288
rect 116144 113288 116492 113364
rect 134640 113288 134852 113424
rect 135456 113364 135668 113424
rect 135456 113358 136892 113364
rect 135456 113294 136822 113358
rect 136886 113294 136892 113358
rect 135456 113288 136892 113294
rect 116144 113228 116220 113288
rect 115192 113086 115404 113228
rect 115192 113022 115198 113086
rect 115262 113022 115404 113086
rect 115192 113016 115404 113022
rect 115600 113086 115812 113228
rect 115600 113022 115606 113086
rect 115670 113022 115812 113086
rect 115600 113016 115812 113022
rect 116008 113152 116628 113228
rect 22168 112880 22788 112956
rect 22304 112820 22380 112880
rect 22712 112820 22788 112880
rect 28288 112956 28364 113016
rect 110432 112956 110508 113016
rect 28288 112950 28636 112956
rect 28288 112886 28294 112950
rect 28358 112886 28636 112950
rect 21760 112814 21972 112820
rect 21760 112750 21902 112814
rect 21966 112750 21972 112814
rect 21760 112678 21972 112750
rect 21760 112614 21766 112678
rect 21830 112614 21972 112678
rect 21760 112608 21972 112614
rect 22168 112678 22380 112820
rect 22168 112614 22174 112678
rect 22238 112614 22380 112678
rect 22168 112608 22380 112614
rect 22576 112608 22788 112820
rect 22984 112814 23196 112820
rect 22984 112750 22990 112814
rect 23054 112750 23196 112814
rect 22984 112678 23196 112750
rect 22984 112614 23126 112678
rect 23190 112614 23196 112678
rect 22984 112608 23196 112614
rect 23392 112814 23604 112820
rect 23392 112750 23398 112814
rect 23462 112750 23604 112814
rect 23392 112678 23604 112750
rect 28288 112744 28636 112886
rect 28560 112684 28636 112744
rect 23392 112614 23534 112678
rect 23598 112614 23604 112678
rect 23392 112608 23604 112614
rect 21760 112406 21972 112412
rect 21760 112342 21766 112406
rect 21830 112342 21972 112406
rect 21760 112270 21972 112342
rect 21760 112206 21902 112270
rect 21966 112206 21972 112270
rect 21760 112200 21972 112206
rect 22168 112406 22380 112412
rect 22168 112342 22174 112406
rect 22238 112342 22380 112406
rect 22168 112270 22380 112342
rect 22168 112206 22310 112270
rect 22374 112206 22380 112270
rect 22168 112200 22380 112206
rect 22576 112200 22788 112412
rect 22984 112406 23196 112412
rect 22984 112342 23126 112406
rect 23190 112342 23196 112406
rect 22984 112270 23196 112342
rect 22984 112206 23126 112270
rect 23190 112206 23196 112270
rect 22984 112200 23196 112206
rect 23392 112406 23604 112412
rect 23392 112342 23534 112406
rect 23598 112342 23604 112406
rect 23392 112270 23604 112342
rect 23392 112206 23398 112270
rect 23462 112206 23604 112270
rect 23392 112200 23604 112206
rect 28288 112406 28636 112684
rect 28288 112342 28430 112406
rect 28494 112342 28636 112406
rect 28288 112200 28636 112342
rect 110160 112744 110508 112956
rect 116008 112880 116220 113152
rect 116144 112820 116220 112880
rect 115192 112814 115404 112820
rect 115192 112750 115198 112814
rect 115262 112750 115404 112814
rect 110160 112684 110236 112744
rect 110160 112406 110508 112684
rect 115192 112678 115404 112750
rect 115192 112614 115198 112678
rect 115262 112614 115404 112678
rect 115192 112608 115404 112614
rect 115600 112814 115812 112820
rect 115600 112750 115606 112814
rect 115670 112750 115812 112814
rect 115600 112678 115812 112750
rect 115600 112614 115742 112678
rect 115806 112614 115812 112678
rect 115600 112608 115812 112614
rect 116008 112678 116220 112820
rect 116008 112614 116150 112678
rect 116214 112614 116220 112678
rect 116008 112608 116220 112614
rect 116416 112880 116628 113152
rect 116824 113222 117036 113228
rect 116824 113158 116830 113222
rect 116894 113158 117036 113222
rect 116824 113086 117036 113158
rect 116824 113022 116966 113086
rect 117030 113022 117036 113086
rect 116824 113016 117036 113022
rect 136816 113086 137028 113092
rect 136816 113022 136822 113086
rect 136886 113022 137028 113086
rect 136816 112968 137028 113022
rect 136816 112912 136944 112968
rect 137000 112956 137028 112968
rect 137000 112950 137572 112956
rect 137000 112912 137502 112950
rect 136816 112886 137502 112912
rect 137566 112886 137572 112950
rect 136816 112880 137572 112886
rect 116416 112820 116492 112880
rect 116416 112608 116628 112820
rect 116824 112814 117036 112820
rect 116824 112750 116966 112814
rect 117030 112750 117036 112814
rect 116824 112678 117036 112750
rect 136192 112683 136258 112684
rect 116824 112614 116830 112678
rect 116894 112614 117036 112678
rect 136150 112619 136193 112683
rect 136257 112619 136300 112683
rect 136192 112618 136258 112619
rect 116824 112608 117036 112614
rect 110160 112342 110302 112406
rect 110366 112342 110508 112406
rect 110160 112200 110508 112342
rect 115192 112406 115404 112412
rect 115192 112342 115198 112406
rect 115262 112342 115404 112406
rect 115192 112270 115404 112342
rect 115192 112206 115198 112270
rect 115262 112206 115404 112270
rect 115192 112200 115404 112206
rect 115600 112406 115812 112412
rect 115600 112342 115742 112406
rect 115806 112342 115812 112406
rect 115600 112270 115812 112342
rect 115600 112206 115742 112270
rect 115806 112206 115812 112270
rect 115600 112200 115812 112206
rect 116008 112406 116220 112412
rect 116008 112342 116150 112406
rect 116214 112342 116220 112406
rect 116008 112270 116220 112342
rect 116008 112206 116014 112270
rect 116078 112206 116220 112270
rect 116008 112200 116220 112206
rect 116416 112270 116628 112412
rect 116416 112206 116422 112270
rect 116486 112206 116628 112270
rect 116416 112200 116628 112206
rect 116824 112406 117036 112412
rect 116824 112342 116830 112406
rect 116894 112342 117036 112406
rect 116824 112270 117036 112342
rect 116824 112206 116830 112270
rect 116894 112206 117036 112270
rect 116824 112200 117036 112206
rect 22576 112140 22652 112200
rect 28560 112140 28636 112200
rect 110432 112140 110508 112200
rect 22304 112064 22652 112140
rect 28288 112134 28636 112140
rect 28288 112070 28430 112134
rect 28494 112070 28636 112134
rect 22304 112004 22380 112064
rect 21760 111998 21972 112004
rect 21760 111934 21902 111998
rect 21966 111934 21972 111998
rect 21760 111862 21972 111934
rect 21760 111798 21902 111862
rect 21966 111798 21972 111862
rect 21760 111792 21972 111798
rect 22168 111998 22788 112004
rect 22168 111934 22310 111998
rect 22374 111934 22788 111998
rect 22168 111928 22788 111934
rect 22168 111862 22380 111928
rect 22168 111798 22174 111862
rect 22238 111798 22380 111862
rect 22168 111792 22380 111798
rect 22576 111862 22788 111928
rect 22576 111798 22718 111862
rect 22782 111798 22788 111862
rect 22576 111792 22788 111798
rect 22984 111998 23196 112004
rect 22984 111934 23126 111998
rect 23190 111934 23196 111998
rect 22984 111862 23196 111934
rect 22984 111798 22990 111862
rect 23054 111798 23196 111862
rect 22984 111792 23196 111798
rect 23392 111998 23604 112004
rect 23392 111934 23398 111998
rect 23462 111934 23604 111998
rect 23392 111862 23604 111934
rect 28288 111928 28636 112070
rect 110160 112134 110508 112140
rect 110160 112070 110302 112134
rect 110366 112070 110508 112134
rect 110160 111928 110508 112070
rect 134640 112134 135396 112140
rect 134640 112070 135326 112134
rect 135390 112070 135396 112134
rect 134640 112064 135396 112070
rect 134640 112004 134852 112064
rect 135456 112004 135668 112140
rect 28560 111868 28636 111928
rect 110432 111868 110508 111928
rect 23392 111798 23398 111862
rect 23462 111798 23604 111862
rect 23392 111792 23604 111798
rect 28288 111656 28636 111868
rect 110160 111656 110508 111868
rect 115192 111998 115404 112004
rect 115192 111934 115198 111998
rect 115262 111934 115404 111998
rect 115192 111862 115404 111934
rect 115192 111798 115334 111862
rect 115398 111798 115404 111862
rect 115192 111792 115404 111798
rect 115600 111998 115812 112004
rect 115600 111934 115742 111998
rect 115806 111934 115812 111998
rect 115600 111862 115812 111934
rect 115600 111798 115606 111862
rect 115670 111798 115812 111862
rect 115600 111792 115812 111798
rect 116008 111998 116220 112004
rect 116008 111934 116014 111998
rect 116078 111934 116220 111998
rect 116008 111868 116220 111934
rect 116416 111998 116628 112004
rect 116416 111934 116422 111998
rect 116486 111934 116628 111998
rect 116416 111868 116628 111934
rect 116008 111862 116628 111868
rect 116008 111798 116014 111862
rect 116078 111798 116628 111862
rect 116008 111792 116628 111798
rect 116824 111998 117036 112004
rect 116824 111934 116830 111998
rect 116894 111934 117036 111998
rect 116824 111862 117036 111934
rect 134640 111928 135668 112004
rect 116824 111798 116966 111862
rect 117030 111798 117036 111862
rect 116824 111792 117036 111798
rect 116144 111732 116220 111792
rect 116144 111656 116492 111732
rect 28424 111596 28500 111656
rect 110160 111596 110236 111656
rect 116416 111596 116492 111656
rect 21760 111590 21972 111596
rect 21760 111526 21902 111590
rect 21966 111526 21972 111590
rect 21760 111454 21972 111526
rect 21760 111390 21766 111454
rect 21830 111390 21972 111454
rect 21760 111384 21972 111390
rect 22168 111590 22380 111596
rect 22168 111526 22174 111590
rect 22238 111526 22380 111590
rect 22168 111384 22380 111526
rect 22576 111590 22788 111596
rect 22576 111526 22718 111590
rect 22782 111526 22788 111590
rect 22576 111454 22788 111526
rect 22576 111390 22582 111454
rect 22646 111390 22788 111454
rect 22576 111384 22788 111390
rect 22984 111590 23196 111596
rect 22984 111526 22990 111590
rect 23054 111526 23196 111590
rect 22984 111454 23196 111526
rect 22984 111390 23126 111454
rect 23190 111390 23196 111454
rect 22984 111384 23196 111390
rect 23392 111590 23604 111596
rect 23392 111526 23398 111590
rect 23462 111526 23604 111590
rect 23392 111454 23604 111526
rect 23392 111390 23534 111454
rect 23598 111390 23604 111454
rect 23392 111384 23604 111390
rect 28288 111384 28636 111596
rect 110160 111384 110508 111596
rect 115192 111590 115404 111596
rect 115192 111526 115334 111590
rect 115398 111526 115404 111590
rect 115192 111454 115404 111526
rect 115192 111390 115334 111454
rect 115398 111390 115404 111454
rect 115192 111384 115404 111390
rect 115600 111590 115812 111596
rect 115600 111526 115606 111590
rect 115670 111526 115812 111590
rect 115600 111454 115812 111526
rect 115600 111390 115742 111454
rect 115806 111390 115812 111454
rect 115600 111384 115812 111390
rect 116008 111590 116220 111596
rect 116008 111526 116014 111590
rect 116078 111526 116220 111590
rect 116008 111384 116220 111526
rect 116416 111454 116628 111596
rect 116416 111390 116422 111454
rect 116486 111390 116628 111454
rect 116416 111384 116628 111390
rect 116824 111590 117036 111596
rect 116824 111526 116966 111590
rect 117030 111526 117036 111590
rect 116824 111454 117036 111526
rect 116824 111390 116830 111454
rect 116894 111390 117036 111454
rect 116824 111384 117036 111390
rect 28424 111324 28500 111384
rect 110432 111324 110508 111384
rect 1224 111318 1980 111324
rect 1224 111254 1230 111318
rect 1294 111288 1980 111318
rect 1294 111254 1798 111288
rect 1224 111248 1798 111254
rect 1768 111232 1798 111248
rect 1854 111232 1980 111288
rect 1768 111112 1980 111232
rect 21760 111182 21972 111188
rect 21760 111118 21766 111182
rect 21830 111118 21972 111182
rect 21760 110976 21972 111118
rect 22168 111182 22788 111188
rect 22168 111118 22582 111182
rect 22646 111118 22788 111182
rect 22168 111112 22788 111118
rect 22168 111052 22380 111112
rect 22168 111046 22516 111052
rect 22168 110982 22310 111046
rect 22374 110982 22446 111046
rect 22510 110982 22516 111046
rect 22168 110976 22516 110982
rect 22576 110976 22788 111112
rect 22984 111182 23196 111188
rect 22984 111118 23126 111182
rect 23190 111118 23196 111182
rect 22984 111046 23196 111118
rect 22984 110982 23126 111046
rect 23190 110982 23196 111046
rect 22984 110976 23196 110982
rect 23392 111182 23604 111188
rect 23392 111118 23534 111182
rect 23598 111118 23604 111182
rect 23392 111046 23604 111118
rect 23392 110982 23398 111046
rect 23462 110982 23604 111046
rect 23392 110976 23604 110982
rect 28288 111112 28636 111324
rect 110160 111112 110508 111324
rect 136816 111318 137572 111324
rect 136816 111288 137502 111318
rect 136816 111232 136944 111288
rect 137000 111254 137502 111288
rect 137566 111254 137572 111318
rect 137000 111248 137572 111254
rect 137000 111232 137028 111248
rect 28288 111052 28364 111112
rect 110432 111052 110508 111112
rect 21896 110916 21972 110976
rect 21760 110568 21972 110916
rect 28288 110910 28636 111052
rect 28288 110846 28294 110910
rect 28358 110846 28636 110910
rect 28288 110840 28636 110846
rect 110160 110840 110508 111052
rect 115192 111182 115404 111188
rect 115192 111118 115334 111182
rect 115398 111118 115404 111182
rect 115192 111046 115404 111118
rect 115192 110982 115198 111046
rect 115262 110982 115404 111046
rect 115192 110976 115404 110982
rect 115600 111182 115812 111188
rect 115600 111118 115742 111182
rect 115806 111118 115812 111182
rect 115600 111046 115812 111118
rect 115600 110982 115606 111046
rect 115670 110982 115812 111046
rect 115600 110976 115812 110982
rect 116008 111182 116628 111188
rect 116008 111118 116422 111182
rect 116486 111118 116628 111182
rect 116008 111112 116628 111118
rect 116008 110976 116220 111112
rect 116416 111046 116628 111112
rect 116416 110982 116558 111046
rect 116622 110982 116628 111046
rect 116416 110976 116628 110982
rect 116824 111182 117036 111188
rect 116824 111118 116830 111182
rect 116894 111118 117036 111182
rect 116824 110976 117036 111118
rect 136816 111112 137028 111232
rect 116824 110916 116900 110976
rect 28424 110780 28500 110840
rect 110296 110780 110372 110840
rect 22168 110774 22380 110780
rect 22478 110774 22788 110780
rect 22168 110710 22310 110774
rect 22374 110710 22380 110774
rect 22440 110710 22446 110774
rect 22510 110710 22788 110774
rect 22168 110644 22380 110710
rect 22478 110704 22788 110710
rect 22168 110568 22516 110644
rect 22576 110568 22788 110704
rect 22984 110774 23196 110780
rect 22984 110710 23126 110774
rect 23190 110710 23196 110774
rect 22984 110638 23196 110710
rect 22984 110574 23126 110638
rect 23190 110574 23196 110638
rect 22984 110568 23196 110574
rect 23392 110774 23604 110780
rect 23392 110710 23398 110774
rect 23462 110710 23604 110774
rect 23392 110638 23604 110710
rect 23392 110574 23398 110638
rect 23462 110574 23604 110638
rect 23392 110568 23604 110574
rect 28288 110638 28636 110780
rect 28288 110574 28294 110638
rect 28358 110574 28636 110638
rect 28288 110568 28636 110574
rect 110160 110568 110508 110780
rect 115192 110774 115404 110780
rect 115192 110710 115198 110774
rect 115262 110710 115404 110774
rect 115192 110638 115404 110710
rect 115192 110574 115198 110638
rect 115262 110574 115404 110638
rect 115192 110568 115404 110574
rect 115600 110774 115812 110780
rect 115600 110710 115606 110774
rect 115670 110710 115812 110774
rect 115600 110638 115812 110710
rect 115600 110574 115742 110638
rect 115806 110574 115812 110638
rect 115600 110568 115812 110574
rect 116008 110644 116220 110780
rect 116416 110774 116628 110780
rect 116416 110710 116558 110774
rect 116622 110710 116628 110774
rect 116008 110568 116356 110644
rect 21760 110508 21836 110568
rect 22304 110508 22380 110568
rect 21760 110160 21972 110508
rect 22168 110160 22380 110508
rect 22440 110508 22516 110568
rect 22440 110432 22788 110508
rect 22576 110236 22788 110432
rect 28406 110372 28504 110568
rect 110294 110372 110392 110568
rect 116144 110508 116220 110568
rect 22478 110230 22788 110236
rect 22440 110166 22446 110230
rect 22510 110166 22788 110230
rect 22478 110160 22788 110166
rect 22984 110366 23196 110372
rect 22984 110302 23126 110366
rect 23190 110302 23196 110366
rect 22984 110230 23196 110302
rect 22984 110166 22990 110230
rect 23054 110166 23196 110230
rect 22984 110160 23196 110166
rect 23392 110366 23604 110372
rect 23392 110302 23398 110366
rect 23462 110302 23604 110366
rect 23392 110230 23604 110302
rect 23392 110166 23534 110230
rect 23598 110166 23604 110230
rect 23392 110160 23604 110166
rect 28288 110296 28636 110372
rect 110160 110296 110508 110372
rect 115192 110366 115404 110372
rect 115192 110302 115198 110366
rect 115262 110302 115404 110366
rect 28288 110236 28364 110296
rect 110160 110236 110236 110296
rect 21896 110100 21972 110160
rect 21760 109958 21972 110100
rect 28288 110094 28636 110236
rect 28288 110030 28566 110094
rect 28630 110030 28636 110094
rect 28288 110024 28636 110030
rect 110160 110094 110508 110236
rect 115192 110230 115404 110302
rect 115192 110166 115198 110230
rect 115262 110166 115404 110230
rect 115192 110160 115404 110166
rect 115600 110366 115812 110372
rect 115600 110302 115742 110366
rect 115806 110302 115812 110366
rect 115600 110230 115812 110302
rect 115600 110166 115742 110230
rect 115806 110166 115812 110230
rect 115600 110160 115812 110166
rect 116008 110230 116220 110508
rect 116280 110508 116356 110568
rect 116416 110568 116628 110710
rect 116824 110568 117036 110916
rect 116416 110508 116492 110568
rect 116960 110508 117036 110568
rect 116280 110432 116628 110508
rect 116008 110166 116014 110230
rect 116078 110166 116220 110230
rect 116008 110160 116220 110166
rect 116416 110160 116628 110432
rect 116824 110160 117036 110508
rect 110160 110030 110166 110094
rect 110230 110030 110508 110094
rect 110160 110024 110508 110030
rect 116824 110100 116900 110160
rect 28424 109964 28500 110024
rect 110296 109964 110372 110024
rect 21760 109894 21902 109958
rect 21966 109894 21972 109958
rect 21760 109888 21972 109894
rect 22168 109958 22516 109964
rect 22168 109894 22446 109958
rect 22510 109894 22516 109958
rect 22168 109888 22516 109894
rect 22168 109828 22380 109888
rect 22576 109828 22788 109964
rect 22168 109822 22788 109828
rect 22168 109758 22310 109822
rect 22374 109758 22788 109822
rect 22168 109752 22788 109758
rect 22984 109958 23196 109964
rect 22984 109894 22990 109958
rect 23054 109894 23196 109958
rect 22984 109752 23196 109894
rect 23392 109958 23604 109964
rect 23392 109894 23534 109958
rect 23598 109894 23604 109958
rect 23392 109752 23604 109894
rect 28288 109822 28636 109964
rect 28288 109758 28566 109822
rect 28630 109758 28636 109822
rect 22304 109692 22380 109752
rect 22984 109692 23060 109752
rect 23392 109692 23468 109752
rect 1224 109686 1980 109692
rect 1224 109622 1230 109686
rect 1294 109622 1980 109686
rect 1224 109616 1980 109622
rect 1768 109608 1980 109616
rect 1768 109552 1798 109608
rect 1854 109552 1980 109608
rect 1768 109480 1980 109552
rect 21760 109686 21972 109692
rect 21760 109622 21902 109686
rect 21966 109622 21972 109686
rect 21760 109550 21972 109622
rect 21760 109486 21766 109550
rect 21830 109486 21972 109550
rect 21760 109480 21972 109486
rect 22168 109556 22380 109692
rect 22478 109686 22788 109692
rect 22440 109622 22446 109686
rect 22510 109622 22788 109686
rect 22478 109616 22788 109622
rect 22168 109550 22516 109556
rect 22168 109486 22446 109550
rect 22510 109486 22516 109550
rect 22168 109480 22516 109486
rect 22576 109480 22788 109616
rect 22984 109344 23196 109692
rect 23392 109344 23604 109692
rect 28288 109686 28636 109758
rect 28288 109622 28294 109686
rect 28358 109622 28636 109686
rect 28288 109616 28636 109622
rect 110160 109822 110508 109964
rect 110160 109758 110166 109822
rect 110230 109758 110508 109822
rect 110160 109686 110508 109758
rect 110160 109622 110166 109686
rect 110230 109622 110302 109686
rect 110366 109622 110508 109686
rect 110160 109616 110508 109622
rect 115192 109958 115404 109964
rect 115192 109894 115198 109958
rect 115262 109894 115404 109958
rect 115192 109752 115404 109894
rect 115600 109958 115812 109964
rect 115600 109894 115742 109958
rect 115806 109894 115812 109958
rect 115600 109752 115812 109894
rect 116008 109958 116220 109964
rect 116008 109894 116014 109958
rect 116078 109894 116220 109958
rect 116008 109752 116220 109894
rect 116416 109828 116628 109964
rect 116824 109958 117036 110100
rect 116824 109894 116966 109958
rect 117030 109894 117036 109958
rect 116824 109888 117036 109894
rect 115192 109692 115268 109752
rect 115600 109692 115676 109752
rect 116144 109692 116220 109752
rect 116280 109752 116628 109828
rect 116280 109692 116356 109752
rect 116552 109692 116628 109752
rect 23120 109284 23196 109344
rect 23528 109284 23604 109344
rect 21760 109278 21972 109284
rect 21760 109214 21766 109278
rect 21830 109214 21972 109278
rect 21760 109142 21972 109214
rect 21760 109078 21902 109142
rect 21966 109078 21972 109142
rect 21760 109072 21972 109078
rect 22168 108936 22380 109284
rect 22478 109278 22788 109284
rect 22440 109214 22446 109278
rect 22510 109214 22788 109278
rect 22478 109208 22788 109214
rect 22576 108936 22788 109208
rect 22984 108936 23196 109284
rect 23392 108936 23604 109284
rect 22304 108876 22380 108936
rect 22712 108876 22788 108936
rect 23120 108876 23196 108936
rect 23528 108876 23604 108936
rect 21760 108870 21972 108876
rect 21760 108806 21902 108870
rect 21966 108806 21972 108870
rect 21760 108734 21972 108806
rect 21760 108670 21902 108734
rect 21966 108670 21972 108734
rect 21760 108664 21972 108670
rect 22168 108740 22380 108876
rect 22576 108740 22788 108876
rect 22168 108734 22788 108740
rect 22168 108670 22310 108734
rect 22374 108670 22788 108734
rect 22168 108664 22788 108670
rect 22984 108734 23196 108876
rect 22984 108670 23126 108734
rect 23190 108670 23196 108734
rect 22984 108664 23196 108670
rect 23392 108734 23604 108876
rect 28288 109414 28636 109420
rect 28288 109350 28294 109414
rect 28358 109350 28636 109414
rect 28288 109278 28636 109350
rect 28288 109214 28294 109278
rect 28358 109214 28636 109278
rect 28288 109006 28636 109214
rect 28288 108942 28294 109006
rect 28358 108942 28636 109006
rect 28288 108870 28636 108942
rect 28288 108806 28430 108870
rect 28494 108806 28636 108870
rect 28288 108800 28636 108806
rect 110160 109414 110508 109420
rect 110160 109350 110166 109414
rect 110230 109350 110508 109414
rect 110160 109278 110508 109350
rect 115192 109344 115404 109692
rect 115328 109284 115404 109344
rect 110160 109214 110302 109278
rect 110366 109214 110438 109278
rect 110502 109214 110508 109278
rect 110160 109006 110508 109214
rect 110160 108942 110438 109006
rect 110502 108942 110508 109006
rect 110160 108800 110508 108942
rect 115192 108936 115404 109284
rect 115328 108876 115404 108936
rect 110160 108740 110236 108800
rect 23392 108670 23398 108734
rect 23462 108670 23604 108734
rect 23392 108664 23604 108670
rect 22304 108604 22380 108664
rect 22304 108528 22652 108604
rect 22576 108468 22652 108528
rect 21760 108462 21972 108468
rect 21760 108398 21902 108462
rect 21966 108398 21972 108462
rect 21760 108326 21972 108398
rect 21760 108262 21766 108326
rect 21830 108262 21972 108326
rect 21760 108256 21972 108262
rect 22168 108462 22380 108468
rect 22168 108398 22310 108462
rect 22374 108398 22380 108462
rect 22168 108326 22380 108398
rect 22168 108262 22174 108326
rect 22238 108262 22380 108326
rect 22168 108256 22380 108262
rect 22576 108256 22788 108468
rect 22984 108462 23196 108468
rect 22984 108398 23126 108462
rect 23190 108398 23196 108462
rect 22984 108326 23196 108398
rect 22984 108262 22990 108326
rect 23054 108262 23196 108326
rect 22984 108256 23196 108262
rect 23392 108462 23604 108468
rect 23392 108398 23398 108462
rect 23462 108398 23604 108462
rect 23392 108326 23604 108398
rect 23392 108262 23534 108326
rect 23598 108262 23604 108326
rect 23392 108256 23604 108262
rect 28288 108462 28636 108740
rect 28288 108398 28430 108462
rect 28494 108398 28566 108462
rect 28630 108398 28636 108462
rect 28288 108256 28636 108398
rect 110160 108256 110508 108740
rect 115192 108734 115404 108876
rect 115192 108670 115198 108734
rect 115262 108670 115404 108734
rect 115192 108664 115404 108670
rect 115600 109344 115812 109692
rect 116008 109616 116356 109692
rect 116008 109556 116220 109616
rect 116008 109550 116356 109556
rect 116008 109486 116150 109550
rect 116214 109486 116286 109550
rect 116350 109486 116356 109550
rect 116008 109480 116356 109486
rect 116416 109480 116628 109692
rect 116824 109686 117036 109692
rect 116824 109622 116966 109686
rect 117030 109622 117036 109686
rect 116824 109550 117036 109622
rect 116824 109486 116966 109550
rect 117030 109486 117036 109550
rect 116824 109480 117036 109486
rect 136816 109686 137572 109692
rect 136816 109622 137502 109686
rect 137566 109622 137572 109686
rect 136816 109616 137572 109622
rect 136816 109608 137028 109616
rect 136816 109552 136944 109608
rect 137000 109552 137028 109608
rect 136816 109480 137028 109552
rect 115600 109284 115676 109344
rect 115600 108936 115812 109284
rect 116008 109278 116220 109284
rect 116318 109278 116628 109284
rect 116008 109214 116150 109278
rect 116214 109214 116220 109278
rect 116280 109214 116286 109278
rect 116350 109214 116628 109278
rect 116008 108936 116220 109214
rect 116318 109208 116628 109214
rect 116416 108936 116628 109208
rect 116824 109278 117036 109284
rect 116824 109214 116966 109278
rect 117030 109214 117036 109278
rect 116824 109142 117036 109214
rect 116824 109078 116966 109142
rect 117030 109078 117036 109142
rect 116824 109072 117036 109078
rect 115600 108876 115676 108936
rect 116008 108876 116084 108936
rect 116552 108876 116628 108936
rect 115600 108734 115812 108876
rect 115600 108670 115606 108734
rect 115670 108670 115812 108734
rect 115600 108664 115812 108670
rect 116008 108734 116220 108876
rect 116008 108670 116014 108734
rect 116078 108670 116220 108734
rect 116008 108664 116220 108670
rect 116416 108664 116628 108876
rect 116824 108870 117036 108876
rect 116824 108806 116966 108870
rect 117030 108806 117036 108870
rect 116824 108734 117036 108806
rect 116824 108670 116966 108734
rect 117030 108670 117036 108734
rect 116824 108664 117036 108670
rect 115192 108462 115404 108468
rect 115192 108398 115198 108462
rect 115262 108398 115404 108462
rect 115192 108326 115404 108398
rect 115192 108262 115334 108326
rect 115398 108262 115404 108326
rect 115192 108256 115404 108262
rect 115600 108462 115812 108468
rect 115600 108398 115606 108462
rect 115670 108398 115812 108462
rect 115600 108326 115812 108398
rect 115600 108262 115742 108326
rect 115806 108262 115812 108326
rect 115600 108256 115812 108262
rect 116008 108462 116628 108468
rect 116008 108398 116014 108462
rect 116078 108398 116628 108462
rect 116008 108392 116628 108398
rect 116008 108332 116220 108392
rect 116008 108326 116356 108332
rect 116008 108262 116286 108326
rect 116350 108262 116356 108326
rect 116008 108256 116356 108262
rect 116416 108256 116628 108392
rect 116824 108462 117036 108468
rect 116824 108398 116966 108462
rect 117030 108398 117036 108462
rect 116824 108326 117036 108398
rect 116824 108262 116830 108326
rect 116894 108262 117036 108326
rect 116824 108256 117036 108262
rect 28560 108196 28636 108256
rect 110296 108196 110372 108256
rect 28288 108190 28636 108196
rect 28288 108126 28566 108190
rect 28630 108126 28636 108190
rect 1224 108054 1980 108060
rect 1224 107990 1230 108054
rect 1294 107990 1980 108054
rect 1224 107984 1980 107990
rect 1768 107928 1980 107984
rect 1768 107872 1798 107928
rect 1854 107872 1980 107928
rect 1768 107848 1980 107872
rect 21760 108054 21972 108060
rect 21760 107990 21766 108054
rect 21830 107990 21972 108054
rect 21760 107918 21972 107990
rect 21760 107854 21902 107918
rect 21966 107854 21972 107918
rect 21760 107848 21972 107854
rect 22168 108054 22380 108060
rect 22168 107990 22174 108054
rect 22238 107990 22380 108054
rect 22168 107918 22380 107990
rect 22168 107854 22310 107918
rect 22374 107854 22380 107918
rect 22168 107848 22380 107854
rect 22576 107918 22788 108060
rect 22576 107854 22582 107918
rect 22646 107854 22788 107918
rect 22576 107848 22788 107854
rect 22984 108054 23196 108060
rect 22984 107990 22990 108054
rect 23054 107990 23196 108054
rect 22984 107918 23196 107990
rect 22984 107854 23126 107918
rect 23190 107854 23196 107918
rect 22984 107848 23196 107854
rect 23392 108054 23604 108060
rect 23392 107990 23534 108054
rect 23598 107990 23604 108054
rect 23392 107918 23604 107990
rect 28288 107984 28636 108126
rect 110160 107984 110508 108196
rect 28424 107924 28500 107984
rect 110432 107924 110508 107984
rect 23392 107854 23398 107918
rect 23462 107854 23604 107918
rect 23392 107848 23604 107854
rect 28288 107712 28636 107924
rect 28560 107652 28636 107712
rect 21760 107646 21972 107652
rect 21760 107582 21902 107646
rect 21966 107582 21972 107646
rect 21760 107510 21972 107582
rect 21760 107446 21902 107510
rect 21966 107446 21972 107510
rect 21760 107440 21972 107446
rect 22168 107646 22788 107652
rect 22168 107582 22310 107646
rect 22374 107582 22582 107646
rect 22646 107582 22788 107646
rect 22168 107576 22788 107582
rect 22168 107440 22380 107576
rect 22576 107516 22788 107576
rect 22478 107510 22788 107516
rect 22440 107446 22446 107510
rect 22510 107446 22582 107510
rect 22646 107446 22788 107510
rect 22478 107440 22788 107446
rect 22984 107646 23196 107652
rect 22984 107582 23126 107646
rect 23190 107582 23196 107646
rect 22984 107510 23196 107582
rect 22984 107446 22990 107510
rect 23054 107446 23196 107510
rect 22984 107440 23196 107446
rect 23392 107646 23604 107652
rect 23392 107582 23398 107646
rect 23462 107582 23604 107646
rect 23392 107510 23604 107582
rect 23392 107446 23534 107510
rect 23598 107446 23604 107510
rect 23392 107440 23604 107446
rect 28288 107440 28636 107652
rect 110160 107712 110508 107924
rect 115192 108054 115404 108060
rect 115192 107990 115334 108054
rect 115398 107990 115404 108054
rect 115192 107918 115404 107990
rect 115192 107854 115198 107918
rect 115262 107854 115404 107918
rect 115192 107848 115404 107854
rect 115600 108054 115812 108060
rect 115600 107990 115742 108054
rect 115806 107990 115812 108054
rect 115600 107918 115812 107990
rect 115600 107854 115606 107918
rect 115670 107854 115812 107918
rect 115600 107848 115812 107854
rect 116008 107924 116220 108060
rect 116318 108054 116628 108060
rect 116280 107990 116286 108054
rect 116350 107990 116628 108054
rect 116318 107984 116628 107990
rect 116416 107924 116628 107984
rect 116008 107918 116628 107924
rect 116008 107854 116150 107918
rect 116214 107854 116422 107918
rect 116486 107854 116628 107918
rect 116008 107848 116628 107854
rect 116824 108054 117036 108060
rect 116824 107990 116830 108054
rect 116894 107990 117036 108054
rect 116824 107918 117036 107990
rect 116824 107854 116966 107918
rect 117030 107854 117036 107918
rect 116824 107848 117036 107854
rect 136816 108054 137572 108060
rect 136816 107990 137502 108054
rect 137566 107990 137572 108054
rect 136816 107984 137572 107990
rect 136816 107928 137028 107984
rect 136816 107872 136944 107928
rect 137000 107872 137028 107928
rect 136816 107848 137028 107872
rect 110160 107652 110236 107712
rect 110160 107440 110508 107652
rect 115192 107646 115404 107652
rect 115192 107582 115198 107646
rect 115262 107582 115404 107646
rect 115192 107510 115404 107582
rect 115192 107446 115198 107510
rect 115262 107446 115404 107510
rect 115192 107440 115404 107446
rect 115600 107646 115812 107652
rect 115600 107582 115606 107646
rect 115670 107582 115812 107646
rect 115600 107510 115812 107582
rect 115600 107446 115606 107510
rect 115670 107446 115812 107510
rect 115600 107440 115812 107446
rect 116008 107646 116220 107652
rect 116008 107582 116150 107646
rect 116214 107582 116220 107646
rect 116008 107510 116220 107582
rect 116008 107446 116014 107510
rect 116078 107446 116220 107510
rect 116008 107440 116220 107446
rect 116416 107646 116628 107652
rect 116416 107582 116422 107646
rect 116486 107582 116628 107646
rect 116416 107440 116628 107582
rect 116824 107646 117036 107652
rect 116824 107582 116966 107646
rect 117030 107582 117036 107646
rect 116824 107510 117036 107582
rect 116824 107446 116966 107510
rect 117030 107446 117036 107510
rect 116824 107440 117036 107446
rect 28424 107380 28500 107440
rect 110432 107380 110508 107440
rect 21760 107238 21972 107244
rect 21760 107174 21902 107238
rect 21966 107174 21972 107238
rect 21760 107032 21972 107174
rect 22168 107238 22516 107244
rect 22168 107174 22446 107238
rect 22510 107174 22516 107238
rect 22168 107168 22516 107174
rect 22576 107238 22788 107244
rect 22576 107174 22582 107238
rect 22646 107174 22788 107238
rect 22168 107102 22380 107168
rect 22168 107038 22174 107102
rect 22238 107038 22380 107102
rect 22168 107032 22380 107038
rect 22576 107102 22788 107174
rect 22576 107038 22582 107102
rect 22646 107038 22788 107102
rect 22576 107032 22788 107038
rect 22984 107238 23196 107244
rect 22984 107174 22990 107238
rect 23054 107174 23196 107238
rect 22984 107102 23196 107174
rect 22984 107038 23126 107102
rect 23190 107038 23196 107102
rect 22984 107032 23196 107038
rect 23392 107238 23604 107244
rect 23392 107174 23534 107238
rect 23598 107174 23604 107238
rect 23392 107102 23604 107174
rect 28288 107168 28636 107380
rect 110160 107168 110508 107380
rect 28424 107108 28500 107168
rect 110432 107108 110508 107168
rect 23392 107038 23534 107102
rect 23598 107038 23604 107102
rect 23392 107032 23604 107038
rect 21896 106972 21972 107032
rect 21760 106694 21972 106972
rect 28288 106896 28636 107108
rect 110160 106896 110508 107108
rect 115192 107238 115404 107244
rect 115192 107174 115198 107238
rect 115262 107174 115404 107238
rect 115192 107102 115404 107174
rect 115192 107038 115198 107102
rect 115262 107038 115404 107102
rect 115192 107032 115404 107038
rect 115600 107238 115812 107244
rect 115600 107174 115606 107238
rect 115670 107174 115812 107238
rect 115600 107102 115812 107174
rect 115600 107038 115742 107102
rect 115806 107038 115812 107102
rect 115600 107032 115812 107038
rect 116008 107238 116220 107244
rect 116008 107174 116014 107238
rect 116078 107174 116220 107238
rect 116008 107102 116220 107174
rect 116008 107038 116014 107102
rect 116078 107038 116220 107102
rect 116008 107032 116220 107038
rect 116416 107032 116628 107244
rect 116824 107238 117036 107244
rect 116824 107174 116966 107238
rect 117030 107174 117036 107238
rect 116824 107032 117036 107174
rect 116416 106972 116492 107032
rect 116144 106896 116492 106972
rect 116824 106972 116900 107032
rect 28288 106836 28364 106896
rect 110296 106836 110372 106896
rect 116144 106836 116220 106896
rect 21760 106630 21902 106694
rect 21966 106630 21972 106694
rect 21760 106624 21972 106630
rect 22168 106830 22380 106836
rect 22168 106766 22174 106830
rect 22238 106766 22380 106830
rect 22168 106624 22380 106766
rect 22576 106830 22788 106836
rect 22576 106766 22582 106830
rect 22646 106766 22788 106830
rect 22576 106694 22788 106766
rect 22576 106630 22718 106694
rect 22782 106630 22788 106694
rect 22576 106624 22788 106630
rect 22984 106830 23196 106836
rect 22984 106766 23126 106830
rect 23190 106766 23196 106830
rect 22984 106694 23196 106766
rect 22984 106630 23126 106694
rect 23190 106630 23196 106694
rect 22984 106624 23196 106630
rect 23392 106830 23604 106836
rect 23392 106766 23534 106830
rect 23598 106766 23604 106830
rect 23392 106694 23604 106766
rect 23392 106630 23398 106694
rect 23462 106630 23604 106694
rect 23392 106624 23604 106630
rect 28288 106624 28636 106836
rect 110160 106624 110508 106836
rect 115192 106830 115404 106836
rect 115192 106766 115198 106830
rect 115262 106766 115404 106830
rect 115192 106694 115404 106766
rect 115192 106630 115198 106694
rect 115262 106630 115404 106694
rect 115192 106624 115404 106630
rect 115600 106830 115812 106836
rect 115600 106766 115742 106830
rect 115806 106766 115812 106830
rect 115600 106694 115812 106766
rect 115600 106630 115606 106694
rect 115670 106630 115812 106694
rect 115600 106624 115812 106630
rect 116008 106830 116628 106836
rect 116008 106766 116014 106830
rect 116078 106766 116628 106830
rect 116008 106760 116628 106766
rect 116008 106624 116220 106760
rect 116416 106694 116628 106760
rect 116416 106630 116558 106694
rect 116622 106630 116628 106694
rect 116416 106624 116628 106630
rect 116824 106694 117036 106972
rect 116824 106630 116966 106694
rect 117030 106630 117036 106694
rect 116824 106624 117036 106630
rect 28288 106564 28364 106624
rect 110432 106564 110508 106624
rect 21760 106422 21972 106428
rect 21760 106358 21902 106422
rect 21966 106358 21972 106422
rect 1768 106248 1980 106292
rect 1768 106192 1798 106248
rect 1854 106192 1980 106248
rect 21760 106216 21972 106358
rect 22168 106422 22788 106428
rect 22168 106358 22718 106422
rect 22782 106358 22788 106422
rect 22168 106352 22788 106358
rect 22168 106292 22380 106352
rect 22168 106286 22516 106292
rect 22168 106222 22446 106286
rect 22510 106222 22516 106286
rect 22168 106216 22516 106222
rect 22576 106216 22788 106352
rect 22984 106422 23196 106428
rect 22984 106358 23126 106422
rect 23190 106358 23196 106422
rect 22984 106286 23196 106358
rect 22984 106222 23126 106286
rect 23190 106222 23196 106286
rect 22984 106216 23196 106222
rect 23392 106422 23604 106428
rect 23392 106358 23398 106422
rect 23462 106358 23604 106422
rect 23392 106286 23604 106358
rect 28288 106352 28636 106564
rect 110160 106352 110508 106564
rect 28424 106292 28500 106352
rect 110432 106292 110508 106352
rect 23392 106222 23534 106286
rect 23598 106222 23604 106286
rect 23392 106216 23604 106222
rect 1768 106156 1980 106192
rect 21896 106156 21972 106216
rect 1224 106150 1980 106156
rect 1224 106086 1230 106150
rect 1294 106086 1980 106150
rect 1224 106080 1980 106086
rect 21760 106014 21972 106156
rect 28288 106080 28636 106292
rect 110160 106150 110508 106292
rect 115192 106422 115404 106428
rect 115192 106358 115198 106422
rect 115262 106358 115404 106422
rect 115192 106286 115404 106358
rect 115192 106222 115334 106286
rect 115398 106222 115404 106286
rect 115192 106216 115404 106222
rect 115600 106422 115812 106428
rect 115600 106358 115606 106422
rect 115670 106358 115812 106422
rect 115600 106286 115812 106358
rect 115600 106222 115742 106286
rect 115806 106222 115812 106286
rect 115600 106216 115812 106222
rect 116008 106292 116220 106428
rect 116416 106422 116628 106428
rect 116416 106358 116558 106422
rect 116622 106358 116628 106422
rect 116416 106292 116628 106358
rect 116008 106216 116628 106292
rect 116824 106422 117036 106428
rect 116824 106358 116966 106422
rect 117030 106358 117036 106422
rect 116824 106216 117036 106358
rect 136816 106286 137572 106292
rect 136816 106248 137502 106286
rect 110160 106086 110302 106150
rect 110366 106086 110508 106150
rect 110160 106080 110508 106086
rect 116144 106156 116220 106216
rect 116824 106156 116900 106216
rect 136816 106192 136944 106248
rect 137000 106222 137502 106248
rect 137566 106222 137572 106286
rect 137000 106216 137572 106222
rect 137000 106192 137028 106216
rect 116144 106080 116492 106156
rect 28288 106020 28364 106080
rect 110296 106020 110372 106080
rect 116416 106020 116492 106080
rect 21760 105950 21766 106014
rect 21830 105950 21972 106014
rect 21760 105944 21972 105950
rect 22168 105808 22380 106020
rect 22478 106014 22788 106020
rect 22440 105950 22446 106014
rect 22510 105950 22788 106014
rect 22478 105944 22788 105950
rect 22576 105808 22788 105944
rect 22984 106014 23196 106020
rect 22984 105950 23126 106014
rect 23190 105950 23196 106014
rect 22984 105878 23196 105950
rect 22984 105814 22990 105878
rect 23054 105814 23196 105878
rect 22984 105808 23196 105814
rect 23392 106014 23604 106020
rect 23392 105950 23534 106014
rect 23598 105950 23604 106014
rect 23392 105878 23604 105950
rect 23392 105814 23534 105878
rect 23598 105814 23604 105878
rect 23392 105808 23604 105814
rect 22168 105748 22244 105808
rect 22576 105748 22652 105808
rect 21760 105742 21972 105748
rect 21760 105678 21766 105742
rect 21830 105678 21972 105742
rect 21760 105400 21972 105678
rect 22168 105612 22380 105748
rect 22576 105612 22788 105748
rect 22168 105536 22788 105612
rect 22168 105476 22380 105536
rect 22168 105470 22516 105476
rect 22168 105406 22310 105470
rect 22374 105406 22446 105470
rect 22510 105406 22516 105470
rect 22168 105400 22516 105406
rect 22576 105400 22788 105536
rect 22984 105606 23196 105612
rect 22984 105542 22990 105606
rect 23054 105542 23196 105606
rect 22984 105400 23196 105542
rect 23392 105606 23604 105612
rect 23392 105542 23534 105606
rect 23598 105542 23604 105606
rect 23392 105400 23604 105542
rect 28288 105536 28636 106020
rect 110160 105878 110508 106020
rect 110160 105814 110302 105878
rect 110366 105814 110508 105878
rect 110160 105536 110508 105814
rect 115192 106014 115404 106020
rect 115192 105950 115334 106014
rect 115398 105950 115404 106014
rect 115192 105878 115404 105950
rect 115192 105814 115334 105878
rect 115398 105814 115404 105878
rect 115192 105808 115404 105814
rect 115600 106014 115812 106020
rect 115600 105950 115742 106014
rect 115806 105950 115812 106014
rect 115600 105878 115812 105950
rect 115600 105814 115742 105878
rect 115806 105814 115812 105878
rect 115600 105808 115812 105814
rect 116008 105808 116220 106020
rect 116416 105808 116628 106020
rect 116824 106014 117036 106156
rect 136816 106080 137028 106192
rect 116824 105950 116830 106014
rect 116894 105950 117036 106014
rect 116824 105944 117036 105950
rect 116144 105748 116220 105808
rect 116552 105748 116628 105808
rect 116008 105672 116628 105748
rect 28424 105476 28500 105536
rect 110432 105476 110508 105536
rect 21760 105340 21836 105400
rect 22984 105340 23060 105400
rect 23392 105340 23468 105400
rect 21760 105198 21972 105340
rect 21760 105134 21902 105198
rect 21966 105134 21972 105198
rect 21760 105128 21972 105134
rect 22168 105198 22380 105204
rect 22478 105198 22788 105204
rect 22168 105134 22310 105198
rect 22374 105134 22380 105198
rect 22440 105134 22446 105198
rect 22510 105134 22788 105198
rect 22168 104992 22380 105134
rect 22478 105128 22788 105134
rect 22576 104992 22788 105128
rect 22984 104992 23196 105340
rect 23392 104992 23604 105340
rect 22168 104932 22244 104992
rect 22576 104932 22652 104992
rect 22984 104932 23060 104992
rect 23528 104932 23604 104992
rect 21760 104926 21972 104932
rect 21760 104862 21902 104926
rect 21966 104862 21972 104926
rect 21760 104790 21972 104862
rect 21760 104726 21902 104790
rect 21966 104726 21972 104790
rect 21760 104720 21972 104726
rect 22168 104720 22380 104932
rect 22576 104790 22788 104932
rect 22576 104726 22582 104790
rect 22646 104726 22788 104790
rect 22576 104720 22788 104726
rect 22984 104790 23196 104932
rect 22984 104726 22990 104790
rect 23054 104726 23196 104790
rect 22984 104720 23196 104726
rect 23392 104790 23604 104932
rect 28288 105062 28636 105476
rect 28288 104998 28294 105062
rect 28358 104998 28636 105062
rect 28288 104926 28636 104998
rect 28288 104862 28566 104926
rect 28630 104862 28636 104926
rect 28288 104856 28636 104862
rect 110160 104856 110508 105476
rect 115192 105606 115404 105612
rect 115192 105542 115334 105606
rect 115398 105542 115404 105606
rect 115192 105400 115404 105542
rect 115600 105606 115812 105612
rect 115600 105542 115742 105606
rect 115806 105542 115812 105606
rect 115600 105400 115812 105542
rect 116008 105400 116220 105672
rect 116416 105470 116628 105672
rect 116416 105406 116422 105470
rect 116486 105406 116628 105470
rect 116416 105400 116628 105406
rect 116824 105742 117036 105748
rect 116824 105678 116830 105742
rect 116894 105678 117036 105742
rect 116824 105400 117036 105678
rect 115192 105340 115268 105400
rect 115600 105340 115676 105400
rect 116960 105340 117036 105400
rect 115192 104992 115404 105340
rect 115600 104992 115812 105340
rect 115328 104932 115404 104992
rect 115736 104932 115812 104992
rect 110296 104796 110372 104856
rect 23392 104726 23534 104790
rect 23598 104726 23604 104790
rect 23392 104720 23604 104726
rect 28288 104790 28636 104796
rect 28288 104726 28294 104790
rect 28358 104726 28636 104790
rect 1224 104654 1980 104660
rect 1224 104590 1230 104654
rect 1294 104590 1980 104654
rect 1224 104584 1980 104590
rect 1768 104568 1980 104584
rect 1768 104512 1798 104568
rect 1854 104512 1980 104568
rect 1768 104448 1980 104512
rect 21760 104518 21972 104524
rect 21760 104454 21902 104518
rect 21966 104454 21972 104518
rect 21760 104382 21972 104454
rect 21760 104318 21902 104382
rect 21966 104318 21972 104382
rect 21760 104312 21972 104318
rect 22168 104388 22380 104524
rect 22576 104518 22788 104524
rect 22576 104454 22582 104518
rect 22646 104454 22788 104518
rect 22576 104388 22788 104454
rect 22168 104312 22788 104388
rect 22984 104518 23196 104524
rect 22984 104454 22990 104518
rect 23054 104454 23196 104518
rect 22984 104382 23196 104454
rect 22984 104318 22990 104382
rect 23054 104318 23196 104382
rect 22984 104312 23196 104318
rect 23392 104518 23604 104524
rect 23392 104454 23534 104518
rect 23598 104454 23604 104518
rect 23392 104382 23604 104454
rect 23392 104318 23398 104382
rect 23462 104318 23604 104382
rect 23392 104312 23604 104318
rect 28288 104518 28636 104726
rect 28288 104454 28430 104518
rect 28494 104454 28566 104518
rect 28630 104454 28636 104518
rect 28288 104312 28636 104454
rect 110160 104312 110508 104796
rect 115192 104790 115404 104932
rect 115192 104726 115198 104790
rect 115262 104726 115404 104790
rect 115192 104720 115404 104726
rect 115600 104790 115812 104932
rect 115600 104726 115606 104790
rect 115670 104726 115812 104790
rect 115600 104720 115812 104726
rect 116008 104992 116220 105204
rect 116416 105198 116628 105204
rect 116416 105134 116422 105198
rect 116486 105134 116628 105198
rect 116416 104992 116628 105134
rect 116824 105198 117036 105340
rect 116824 105134 116966 105198
rect 117030 105134 117036 105198
rect 116824 105128 117036 105134
rect 116008 104932 116084 104992
rect 116416 104932 116492 104992
rect 116008 104856 116628 104932
rect 116008 104790 116220 104856
rect 116008 104726 116014 104790
rect 116078 104726 116220 104790
rect 116008 104720 116220 104726
rect 116416 104720 116628 104856
rect 116824 104926 117036 104932
rect 116824 104862 116966 104926
rect 117030 104862 117036 104926
rect 116824 104790 117036 104862
rect 116824 104726 116966 104790
rect 117030 104726 117036 104790
rect 116824 104720 117036 104726
rect 136816 104568 137028 104660
rect 115192 104518 115404 104524
rect 115192 104454 115198 104518
rect 115262 104454 115404 104518
rect 115192 104382 115404 104454
rect 115192 104318 115198 104382
rect 115262 104318 115404 104382
rect 115192 104312 115404 104318
rect 115600 104518 115812 104524
rect 115600 104454 115606 104518
rect 115670 104454 115812 104518
rect 115600 104382 115812 104454
rect 115600 104318 115606 104382
rect 115670 104318 115812 104382
rect 115600 104312 115812 104318
rect 116008 104518 116220 104524
rect 116008 104454 116014 104518
rect 116078 104454 116220 104518
rect 116008 104388 116220 104454
rect 116416 104388 116628 104524
rect 116008 104382 116628 104388
rect 116008 104318 116150 104382
rect 116214 104318 116628 104382
rect 116008 104312 116628 104318
rect 116824 104518 117036 104524
rect 116824 104454 116966 104518
rect 117030 104454 117036 104518
rect 116824 104382 117036 104454
rect 136816 104512 136944 104568
rect 137000 104524 137028 104568
rect 137000 104518 137572 104524
rect 137000 104512 137502 104518
rect 136816 104454 137502 104512
rect 137566 104454 137572 104518
rect 136816 104448 137572 104454
rect 116824 104318 116966 104382
rect 117030 104318 117036 104382
rect 116824 104312 117036 104318
rect 22304 104252 22380 104312
rect 28288 104252 28364 104312
rect 110432 104252 110508 104312
rect 22304 104176 22652 104252
rect 22576 104116 22652 104176
rect 28288 104246 28636 104252
rect 28288 104182 28430 104246
rect 28494 104182 28636 104246
rect 21760 104110 21972 104116
rect 21760 104046 21902 104110
rect 21966 104046 21972 104110
rect 21760 103974 21972 104046
rect 21760 103910 21766 103974
rect 21830 103910 21972 103974
rect 21760 103904 21972 103910
rect 22168 103980 22380 104116
rect 22576 103980 22788 104116
rect 22168 103974 22788 103980
rect 22168 103910 22174 103974
rect 22238 103910 22788 103974
rect 22168 103904 22788 103910
rect 22984 104110 23196 104116
rect 22984 104046 22990 104110
rect 23054 104046 23196 104110
rect 22984 103974 23196 104046
rect 22984 103910 23126 103974
rect 23190 103910 23196 103974
rect 22984 103904 23196 103910
rect 23392 104110 23604 104116
rect 23392 104046 23398 104110
rect 23462 104046 23604 104110
rect 23392 103974 23604 104046
rect 28288 104040 28636 104182
rect 110160 104040 110508 104252
rect 115192 104110 115404 104116
rect 115192 104046 115198 104110
rect 115262 104046 115404 104110
rect 28560 103980 28636 104040
rect 110296 103980 110372 104040
rect 23392 103910 23534 103974
rect 23598 103910 23604 103974
rect 23392 103904 23604 103910
rect 28288 103768 28636 103980
rect 110160 103768 110508 103980
rect 115192 103974 115404 104046
rect 115192 103910 115334 103974
rect 115398 103910 115404 103974
rect 115192 103904 115404 103910
rect 115600 104110 115812 104116
rect 115600 104046 115606 104110
rect 115670 104046 115812 104110
rect 115600 103974 115812 104046
rect 115600 103910 115742 103974
rect 115806 103910 115812 103974
rect 115600 103904 115812 103910
rect 116008 104110 116220 104116
rect 116008 104046 116150 104110
rect 116214 104046 116220 104110
rect 116008 103980 116220 104046
rect 116416 103980 116628 104116
rect 116008 103974 116628 103980
rect 116008 103910 116014 103974
rect 116078 103910 116628 103974
rect 116008 103904 116628 103910
rect 116824 104110 117036 104116
rect 116824 104046 116966 104110
rect 117030 104046 117036 104110
rect 116824 103974 117036 104046
rect 116824 103910 116830 103974
rect 116894 103910 117036 103974
rect 116824 103904 117036 103910
rect 28424 103708 28500 103768
rect 110296 103708 110372 103768
rect 21760 103702 21972 103708
rect 21760 103638 21766 103702
rect 21830 103638 21972 103702
rect 21760 103566 21972 103638
rect 21760 103502 21766 103566
rect 21830 103502 21972 103566
rect 21760 103496 21972 103502
rect 22168 103702 22380 103708
rect 22168 103638 22174 103702
rect 22238 103638 22380 103702
rect 22168 103566 22380 103638
rect 22168 103502 22310 103566
rect 22374 103502 22380 103566
rect 22168 103496 22380 103502
rect 22576 103496 22788 103708
rect 22984 103702 23196 103708
rect 22984 103638 23126 103702
rect 23190 103638 23196 103702
rect 22984 103566 23196 103638
rect 22984 103502 23126 103566
rect 23190 103502 23196 103566
rect 22984 103496 23196 103502
rect 23392 103702 23604 103708
rect 23392 103638 23534 103702
rect 23598 103638 23604 103702
rect 23392 103566 23604 103638
rect 23392 103502 23398 103566
rect 23462 103502 23604 103566
rect 23392 103496 23604 103502
rect 28288 103496 28636 103708
rect 110160 103496 110508 103708
rect 115192 103702 115404 103708
rect 115192 103638 115334 103702
rect 115398 103638 115404 103702
rect 115192 103566 115404 103638
rect 115192 103502 115334 103566
rect 115398 103502 115404 103566
rect 115192 103496 115404 103502
rect 115600 103702 115812 103708
rect 115600 103638 115742 103702
rect 115806 103638 115812 103702
rect 115600 103566 115812 103638
rect 115600 103502 115742 103566
rect 115806 103502 115812 103566
rect 115600 103496 115812 103502
rect 116008 103702 116628 103708
rect 116008 103638 116014 103702
rect 116078 103638 116628 103702
rect 116008 103632 116628 103638
rect 116008 103572 116220 103632
rect 116008 103566 116356 103572
rect 116008 103502 116286 103566
rect 116350 103502 116356 103566
rect 116008 103496 116356 103502
rect 116416 103496 116628 103632
rect 116824 103702 117036 103708
rect 116824 103638 116830 103702
rect 116894 103638 117036 103702
rect 116824 103566 117036 103638
rect 116824 103502 116830 103566
rect 116894 103502 117036 103566
rect 116824 103496 117036 103502
rect 22576 103436 22652 103496
rect 22304 103360 22652 103436
rect 28288 103436 28364 103496
rect 110160 103436 110236 103496
rect 22304 103300 22380 103360
rect 21760 103294 21972 103300
rect 21760 103230 21766 103294
rect 21830 103230 21972 103294
rect 21760 103158 21972 103230
rect 21760 103094 21902 103158
rect 21966 103094 21972 103158
rect 21760 103088 21972 103094
rect 22168 103294 22788 103300
rect 22168 103230 22310 103294
rect 22374 103230 22788 103294
rect 22168 103224 22788 103230
rect 22168 103164 22380 103224
rect 22168 103158 22516 103164
rect 22168 103094 22174 103158
rect 22238 103094 22446 103158
rect 22510 103094 22516 103158
rect 22168 103088 22516 103094
rect 22576 103088 22788 103224
rect 22984 103294 23196 103300
rect 22984 103230 23126 103294
rect 23190 103230 23196 103294
rect 22984 103158 23196 103230
rect 22984 103094 22990 103158
rect 23054 103094 23196 103158
rect 22984 103088 23196 103094
rect 23392 103294 23604 103300
rect 23392 103230 23398 103294
rect 23462 103230 23604 103294
rect 23392 103158 23604 103230
rect 28288 103224 28636 103436
rect 110160 103224 110508 103436
rect 115192 103294 115404 103300
rect 115192 103230 115334 103294
rect 115398 103230 115404 103294
rect 28424 103164 28500 103224
rect 110296 103164 110372 103224
rect 23392 103094 23398 103158
rect 23462 103094 23604 103158
rect 23392 103088 23604 103094
rect 1768 102888 1980 103028
rect 28288 102952 28636 103164
rect 110160 102952 110508 103164
rect 115192 103158 115404 103230
rect 115192 103094 115334 103158
rect 115398 103094 115404 103158
rect 115192 103088 115404 103094
rect 115600 103294 115812 103300
rect 115600 103230 115742 103294
rect 115806 103230 115812 103294
rect 115600 103158 115812 103230
rect 115600 103094 115742 103158
rect 115806 103094 115812 103158
rect 115600 103088 115812 103094
rect 116008 103164 116220 103300
rect 116318 103294 116628 103300
rect 116280 103230 116286 103294
rect 116350 103230 116628 103294
rect 116318 103224 116628 103230
rect 116416 103164 116628 103224
rect 116008 103088 116628 103164
rect 116824 103294 117036 103300
rect 116824 103230 116830 103294
rect 116894 103230 117036 103294
rect 116824 103158 117036 103230
rect 116824 103094 116966 103158
rect 117030 103094 117036 103158
rect 116824 103088 117036 103094
rect 116144 103028 116220 103088
rect 116144 102952 116492 103028
rect 28424 102892 28500 102952
rect 110432 102892 110508 102952
rect 116416 102892 116492 102952
rect 136816 102892 137028 103028
rect 1768 102832 1798 102888
rect 1854 102832 1980 102888
rect 1768 102756 1980 102832
rect 1224 102750 1980 102756
rect 1224 102686 1230 102750
rect 1294 102686 1980 102750
rect 1224 102680 1980 102686
rect 21760 102886 21972 102892
rect 21760 102822 21902 102886
rect 21966 102822 21972 102886
rect 21760 102750 21972 102822
rect 21760 102686 21766 102750
rect 21830 102686 21972 102750
rect 21760 102680 21972 102686
rect 22168 102886 22380 102892
rect 22478 102886 22788 102892
rect 22168 102822 22174 102886
rect 22238 102822 22380 102886
rect 22440 102822 22446 102886
rect 22510 102822 22788 102886
rect 22168 102680 22380 102822
rect 22478 102816 22788 102822
rect 22576 102750 22788 102816
rect 22576 102686 22582 102750
rect 22646 102686 22788 102750
rect 22576 102680 22788 102686
rect 22984 102886 23196 102892
rect 22984 102822 22990 102886
rect 23054 102822 23196 102886
rect 22984 102750 23196 102822
rect 22984 102686 23126 102750
rect 23190 102686 23196 102750
rect 22984 102680 23196 102686
rect 23392 102886 23604 102892
rect 23392 102822 23398 102886
rect 23462 102822 23604 102886
rect 23392 102750 23604 102822
rect 23392 102686 23534 102750
rect 23598 102686 23604 102750
rect 23392 102680 23604 102686
rect 28288 102680 28636 102892
rect 110160 102680 110508 102892
rect 115192 102886 115404 102892
rect 115192 102822 115334 102886
rect 115398 102822 115404 102886
rect 115192 102750 115404 102822
rect 115192 102686 115198 102750
rect 115262 102686 115404 102750
rect 115192 102680 115404 102686
rect 115600 102886 115812 102892
rect 115600 102822 115742 102886
rect 115806 102822 115812 102886
rect 115600 102750 115812 102822
rect 115600 102686 115742 102750
rect 115806 102686 115812 102750
rect 115600 102680 115812 102686
rect 116008 102750 116220 102892
rect 116008 102686 116150 102750
rect 116214 102686 116220 102750
rect 116008 102680 116220 102686
rect 116416 102750 116628 102892
rect 116416 102686 116422 102750
rect 116486 102686 116628 102750
rect 116416 102680 116628 102686
rect 116824 102886 117036 102892
rect 116824 102822 116966 102886
rect 117030 102822 117036 102886
rect 116824 102750 117036 102822
rect 116824 102686 116830 102750
rect 116894 102686 117036 102750
rect 116824 102680 117036 102686
rect 136816 102888 137572 102892
rect 136816 102832 136944 102888
rect 137000 102886 137572 102888
rect 137000 102832 137502 102886
rect 136816 102822 137502 102832
rect 137566 102822 137572 102886
rect 136816 102816 137572 102822
rect 136816 102680 137028 102816
rect 28288 102620 28364 102680
rect 110296 102620 110372 102680
rect 21760 102478 21972 102484
rect 21760 102414 21766 102478
rect 21830 102414 21972 102478
rect 21760 102272 21972 102414
rect 22168 102342 22380 102484
rect 22168 102278 22310 102342
rect 22374 102278 22380 102342
rect 22168 102272 22380 102278
rect 22576 102478 22788 102484
rect 22576 102414 22582 102478
rect 22646 102414 22788 102478
rect 22576 102342 22788 102414
rect 22576 102278 22718 102342
rect 22782 102278 22788 102342
rect 22576 102272 22788 102278
rect 22984 102478 23196 102484
rect 22984 102414 23126 102478
rect 23190 102414 23196 102478
rect 22984 102342 23196 102414
rect 22984 102278 22990 102342
rect 23054 102278 23196 102342
rect 22984 102272 23196 102278
rect 23392 102478 23604 102484
rect 23392 102414 23534 102478
rect 23598 102414 23604 102478
rect 23392 102342 23604 102414
rect 23392 102278 23398 102342
rect 23462 102278 23604 102342
rect 23392 102272 23604 102278
rect 28288 102408 28636 102620
rect 110160 102408 110508 102620
rect 115192 102478 115404 102484
rect 115192 102414 115198 102478
rect 115262 102414 115404 102478
rect 28288 102348 28364 102408
rect 110296 102348 110372 102408
rect 21896 102212 21972 102272
rect 21760 102070 21972 102212
rect 28288 102136 28636 102348
rect 110160 102136 110508 102348
rect 115192 102342 115404 102414
rect 115192 102278 115198 102342
rect 115262 102278 115404 102342
rect 115192 102272 115404 102278
rect 115600 102478 115812 102484
rect 115600 102414 115742 102478
rect 115806 102414 115812 102478
rect 115600 102342 115812 102414
rect 115600 102278 115606 102342
rect 115670 102278 115812 102342
rect 115600 102272 115812 102278
rect 116008 102478 116628 102484
rect 116008 102414 116150 102478
rect 116214 102414 116422 102478
rect 116486 102414 116628 102478
rect 116008 102408 116628 102414
rect 116008 102272 116220 102408
rect 116416 102342 116628 102408
rect 116416 102278 116558 102342
rect 116622 102278 116628 102342
rect 116416 102272 116628 102278
rect 116824 102478 117036 102484
rect 116824 102414 116830 102478
rect 116894 102414 117036 102478
rect 116824 102272 117036 102414
rect 116960 102212 117036 102272
rect 28424 102076 28500 102136
rect 110160 102076 110236 102136
rect 21760 102006 21766 102070
rect 21830 102006 21972 102070
rect 21760 102000 21972 102006
rect 22168 102070 22516 102076
rect 22168 102006 22310 102070
rect 22374 102006 22446 102070
rect 22510 102006 22516 102070
rect 22168 102000 22516 102006
rect 22576 102070 22788 102076
rect 22576 102006 22718 102070
rect 22782 102006 22788 102070
rect 22168 101940 22380 102000
rect 22576 101940 22788 102006
rect 22168 101864 22788 101940
rect 22984 102070 23196 102076
rect 22984 102006 22990 102070
rect 23054 102006 23196 102070
rect 22984 101934 23196 102006
rect 22984 101870 23126 101934
rect 23190 101870 23196 101934
rect 22984 101864 23196 101870
rect 23392 102070 23604 102076
rect 23392 102006 23398 102070
rect 23462 102006 23604 102070
rect 23392 101934 23604 102006
rect 23392 101870 23534 101934
rect 23598 101870 23604 101934
rect 23392 101864 23604 101870
rect 22304 101804 22380 101864
rect 21760 101798 21972 101804
rect 21760 101734 21766 101798
rect 21830 101734 21972 101798
rect 21760 101456 21972 101734
rect 22168 101456 22380 101804
rect 22478 101798 22788 101804
rect 22440 101734 22446 101798
rect 22510 101734 22788 101798
rect 22478 101728 22788 101734
rect 22576 101526 22788 101728
rect 22576 101462 22718 101526
rect 22782 101462 22788 101526
rect 22576 101456 22788 101462
rect 22984 101662 23196 101668
rect 22984 101598 23126 101662
rect 23190 101598 23196 101662
rect 22984 101456 23196 101598
rect 23392 101662 23604 101668
rect 23392 101598 23534 101662
rect 23598 101598 23604 101662
rect 23392 101456 23604 101598
rect 21896 101396 21972 101456
rect 23120 101396 23196 101456
rect 23528 101396 23604 101456
rect 1224 101254 1980 101260
rect 1224 101190 1230 101254
rect 1294 101208 1980 101254
rect 1294 101190 1798 101208
rect 1224 101184 1798 101190
rect 1768 101152 1798 101184
rect 1854 101152 1980 101208
rect 21760 101254 21972 101396
rect 21760 101190 21902 101254
rect 21966 101190 21972 101254
rect 21760 101184 21972 101190
rect 1768 101048 1980 101152
rect 22168 101048 22380 101260
rect 22576 101254 22788 101260
rect 22576 101190 22718 101254
rect 22782 101190 22788 101254
rect 22576 101124 22788 101190
rect 22304 100988 22380 101048
rect 22440 101048 22788 101124
rect 22984 101048 23196 101396
rect 22440 100988 22516 101048
rect 23120 100988 23196 101048
rect 21760 100982 21972 100988
rect 21760 100918 21902 100982
rect 21966 100918 21972 100982
rect 21760 100846 21972 100918
rect 21760 100782 21766 100846
rect 21830 100782 21972 100846
rect 21760 100776 21972 100782
rect 22168 100912 22516 100988
rect 22168 100852 22380 100912
rect 22168 100846 22516 100852
rect 22168 100782 22446 100846
rect 22510 100782 22516 100846
rect 22168 100776 22516 100782
rect 22576 100776 22788 100988
rect 22304 100716 22380 100776
rect 22576 100716 22652 100776
rect 22304 100640 22652 100716
rect 22984 100640 23196 100988
rect 23392 101048 23604 101396
rect 28288 101662 28636 102076
rect 28288 101598 28294 101662
rect 28358 101598 28636 101662
rect 28288 101592 28636 101598
rect 110160 101592 110508 102076
rect 115192 102070 115404 102076
rect 115192 102006 115198 102070
rect 115262 102006 115404 102070
rect 115192 101934 115404 102006
rect 115192 101870 115198 101934
rect 115262 101870 115404 101934
rect 115192 101864 115404 101870
rect 115600 102070 115812 102076
rect 115600 102006 115606 102070
rect 115670 102006 115812 102070
rect 115600 101934 115812 102006
rect 115600 101870 115606 101934
rect 115670 101870 115812 101934
rect 115600 101864 115812 101870
rect 116008 101940 116220 102076
rect 116416 102070 116628 102076
rect 116416 102006 116558 102070
rect 116622 102006 116628 102070
rect 116416 101940 116628 102006
rect 116824 102070 117036 102212
rect 116824 102006 116966 102070
rect 117030 102006 117036 102070
rect 116824 102000 117036 102006
rect 116008 101864 116628 101940
rect 116008 101804 116084 101864
rect 116416 101804 116492 101864
rect 28288 101532 28364 101592
rect 110432 101532 110508 101592
rect 28288 101390 28636 101532
rect 28288 101326 28294 101390
rect 28358 101326 28566 101390
rect 28630 101326 28636 101390
rect 28288 101118 28636 101326
rect 28288 101054 28566 101118
rect 28630 101054 28636 101118
rect 23392 100988 23468 101048
rect 23392 100640 23604 100988
rect 28288 100982 28636 101054
rect 28288 100918 28294 100982
rect 28358 100918 28636 100982
rect 28288 100912 28636 100918
rect 110160 101390 110508 101532
rect 115192 101662 115404 101668
rect 115192 101598 115198 101662
rect 115262 101598 115404 101662
rect 115192 101456 115404 101598
rect 115600 101662 115812 101668
rect 115600 101598 115606 101662
rect 115670 101598 115812 101662
rect 115600 101456 115812 101598
rect 116008 101456 116220 101804
rect 116416 101532 116628 101804
rect 116318 101526 116628 101532
rect 116280 101462 116286 101526
rect 116350 101462 116628 101526
rect 116318 101456 116628 101462
rect 116824 101798 117036 101804
rect 116824 101734 116966 101798
rect 117030 101734 117036 101798
rect 116824 101456 117036 101734
rect 115328 101396 115404 101456
rect 115736 101396 115812 101456
rect 110160 101326 110166 101390
rect 110230 101326 110508 101390
rect 110160 101118 110508 101326
rect 110160 101054 110166 101118
rect 110230 101054 110508 101118
rect 110160 100982 110508 101054
rect 110160 100918 110302 100982
rect 110366 100918 110508 100982
rect 110160 100912 110508 100918
rect 115192 101048 115404 101396
rect 115600 101048 115812 101396
rect 116824 101396 116900 101456
rect 116008 101254 116356 101260
rect 116008 101190 116286 101254
rect 116350 101190 116356 101254
rect 116008 101184 116356 101190
rect 116008 101048 116220 101184
rect 116416 101124 116628 101260
rect 116824 101254 117036 101396
rect 116824 101190 116966 101254
rect 117030 101190 117036 101254
rect 116824 101184 117036 101190
rect 136816 101254 137572 101260
rect 136816 101208 137502 101254
rect 115192 100988 115268 101048
rect 115736 100988 115812 101048
rect 116144 100988 116220 101048
rect 116280 101048 116628 101124
rect 136816 101152 136944 101208
rect 137000 101190 137502 101208
rect 137566 101190 137572 101254
rect 137000 101184 137572 101190
rect 137000 101152 137028 101184
rect 136816 101048 137028 101152
rect 116280 100988 116356 101048
rect 22984 100580 23060 100640
rect 23528 100580 23604 100640
rect 21760 100574 21972 100580
rect 21760 100510 21766 100574
rect 21830 100510 21972 100574
rect 21760 100438 21972 100510
rect 21760 100374 21766 100438
rect 21830 100374 21972 100438
rect 21760 100368 21972 100374
rect 22168 100232 22380 100580
rect 22478 100574 22788 100580
rect 22440 100510 22446 100574
rect 22510 100510 22788 100574
rect 22478 100504 22788 100510
rect 22576 100308 22788 100504
rect 22984 100438 23196 100580
rect 22984 100374 22990 100438
rect 23054 100374 23196 100438
rect 22984 100368 23196 100374
rect 23392 100438 23604 100580
rect 23392 100374 23398 100438
rect 23462 100374 23604 100438
rect 23392 100368 23604 100374
rect 28288 100710 28636 100716
rect 28288 100646 28294 100710
rect 28358 100646 28636 100710
rect 28288 100438 28636 100646
rect 28288 100374 28430 100438
rect 28494 100374 28636 100438
rect 28288 100368 28636 100374
rect 110160 100710 110508 100716
rect 110160 100646 110302 100710
rect 110366 100646 110508 100710
rect 110160 100574 110508 100646
rect 115192 100640 115404 100988
rect 115328 100580 115404 100640
rect 110160 100510 110302 100574
rect 110366 100510 110508 100574
rect 110160 100368 110508 100510
rect 115192 100438 115404 100580
rect 115192 100374 115334 100438
rect 115398 100374 115404 100438
rect 115192 100368 115404 100374
rect 115600 100640 115812 100988
rect 116008 100912 116356 100988
rect 116008 100852 116220 100912
rect 116416 100852 116628 100988
rect 116008 100846 116628 100852
rect 116008 100782 116150 100846
rect 116214 100782 116422 100846
rect 116486 100782 116628 100846
rect 116008 100776 116628 100782
rect 116824 100982 117036 100988
rect 116824 100918 116966 100982
rect 117030 100918 117036 100982
rect 116824 100846 117036 100918
rect 116824 100782 116966 100846
rect 117030 100782 117036 100846
rect 116824 100776 117036 100782
rect 115600 100580 115676 100640
rect 115600 100438 115812 100580
rect 115600 100374 115742 100438
rect 115806 100374 115812 100438
rect 115600 100368 115812 100374
rect 116008 100574 116220 100580
rect 116008 100510 116150 100574
rect 116214 100510 116220 100574
rect 28424 100308 28500 100368
rect 110432 100308 110508 100368
rect 22304 100172 22380 100232
rect 22440 100232 22788 100308
rect 22440 100172 22516 100232
rect 21760 100166 21972 100172
rect 21760 100102 21766 100166
rect 21830 100102 21972 100166
rect 21760 100030 21972 100102
rect 21760 99966 21902 100030
rect 21966 99966 21972 100030
rect 21760 99960 21972 99966
rect 22168 100096 22516 100172
rect 22168 100036 22380 100096
rect 22576 100036 22788 100172
rect 22168 100030 22788 100036
rect 22168 99966 22174 100030
rect 22238 99966 22788 100030
rect 22168 99960 22788 99966
rect 22984 100166 23196 100172
rect 22984 100102 22990 100166
rect 23054 100102 23196 100166
rect 22984 100030 23196 100102
rect 22984 99966 22990 100030
rect 23054 99966 23196 100030
rect 22984 99960 23196 99966
rect 23392 100166 23604 100172
rect 23392 100102 23398 100166
rect 23462 100102 23604 100166
rect 23392 100030 23604 100102
rect 28288 100096 28636 100308
rect 110160 100302 110508 100308
rect 110160 100238 110302 100302
rect 110366 100238 110508 100302
rect 110160 100096 110508 100238
rect 116008 100232 116220 100510
rect 116416 100574 116628 100580
rect 116416 100510 116422 100574
rect 116486 100510 116628 100574
rect 116416 100232 116628 100510
rect 116824 100574 117036 100580
rect 116824 100510 116966 100574
rect 117030 100510 117036 100574
rect 116824 100438 117036 100510
rect 116824 100374 116966 100438
rect 117030 100374 117036 100438
rect 116824 100368 117036 100374
rect 116008 100172 116084 100232
rect 116552 100172 116628 100232
rect 110432 100036 110508 100096
rect 23392 99966 23398 100030
rect 23462 99966 23604 100030
rect 23392 99960 23604 99966
rect 28288 100030 28636 100036
rect 28288 99966 28430 100030
rect 28494 99966 28636 100030
rect 28288 99960 28636 99966
rect 110160 99960 110508 100036
rect 115192 100166 115404 100172
rect 115192 100102 115334 100166
rect 115398 100102 115404 100166
rect 115192 100030 115404 100102
rect 115192 99966 115198 100030
rect 115262 99966 115404 100030
rect 115192 99960 115404 99966
rect 115600 100166 115812 100172
rect 115600 100102 115742 100166
rect 115806 100102 115812 100166
rect 115600 100030 115812 100102
rect 115600 99966 115606 100030
rect 115670 99966 115812 100030
rect 115600 99960 115812 99966
rect 116008 100030 116220 100172
rect 116008 99966 116014 100030
rect 116078 99966 116220 100030
rect 116008 99960 116220 99966
rect 116416 99960 116628 100172
rect 116824 100166 117036 100172
rect 116824 100102 116966 100166
rect 117030 100102 117036 100166
rect 116824 100030 117036 100102
rect 116824 99966 116830 100030
rect 116894 99966 117036 100030
rect 116824 99960 117036 99966
rect 22304 99900 22380 99960
rect 22304 99824 22652 99900
rect 22576 99764 22652 99824
rect 28406 99764 28504 99960
rect 110294 99764 110392 99960
rect 21760 99758 21972 99764
rect 21760 99694 21902 99758
rect 21966 99694 21972 99758
rect 1224 99622 1980 99628
rect 1224 99558 1230 99622
rect 1294 99558 1980 99622
rect 1224 99552 1980 99558
rect 21760 99622 21972 99694
rect 21760 99558 21766 99622
rect 21830 99558 21972 99622
rect 21760 99552 21972 99558
rect 22168 99758 22380 99764
rect 22168 99694 22174 99758
rect 22238 99694 22380 99758
rect 22168 99628 22380 99694
rect 22168 99622 22516 99628
rect 22168 99558 22174 99622
rect 22238 99558 22446 99622
rect 22510 99558 22516 99622
rect 22168 99552 22516 99558
rect 22576 99552 22788 99764
rect 22984 99758 23196 99764
rect 22984 99694 22990 99758
rect 23054 99694 23196 99758
rect 22984 99622 23196 99694
rect 22984 99558 22990 99622
rect 23054 99558 23196 99622
rect 22984 99552 23196 99558
rect 23392 99758 23604 99764
rect 23392 99694 23398 99758
rect 23462 99694 23604 99758
rect 23392 99622 23604 99694
rect 23392 99558 23534 99622
rect 23598 99558 23604 99622
rect 23392 99552 23604 99558
rect 28288 99758 28636 99764
rect 28288 99694 28566 99758
rect 28630 99694 28636 99758
rect 28288 99552 28636 99694
rect 110160 99552 110508 99764
rect 115192 99758 115404 99764
rect 115192 99694 115198 99758
rect 115262 99694 115404 99758
rect 115192 99622 115404 99694
rect 115192 99558 115198 99622
rect 115262 99558 115404 99622
rect 115192 99552 115404 99558
rect 115600 99758 115812 99764
rect 115600 99694 115606 99758
rect 115670 99694 115812 99758
rect 115600 99622 115812 99694
rect 115600 99558 115742 99622
rect 115806 99558 115812 99622
rect 115600 99552 115812 99558
rect 116008 99758 116220 99764
rect 116008 99694 116014 99758
rect 116078 99694 116220 99758
rect 116008 99628 116220 99694
rect 116008 99622 116356 99628
rect 116008 99558 116286 99622
rect 116350 99558 116356 99622
rect 116008 99552 116356 99558
rect 116416 99622 116628 99764
rect 116416 99558 116422 99622
rect 116486 99558 116628 99622
rect 116416 99552 116628 99558
rect 116824 99758 117036 99764
rect 116824 99694 116830 99758
rect 116894 99694 117036 99758
rect 116824 99622 117036 99694
rect 116824 99558 116830 99622
rect 116894 99558 117036 99622
rect 116824 99552 117036 99558
rect 136816 99622 137572 99628
rect 136816 99558 137502 99622
rect 137566 99558 137572 99622
rect 136816 99552 137572 99558
rect 1768 99528 1980 99552
rect 1768 99472 1798 99528
rect 1854 99472 1980 99528
rect 1768 99416 1980 99472
rect 28288 99492 28364 99552
rect 110296 99492 110372 99552
rect 136816 99528 137028 99552
rect 28288 99486 28636 99492
rect 28288 99422 28566 99486
rect 28630 99422 28636 99486
rect 21760 99350 21972 99356
rect 21760 99286 21766 99350
rect 21830 99286 21972 99350
rect 21760 99214 21972 99286
rect 21760 99150 21902 99214
rect 21966 99150 21972 99214
rect 21760 99144 21972 99150
rect 22168 99350 22380 99356
rect 22478 99350 22788 99356
rect 22168 99286 22174 99350
rect 22238 99286 22380 99350
rect 22440 99286 22446 99350
rect 22510 99286 22788 99350
rect 22168 99144 22380 99286
rect 22478 99280 22788 99286
rect 22576 99214 22788 99280
rect 22576 99150 22582 99214
rect 22646 99150 22788 99214
rect 22576 99144 22788 99150
rect 22984 99350 23196 99356
rect 22984 99286 22990 99350
rect 23054 99286 23196 99350
rect 22984 99214 23196 99286
rect 22984 99150 22990 99214
rect 23054 99150 23196 99214
rect 22984 99144 23196 99150
rect 23392 99350 23604 99356
rect 23392 99286 23534 99350
rect 23598 99286 23604 99350
rect 23392 99214 23604 99286
rect 23392 99150 23398 99214
rect 23462 99150 23604 99214
rect 23392 99144 23604 99150
rect 28288 99280 28636 99422
rect 110160 99280 110508 99492
rect 136816 99472 136944 99528
rect 137000 99472 137028 99528
rect 136816 99416 137028 99472
rect 115192 99350 115404 99356
rect 115192 99286 115198 99350
rect 115262 99286 115404 99350
rect 28288 99220 28364 99280
rect 110296 99220 110372 99280
rect 28288 99008 28636 99220
rect 110160 99008 110508 99220
rect 115192 99214 115404 99286
rect 115192 99150 115198 99214
rect 115262 99150 115404 99214
rect 115192 99144 115404 99150
rect 115600 99350 115812 99356
rect 115600 99286 115742 99350
rect 115806 99286 115812 99350
rect 115600 99214 115812 99286
rect 115600 99150 115606 99214
rect 115670 99150 115812 99214
rect 115600 99144 115812 99150
rect 116008 99214 116220 99356
rect 116318 99350 116628 99356
rect 116280 99286 116286 99350
rect 116350 99286 116422 99350
rect 116486 99286 116628 99350
rect 116318 99280 116628 99286
rect 116008 99150 116150 99214
rect 116214 99150 116220 99214
rect 116008 99144 116220 99150
rect 116416 99214 116628 99280
rect 116416 99150 116558 99214
rect 116622 99150 116628 99214
rect 116416 99144 116628 99150
rect 116824 99350 117036 99356
rect 116824 99286 116830 99350
rect 116894 99286 117036 99350
rect 116824 99214 117036 99286
rect 116824 99150 116966 99214
rect 117030 99150 117036 99214
rect 116824 99144 117036 99150
rect 28560 98948 28636 99008
rect 110296 98948 110372 99008
rect 21760 98942 21972 98948
rect 21760 98878 21902 98942
rect 21966 98878 21972 98942
rect 21760 98806 21972 98878
rect 21760 98742 21902 98806
rect 21966 98742 21972 98806
rect 21760 98736 21972 98742
rect 22168 98942 22788 98948
rect 22168 98878 22582 98942
rect 22646 98878 22788 98942
rect 22168 98872 22788 98878
rect 22168 98806 22380 98872
rect 22168 98742 22174 98806
rect 22238 98742 22380 98806
rect 22168 98736 22380 98742
rect 22576 98736 22788 98872
rect 22984 98942 23196 98948
rect 22984 98878 22990 98942
rect 23054 98878 23196 98942
rect 22984 98806 23196 98878
rect 22984 98742 23126 98806
rect 23190 98742 23196 98806
rect 22984 98736 23196 98742
rect 23392 98942 23604 98948
rect 23392 98878 23398 98942
rect 23462 98878 23604 98942
rect 23392 98806 23604 98878
rect 23392 98742 23398 98806
rect 23462 98742 23604 98806
rect 23392 98736 23604 98742
rect 28288 98736 28636 98948
rect 110160 98736 110508 98948
rect 115192 98942 115404 98948
rect 115192 98878 115198 98942
rect 115262 98878 115404 98942
rect 115192 98806 115404 98878
rect 115192 98742 115198 98806
rect 115262 98742 115404 98806
rect 115192 98736 115404 98742
rect 115600 98942 115812 98948
rect 115600 98878 115606 98942
rect 115670 98878 115812 98942
rect 115600 98806 115812 98878
rect 115600 98742 115606 98806
rect 115670 98742 115812 98806
rect 115600 98736 115812 98742
rect 116008 98942 116220 98948
rect 116008 98878 116150 98942
rect 116214 98878 116220 98942
rect 116008 98812 116220 98878
rect 116416 98942 116628 98948
rect 116416 98878 116558 98942
rect 116622 98878 116628 98942
rect 116416 98812 116628 98878
rect 116008 98806 116628 98812
rect 116008 98742 116014 98806
rect 116078 98742 116628 98806
rect 116008 98736 116628 98742
rect 116824 98942 117036 98948
rect 116824 98878 116966 98942
rect 117030 98878 117036 98942
rect 116824 98806 117036 98878
rect 116824 98742 116966 98806
rect 117030 98742 117036 98806
rect 116824 98736 117036 98742
rect 28424 98676 28500 98736
rect 110160 98676 110236 98736
rect 21760 98534 21972 98540
rect 21760 98470 21902 98534
rect 21966 98470 21972 98534
rect 21760 98328 21972 98470
rect 22168 98534 22380 98540
rect 22168 98470 22174 98534
rect 22238 98470 22380 98534
rect 22168 98398 22380 98470
rect 22168 98334 22174 98398
rect 22238 98334 22380 98398
rect 22168 98328 22380 98334
rect 22576 98398 22788 98540
rect 22576 98334 22582 98398
rect 22646 98334 22788 98398
rect 22576 98328 22788 98334
rect 22984 98534 23196 98540
rect 22984 98470 23126 98534
rect 23190 98470 23196 98534
rect 22984 98398 23196 98470
rect 22984 98334 22990 98398
rect 23054 98334 23196 98398
rect 22984 98328 23196 98334
rect 23392 98534 23604 98540
rect 23392 98470 23398 98534
rect 23462 98470 23604 98534
rect 23392 98398 23604 98470
rect 28288 98464 28636 98676
rect 110160 98464 110508 98676
rect 28424 98404 28500 98464
rect 110432 98404 110508 98464
rect 23392 98334 23534 98398
rect 23598 98334 23604 98398
rect 23392 98328 23604 98334
rect 21896 98268 21972 98328
rect 1768 97860 1980 97996
rect 21760 97920 21972 98268
rect 28288 98192 28636 98404
rect 110160 98192 110508 98404
rect 115192 98534 115404 98540
rect 115192 98470 115198 98534
rect 115262 98470 115404 98534
rect 115192 98398 115404 98470
rect 115192 98334 115334 98398
rect 115398 98334 115404 98398
rect 115192 98328 115404 98334
rect 115600 98534 115812 98540
rect 115600 98470 115606 98534
rect 115670 98470 115812 98534
rect 115600 98398 115812 98470
rect 115600 98334 115742 98398
rect 115806 98334 115812 98398
rect 115600 98328 115812 98334
rect 116008 98534 116220 98540
rect 116008 98470 116014 98534
rect 116078 98470 116220 98534
rect 116008 98398 116220 98470
rect 116008 98334 116014 98398
rect 116078 98334 116220 98398
rect 116008 98328 116220 98334
rect 116416 98398 116628 98540
rect 116416 98334 116422 98398
rect 116486 98334 116628 98398
rect 116416 98328 116628 98334
rect 116824 98534 117036 98540
rect 116824 98470 116966 98534
rect 117030 98470 117036 98534
rect 116824 98328 117036 98470
rect 116824 98268 116900 98328
rect 28288 98132 28364 98192
rect 110296 98132 110372 98192
rect 21896 97860 21972 97920
rect 1224 97854 1980 97860
rect 1224 97790 1230 97854
rect 1294 97848 1980 97854
rect 1294 97792 1798 97848
rect 1854 97792 1980 97848
rect 1294 97790 1980 97792
rect 1224 97784 1980 97790
rect 1768 97648 1980 97784
rect 21760 97512 21972 97860
rect 22168 98126 22380 98132
rect 22168 98062 22174 98126
rect 22238 98062 22380 98126
rect 22168 97920 22380 98062
rect 22576 98126 22788 98132
rect 22576 98062 22582 98126
rect 22646 98062 22788 98126
rect 22576 97920 22788 98062
rect 22984 98126 23196 98132
rect 22984 98062 22990 98126
rect 23054 98062 23196 98126
rect 22984 97990 23196 98062
rect 22984 97926 23126 97990
rect 23190 97926 23196 97990
rect 22984 97920 23196 97926
rect 23392 98126 23604 98132
rect 23392 98062 23534 98126
rect 23598 98062 23604 98126
rect 23392 97990 23604 98062
rect 23392 97926 23398 97990
rect 23462 97926 23604 97990
rect 23392 97920 23604 97926
rect 28288 97990 28636 98132
rect 28288 97926 28294 97990
rect 28358 97926 28636 97990
rect 22168 97860 22244 97920
rect 22712 97860 22788 97920
rect 22168 97784 22788 97860
rect 22168 97512 22380 97784
rect 22576 97582 22788 97784
rect 22576 97518 22582 97582
rect 22646 97518 22788 97582
rect 22576 97512 22788 97518
rect 22984 97718 23196 97724
rect 22984 97654 23126 97718
rect 23190 97654 23196 97718
rect 22984 97582 23196 97654
rect 22984 97518 23126 97582
rect 23190 97518 23196 97582
rect 22984 97512 23196 97518
rect 23392 97718 23604 97724
rect 23392 97654 23398 97718
rect 23462 97654 23604 97718
rect 23392 97582 23604 97654
rect 23392 97518 23398 97582
rect 23462 97518 23604 97582
rect 23392 97512 23604 97518
rect 28288 97648 28636 97926
rect 110160 97648 110508 98132
rect 115192 98126 115404 98132
rect 115192 98062 115334 98126
rect 115398 98062 115404 98126
rect 115192 97990 115404 98062
rect 115192 97926 115198 97990
rect 115262 97926 115404 97990
rect 115192 97920 115404 97926
rect 115600 98126 115812 98132
rect 115600 98062 115742 98126
rect 115806 98062 115812 98126
rect 115600 97990 115812 98062
rect 115600 97926 115606 97990
rect 115670 97926 115812 97990
rect 115600 97920 115812 97926
rect 116008 98126 116628 98132
rect 116008 98062 116014 98126
rect 116078 98062 116422 98126
rect 116486 98062 116628 98126
rect 116008 98056 116628 98062
rect 116008 97920 116220 98056
rect 116416 97920 116628 98056
rect 116824 97920 117036 98268
rect 116552 97860 116628 97920
rect 116960 97860 117036 97920
rect 116008 97784 116628 97860
rect 115192 97718 115404 97724
rect 115192 97654 115198 97718
rect 115262 97654 115404 97718
rect 28288 97588 28364 97648
rect 110160 97588 110236 97648
rect 28288 97582 28636 97588
rect 28288 97518 28294 97582
rect 28358 97518 28636 97582
rect 21760 97452 21836 97512
rect 21760 97310 21972 97452
rect 28288 97376 28636 97518
rect 110160 97446 110508 97588
rect 115192 97582 115404 97654
rect 115192 97518 115334 97582
rect 115398 97518 115404 97582
rect 115192 97512 115404 97518
rect 115600 97718 115812 97724
rect 115600 97654 115606 97718
rect 115670 97654 115812 97718
rect 115600 97582 115812 97654
rect 115600 97518 115742 97582
rect 115806 97518 115812 97582
rect 115600 97512 115812 97518
rect 116008 97588 116220 97784
rect 116008 97582 116356 97588
rect 116008 97518 116286 97582
rect 116350 97518 116356 97582
rect 116008 97512 116356 97518
rect 116416 97512 116628 97784
rect 116824 97512 117036 97860
rect 136816 97860 137028 97996
rect 136816 97854 137572 97860
rect 136816 97848 137502 97854
rect 136816 97792 136944 97848
rect 137000 97792 137502 97848
rect 136816 97790 137502 97792
rect 137566 97790 137572 97854
rect 136816 97784 137572 97790
rect 136816 97648 137028 97784
rect 110160 97382 110166 97446
rect 110230 97382 110508 97446
rect 110160 97376 110508 97382
rect 28424 97316 28500 97376
rect 110432 97316 110508 97376
rect 116824 97452 116900 97512
rect 21760 97246 21766 97310
rect 21830 97246 21972 97310
rect 21760 97240 21972 97246
rect 22168 97310 22788 97316
rect 22168 97246 22582 97310
rect 22646 97246 22788 97310
rect 22168 97240 22788 97246
rect 22168 97104 22380 97240
rect 22576 97104 22788 97240
rect 22984 97310 23196 97316
rect 22984 97246 23126 97310
rect 23190 97246 23196 97310
rect 22984 97104 23196 97246
rect 23392 97310 23604 97316
rect 23392 97246 23398 97310
rect 23462 97246 23604 97310
rect 23392 97104 23604 97246
rect 22168 97044 22244 97104
rect 22576 97044 22652 97104
rect 22984 97044 23060 97104
rect 23528 97044 23604 97104
rect 21760 97038 21972 97044
rect 21760 96974 21766 97038
rect 21830 96974 21972 97038
rect 21760 96902 21972 96974
rect 21760 96838 21902 96902
rect 21966 96838 21972 96902
rect 21760 96832 21972 96838
rect 22168 96832 22380 97044
rect 22576 96902 22788 97044
rect 22576 96838 22718 96902
rect 22782 96838 22788 96902
rect 22576 96832 22788 96838
rect 22984 96696 23196 97044
rect 23120 96636 23196 96696
rect 21760 96630 21972 96636
rect 21760 96566 21902 96630
rect 21966 96566 21972 96630
rect 21760 96494 21972 96566
rect 21760 96430 21766 96494
rect 21830 96430 21972 96494
rect 21760 96424 21972 96430
rect 22168 96500 22380 96636
rect 22576 96630 22788 96636
rect 22576 96566 22718 96630
rect 22782 96566 22788 96630
rect 22576 96500 22788 96566
rect 22168 96424 22788 96500
rect 22984 96494 23196 96636
rect 22984 96430 22990 96494
rect 23054 96430 23196 96494
rect 22984 96424 23196 96430
rect 23392 96696 23604 97044
rect 28288 97038 28636 97316
rect 28288 96974 28430 97038
rect 28494 96974 28636 97038
rect 28288 96968 28636 96974
rect 110160 97174 110508 97316
rect 110160 97110 110166 97174
rect 110230 97110 110508 97174
rect 110160 97038 110508 97110
rect 115192 97310 115404 97316
rect 115192 97246 115334 97310
rect 115398 97246 115404 97310
rect 115192 97104 115404 97246
rect 115600 97310 115812 97316
rect 115600 97246 115742 97310
rect 115806 97246 115812 97310
rect 115600 97104 115812 97246
rect 115328 97044 115404 97104
rect 115736 97044 115812 97104
rect 110160 96974 110302 97038
rect 110366 96974 110508 97038
rect 110160 96968 110508 96974
rect 28288 96766 28636 96772
rect 28288 96702 28430 96766
rect 28494 96702 28636 96766
rect 23392 96636 23468 96696
rect 23392 96494 23604 96636
rect 23392 96430 23534 96494
rect 23598 96430 23604 96494
rect 23392 96424 23604 96430
rect 28288 96424 28636 96702
rect 110160 96766 110508 96772
rect 110160 96702 110302 96766
rect 110366 96702 110508 96766
rect 110160 96424 110508 96702
rect 115192 96696 115404 97044
rect 115600 96696 115812 97044
rect 116008 97104 116220 97316
rect 116318 97310 116628 97316
rect 116280 97246 116286 97310
rect 116350 97246 116628 97310
rect 116318 97240 116628 97246
rect 116824 97310 117036 97452
rect 116824 97246 116830 97310
rect 116894 97246 117036 97310
rect 116824 97240 117036 97246
rect 116416 97104 116628 97240
rect 116008 97044 116084 97104
rect 116416 97044 116492 97104
rect 116008 96968 116628 97044
rect 116008 96832 116220 96968
rect 116416 96902 116628 96968
rect 116416 96838 116558 96902
rect 116622 96838 116628 96902
rect 116416 96832 116628 96838
rect 116824 97038 117036 97044
rect 116824 96974 116830 97038
rect 116894 96974 117036 97038
rect 116824 96902 117036 96974
rect 116824 96838 116966 96902
rect 117030 96838 117036 96902
rect 116824 96832 117036 96838
rect 115192 96636 115268 96696
rect 115736 96636 115812 96696
rect 115192 96494 115404 96636
rect 115192 96430 115334 96494
rect 115398 96430 115404 96494
rect 115192 96424 115404 96430
rect 115600 96494 115812 96636
rect 115600 96430 115742 96494
rect 115806 96430 115812 96494
rect 115600 96424 115812 96430
rect 116008 96500 116220 96636
rect 116416 96630 116628 96636
rect 116416 96566 116558 96630
rect 116622 96566 116628 96630
rect 116008 96494 116356 96500
rect 116008 96430 116286 96494
rect 116350 96430 116356 96494
rect 116008 96424 116356 96430
rect 22168 96288 22380 96424
rect 22576 96288 22788 96424
rect 28560 96364 28636 96424
rect 110296 96364 110372 96424
rect 116008 96364 116220 96424
rect 116416 96364 116628 96566
rect 116824 96630 117036 96636
rect 116824 96566 116966 96630
rect 117030 96566 117036 96630
rect 116824 96494 117036 96566
rect 116824 96430 116966 96494
rect 117030 96430 117036 96494
rect 116824 96424 117036 96430
rect 22576 96228 22652 96288
rect 1224 96222 1980 96228
rect 1224 96158 1230 96222
rect 1294 96168 1980 96222
rect 1294 96158 1798 96168
rect 1224 96152 1798 96158
rect 1768 96112 1798 96152
rect 1854 96112 1980 96168
rect 1768 96016 1980 96112
rect 21760 96222 21972 96228
rect 21760 96158 21766 96222
rect 21830 96158 21972 96222
rect 21760 96086 21972 96158
rect 21760 96022 21902 96086
rect 21966 96022 21972 96086
rect 21760 96016 21972 96022
rect 22168 96086 22380 96228
rect 22168 96022 22174 96086
rect 22238 96022 22380 96086
rect 22168 96016 22380 96022
rect 22576 96086 22788 96228
rect 22576 96022 22718 96086
rect 22782 96022 22788 96086
rect 22576 96016 22788 96022
rect 22984 96222 23196 96228
rect 22984 96158 22990 96222
rect 23054 96158 23196 96222
rect 22984 96086 23196 96158
rect 22984 96022 22990 96086
rect 23054 96022 23196 96086
rect 22984 96016 23196 96022
rect 23392 96222 23604 96228
rect 23392 96158 23534 96222
rect 23598 96158 23604 96222
rect 23392 96086 23604 96158
rect 28288 96152 28636 96364
rect 110160 96152 110508 96364
rect 116008 96288 116628 96364
rect 116008 96228 116084 96288
rect 28424 96092 28500 96152
rect 110432 96092 110508 96152
rect 23392 96022 23398 96086
rect 23462 96022 23604 96086
rect 23392 96016 23604 96022
rect 21760 95814 21972 95820
rect 21760 95750 21902 95814
rect 21966 95750 21972 95814
rect 21760 95678 21972 95750
rect 21760 95614 21902 95678
rect 21966 95614 21972 95678
rect 21760 95608 21972 95614
rect 22168 95814 22380 95820
rect 22168 95750 22174 95814
rect 22238 95750 22380 95814
rect 22168 95684 22380 95750
rect 22576 95814 22788 95820
rect 22576 95750 22718 95814
rect 22782 95750 22788 95814
rect 22576 95684 22788 95750
rect 22168 95608 22788 95684
rect 22984 95814 23196 95820
rect 22984 95750 22990 95814
rect 23054 95750 23196 95814
rect 22984 95678 23196 95750
rect 22984 95614 22990 95678
rect 23054 95614 23196 95678
rect 22984 95608 23196 95614
rect 23392 95814 23604 95820
rect 23392 95750 23398 95814
rect 23462 95750 23604 95814
rect 23392 95678 23604 95750
rect 23392 95614 23398 95678
rect 23462 95614 23604 95678
rect 23392 95608 23604 95614
rect 28288 95814 28636 96092
rect 28288 95750 28430 95814
rect 28494 95750 28636 95814
rect 28288 95608 28636 95750
rect 110160 95814 110508 96092
rect 115192 96222 115404 96228
rect 115192 96158 115334 96222
rect 115398 96158 115404 96222
rect 115192 96086 115404 96158
rect 115192 96022 115334 96086
rect 115398 96022 115404 96086
rect 115192 96016 115404 96022
rect 115600 96222 115812 96228
rect 115600 96158 115742 96222
rect 115806 96158 115812 96222
rect 115600 96086 115812 96158
rect 115600 96022 115742 96086
rect 115806 96022 115812 96086
rect 115600 96016 115812 96022
rect 116008 96016 116220 96228
rect 116318 96222 116628 96228
rect 116280 96158 116286 96222
rect 116350 96158 116628 96222
rect 116318 96152 116628 96158
rect 116416 96086 116628 96152
rect 116416 96022 116558 96086
rect 116622 96022 116628 96086
rect 116416 96016 116628 96022
rect 116824 96222 117036 96228
rect 116824 96158 116966 96222
rect 117030 96158 117036 96222
rect 116824 96086 117036 96158
rect 116824 96022 116966 96086
rect 117030 96022 117036 96086
rect 116824 96016 117036 96022
rect 136816 96168 137028 96228
rect 136816 96112 136944 96168
rect 137000 96112 137028 96168
rect 136816 96092 137028 96112
rect 136816 96086 137572 96092
rect 136816 96022 137502 96086
rect 137566 96022 137572 96086
rect 136816 96016 137572 96022
rect 110160 95750 110166 95814
rect 110230 95750 110508 95814
rect 110160 95608 110508 95750
rect 115192 95814 115404 95820
rect 115192 95750 115334 95814
rect 115398 95750 115404 95814
rect 115192 95678 115404 95750
rect 115192 95614 115198 95678
rect 115262 95614 115404 95678
rect 115192 95608 115404 95614
rect 115600 95814 115812 95820
rect 115600 95750 115742 95814
rect 115806 95750 115812 95814
rect 115600 95678 115812 95750
rect 115600 95614 115606 95678
rect 115670 95614 115812 95678
rect 115600 95608 115812 95614
rect 116008 95684 116220 95820
rect 116416 95814 116628 95820
rect 116416 95750 116558 95814
rect 116622 95750 116628 95814
rect 116416 95684 116628 95750
rect 116008 95678 116628 95684
rect 116008 95614 116150 95678
rect 116214 95614 116628 95678
rect 116008 95608 116628 95614
rect 116824 95814 117036 95820
rect 116824 95750 116966 95814
rect 117030 95750 117036 95814
rect 116824 95678 117036 95750
rect 116824 95614 116966 95678
rect 117030 95614 117036 95678
rect 116824 95608 117036 95614
rect 22304 95548 22380 95608
rect 28288 95548 28364 95608
rect 110432 95548 110508 95608
rect 22304 95472 22652 95548
rect 22576 95412 22652 95472
rect 28288 95542 28636 95548
rect 28288 95478 28430 95542
rect 28494 95478 28636 95542
rect 21760 95406 21972 95412
rect 21760 95342 21902 95406
rect 21966 95342 21972 95406
rect 21760 95270 21972 95342
rect 21760 95206 21766 95270
rect 21830 95206 21972 95270
rect 21760 95200 21972 95206
rect 22168 95270 22380 95412
rect 22168 95206 22174 95270
rect 22238 95206 22380 95270
rect 22168 95200 22380 95206
rect 22576 95270 22788 95412
rect 22576 95206 22582 95270
rect 22646 95206 22788 95270
rect 22576 95200 22788 95206
rect 22984 95406 23196 95412
rect 22984 95342 22990 95406
rect 23054 95342 23196 95406
rect 22984 95270 23196 95342
rect 22984 95206 23126 95270
rect 23190 95206 23196 95270
rect 22984 95200 23196 95206
rect 23392 95406 23604 95412
rect 23392 95342 23398 95406
rect 23462 95342 23604 95406
rect 23392 95270 23604 95342
rect 28288 95336 28636 95478
rect 28560 95276 28636 95336
rect 23392 95206 23534 95270
rect 23598 95206 23604 95270
rect 23392 95200 23604 95206
rect 28288 95064 28636 95276
rect 110160 95542 110508 95548
rect 110160 95478 110166 95542
rect 110230 95478 110508 95542
rect 110160 95336 110508 95478
rect 115192 95406 115404 95412
rect 115192 95342 115198 95406
rect 115262 95342 115404 95406
rect 110160 95276 110236 95336
rect 110160 95064 110508 95276
rect 115192 95270 115404 95342
rect 115192 95206 115334 95270
rect 115398 95206 115404 95270
rect 115192 95200 115404 95206
rect 115600 95406 115812 95412
rect 115600 95342 115606 95406
rect 115670 95342 115812 95406
rect 115600 95270 115812 95342
rect 115600 95206 115742 95270
rect 115806 95206 115812 95270
rect 115600 95200 115812 95206
rect 116008 95406 116220 95412
rect 116008 95342 116150 95406
rect 116214 95342 116220 95406
rect 116008 95270 116220 95342
rect 116008 95206 116014 95270
rect 116078 95206 116220 95270
rect 116008 95200 116220 95206
rect 116416 95270 116628 95412
rect 116416 95206 116422 95270
rect 116486 95206 116628 95270
rect 116416 95200 116628 95206
rect 116824 95406 117036 95412
rect 116824 95342 116966 95406
rect 117030 95342 117036 95406
rect 116824 95270 117036 95342
rect 116824 95206 116830 95270
rect 116894 95206 117036 95270
rect 116824 95200 117036 95206
rect 28424 95004 28500 95064
rect 110296 95004 110372 95064
rect 21760 94998 21972 95004
rect 21760 94934 21766 94998
rect 21830 94934 21972 94998
rect 21760 94862 21972 94934
rect 21760 94798 21902 94862
rect 21966 94798 21972 94862
rect 21760 94792 21972 94798
rect 22168 94998 22380 95004
rect 22168 94934 22174 94998
rect 22238 94934 22380 94998
rect 22168 94862 22380 94934
rect 22168 94798 22310 94862
rect 22374 94798 22380 94862
rect 22168 94792 22380 94798
rect 22576 94998 22788 95004
rect 22576 94934 22582 94998
rect 22646 94934 22788 94998
rect 22576 94792 22788 94934
rect 22984 94998 23196 95004
rect 22984 94934 23126 94998
rect 23190 94934 23196 94998
rect 22984 94862 23196 94934
rect 22984 94798 23126 94862
rect 23190 94798 23196 94862
rect 22984 94792 23196 94798
rect 23392 94998 23604 95004
rect 23392 94934 23534 94998
rect 23598 94934 23604 94998
rect 23392 94862 23604 94934
rect 23392 94798 23534 94862
rect 23598 94798 23604 94862
rect 23392 94792 23604 94798
rect 28288 94792 28636 95004
rect 110160 94792 110508 95004
rect 115192 94998 115404 95004
rect 115192 94934 115334 94998
rect 115398 94934 115404 94998
rect 115192 94862 115404 94934
rect 115192 94798 115198 94862
rect 115262 94798 115404 94862
rect 115192 94792 115404 94798
rect 115600 94998 115812 95004
rect 115600 94934 115742 94998
rect 115806 94934 115812 94998
rect 115600 94862 115812 94934
rect 115600 94798 115606 94862
rect 115670 94798 115812 94862
rect 115600 94792 115812 94798
rect 116008 94998 116628 95004
rect 116008 94934 116014 94998
rect 116078 94934 116422 94998
rect 116486 94934 116628 94998
rect 116008 94928 116628 94934
rect 116008 94868 116220 94928
rect 116008 94792 116356 94868
rect 116416 94792 116628 94928
rect 116824 94998 117036 95004
rect 116824 94934 116830 94998
rect 116894 94934 117036 94998
rect 116824 94862 117036 94934
rect 116824 94798 116830 94862
rect 116894 94798 117036 94862
rect 116824 94792 117036 94798
rect 22576 94732 22652 94792
rect 22304 94656 22652 94732
rect 28288 94732 28364 94792
rect 110432 94732 110508 94792
rect 22304 94596 22380 94656
rect 1224 94590 1980 94596
rect 1224 94526 1230 94590
rect 1294 94526 1980 94590
rect 1224 94520 1980 94526
rect 1768 94488 1980 94520
rect 1768 94432 1798 94488
rect 1854 94432 1980 94488
rect 1768 94384 1980 94432
rect 21760 94590 21972 94596
rect 21760 94526 21902 94590
rect 21966 94526 21972 94590
rect 21760 94384 21972 94526
rect 22168 94590 22788 94596
rect 22168 94526 22310 94590
rect 22374 94526 22788 94590
rect 22168 94520 22788 94526
rect 22168 94384 22380 94520
rect 22576 94454 22788 94520
rect 22576 94390 22582 94454
rect 22646 94390 22788 94454
rect 22576 94384 22788 94390
rect 22984 94590 23196 94596
rect 22984 94526 23126 94590
rect 23190 94526 23196 94590
rect 22984 94454 23196 94526
rect 22984 94390 23126 94454
rect 23190 94390 23196 94454
rect 22984 94384 23196 94390
rect 23392 94590 23604 94596
rect 23392 94526 23534 94590
rect 23598 94526 23604 94590
rect 23392 94454 23604 94526
rect 28288 94520 28636 94732
rect 110160 94520 110508 94732
rect 116280 94732 116356 94792
rect 116280 94656 116492 94732
rect 116416 94596 116492 94656
rect 115192 94590 115404 94596
rect 115192 94526 115198 94590
rect 115262 94526 115404 94590
rect 28424 94460 28500 94520
rect 110296 94460 110372 94520
rect 23392 94390 23398 94454
rect 23462 94390 23604 94454
rect 23392 94384 23604 94390
rect 21896 94324 21972 94384
rect 21760 93976 21972 94324
rect 28288 94248 28636 94460
rect 110160 94318 110508 94460
rect 115192 94454 115404 94526
rect 115192 94390 115334 94454
rect 115398 94390 115404 94454
rect 115192 94384 115404 94390
rect 115600 94590 115812 94596
rect 115600 94526 115606 94590
rect 115670 94526 115812 94590
rect 115600 94454 115812 94526
rect 115600 94390 115606 94454
rect 115670 94390 115812 94454
rect 115600 94384 115812 94390
rect 116008 94520 116628 94596
rect 116008 94460 116220 94520
rect 116008 94454 116356 94460
rect 116008 94390 116014 94454
rect 116078 94390 116286 94454
rect 116350 94390 116356 94454
rect 116008 94384 116356 94390
rect 116416 94384 116628 94520
rect 116824 94590 117036 94596
rect 116824 94526 116830 94590
rect 116894 94526 117036 94590
rect 116824 94384 117036 94526
rect 136816 94488 137028 94596
rect 136816 94432 136944 94488
rect 137000 94460 137028 94488
rect 137000 94454 137572 94460
rect 137000 94432 137502 94454
rect 136816 94390 137502 94432
rect 137566 94390 137572 94454
rect 136816 94384 137572 94390
rect 116960 94324 117036 94384
rect 110160 94254 110166 94318
rect 110230 94254 110508 94318
rect 110160 94248 110508 94254
rect 28424 94188 28500 94248
rect 110432 94188 110508 94248
rect 21896 93916 21972 93976
rect 21760 93568 21972 93916
rect 22168 93976 22380 94188
rect 22576 94182 22788 94188
rect 22576 94118 22582 94182
rect 22646 94118 22788 94182
rect 22576 94052 22788 94118
rect 22440 93976 22788 94052
rect 22984 94182 23196 94188
rect 22984 94118 23126 94182
rect 23190 94118 23196 94182
rect 22984 94046 23196 94118
rect 22984 93982 23126 94046
rect 23190 93982 23196 94046
rect 22984 93976 23196 93982
rect 23392 94182 23604 94188
rect 23392 94118 23398 94182
rect 23462 94118 23604 94182
rect 23392 94046 23604 94118
rect 23392 93982 23534 94046
rect 23598 93982 23604 94046
rect 23392 93976 23604 93982
rect 22168 93916 22244 93976
rect 22440 93916 22516 93976
rect 22168 93840 22516 93916
rect 22576 93916 22652 93976
rect 22168 93568 22380 93840
rect 22576 93644 22788 93916
rect 22478 93638 22788 93644
rect 22440 93574 22446 93638
rect 22510 93574 22788 93638
rect 22478 93568 22788 93574
rect 22984 93774 23196 93780
rect 22984 93710 23126 93774
rect 23190 93710 23196 93774
rect 22984 93638 23196 93710
rect 22984 93574 22990 93638
rect 23054 93574 23196 93638
rect 22984 93568 23196 93574
rect 23392 93774 23604 93780
rect 23392 93710 23534 93774
rect 23598 93710 23604 93774
rect 23392 93638 23604 93710
rect 23392 93574 23398 93638
rect 23462 93574 23604 93638
rect 23392 93568 23604 93574
rect 28288 93704 28636 94188
rect 110160 94046 110508 94188
rect 110160 93982 110166 94046
rect 110230 93982 110508 94046
rect 110160 93704 110508 93982
rect 115192 94182 115404 94188
rect 115192 94118 115334 94182
rect 115398 94118 115404 94182
rect 115192 94046 115404 94118
rect 115192 93982 115334 94046
rect 115398 93982 115404 94046
rect 115192 93976 115404 93982
rect 115600 94182 115812 94188
rect 115600 94118 115606 94182
rect 115670 94118 115812 94182
rect 115600 94046 115812 94118
rect 115600 93982 115742 94046
rect 115806 93982 115812 94046
rect 115600 93976 115812 93982
rect 116008 94182 116220 94188
rect 116318 94182 116628 94188
rect 116008 94118 116014 94182
rect 116078 94118 116220 94182
rect 116280 94118 116286 94182
rect 116350 94118 116628 94182
rect 116008 93976 116220 94118
rect 116318 94112 116628 94118
rect 116416 94052 116628 94112
rect 116280 93976 116628 94052
rect 116824 93976 117036 94324
rect 116280 93916 116356 93976
rect 116552 93916 116628 93976
rect 116960 93916 117036 93976
rect 116008 93840 116356 93916
rect 28288 93644 28364 93704
rect 110432 93644 110508 93704
rect 21896 93508 21972 93568
rect 21760 93366 21972 93508
rect 22304 93432 22652 93508
rect 28288 93502 28636 93644
rect 28288 93438 28566 93502
rect 28630 93438 28636 93502
rect 28288 93432 28636 93438
rect 110160 93432 110508 93644
rect 115192 93774 115404 93780
rect 115192 93710 115334 93774
rect 115398 93710 115404 93774
rect 115192 93638 115404 93710
rect 115192 93574 115198 93638
rect 115262 93574 115404 93638
rect 115192 93568 115404 93574
rect 115600 93774 115812 93780
rect 115600 93710 115742 93774
rect 115806 93710 115812 93774
rect 115600 93638 115812 93710
rect 115600 93574 115606 93638
rect 115670 93574 115812 93638
rect 115600 93568 115812 93574
rect 116008 93568 116220 93840
rect 116416 93638 116628 93916
rect 116416 93574 116422 93638
rect 116486 93574 116628 93638
rect 116416 93568 116628 93574
rect 116824 93568 117036 93916
rect 116960 93508 117036 93568
rect 22304 93372 22380 93432
rect 22576 93372 22652 93432
rect 28560 93372 28636 93432
rect 110296 93372 110372 93432
rect 21760 93302 21902 93366
rect 21966 93302 21972 93366
rect 21760 93296 21972 93302
rect 22168 93366 22516 93372
rect 22168 93302 22446 93366
rect 22510 93302 22516 93366
rect 22168 93296 22516 93302
rect 22168 93236 22380 93296
rect 22168 93160 22516 93236
rect 22576 93160 22788 93372
rect 22984 93366 23196 93372
rect 22984 93302 22990 93366
rect 23054 93302 23196 93366
rect 22984 93160 23196 93302
rect 23392 93366 23604 93372
rect 23392 93302 23398 93366
rect 23462 93302 23604 93366
rect 23392 93160 23604 93302
rect 22304 93100 22380 93160
rect 21760 93094 21972 93100
rect 21760 93030 21902 93094
rect 21966 93030 21972 93094
rect 1224 92958 1980 92964
rect 1224 92894 1230 92958
rect 1294 92894 1980 92958
rect 1224 92888 1980 92894
rect 21760 92958 21972 93030
rect 21760 92894 21766 92958
rect 21830 92894 21972 92958
rect 21760 92888 21972 92894
rect 22168 92888 22380 93100
rect 22440 93100 22516 93160
rect 23120 93100 23196 93160
rect 23528 93100 23604 93160
rect 22440 93024 22788 93100
rect 22576 92958 22788 93024
rect 22576 92894 22582 92958
rect 22646 92894 22788 92958
rect 22576 92888 22788 92894
rect 1768 92808 1980 92888
rect 1768 92752 1798 92808
rect 1854 92752 1980 92808
rect 22984 92752 23196 93100
rect 23392 92752 23604 93100
rect 28288 93230 28636 93372
rect 28288 93166 28566 93230
rect 28630 93166 28636 93230
rect 28288 93094 28636 93166
rect 28288 93030 28294 93094
rect 28358 93030 28636 93094
rect 28288 93024 28636 93030
rect 110160 93094 110508 93372
rect 110160 93030 110302 93094
rect 110366 93030 110508 93094
rect 110160 93024 110508 93030
rect 115192 93366 115404 93372
rect 115192 93302 115198 93366
rect 115262 93302 115404 93366
rect 115192 93160 115404 93302
rect 115600 93366 115812 93372
rect 115600 93302 115606 93366
rect 115670 93302 115812 93366
rect 115600 93160 115812 93302
rect 116008 93366 116628 93372
rect 116008 93302 116422 93366
rect 116486 93302 116628 93366
rect 116008 93296 116628 93302
rect 116824 93366 117036 93508
rect 116824 93302 116830 93366
rect 116894 93302 117036 93366
rect 116824 93296 117036 93302
rect 116008 93236 116220 93296
rect 116008 93160 116356 93236
rect 116416 93160 116628 93296
rect 115192 93100 115268 93160
rect 115600 93100 115676 93160
rect 116144 93100 116220 93160
rect 1768 92616 1980 92752
rect 23120 92692 23196 92752
rect 23528 92692 23604 92752
rect 21760 92686 21972 92692
rect 21760 92622 21766 92686
rect 21830 92622 21972 92686
rect 21760 92550 21972 92622
rect 21760 92486 21902 92550
rect 21966 92486 21972 92550
rect 21760 92480 21972 92486
rect 22168 92344 22380 92692
rect 22576 92686 22788 92692
rect 22576 92622 22582 92686
rect 22646 92622 22788 92686
rect 22576 92420 22788 92622
rect 22304 92284 22380 92344
rect 22440 92344 22788 92420
rect 22984 92344 23196 92692
rect 22440 92284 22516 92344
rect 22712 92284 22788 92344
rect 23120 92284 23196 92344
rect 21760 92278 21972 92284
rect 21760 92214 21902 92278
rect 21966 92214 21972 92278
rect 21760 92142 21972 92214
rect 21760 92078 21766 92142
rect 21830 92078 21972 92142
rect 21760 92072 21972 92078
rect 22168 92208 22516 92284
rect 22168 92148 22380 92208
rect 22168 92142 22516 92148
rect 22168 92078 22446 92142
rect 22510 92078 22516 92142
rect 22168 92072 22516 92078
rect 22576 92072 22788 92284
rect 22984 92142 23196 92284
rect 22984 92078 23126 92142
rect 23190 92078 23196 92142
rect 22984 92072 23196 92078
rect 23392 92344 23604 92692
rect 28288 92822 28636 92828
rect 28288 92758 28294 92822
rect 28358 92758 28636 92822
rect 28288 92686 28636 92758
rect 28288 92622 28566 92686
rect 28630 92622 28636 92686
rect 28288 92414 28636 92622
rect 28288 92350 28430 92414
rect 28494 92350 28566 92414
rect 28630 92350 28636 92414
rect 23392 92284 23468 92344
rect 23392 92142 23604 92284
rect 28288 92208 28636 92350
rect 28560 92148 28636 92208
rect 23392 92078 23534 92142
rect 23598 92078 23604 92142
rect 23392 92072 23604 92078
rect 28288 92142 28636 92148
rect 28288 92078 28430 92142
rect 28494 92078 28636 92142
rect 21760 91870 21972 91876
rect 21760 91806 21766 91870
rect 21830 91806 21972 91870
rect 21760 91734 21972 91806
rect 21760 91670 21766 91734
rect 21830 91670 21972 91734
rect 21760 91664 21972 91670
rect 22168 91734 22380 91876
rect 22478 91870 22788 91876
rect 22440 91806 22446 91870
rect 22510 91806 22788 91870
rect 22478 91800 22788 91806
rect 22168 91670 22310 91734
rect 22374 91670 22380 91734
rect 22168 91664 22380 91670
rect 22576 91734 22788 91800
rect 22576 91670 22718 91734
rect 22782 91670 22788 91734
rect 22576 91664 22788 91670
rect 22984 91870 23196 91876
rect 22984 91806 23126 91870
rect 23190 91806 23196 91870
rect 22984 91734 23196 91806
rect 22984 91670 22990 91734
rect 23054 91670 23196 91734
rect 22984 91664 23196 91670
rect 23392 91870 23604 91876
rect 23392 91806 23534 91870
rect 23598 91806 23604 91870
rect 23392 91734 23604 91806
rect 23392 91670 23534 91734
rect 23598 91670 23604 91734
rect 23392 91664 23604 91670
rect 28288 91664 28636 92078
rect 110160 92822 110508 92828
rect 110160 92758 110302 92822
rect 110366 92758 110508 92822
rect 110160 92686 110508 92758
rect 115192 92752 115404 93100
rect 115600 92752 115812 93100
rect 116008 92888 116220 93100
rect 116280 93100 116356 93160
rect 116280 93024 116628 93100
rect 116416 92958 116628 93024
rect 116416 92894 116422 92958
rect 116486 92894 116628 92958
rect 116416 92888 116628 92894
rect 116824 93094 117036 93100
rect 116824 93030 116830 93094
rect 116894 93030 117036 93094
rect 116824 92958 117036 93030
rect 116824 92894 116830 92958
rect 116894 92894 117036 92958
rect 116824 92888 117036 92894
rect 136816 92958 137572 92964
rect 136816 92894 137502 92958
rect 137566 92894 137572 92958
rect 136816 92888 137572 92894
rect 115328 92692 115404 92752
rect 115736 92692 115812 92752
rect 136816 92808 137028 92888
rect 136816 92752 136944 92808
rect 137000 92752 137028 92808
rect 110160 92622 110302 92686
rect 110366 92622 110508 92686
rect 110160 92414 110508 92622
rect 110160 92350 110302 92414
rect 110366 92350 110508 92414
rect 110160 92208 110508 92350
rect 115192 92344 115404 92692
rect 115600 92344 115812 92692
rect 116008 92686 116628 92692
rect 116008 92622 116422 92686
rect 116486 92622 116628 92686
rect 116008 92616 116628 92622
rect 116008 92344 116220 92616
rect 116416 92420 116628 92616
rect 116824 92686 117036 92692
rect 116824 92622 116830 92686
rect 116894 92622 117036 92686
rect 116824 92550 117036 92622
rect 136816 92616 137028 92752
rect 116824 92486 116966 92550
rect 117030 92486 117036 92550
rect 116824 92480 117036 92486
rect 116280 92344 116628 92420
rect 115192 92284 115268 92344
rect 115600 92284 115676 92344
rect 116280 92284 116356 92344
rect 110160 92148 110236 92208
rect 110160 91870 110508 92148
rect 115192 92142 115404 92284
rect 115192 92078 115334 92142
rect 115398 92078 115404 92142
rect 115192 92072 115404 92078
rect 115600 92142 115812 92284
rect 115600 92078 115606 92142
rect 115670 92078 115812 92142
rect 115600 92072 115812 92078
rect 116008 92208 116356 92284
rect 116008 92148 116220 92208
rect 116008 92142 116356 92148
rect 116008 92078 116286 92142
rect 116350 92078 116356 92142
rect 116008 92072 116356 92078
rect 116416 92072 116628 92284
rect 116824 92278 117036 92284
rect 116824 92214 116966 92278
rect 117030 92214 117036 92278
rect 116824 92142 117036 92214
rect 116824 92078 116966 92142
rect 117030 92078 117036 92142
rect 116824 92072 117036 92078
rect 116144 92012 116220 92072
rect 116416 92012 116492 92072
rect 116144 91936 116492 92012
rect 110160 91806 110438 91870
rect 110502 91806 110508 91870
rect 110160 91664 110508 91806
rect 115192 91870 115404 91876
rect 115192 91806 115334 91870
rect 115398 91806 115404 91870
rect 115192 91734 115404 91806
rect 115192 91670 115334 91734
rect 115398 91670 115404 91734
rect 115192 91664 115404 91670
rect 115600 91870 115812 91876
rect 115600 91806 115606 91870
rect 115670 91806 115812 91870
rect 115600 91734 115812 91806
rect 115600 91670 115606 91734
rect 115670 91670 115812 91734
rect 115600 91664 115812 91670
rect 116008 91740 116220 91876
rect 116318 91870 116628 91876
rect 116280 91806 116286 91870
rect 116350 91806 116628 91870
rect 116318 91800 116628 91806
rect 116416 91740 116628 91800
rect 116008 91734 116628 91740
rect 116008 91670 116150 91734
rect 116214 91670 116628 91734
rect 116008 91664 116628 91670
rect 116824 91870 117036 91876
rect 116824 91806 116966 91870
rect 117030 91806 117036 91870
rect 116824 91734 117036 91806
rect 116824 91670 116966 91734
rect 117030 91670 117036 91734
rect 116824 91664 117036 91670
rect 28424 91604 28500 91664
rect 110432 91604 110508 91664
rect 21760 91462 21972 91468
rect 21760 91398 21766 91462
rect 21830 91398 21972 91462
rect 21760 91326 21972 91398
rect 21760 91262 21902 91326
rect 21966 91262 21972 91326
rect 21760 91256 21972 91262
rect 22168 91462 22380 91468
rect 22168 91398 22310 91462
rect 22374 91398 22380 91462
rect 22168 91332 22380 91398
rect 22576 91462 22788 91468
rect 22576 91398 22718 91462
rect 22782 91398 22788 91462
rect 22576 91332 22788 91398
rect 22168 91326 22788 91332
rect 22168 91262 22174 91326
rect 22238 91262 22718 91326
rect 22782 91262 22788 91326
rect 22168 91256 22788 91262
rect 22984 91462 23196 91468
rect 22984 91398 22990 91462
rect 23054 91398 23196 91462
rect 22984 91326 23196 91398
rect 22984 91262 22990 91326
rect 23054 91262 23196 91326
rect 22984 91256 23196 91262
rect 23392 91462 23604 91468
rect 23392 91398 23534 91462
rect 23598 91398 23604 91462
rect 23392 91326 23604 91398
rect 23392 91262 23398 91326
rect 23462 91262 23604 91326
rect 23392 91256 23604 91262
rect 28288 91392 28636 91604
rect 110160 91598 110508 91604
rect 110160 91534 110438 91598
rect 110502 91534 110508 91598
rect 110160 91392 110508 91534
rect 116144 91604 116220 91664
rect 116144 91528 116492 91604
rect 116416 91468 116492 91528
rect 28288 91332 28364 91392
rect 110432 91332 110508 91392
rect 1224 91190 1980 91196
rect 1224 91126 1230 91190
rect 1294 91128 1980 91190
rect 1294 91126 1798 91128
rect 1224 91120 1798 91126
rect 1768 91072 1798 91120
rect 1854 91072 1980 91128
rect 28288 91120 28636 91332
rect 110160 91120 110508 91332
rect 115192 91462 115404 91468
rect 115192 91398 115334 91462
rect 115398 91398 115404 91462
rect 115192 91326 115404 91398
rect 115192 91262 115198 91326
rect 115262 91262 115404 91326
rect 115192 91256 115404 91262
rect 115600 91462 115812 91468
rect 115600 91398 115606 91462
rect 115670 91398 115812 91462
rect 115600 91326 115812 91398
rect 115600 91262 115606 91326
rect 115670 91262 115812 91326
rect 115600 91256 115812 91262
rect 116008 91462 116220 91468
rect 116008 91398 116150 91462
rect 116214 91398 116220 91462
rect 116008 91326 116220 91398
rect 116008 91262 116150 91326
rect 116214 91262 116220 91326
rect 116008 91256 116220 91262
rect 116416 91256 116628 91468
rect 116824 91462 117036 91468
rect 116824 91398 116966 91462
rect 117030 91398 117036 91462
rect 116824 91326 117036 91398
rect 116824 91262 116966 91326
rect 117030 91262 117036 91326
rect 116824 91256 117036 91262
rect 1768 90984 1980 91072
rect 28560 91060 28636 91120
rect 110432 91060 110508 91120
rect 136816 91190 137572 91196
rect 136816 91128 137502 91190
rect 136816 91072 136944 91128
rect 137000 91126 137502 91128
rect 137566 91126 137572 91190
rect 137000 91120 137572 91126
rect 137000 91072 137028 91120
rect 21760 91054 21972 91060
rect 21760 90990 21902 91054
rect 21966 90990 21972 91054
rect 21760 90918 21972 90990
rect 21760 90854 21766 90918
rect 21830 90854 21972 90918
rect 21760 90848 21972 90854
rect 22168 91054 22380 91060
rect 22168 90990 22174 91054
rect 22238 90990 22380 91054
rect 22168 90918 22380 90990
rect 22168 90854 22174 90918
rect 22238 90854 22380 90918
rect 22168 90848 22380 90854
rect 22576 91054 22788 91060
rect 22576 90990 22718 91054
rect 22782 90990 22788 91054
rect 22576 90918 22788 90990
rect 22576 90854 22582 90918
rect 22646 90854 22788 90918
rect 22576 90848 22788 90854
rect 22984 91054 23196 91060
rect 22984 90990 22990 91054
rect 23054 90990 23196 91054
rect 22984 90918 23196 90990
rect 22984 90854 22990 90918
rect 23054 90854 23196 90918
rect 22984 90848 23196 90854
rect 23392 91054 23604 91060
rect 23392 90990 23398 91054
rect 23462 90990 23604 91054
rect 23392 90918 23604 90990
rect 23392 90854 23534 90918
rect 23598 90854 23604 90918
rect 23392 90848 23604 90854
rect 28288 90848 28636 91060
rect 110160 90848 110508 91060
rect 115192 91054 115404 91060
rect 115192 90990 115198 91054
rect 115262 90990 115404 91054
rect 115192 90918 115404 90990
rect 115192 90854 115334 90918
rect 115398 90854 115404 90918
rect 115192 90848 115404 90854
rect 115600 91054 115812 91060
rect 115600 90990 115606 91054
rect 115670 90990 115812 91054
rect 115600 90918 115812 90990
rect 115600 90854 115742 90918
rect 115806 90854 115812 90918
rect 115600 90848 115812 90854
rect 116008 91054 116220 91060
rect 116008 90990 116150 91054
rect 116214 90990 116220 91054
rect 116008 90924 116220 90990
rect 116416 90924 116628 91060
rect 116008 90918 116628 90924
rect 116008 90854 116422 90918
rect 116486 90854 116628 90918
rect 116008 90848 116628 90854
rect 116824 91054 117036 91060
rect 116824 90990 116966 91054
rect 117030 90990 117036 91054
rect 116824 90918 117036 90990
rect 136816 90984 137028 91072
rect 116824 90854 116830 90918
rect 116894 90854 117036 90918
rect 116824 90848 117036 90854
rect 28560 90788 28636 90848
rect 110296 90788 110372 90848
rect 21760 90646 21972 90652
rect 21760 90582 21766 90646
rect 21830 90582 21972 90646
rect 21760 90440 21972 90582
rect 22168 90646 22380 90652
rect 22168 90582 22174 90646
rect 22238 90582 22380 90646
rect 22168 90440 22380 90582
rect 22576 90646 22788 90652
rect 22576 90582 22582 90646
rect 22646 90582 22788 90646
rect 22576 90516 22788 90582
rect 22478 90510 22788 90516
rect 22440 90446 22446 90510
rect 22510 90446 22788 90510
rect 22478 90440 22788 90446
rect 22984 90646 23196 90652
rect 22984 90582 22990 90646
rect 23054 90582 23196 90646
rect 22984 90510 23196 90582
rect 22984 90446 23126 90510
rect 23190 90446 23196 90510
rect 22984 90440 23196 90446
rect 23392 90646 23604 90652
rect 23392 90582 23534 90646
rect 23598 90582 23604 90646
rect 23392 90510 23604 90582
rect 28288 90576 28636 90788
rect 110160 90576 110508 90788
rect 115192 90646 115404 90652
rect 115192 90582 115334 90646
rect 115398 90582 115404 90646
rect 28424 90516 28500 90576
rect 110296 90516 110372 90576
rect 23392 90446 23534 90510
rect 23598 90446 23604 90510
rect 23392 90440 23604 90446
rect 21896 90380 21972 90440
rect 21760 90102 21972 90380
rect 28288 90304 28636 90516
rect 110160 90304 110508 90516
rect 115192 90510 115404 90582
rect 115192 90446 115334 90510
rect 115398 90446 115404 90510
rect 115192 90440 115404 90446
rect 115600 90646 115812 90652
rect 115600 90582 115742 90646
rect 115806 90582 115812 90646
rect 115600 90510 115812 90582
rect 115600 90446 115742 90510
rect 115806 90446 115812 90510
rect 115600 90440 115812 90446
rect 116008 90510 116220 90652
rect 116416 90646 116628 90652
rect 116416 90582 116422 90646
rect 116486 90582 116628 90646
rect 116416 90516 116628 90582
rect 116318 90510 116628 90516
rect 116008 90446 116150 90510
rect 116214 90446 116220 90510
rect 116280 90446 116286 90510
rect 116350 90446 116628 90510
rect 116008 90440 116220 90446
rect 116318 90440 116628 90446
rect 116824 90646 117036 90652
rect 116824 90582 116830 90646
rect 116894 90582 117036 90646
rect 116824 90440 117036 90582
rect 116824 90380 116900 90440
rect 116144 90304 116492 90380
rect 28560 90244 28636 90304
rect 110296 90244 110372 90304
rect 116144 90244 116220 90304
rect 116416 90244 116492 90304
rect 21760 90038 21766 90102
rect 21830 90038 21972 90102
rect 21760 90032 21972 90038
rect 22168 90238 22516 90244
rect 22168 90174 22446 90238
rect 22510 90174 22516 90238
rect 22168 90168 22516 90174
rect 22168 90108 22380 90168
rect 22576 90108 22788 90244
rect 22168 90102 22788 90108
rect 22168 90038 22174 90102
rect 22238 90038 22788 90102
rect 22168 90032 22788 90038
rect 22984 90238 23196 90244
rect 22984 90174 23126 90238
rect 23190 90174 23196 90238
rect 22984 90102 23196 90174
rect 22984 90038 22990 90102
rect 23054 90038 23196 90102
rect 22984 90032 23196 90038
rect 23392 90238 23604 90244
rect 23392 90174 23534 90238
rect 23598 90174 23604 90238
rect 23392 90102 23604 90174
rect 23392 90038 23534 90102
rect 23598 90038 23604 90102
rect 23392 90032 23604 90038
rect 28288 90032 28636 90244
rect 110160 90032 110508 90244
rect 115192 90238 115404 90244
rect 115192 90174 115334 90238
rect 115398 90174 115404 90238
rect 115192 90102 115404 90174
rect 115192 90038 115198 90102
rect 115262 90038 115404 90102
rect 115192 90032 115404 90038
rect 115600 90238 115812 90244
rect 115600 90174 115742 90238
rect 115806 90174 115812 90238
rect 115600 90102 115812 90174
rect 115600 90038 115742 90102
rect 115806 90038 115812 90102
rect 115600 90032 115812 90038
rect 116008 90238 116356 90244
rect 116008 90174 116150 90238
rect 116214 90174 116286 90238
rect 116350 90174 116356 90238
rect 116008 90168 116356 90174
rect 116008 90108 116220 90168
rect 116008 90102 116356 90108
rect 116008 90038 116014 90102
rect 116078 90038 116286 90102
rect 116350 90038 116356 90102
rect 116008 90032 116356 90038
rect 116416 90032 116628 90244
rect 116824 90102 117036 90380
rect 116824 90038 116830 90102
rect 116894 90038 117036 90102
rect 116824 90032 117036 90038
rect 28424 89972 28500 90032
rect 110160 89972 110236 90032
rect 21760 89830 21972 89836
rect 21760 89766 21766 89830
rect 21830 89766 21972 89830
rect 21760 89624 21972 89766
rect 22168 89830 22380 89836
rect 22168 89766 22174 89830
rect 22238 89766 22380 89830
rect 22168 89700 22380 89766
rect 22576 89700 22788 89836
rect 22168 89694 22788 89700
rect 22168 89630 22582 89694
rect 22646 89630 22788 89694
rect 22168 89624 22788 89630
rect 22984 89830 23196 89836
rect 22984 89766 22990 89830
rect 23054 89766 23196 89830
rect 22984 89694 23196 89766
rect 22984 89630 22990 89694
rect 23054 89630 23196 89694
rect 22984 89624 23196 89630
rect 23392 89830 23604 89836
rect 23392 89766 23534 89830
rect 23598 89766 23604 89830
rect 23392 89694 23604 89766
rect 28288 89760 28636 89972
rect 110160 89760 110508 89972
rect 28424 89700 28500 89760
rect 110432 89700 110508 89760
rect 23392 89630 23534 89694
rect 23598 89630 23604 89694
rect 23392 89624 23604 89630
rect 21760 89564 21836 89624
rect 1224 89558 1980 89564
rect 1224 89494 1230 89558
rect 1294 89494 1980 89558
rect 1224 89488 1980 89494
rect 1768 89448 1980 89488
rect 1768 89392 1798 89448
rect 1854 89392 1980 89448
rect 1768 89352 1980 89392
rect 21760 89422 21972 89564
rect 28288 89558 28636 89700
rect 28288 89494 28294 89558
rect 28358 89494 28636 89558
rect 28288 89488 28636 89494
rect 110160 89488 110508 89700
rect 115192 89830 115404 89836
rect 115192 89766 115198 89830
rect 115262 89766 115404 89830
rect 115192 89694 115404 89766
rect 115192 89630 115198 89694
rect 115262 89630 115404 89694
rect 115192 89624 115404 89630
rect 115600 89830 115812 89836
rect 115600 89766 115742 89830
rect 115806 89766 115812 89830
rect 115600 89694 115812 89766
rect 115600 89630 115742 89694
rect 115806 89630 115812 89694
rect 115600 89624 115812 89630
rect 116008 89830 116220 89836
rect 116318 89830 116628 89836
rect 116008 89766 116014 89830
rect 116078 89766 116220 89830
rect 116280 89766 116286 89830
rect 116350 89766 116628 89830
rect 116008 89624 116220 89766
rect 116318 89760 116628 89766
rect 116416 89624 116628 89760
rect 116824 89830 117036 89836
rect 116824 89766 116830 89830
rect 116894 89766 117036 89830
rect 116824 89624 117036 89766
rect 116416 89564 116492 89624
rect 116144 89488 116492 89564
rect 116824 89564 116900 89624
rect 28288 89428 28364 89488
rect 110296 89428 110372 89488
rect 116144 89428 116220 89488
rect 21760 89358 21766 89422
rect 21830 89358 21972 89422
rect 21760 89352 21972 89358
rect 22168 89216 22380 89428
rect 22576 89422 22788 89428
rect 22576 89358 22582 89422
rect 22646 89358 22788 89422
rect 22576 89292 22788 89358
rect 22478 89286 22788 89292
rect 22440 89222 22446 89286
rect 22510 89222 22788 89286
rect 22478 89216 22788 89222
rect 22984 89422 23196 89428
rect 22984 89358 22990 89422
rect 23054 89358 23196 89422
rect 22984 89216 23196 89358
rect 23392 89422 23604 89428
rect 23392 89358 23534 89422
rect 23598 89358 23604 89422
rect 23392 89216 23604 89358
rect 28288 89286 28636 89428
rect 28288 89222 28294 89286
rect 28358 89222 28636 89286
rect 28288 89216 28636 89222
rect 110160 89216 110508 89428
rect 115192 89422 115404 89428
rect 115192 89358 115198 89422
rect 115262 89358 115404 89422
rect 115192 89216 115404 89358
rect 115600 89422 115812 89428
rect 115600 89358 115742 89422
rect 115806 89358 115812 89422
rect 115600 89216 115812 89358
rect 116008 89352 116628 89428
rect 116824 89422 117036 89564
rect 116824 89358 116966 89422
rect 117030 89358 117036 89422
rect 116824 89352 117036 89358
rect 136816 89558 137572 89564
rect 136816 89494 137502 89558
rect 137566 89494 137572 89558
rect 136816 89488 137572 89494
rect 136816 89448 137028 89488
rect 136816 89392 136944 89448
rect 137000 89392 137028 89448
rect 136816 89352 137028 89392
rect 116008 89216 116220 89352
rect 116416 89216 116628 89352
rect 22304 89156 22380 89216
rect 22984 89156 23060 89216
rect 23392 89156 23468 89216
rect 21760 89150 21972 89156
rect 21760 89086 21766 89150
rect 21830 89086 21972 89150
rect 21760 89014 21972 89086
rect 21760 88950 21902 89014
rect 21966 88950 21972 89014
rect 21760 88944 21972 88950
rect 22168 89080 22788 89156
rect 22168 89020 22380 89080
rect 22168 89014 22516 89020
rect 22168 88950 22174 89014
rect 22238 88950 22446 89014
rect 22510 88950 22516 89014
rect 22168 88944 22516 88950
rect 22576 88944 22788 89080
rect 22984 88808 23196 89156
rect 23392 88808 23604 89156
rect 28406 89020 28504 89216
rect 110294 89020 110392 89216
rect 115192 89156 115268 89216
rect 115600 89156 115676 89216
rect 116008 89156 116084 89216
rect 116552 89156 116628 89216
rect 28288 88944 28636 89020
rect 110160 89014 110508 89020
rect 110160 88950 110166 89014
rect 110230 88950 110508 89014
rect 110160 88944 110508 88950
rect 28424 88884 28500 88944
rect 22984 88748 23060 88808
rect 23392 88748 23468 88808
rect 21760 88742 21972 88748
rect 21760 88678 21902 88742
rect 21966 88678 21972 88742
rect 21760 88606 21972 88678
rect 21760 88542 21766 88606
rect 21830 88542 21972 88606
rect 21760 88536 21972 88542
rect 22168 88606 22380 88612
rect 22168 88542 22174 88606
rect 22238 88542 22380 88606
rect 22168 88400 22380 88542
rect 22576 88476 22788 88612
rect 22440 88400 22788 88476
rect 22984 88400 23196 88748
rect 22168 88340 22244 88400
rect 22440 88340 22516 88400
rect 21760 88334 21972 88340
rect 21760 88270 21766 88334
rect 21830 88270 21972 88334
rect 21760 88198 21972 88270
rect 21760 88134 21902 88198
rect 21966 88134 21972 88198
rect 21760 88128 21972 88134
rect 22168 88264 22516 88340
rect 22576 88340 22652 88400
rect 23120 88340 23196 88400
rect 22168 88128 22380 88264
rect 22576 88198 22788 88340
rect 22576 88134 22718 88198
rect 22782 88134 22788 88198
rect 22576 88128 22788 88134
rect 22984 88198 23196 88340
rect 22984 88134 23126 88198
rect 23190 88134 23196 88198
rect 22984 88128 23196 88134
rect 23392 88400 23604 88748
rect 23392 88340 23468 88400
rect 23392 88198 23604 88340
rect 28288 88264 28636 88884
rect 110160 88742 110508 88884
rect 115192 88808 115404 89156
rect 115600 88808 115812 89156
rect 116008 88944 116220 89156
rect 116416 89014 116628 89156
rect 116416 88950 116558 89014
rect 116622 88950 116628 89014
rect 116416 88944 116628 88950
rect 116824 89150 117036 89156
rect 116824 89086 116966 89150
rect 117030 89086 117036 89150
rect 116824 89014 117036 89086
rect 116824 88950 116830 89014
rect 116894 88950 117036 89014
rect 116824 88944 117036 88950
rect 115328 88748 115404 88808
rect 115736 88748 115812 88808
rect 110160 88678 110166 88742
rect 110230 88678 110302 88742
rect 110366 88678 110508 88742
rect 110160 88470 110508 88678
rect 110160 88406 110302 88470
rect 110366 88406 110438 88470
rect 110502 88406 110508 88470
rect 110160 88264 110508 88406
rect 115192 88400 115404 88748
rect 115600 88400 115812 88748
rect 116824 88742 117036 88748
rect 116824 88678 116830 88742
rect 116894 88678 117036 88742
rect 116008 88400 116220 88612
rect 116416 88606 116628 88612
rect 116416 88542 116558 88606
rect 116622 88542 116628 88606
rect 116416 88476 116628 88542
rect 116824 88606 117036 88678
rect 116824 88542 116830 88606
rect 116894 88542 117036 88606
rect 116824 88536 117036 88542
rect 116318 88470 116628 88476
rect 116280 88406 116286 88470
rect 116350 88406 116628 88470
rect 116318 88400 116628 88406
rect 115328 88340 115404 88400
rect 115736 88340 115812 88400
rect 116144 88340 116220 88400
rect 28424 88204 28500 88264
rect 110432 88204 110508 88264
rect 23392 88134 23398 88198
rect 23462 88134 23604 88198
rect 23392 88128 23604 88134
rect 21760 87926 21972 87932
rect 21760 87862 21902 87926
rect 21966 87862 21972 87926
rect 1768 87768 1980 87796
rect 1768 87712 1798 87768
rect 1854 87712 1980 87768
rect 21760 87790 21972 87862
rect 21760 87726 21766 87790
rect 21830 87726 21972 87790
rect 21760 87720 21972 87726
rect 22168 87796 22380 87932
rect 22576 87926 22788 87932
rect 22576 87862 22718 87926
rect 22782 87862 22788 87926
rect 22576 87796 22788 87862
rect 22168 87720 22788 87796
rect 22984 87926 23196 87932
rect 22984 87862 23126 87926
rect 23190 87862 23196 87926
rect 22984 87790 23196 87862
rect 22984 87726 23126 87790
rect 23190 87726 23196 87790
rect 22984 87720 23196 87726
rect 23392 87926 23604 87932
rect 23392 87862 23398 87926
rect 23462 87862 23604 87926
rect 23392 87790 23604 87862
rect 23392 87726 23534 87790
rect 23598 87726 23604 87790
rect 23392 87720 23604 87726
rect 28288 87926 28636 88204
rect 28288 87862 28294 87926
rect 28358 87862 28636 87926
rect 28288 87720 28636 87862
rect 110160 88198 110508 88204
rect 110160 88134 110438 88198
rect 110502 88134 110508 88198
rect 110160 87720 110508 88134
rect 115192 88198 115404 88340
rect 115192 88134 115198 88198
rect 115262 88134 115404 88198
rect 115192 88128 115404 88134
rect 115600 88198 115812 88340
rect 115600 88134 115606 88198
rect 115670 88134 115812 88198
rect 115600 88128 115812 88134
rect 116008 88264 116628 88340
rect 116008 88204 116220 88264
rect 116008 88198 116356 88204
rect 116008 88134 116286 88198
rect 116350 88134 116356 88198
rect 116008 88128 116356 88134
rect 116416 88198 116628 88264
rect 116416 88134 116558 88198
rect 116622 88134 116628 88198
rect 116416 88128 116628 88134
rect 116824 88334 117036 88340
rect 116824 88270 116830 88334
rect 116894 88270 117036 88334
rect 116824 88198 117036 88270
rect 116824 88134 116966 88198
rect 117030 88134 117036 88198
rect 116824 88128 117036 88134
rect 115192 87926 115404 87932
rect 115192 87862 115198 87926
rect 115262 87862 115404 87926
rect 115192 87790 115404 87862
rect 115192 87726 115334 87790
rect 115398 87726 115404 87790
rect 115192 87720 115404 87726
rect 115600 87926 115812 87932
rect 115600 87862 115606 87926
rect 115670 87862 115812 87926
rect 115600 87790 115812 87862
rect 115600 87726 115742 87790
rect 115806 87726 115812 87790
rect 115600 87720 115812 87726
rect 116008 87790 116220 87932
rect 116416 87926 116628 87932
rect 116416 87862 116558 87926
rect 116622 87862 116628 87926
rect 116416 87796 116628 87862
rect 116318 87790 116628 87796
rect 116008 87726 116150 87790
rect 116214 87726 116220 87790
rect 116280 87726 116286 87790
rect 116350 87726 116422 87790
rect 116486 87726 116628 87790
rect 116008 87720 116220 87726
rect 116318 87720 116628 87726
rect 116824 87926 117036 87932
rect 116824 87862 116966 87926
rect 117030 87862 117036 87926
rect 116824 87790 117036 87862
rect 116824 87726 116966 87790
rect 117030 87726 117036 87790
rect 116824 87720 117036 87726
rect 136816 87790 137572 87796
rect 136816 87768 137502 87790
rect 1768 87660 1980 87712
rect 1224 87654 1980 87660
rect 1224 87590 1230 87654
rect 1294 87590 1980 87654
rect 1224 87584 1980 87590
rect 22304 87660 22380 87720
rect 28288 87660 28364 87720
rect 110296 87660 110372 87720
rect 136816 87712 136944 87768
rect 137000 87726 137502 87768
rect 137566 87726 137572 87790
rect 137000 87720 137572 87726
rect 137000 87712 137028 87720
rect 22304 87584 22652 87660
rect 22576 87524 22652 87584
rect 28288 87654 28636 87660
rect 28288 87590 28294 87654
rect 28358 87590 28636 87654
rect 21760 87518 21972 87524
rect 21760 87454 21766 87518
rect 21830 87454 21972 87518
rect 21760 87382 21972 87454
rect 21760 87318 21766 87382
rect 21830 87318 21972 87382
rect 21760 87312 21972 87318
rect 22168 87382 22380 87524
rect 22168 87318 22174 87382
rect 22238 87318 22380 87382
rect 22168 87312 22380 87318
rect 22576 87382 22788 87524
rect 22576 87318 22582 87382
rect 22646 87318 22788 87382
rect 22576 87312 22788 87318
rect 22984 87518 23196 87524
rect 22984 87454 23126 87518
rect 23190 87454 23196 87518
rect 22984 87382 23196 87454
rect 22984 87318 22990 87382
rect 23054 87318 23196 87382
rect 22984 87312 23196 87318
rect 23392 87518 23604 87524
rect 23392 87454 23534 87518
rect 23598 87454 23604 87518
rect 23392 87382 23604 87454
rect 23392 87318 23534 87382
rect 23598 87318 23604 87382
rect 23392 87312 23604 87318
rect 28288 87448 28636 87590
rect 110160 87448 110508 87660
rect 136816 87584 137028 87712
rect 28288 87388 28364 87448
rect 110432 87388 110508 87448
rect 28288 87176 28636 87388
rect 110160 87176 110508 87388
rect 115192 87518 115404 87524
rect 115192 87454 115334 87518
rect 115398 87454 115404 87518
rect 115192 87382 115404 87454
rect 115192 87318 115198 87382
rect 115262 87318 115404 87382
rect 115192 87312 115404 87318
rect 115600 87518 115812 87524
rect 115600 87454 115742 87518
rect 115806 87454 115812 87518
rect 115600 87382 115812 87454
rect 115600 87318 115742 87382
rect 115806 87318 115812 87382
rect 115600 87312 115812 87318
rect 116008 87518 116356 87524
rect 116008 87454 116150 87518
rect 116214 87454 116286 87518
rect 116350 87454 116356 87518
rect 116008 87448 116356 87454
rect 116416 87518 116628 87524
rect 116416 87454 116422 87518
rect 116486 87454 116628 87518
rect 116008 87388 116220 87448
rect 116008 87382 116356 87388
rect 116008 87318 116014 87382
rect 116078 87318 116286 87382
rect 116350 87318 116356 87382
rect 116008 87312 116356 87318
rect 116416 87312 116628 87454
rect 116824 87518 117036 87524
rect 116824 87454 116966 87518
rect 117030 87454 117036 87518
rect 116824 87382 117036 87454
rect 116824 87318 116966 87382
rect 117030 87318 117036 87382
rect 116824 87312 117036 87318
rect 28424 87116 28500 87176
rect 110432 87116 110508 87176
rect 21760 87110 21972 87116
rect 21760 87046 21766 87110
rect 21830 87046 21972 87110
rect 21760 86974 21972 87046
rect 21760 86910 21902 86974
rect 21966 86910 21972 86974
rect 21760 86904 21972 86910
rect 22168 87110 22788 87116
rect 22168 87046 22174 87110
rect 22238 87046 22582 87110
rect 22646 87046 22788 87110
rect 22168 87040 22788 87046
rect 22168 86980 22380 87040
rect 22168 86904 22516 86980
rect 22576 86904 22788 87040
rect 22984 87110 23196 87116
rect 22984 87046 22990 87110
rect 23054 87046 23196 87110
rect 22984 86974 23196 87046
rect 22984 86910 23126 86974
rect 23190 86910 23196 86974
rect 22984 86904 23196 86910
rect 23392 87110 23604 87116
rect 23392 87046 23534 87110
rect 23598 87046 23604 87110
rect 23392 86974 23604 87046
rect 23392 86910 23398 86974
rect 23462 86910 23604 86974
rect 23392 86904 23604 86910
rect 28288 86904 28636 87116
rect 110160 86904 110508 87116
rect 115192 87110 115404 87116
rect 115192 87046 115198 87110
rect 115262 87046 115404 87110
rect 115192 86974 115404 87046
rect 115192 86910 115198 86974
rect 115262 86910 115404 86974
rect 115192 86904 115404 86910
rect 115600 87110 115812 87116
rect 115600 87046 115742 87110
rect 115806 87046 115812 87110
rect 115600 86974 115812 87046
rect 115600 86910 115606 86974
rect 115670 86910 115812 86974
rect 115600 86904 115812 86910
rect 116008 87110 116220 87116
rect 116318 87110 116628 87116
rect 116008 87046 116014 87110
rect 116078 87046 116220 87110
rect 116280 87046 116286 87110
rect 116350 87046 116628 87110
rect 116008 86974 116220 87046
rect 116318 87040 116628 87046
rect 116008 86910 116150 86974
rect 116214 86910 116220 86974
rect 116008 86904 116220 86910
rect 116416 86904 116628 87040
rect 116824 87110 117036 87116
rect 116824 87046 116966 87110
rect 117030 87046 117036 87110
rect 116824 86974 117036 87046
rect 116824 86910 116966 86974
rect 117030 86910 117036 86974
rect 116824 86904 117036 86910
rect 22440 86844 22516 86904
rect 28288 86844 28364 86904
rect 110432 86844 110508 86904
rect 22440 86768 22652 86844
rect 22576 86708 22652 86768
rect 21760 86702 21972 86708
rect 21760 86638 21902 86702
rect 21966 86638 21972 86702
rect 21760 86566 21972 86638
rect 21760 86502 21766 86566
rect 21830 86502 21972 86566
rect 21760 86496 21972 86502
rect 22168 86632 22788 86708
rect 22168 86572 22380 86632
rect 22168 86566 22516 86572
rect 22168 86502 22446 86566
rect 22510 86502 22516 86566
rect 22168 86496 22516 86502
rect 22576 86496 22788 86632
rect 22984 86702 23196 86708
rect 22984 86638 23126 86702
rect 23190 86638 23196 86702
rect 22984 86566 23196 86638
rect 22984 86502 22990 86566
rect 23054 86502 23196 86566
rect 22984 86496 23196 86502
rect 23392 86702 23604 86708
rect 23392 86638 23398 86702
rect 23462 86638 23604 86702
rect 23392 86566 23604 86638
rect 23392 86502 23534 86566
rect 23598 86502 23604 86566
rect 23392 86496 23604 86502
rect 28288 86632 28636 86844
rect 110160 86632 110508 86844
rect 115192 86702 115404 86708
rect 115192 86638 115198 86702
rect 115262 86638 115404 86702
rect 28288 86572 28364 86632
rect 110296 86572 110372 86632
rect 28288 86360 28636 86572
rect 110160 86360 110508 86572
rect 115192 86566 115404 86638
rect 115192 86502 115334 86566
rect 115398 86502 115404 86566
rect 115192 86496 115404 86502
rect 115600 86702 115812 86708
rect 115600 86638 115606 86702
rect 115670 86638 115812 86702
rect 115600 86566 115812 86638
rect 115600 86502 115742 86566
rect 115806 86502 115812 86566
rect 115600 86496 115812 86502
rect 116008 86702 116220 86708
rect 116008 86638 116150 86702
rect 116214 86638 116220 86702
rect 116008 86566 116220 86638
rect 116008 86502 116014 86566
rect 116078 86502 116220 86566
rect 116008 86496 116220 86502
rect 116416 86566 116628 86708
rect 116416 86502 116422 86566
rect 116486 86502 116628 86566
rect 116416 86496 116628 86502
rect 116824 86702 117036 86708
rect 116824 86638 116966 86702
rect 117030 86638 117036 86702
rect 116824 86566 117036 86638
rect 116824 86502 116830 86566
rect 116894 86502 117036 86566
rect 116824 86496 117036 86502
rect 28560 86300 28636 86360
rect 110296 86300 110372 86360
rect 21760 86294 21972 86300
rect 21760 86230 21766 86294
rect 21830 86230 21972 86294
rect 1224 86158 1980 86164
rect 1224 86094 1230 86158
rect 1294 86094 1980 86158
rect 1224 86088 1980 86094
rect 21760 86158 21972 86230
rect 21760 86094 21766 86158
rect 21830 86094 21972 86158
rect 21760 86088 21972 86094
rect 22168 86158 22380 86300
rect 22478 86294 22788 86300
rect 22440 86230 22446 86294
rect 22510 86230 22788 86294
rect 22478 86224 22788 86230
rect 22168 86094 22310 86158
rect 22374 86094 22380 86158
rect 22168 86088 22380 86094
rect 22576 86088 22788 86224
rect 22984 86294 23196 86300
rect 22984 86230 22990 86294
rect 23054 86230 23196 86294
rect 22984 86158 23196 86230
rect 22984 86094 22990 86158
rect 23054 86094 23196 86158
rect 22984 86088 23196 86094
rect 23392 86294 23604 86300
rect 23392 86230 23534 86294
rect 23598 86230 23604 86294
rect 23392 86158 23604 86230
rect 23392 86094 23534 86158
rect 23598 86094 23604 86158
rect 23392 86088 23604 86094
rect 28288 86088 28636 86300
rect 1768 86032 1798 86088
rect 1854 86032 1980 86088
rect 1768 85952 1980 86032
rect 22576 86028 22652 86088
rect 28560 86028 28636 86088
rect 22304 85952 22652 86028
rect 22304 85892 22380 85952
rect 21760 85886 21972 85892
rect 21760 85822 21766 85886
rect 21830 85822 21972 85886
rect 21760 85680 21972 85822
rect 22168 85886 22788 85892
rect 22168 85822 22310 85886
rect 22374 85822 22788 85886
rect 22168 85816 22788 85822
rect 22168 85680 22380 85816
rect 22576 85756 22788 85816
rect 22478 85750 22788 85756
rect 22440 85686 22446 85750
rect 22510 85686 22718 85750
rect 22782 85686 22788 85750
rect 22478 85680 22788 85686
rect 22984 85886 23196 85892
rect 22984 85822 22990 85886
rect 23054 85822 23196 85886
rect 22984 85750 23196 85822
rect 22984 85686 22990 85750
rect 23054 85686 23196 85750
rect 22984 85680 23196 85686
rect 23392 85886 23604 85892
rect 23392 85822 23534 85886
rect 23598 85822 23604 85886
rect 23392 85750 23604 85822
rect 28288 85816 28636 86028
rect 110160 86088 110508 86300
rect 115192 86294 115404 86300
rect 115192 86230 115334 86294
rect 115398 86230 115404 86294
rect 115192 86158 115404 86230
rect 115192 86094 115334 86158
rect 115398 86094 115404 86158
rect 115192 86088 115404 86094
rect 115600 86294 115812 86300
rect 115600 86230 115742 86294
rect 115806 86230 115812 86294
rect 115600 86158 115812 86230
rect 115600 86094 115606 86158
rect 115670 86094 115812 86158
rect 115600 86088 115812 86094
rect 116008 86294 116220 86300
rect 116008 86230 116014 86294
rect 116078 86230 116220 86294
rect 116008 86164 116220 86230
rect 116416 86294 116628 86300
rect 116416 86230 116422 86294
rect 116486 86230 116628 86294
rect 116416 86164 116628 86230
rect 116008 86088 116628 86164
rect 116824 86294 117036 86300
rect 116824 86230 116830 86294
rect 116894 86230 117036 86294
rect 116824 86158 117036 86230
rect 116824 86094 116830 86158
rect 116894 86094 117036 86158
rect 116824 86088 117036 86094
rect 136816 86088 137028 86164
rect 110160 86028 110236 86088
rect 116144 86028 116220 86088
rect 136816 86032 136944 86088
rect 137000 86032 137028 86088
rect 136816 86028 137028 86032
rect 110160 85816 110508 86028
rect 116144 85952 116492 86028
rect 136816 86022 137572 86028
rect 136816 85958 137502 86022
rect 137566 85958 137572 86022
rect 136816 85952 137572 85958
rect 116416 85892 116492 85952
rect 28560 85756 28636 85816
rect 110432 85756 110508 85816
rect 23392 85686 23534 85750
rect 23598 85686 23604 85750
rect 23392 85680 23604 85686
rect 21896 85620 21972 85680
rect 21760 85478 21972 85620
rect 28288 85544 28636 85756
rect 110160 85614 110508 85756
rect 115192 85886 115404 85892
rect 115192 85822 115334 85886
rect 115398 85822 115404 85886
rect 115192 85750 115404 85822
rect 115192 85686 115334 85750
rect 115398 85686 115404 85750
rect 115192 85680 115404 85686
rect 115600 85886 115812 85892
rect 115600 85822 115606 85886
rect 115670 85822 115812 85886
rect 115600 85750 115812 85822
rect 115600 85686 115606 85750
rect 115670 85686 115812 85750
rect 115600 85680 115812 85686
rect 116008 85756 116220 85892
rect 116416 85756 116628 85892
rect 116008 85750 116628 85756
rect 116008 85686 116014 85750
rect 116078 85686 116628 85750
rect 116008 85680 116628 85686
rect 116824 85886 117036 85892
rect 116824 85822 116830 85886
rect 116894 85822 117036 85886
rect 116824 85680 117036 85822
rect 110160 85550 110166 85614
rect 110230 85550 110508 85614
rect 110160 85544 110508 85550
rect 116824 85620 116900 85680
rect 28424 85484 28500 85544
rect 110160 85484 110236 85544
rect 21760 85414 21766 85478
rect 21830 85414 21972 85478
rect 21760 85408 21972 85414
rect 22168 85478 22516 85484
rect 22168 85414 22446 85478
rect 22510 85414 22516 85478
rect 22168 85408 22516 85414
rect 22576 85478 22788 85484
rect 22576 85414 22718 85478
rect 22782 85414 22788 85478
rect 22168 85272 22380 85408
rect 22576 85272 22788 85414
rect 22984 85478 23196 85484
rect 22984 85414 22990 85478
rect 23054 85414 23196 85478
rect 22984 85342 23196 85414
rect 22984 85278 22990 85342
rect 23054 85278 23196 85342
rect 22984 85272 23196 85278
rect 23392 85478 23604 85484
rect 23392 85414 23534 85478
rect 23598 85414 23604 85478
rect 23392 85342 23604 85414
rect 23392 85278 23534 85342
rect 23598 85278 23604 85342
rect 23392 85272 23604 85278
rect 22168 85212 22244 85272
rect 22576 85212 22652 85272
rect 21760 85206 21972 85212
rect 21760 85142 21766 85206
rect 21830 85142 21972 85206
rect 21760 84864 21972 85142
rect 22168 84864 22380 85212
rect 22576 84934 22788 85212
rect 22576 84870 22718 84934
rect 22782 84870 22788 84934
rect 22576 84864 22788 84870
rect 22984 85070 23196 85076
rect 22984 85006 22990 85070
rect 23054 85006 23196 85070
rect 22984 84864 23196 85006
rect 23392 85070 23604 85076
rect 23392 85006 23534 85070
rect 23598 85006 23604 85070
rect 23392 84864 23604 85006
rect 28288 85000 28636 85484
rect 110160 85342 110508 85484
rect 110160 85278 110166 85342
rect 110230 85278 110508 85342
rect 110160 85000 110508 85278
rect 115192 85478 115404 85484
rect 115192 85414 115334 85478
rect 115398 85414 115404 85478
rect 115192 85342 115404 85414
rect 115192 85278 115334 85342
rect 115398 85278 115404 85342
rect 115192 85272 115404 85278
rect 115600 85478 115812 85484
rect 115600 85414 115606 85478
rect 115670 85414 115812 85478
rect 115600 85342 115812 85414
rect 115600 85278 115742 85342
rect 115806 85278 115812 85342
rect 115600 85272 115812 85278
rect 116008 85478 116220 85484
rect 116008 85414 116014 85478
rect 116078 85414 116220 85478
rect 116008 85272 116220 85414
rect 116416 85348 116628 85484
rect 116824 85478 117036 85620
rect 116824 85414 116966 85478
rect 117030 85414 117036 85478
rect 116824 85408 117036 85414
rect 116280 85272 116628 85348
rect 116008 85212 116084 85272
rect 116280 85212 116356 85272
rect 116008 85136 116356 85212
rect 116416 85212 116492 85272
rect 28288 84940 28364 85000
rect 110432 84940 110508 85000
rect 21896 84804 21972 84864
rect 21760 84662 21972 84804
rect 22984 84804 23060 84864
rect 23392 84804 23468 84864
rect 21760 84598 21902 84662
rect 21966 84598 21972 84662
rect 21760 84592 21972 84598
rect 22168 84662 22788 84668
rect 22168 84598 22718 84662
rect 22782 84598 22788 84662
rect 22168 84592 22788 84598
rect 22168 84532 22380 84592
rect 1768 84408 1980 84532
rect 1768 84396 1798 84408
rect 1224 84390 1798 84396
rect 1224 84326 1230 84390
rect 1294 84352 1798 84390
rect 1854 84352 1980 84408
rect 22168 84456 22516 84532
rect 22576 84456 22788 84592
rect 22984 84456 23196 84804
rect 23392 84456 23604 84804
rect 28288 84798 28636 84940
rect 28288 84734 28566 84798
rect 28630 84734 28636 84798
rect 28288 84526 28636 84734
rect 28288 84462 28566 84526
rect 28630 84462 28636 84526
rect 22168 84396 22244 84456
rect 22440 84396 22516 84456
rect 22984 84396 23060 84456
rect 23392 84396 23468 84456
rect 1294 84326 1980 84352
rect 1224 84320 1980 84326
rect 21760 84390 21972 84396
rect 21760 84326 21902 84390
rect 21966 84326 21972 84390
rect 21760 84254 21972 84326
rect 21760 84190 21766 84254
rect 21830 84190 21972 84254
rect 21760 84184 21972 84190
rect 22168 84184 22380 84396
rect 22440 84320 22788 84396
rect 22576 84254 22788 84320
rect 22576 84190 22582 84254
rect 22646 84190 22788 84254
rect 22576 84184 22788 84190
rect 22984 84048 23196 84396
rect 23392 84048 23604 84396
rect 28288 84390 28636 84462
rect 28288 84326 28430 84390
rect 28494 84326 28636 84390
rect 28288 84320 28636 84326
rect 110160 84390 110508 84940
rect 110160 84326 110166 84390
rect 110230 84326 110508 84390
rect 110160 84320 110508 84326
rect 115192 85070 115404 85076
rect 115192 85006 115334 85070
rect 115398 85006 115404 85070
rect 115192 84864 115404 85006
rect 115600 85070 115812 85076
rect 115600 85006 115742 85070
rect 115806 85006 115812 85070
rect 115600 84864 115812 85006
rect 116008 84864 116220 85136
rect 116416 84934 116628 85212
rect 116416 84870 116558 84934
rect 116622 84870 116628 84934
rect 116416 84864 116628 84870
rect 116824 85206 117036 85212
rect 116824 85142 116966 85206
rect 117030 85142 117036 85206
rect 116824 84864 117036 85142
rect 115192 84804 115268 84864
rect 115600 84804 115676 84864
rect 116824 84804 116900 84864
rect 115192 84456 115404 84804
rect 115600 84456 115812 84804
rect 116008 84532 116220 84668
rect 116416 84662 116628 84668
rect 116416 84598 116558 84662
rect 116622 84598 116628 84662
rect 116416 84532 116628 84598
rect 116824 84662 117036 84804
rect 116824 84598 116966 84662
rect 117030 84598 117036 84662
rect 116824 84592 117036 84598
rect 116008 84456 116628 84532
rect 115192 84396 115268 84456
rect 115600 84396 115676 84456
rect 116144 84396 116220 84456
rect 116552 84396 116628 84456
rect 136816 84526 137572 84532
rect 136816 84462 137502 84526
rect 137566 84462 137572 84526
rect 136816 84456 137572 84462
rect 136816 84408 137028 84456
rect 23120 83988 23196 84048
rect 23528 83988 23604 84048
rect 21760 83982 21972 83988
rect 21760 83918 21766 83982
rect 21830 83918 21972 83982
rect 21760 83846 21972 83918
rect 21760 83782 21902 83846
rect 21966 83782 21972 83846
rect 21760 83776 21972 83782
rect 22168 83852 22380 83988
rect 22576 83982 22788 83988
rect 22576 83918 22582 83982
rect 22646 83918 22788 83982
rect 22576 83852 22788 83918
rect 22168 83776 22788 83852
rect 22984 83846 23196 83988
rect 22984 83782 23126 83846
rect 23190 83782 23196 83846
rect 22984 83776 23196 83782
rect 23392 83846 23604 83988
rect 23392 83782 23398 83846
rect 23462 83782 23604 83846
rect 23392 83776 23604 83782
rect 28288 84118 28636 84124
rect 28288 84054 28430 84118
rect 28494 84054 28636 84118
rect 28288 83982 28636 84054
rect 28288 83918 28430 83982
rect 28494 83918 28636 83982
rect 28288 83776 28636 83918
rect 110160 84118 110508 84124
rect 110160 84054 110166 84118
rect 110230 84054 110508 84118
rect 110160 83776 110508 84054
rect 115192 84048 115404 84396
rect 115600 84048 115812 84396
rect 116008 84184 116220 84396
rect 116416 84184 116628 84396
rect 116824 84390 117036 84396
rect 116824 84326 116966 84390
rect 117030 84326 117036 84390
rect 116824 84254 117036 84326
rect 136816 84352 136944 84408
rect 137000 84352 137028 84408
rect 136816 84320 137028 84352
rect 116824 84190 116830 84254
rect 116894 84190 117036 84254
rect 116824 84184 117036 84190
rect 116416 84124 116492 84184
rect 115192 83988 115268 84048
rect 115736 83988 115812 84048
rect 116144 84048 116492 84124
rect 116144 83988 116220 84048
rect 115192 83846 115404 83988
rect 115192 83782 115198 83846
rect 115262 83782 115404 83846
rect 115192 83776 115404 83782
rect 115600 83846 115812 83988
rect 115600 83782 115606 83846
rect 115670 83782 115812 83846
rect 115600 83776 115812 83782
rect 116008 83912 116628 83988
rect 22168 83640 22380 83776
rect 22576 83640 22788 83776
rect 28424 83716 28500 83776
rect 110432 83716 110508 83776
rect 22712 83580 22788 83640
rect 28288 83710 28636 83716
rect 28288 83646 28430 83710
rect 28494 83646 28636 83710
rect 21760 83574 21972 83580
rect 21760 83510 21902 83574
rect 21966 83510 21972 83574
rect 21760 83438 21972 83510
rect 21760 83374 21766 83438
rect 21830 83374 21972 83438
rect 21760 83368 21972 83374
rect 22168 83444 22380 83580
rect 22576 83444 22788 83580
rect 22168 83438 22788 83444
rect 22168 83374 22310 83438
rect 22374 83374 22788 83438
rect 22168 83368 22788 83374
rect 22984 83574 23196 83580
rect 22984 83510 23126 83574
rect 23190 83510 23196 83574
rect 22984 83438 23196 83510
rect 22984 83374 22990 83438
rect 23054 83374 23196 83438
rect 22984 83368 23196 83374
rect 23392 83574 23604 83580
rect 23392 83510 23398 83574
rect 23462 83510 23604 83574
rect 23392 83438 23604 83510
rect 28288 83504 28636 83646
rect 110160 83504 110508 83716
rect 116008 83640 116220 83912
rect 116416 83640 116628 83912
rect 116824 83982 117036 83988
rect 116824 83918 116830 83982
rect 116894 83918 117036 83982
rect 116824 83846 117036 83918
rect 116824 83782 116966 83846
rect 117030 83782 117036 83846
rect 116824 83776 117036 83782
rect 116416 83580 116492 83640
rect 115192 83574 115404 83580
rect 115192 83510 115198 83574
rect 115262 83510 115404 83574
rect 28560 83444 28636 83504
rect 110296 83444 110372 83504
rect 23392 83374 23398 83438
rect 23462 83374 23604 83438
rect 23392 83368 23604 83374
rect 28288 83232 28636 83444
rect 110160 83232 110508 83444
rect 115192 83438 115404 83510
rect 115192 83374 115198 83438
rect 115262 83374 115404 83438
rect 115192 83368 115404 83374
rect 115600 83574 115812 83580
rect 115600 83510 115606 83574
rect 115670 83510 115812 83574
rect 115600 83438 115812 83510
rect 115600 83374 115742 83438
rect 115806 83374 115812 83438
rect 115600 83368 115812 83374
rect 116008 83444 116220 83580
rect 116416 83444 116628 83580
rect 116008 83438 116628 83444
rect 116008 83374 116014 83438
rect 116078 83374 116422 83438
rect 116486 83374 116628 83438
rect 116008 83368 116628 83374
rect 116824 83574 117036 83580
rect 116824 83510 116966 83574
rect 117030 83510 117036 83574
rect 116824 83438 117036 83510
rect 116824 83374 116966 83438
rect 117030 83374 117036 83438
rect 116824 83368 117036 83374
rect 28288 83172 28364 83232
rect 110296 83172 110372 83232
rect 21760 83166 21972 83172
rect 21760 83102 21766 83166
rect 21830 83102 21972 83166
rect 21760 83030 21972 83102
rect 21760 82966 21766 83030
rect 21830 82966 21972 83030
rect 21760 82960 21972 82966
rect 22168 83166 22380 83172
rect 22168 83102 22310 83166
rect 22374 83102 22380 83166
rect 22168 83030 22380 83102
rect 22168 82966 22174 83030
rect 22238 82966 22380 83030
rect 22168 82960 22380 82966
rect 22576 83030 22788 83172
rect 22576 82966 22582 83030
rect 22646 82966 22788 83030
rect 22576 82960 22788 82966
rect 22984 83166 23196 83172
rect 22984 83102 22990 83166
rect 23054 83102 23196 83166
rect 22984 83030 23196 83102
rect 22984 82966 22990 83030
rect 23054 82966 23196 83030
rect 22984 82960 23196 82966
rect 23392 83166 23604 83172
rect 23392 83102 23398 83166
rect 23462 83102 23604 83166
rect 23392 83030 23604 83102
rect 23392 82966 23398 83030
rect 23462 82966 23604 83030
rect 23392 82960 23604 82966
rect 28288 82960 28636 83172
rect 110160 82960 110508 83172
rect 115192 83166 115404 83172
rect 115192 83102 115198 83166
rect 115262 83102 115404 83166
rect 115192 83030 115404 83102
rect 115192 82966 115198 83030
rect 115262 82966 115404 83030
rect 115192 82960 115404 82966
rect 115600 83166 115812 83172
rect 115600 83102 115742 83166
rect 115806 83102 115812 83166
rect 115600 83030 115812 83102
rect 115600 82966 115742 83030
rect 115806 82966 115812 83030
rect 115600 82960 115812 82966
rect 116008 83166 116220 83172
rect 116008 83102 116014 83166
rect 116078 83102 116220 83166
rect 116008 83030 116220 83102
rect 116008 82966 116014 83030
rect 116078 82966 116220 83030
rect 116008 82960 116220 82966
rect 116416 83166 116628 83172
rect 116416 83102 116422 83166
rect 116486 83102 116628 83166
rect 116416 82960 116628 83102
rect 116824 83166 117036 83172
rect 116824 83102 116966 83166
rect 117030 83102 117036 83166
rect 116824 83030 117036 83102
rect 116824 82966 116830 83030
rect 116894 82966 117036 83030
rect 116824 82960 117036 82966
rect 28424 82900 28500 82960
rect 110432 82900 110508 82960
rect 1224 82758 1980 82764
rect 1224 82694 1230 82758
rect 1294 82728 1980 82758
rect 1294 82694 1798 82728
rect 1224 82688 1798 82694
rect 1768 82672 1798 82688
rect 1854 82672 1980 82728
rect 1768 82552 1980 82672
rect 21760 82758 21972 82764
rect 21760 82694 21766 82758
rect 21830 82694 21972 82758
rect 21760 82622 21972 82694
rect 21760 82558 21902 82622
rect 21966 82558 21972 82622
rect 21760 82552 21972 82558
rect 22168 82758 22788 82764
rect 22168 82694 22174 82758
rect 22238 82694 22582 82758
rect 22646 82694 22788 82758
rect 22168 82688 22788 82694
rect 22168 82552 22380 82688
rect 22576 82628 22788 82688
rect 22478 82622 22788 82628
rect 22440 82558 22446 82622
rect 22510 82558 22788 82622
rect 22478 82552 22788 82558
rect 22984 82758 23196 82764
rect 22984 82694 22990 82758
rect 23054 82694 23196 82758
rect 22984 82622 23196 82694
rect 22984 82558 23126 82622
rect 23190 82558 23196 82622
rect 22984 82552 23196 82558
rect 23392 82758 23604 82764
rect 23392 82694 23398 82758
rect 23462 82694 23604 82758
rect 23392 82622 23604 82694
rect 28288 82688 28636 82900
rect 110160 82688 110508 82900
rect 115192 82758 115404 82764
rect 115192 82694 115198 82758
rect 115262 82694 115404 82758
rect 28424 82628 28500 82688
rect 110160 82628 110236 82688
rect 23392 82558 23398 82622
rect 23462 82558 23604 82622
rect 23392 82552 23604 82558
rect 22304 82492 22380 82552
rect 22304 82416 22652 82492
rect 22576 82356 22652 82416
rect 28288 82416 28636 82628
rect 110160 82416 110508 82628
rect 115192 82622 115404 82694
rect 115192 82558 115198 82622
rect 115262 82558 115404 82622
rect 115192 82552 115404 82558
rect 115600 82758 115812 82764
rect 115600 82694 115742 82758
rect 115806 82694 115812 82758
rect 115600 82622 115812 82694
rect 115600 82558 115606 82622
rect 115670 82558 115812 82622
rect 115600 82552 115812 82558
rect 116008 82758 116220 82764
rect 116008 82694 116014 82758
rect 116078 82694 116220 82758
rect 116008 82628 116220 82694
rect 116416 82628 116628 82764
rect 116008 82622 116628 82628
rect 116008 82558 116014 82622
rect 116078 82558 116628 82622
rect 116008 82552 116628 82558
rect 116824 82758 117036 82764
rect 116824 82694 116830 82758
rect 116894 82694 117036 82758
rect 116824 82622 117036 82694
rect 116824 82558 116966 82622
rect 117030 82558 117036 82622
rect 116824 82552 117036 82558
rect 136816 82758 137572 82764
rect 136816 82728 137502 82758
rect 136816 82672 136944 82728
rect 137000 82694 137502 82728
rect 137566 82694 137572 82758
rect 137000 82688 137572 82694
rect 137000 82672 137028 82688
rect 136816 82552 137028 82672
rect 28288 82356 28364 82416
rect 110296 82356 110372 82416
rect 21760 82350 21972 82356
rect 21760 82286 21902 82350
rect 21966 82286 21972 82350
rect 21760 82214 21972 82286
rect 21760 82150 21766 82214
rect 21830 82150 21972 82214
rect 21760 82144 21972 82150
rect 22168 82350 22516 82356
rect 22168 82286 22446 82350
rect 22510 82286 22516 82350
rect 22168 82280 22516 82286
rect 22168 82144 22380 82280
rect 22576 82214 22788 82356
rect 22576 82150 22582 82214
rect 22646 82150 22788 82214
rect 22576 82144 22788 82150
rect 22984 82350 23196 82356
rect 22984 82286 23126 82350
rect 23190 82286 23196 82350
rect 22984 82214 23196 82286
rect 22984 82150 23126 82214
rect 23190 82150 23196 82214
rect 22984 82144 23196 82150
rect 23392 82350 23604 82356
rect 23392 82286 23398 82350
rect 23462 82286 23604 82350
rect 23392 82214 23604 82286
rect 23392 82150 23534 82214
rect 23598 82150 23604 82214
rect 23392 82144 23604 82150
rect 28288 82144 28636 82356
rect 28560 82084 28636 82144
rect 21760 81942 21972 81948
rect 21760 81878 21766 81942
rect 21830 81878 21972 81942
rect 21760 81736 21972 81878
rect 22168 81806 22380 81948
rect 22168 81742 22310 81806
rect 22374 81742 22380 81806
rect 22168 81736 22380 81742
rect 22576 81942 22788 81948
rect 22576 81878 22582 81942
rect 22646 81878 22788 81942
rect 22576 81806 22788 81878
rect 22576 81742 22582 81806
rect 22646 81742 22788 81806
rect 22576 81736 22788 81742
rect 22984 81942 23196 81948
rect 22984 81878 23126 81942
rect 23190 81878 23196 81942
rect 22984 81806 23196 81878
rect 22984 81742 23126 81806
rect 23190 81742 23196 81806
rect 22984 81736 23196 81742
rect 23392 81942 23604 81948
rect 23392 81878 23534 81942
rect 23598 81878 23604 81942
rect 23392 81806 23604 81878
rect 28288 81872 28636 82084
rect 110160 82144 110508 82356
rect 115192 82350 115404 82356
rect 115192 82286 115198 82350
rect 115262 82286 115404 82350
rect 115192 82214 115404 82286
rect 115192 82150 115334 82214
rect 115398 82150 115404 82214
rect 115192 82144 115404 82150
rect 115600 82350 115812 82356
rect 115600 82286 115606 82350
rect 115670 82286 115812 82350
rect 115600 82214 115812 82286
rect 115600 82150 115742 82214
rect 115806 82150 115812 82214
rect 115600 82144 115812 82150
rect 116008 82350 116220 82356
rect 116008 82286 116014 82350
rect 116078 82286 116220 82350
rect 116008 82214 116220 82286
rect 116008 82150 116014 82214
rect 116078 82150 116220 82214
rect 116008 82144 116220 82150
rect 116416 82214 116628 82356
rect 116416 82150 116422 82214
rect 116486 82150 116628 82214
rect 116416 82144 116628 82150
rect 116824 82350 117036 82356
rect 116824 82286 116966 82350
rect 117030 82286 117036 82350
rect 116824 82214 117036 82286
rect 116824 82150 116830 82214
rect 116894 82150 117036 82214
rect 116824 82144 117036 82150
rect 110160 82084 110236 82144
rect 110160 81872 110508 82084
rect 115192 81942 115404 81948
rect 115192 81878 115334 81942
rect 115398 81878 115404 81942
rect 28424 81812 28500 81872
rect 110296 81812 110372 81872
rect 23392 81742 23534 81806
rect 23598 81742 23604 81806
rect 23392 81736 23604 81742
rect 21896 81676 21972 81736
rect 21760 81328 21972 81676
rect 28288 81600 28636 81812
rect 110160 81600 110508 81812
rect 115192 81806 115404 81878
rect 115192 81742 115198 81806
rect 115262 81742 115404 81806
rect 115192 81736 115404 81742
rect 115600 81942 115812 81948
rect 115600 81878 115742 81942
rect 115806 81878 115812 81942
rect 115600 81806 115812 81878
rect 115600 81742 115606 81806
rect 115670 81742 115812 81806
rect 115600 81736 115812 81742
rect 116008 81942 116628 81948
rect 116008 81878 116014 81942
rect 116078 81878 116422 81942
rect 116486 81878 116628 81942
rect 116008 81872 116628 81878
rect 116008 81812 116220 81872
rect 116008 81806 116356 81812
rect 116008 81742 116286 81806
rect 116350 81742 116356 81806
rect 116008 81736 116356 81742
rect 116416 81736 116628 81872
rect 116824 81942 117036 81948
rect 116824 81878 116830 81942
rect 116894 81878 117036 81942
rect 116824 81736 117036 81878
rect 116960 81676 117036 81736
rect 28560 81540 28636 81600
rect 110296 81540 110372 81600
rect 22168 81534 22788 81540
rect 22168 81470 22310 81534
rect 22374 81470 22582 81534
rect 22646 81470 22788 81534
rect 22168 81464 22788 81470
rect 22168 81328 22380 81464
rect 22576 81328 22788 81464
rect 22984 81534 23196 81540
rect 22984 81470 23126 81534
rect 23190 81470 23196 81534
rect 22984 81398 23196 81470
rect 22984 81334 22990 81398
rect 23054 81334 23196 81398
rect 22984 81328 23196 81334
rect 23392 81534 23604 81540
rect 23392 81470 23534 81534
rect 23598 81470 23604 81534
rect 23392 81398 23604 81470
rect 23392 81334 23534 81398
rect 23598 81334 23604 81398
rect 23392 81328 23604 81334
rect 21760 81268 21836 81328
rect 22304 81268 22380 81328
rect 22712 81268 22788 81328
rect 1224 81126 1980 81132
rect 1224 81062 1230 81126
rect 1294 81062 1980 81126
rect 1224 81056 1980 81062
rect 1768 81048 1980 81056
rect 1768 80992 1798 81048
rect 1854 80992 1980 81048
rect 1768 80920 1980 80992
rect 21760 80920 21972 81268
rect 22168 80990 22380 81268
rect 22168 80926 22174 80990
rect 22238 80926 22380 80990
rect 22168 80920 22380 80926
rect 22576 80920 22788 81268
rect 22984 81126 23196 81132
rect 22984 81062 22990 81126
rect 23054 81062 23196 81126
rect 22984 80920 23196 81062
rect 23392 81126 23604 81132
rect 23392 81062 23534 81126
rect 23598 81062 23604 81126
rect 23392 80920 23604 81062
rect 28288 81126 28636 81540
rect 28288 81062 28294 81126
rect 28358 81062 28636 81126
rect 28288 81056 28636 81062
rect 110160 81056 110508 81540
rect 115192 81534 115404 81540
rect 115192 81470 115198 81534
rect 115262 81470 115404 81534
rect 115192 81398 115404 81470
rect 115192 81334 115198 81398
rect 115262 81334 115404 81398
rect 115192 81328 115404 81334
rect 115600 81534 115812 81540
rect 115600 81470 115606 81534
rect 115670 81470 115812 81534
rect 115600 81398 115812 81470
rect 115600 81334 115606 81398
rect 115670 81334 115812 81398
rect 115600 81328 115812 81334
rect 116008 81404 116220 81540
rect 116318 81534 116628 81540
rect 116280 81470 116286 81534
rect 116350 81470 116628 81534
rect 116318 81464 116628 81470
rect 116416 81404 116628 81464
rect 116008 81328 116628 81404
rect 116008 81268 116084 81328
rect 116552 81268 116628 81328
rect 110432 80996 110508 81056
rect 21760 80860 21836 80920
rect 22984 80860 23060 80920
rect 23528 80860 23604 80920
rect 21760 80718 21972 80860
rect 21760 80654 21902 80718
rect 21966 80654 21972 80718
rect 21760 80648 21972 80654
rect 22168 80718 22380 80724
rect 22168 80654 22174 80718
rect 22238 80654 22380 80718
rect 22168 80512 22380 80654
rect 22576 80588 22788 80724
rect 22478 80582 22788 80588
rect 22440 80518 22446 80582
rect 22510 80518 22788 80582
rect 22478 80512 22788 80518
rect 22984 80512 23196 80860
rect 23392 80512 23604 80860
rect 22168 80452 22244 80512
rect 22984 80452 23060 80512
rect 23528 80452 23604 80512
rect 21760 80446 21972 80452
rect 21760 80382 21902 80446
rect 21966 80382 21972 80446
rect 21760 80310 21972 80382
rect 21760 80246 21902 80310
rect 21966 80246 21972 80310
rect 21760 80240 21972 80246
rect 22168 80376 22788 80452
rect 22168 80316 22380 80376
rect 22168 80310 22516 80316
rect 22168 80246 22446 80310
rect 22510 80246 22516 80310
rect 22168 80240 22516 80246
rect 22576 80310 22788 80376
rect 22576 80246 22718 80310
rect 22782 80246 22788 80310
rect 22576 80240 22788 80246
rect 22984 80104 23196 80452
rect 23392 80104 23604 80452
rect 28288 80854 28636 80996
rect 28288 80790 28294 80854
rect 28358 80790 28566 80854
rect 28630 80790 28636 80854
rect 28288 80582 28636 80790
rect 28288 80518 28566 80582
rect 28630 80518 28636 80582
rect 28288 80446 28636 80518
rect 28288 80382 28294 80446
rect 28358 80382 28636 80446
rect 28288 80376 28636 80382
rect 110160 80446 110508 80996
rect 115192 81126 115404 81132
rect 115192 81062 115198 81126
rect 115262 81062 115404 81126
rect 115192 80920 115404 81062
rect 115600 81126 115812 81132
rect 115600 81062 115606 81126
rect 115670 81062 115812 81126
rect 115600 80920 115812 81062
rect 116008 80990 116220 81268
rect 116008 80926 116150 80990
rect 116214 80926 116220 80990
rect 116008 80920 116220 80926
rect 116416 80920 116628 81268
rect 116824 81328 117036 81676
rect 116824 81268 116900 81328
rect 116824 80920 117036 81268
rect 136816 81126 137572 81132
rect 136816 81062 137502 81126
rect 137566 81062 137572 81126
rect 136816 81056 137572 81062
rect 136816 81048 137028 81056
rect 136816 80992 136944 81048
rect 137000 80992 137028 81048
rect 136816 80920 137028 80992
rect 115328 80860 115404 80920
rect 115736 80860 115812 80920
rect 110160 80382 110438 80446
rect 110502 80382 110508 80446
rect 110160 80376 110508 80382
rect 115192 80512 115404 80860
rect 115600 80512 115812 80860
rect 116824 80860 116900 80920
rect 116008 80718 116220 80724
rect 116008 80654 116150 80718
rect 116214 80654 116220 80718
rect 116008 80512 116220 80654
rect 116416 80588 116628 80724
rect 116824 80718 117036 80860
rect 116824 80654 116830 80718
rect 116894 80654 117036 80718
rect 116824 80648 117036 80654
rect 116280 80512 116628 80588
rect 115192 80452 115268 80512
rect 115600 80452 115676 80512
rect 116008 80452 116084 80512
rect 116280 80452 116356 80512
rect 116552 80452 116628 80512
rect 22984 80044 23060 80104
rect 23528 80044 23604 80104
rect 21760 80038 21972 80044
rect 21760 79974 21902 80038
rect 21966 79974 21972 80038
rect 21760 79902 21972 79974
rect 21760 79838 21766 79902
rect 21830 79838 21972 79902
rect 21760 79832 21972 79838
rect 22168 80038 22788 80044
rect 22168 79974 22718 80038
rect 22782 79974 22788 80038
rect 22168 79968 22788 79974
rect 22168 79696 22380 79968
rect 22304 79636 22380 79696
rect 21760 79630 21972 79636
rect 21760 79566 21766 79630
rect 21830 79566 21972 79630
rect 1224 79494 1980 79500
rect 1224 79430 1230 79494
rect 1294 79430 1980 79494
rect 1224 79424 1980 79430
rect 21760 79494 21972 79566
rect 21760 79430 21902 79494
rect 21966 79430 21972 79494
rect 21760 79424 21972 79430
rect 22168 79424 22380 79636
rect 22576 79696 22788 79968
rect 22984 79902 23196 80044
rect 22984 79838 22990 79902
rect 23054 79838 23196 79902
rect 22984 79832 23196 79838
rect 23392 79902 23604 80044
rect 23392 79838 23534 79902
rect 23598 79838 23604 79902
rect 23392 79832 23604 79838
rect 28288 80174 28636 80180
rect 28288 80110 28294 80174
rect 28358 80110 28636 80174
rect 28288 79832 28636 80110
rect 110160 80174 110508 80180
rect 110160 80110 110438 80174
rect 110502 80110 110508 80174
rect 110160 80038 110508 80110
rect 115192 80104 115404 80452
rect 115600 80104 115812 80452
rect 116008 80376 116356 80452
rect 116008 80316 116220 80376
rect 116008 80310 116356 80316
rect 116008 80246 116014 80310
rect 116078 80246 116286 80310
rect 116350 80246 116356 80310
rect 116008 80240 116356 80246
rect 116416 80240 116628 80452
rect 116824 80446 117036 80452
rect 116824 80382 116830 80446
rect 116894 80382 117036 80446
rect 116824 80310 117036 80382
rect 116824 80246 116830 80310
rect 116894 80246 117036 80310
rect 116824 80240 117036 80246
rect 115328 80044 115404 80104
rect 115736 80044 115812 80104
rect 110160 79974 110166 80038
rect 110230 79974 110508 80038
rect 110160 79832 110508 79974
rect 115192 79902 115404 80044
rect 115192 79838 115334 79902
rect 115398 79838 115404 79902
rect 115192 79832 115404 79838
rect 115600 79902 115812 80044
rect 115600 79838 115742 79902
rect 115806 79838 115812 79902
rect 115600 79832 115812 79838
rect 116008 80038 116220 80044
rect 116318 80038 116628 80044
rect 116008 79974 116014 80038
rect 116078 79974 116220 80038
rect 116280 79974 116286 80038
rect 116350 79974 116628 80038
rect 28288 79772 28364 79832
rect 110432 79772 110508 79832
rect 22576 79636 22652 79696
rect 22576 79494 22788 79636
rect 22576 79430 22718 79494
rect 22782 79430 22788 79494
rect 22576 79424 22788 79430
rect 22984 79630 23196 79636
rect 22984 79566 22990 79630
rect 23054 79566 23196 79630
rect 22984 79494 23196 79566
rect 22984 79430 23126 79494
rect 23190 79430 23196 79494
rect 22984 79424 23196 79430
rect 23392 79630 23604 79636
rect 23392 79566 23534 79630
rect 23598 79566 23604 79630
rect 23392 79494 23604 79566
rect 28288 79560 28636 79772
rect 110160 79766 110508 79772
rect 110160 79702 110166 79766
rect 110230 79702 110508 79766
rect 110160 79560 110508 79702
rect 116008 79696 116220 79974
rect 116318 79968 116628 79974
rect 116416 79772 116628 79968
rect 116824 80038 117036 80044
rect 116824 79974 116830 80038
rect 116894 79974 117036 80038
rect 116824 79902 117036 79974
rect 116824 79838 116830 79902
rect 116894 79838 117036 79902
rect 116824 79832 117036 79838
rect 116318 79766 116628 79772
rect 116280 79702 116286 79766
rect 116350 79702 116628 79766
rect 116318 79696 116628 79702
rect 115192 79630 115404 79636
rect 115192 79566 115334 79630
rect 115398 79566 115404 79630
rect 28560 79500 28636 79560
rect 110296 79500 110372 79560
rect 23392 79430 23398 79494
rect 23462 79430 23604 79494
rect 23392 79424 23604 79430
rect 1768 79368 1980 79424
rect 1768 79312 1798 79368
rect 1854 79312 1980 79368
rect 1768 79288 1980 79312
rect 21760 79222 21972 79228
rect 21760 79158 21902 79222
rect 21966 79158 21972 79222
rect 21760 79086 21972 79158
rect 21760 79022 21766 79086
rect 21830 79022 21972 79086
rect 21760 79016 21972 79022
rect 22168 79092 22380 79228
rect 22576 79222 22788 79228
rect 22576 79158 22718 79222
rect 22782 79158 22788 79222
rect 22576 79092 22788 79158
rect 22168 79016 22788 79092
rect 22984 79222 23196 79228
rect 22984 79158 23126 79222
rect 23190 79158 23196 79222
rect 22984 79086 23196 79158
rect 22984 79022 23126 79086
rect 23190 79022 23196 79086
rect 22984 79016 23196 79022
rect 23392 79222 23604 79228
rect 23392 79158 23398 79222
rect 23462 79158 23604 79222
rect 23392 79086 23604 79158
rect 23392 79022 23398 79086
rect 23462 79022 23604 79086
rect 23392 79016 23604 79022
rect 28288 79222 28636 79500
rect 28288 79158 28294 79222
rect 28358 79158 28636 79222
rect 28288 79016 28636 79158
rect 110160 79016 110508 79500
rect 115192 79494 115404 79566
rect 115192 79430 115198 79494
rect 115262 79430 115404 79494
rect 115192 79424 115404 79430
rect 115600 79630 115812 79636
rect 115600 79566 115742 79630
rect 115806 79566 115812 79630
rect 115600 79494 115812 79566
rect 115600 79430 115606 79494
rect 115670 79430 115812 79494
rect 115600 79424 115812 79430
rect 116008 79560 116628 79636
rect 116008 79500 116220 79560
rect 116008 79494 116356 79500
rect 116008 79430 116286 79494
rect 116350 79430 116356 79494
rect 116008 79424 116356 79430
rect 116416 79494 116628 79560
rect 116416 79430 116558 79494
rect 116622 79430 116628 79494
rect 116416 79424 116628 79430
rect 116824 79630 117036 79636
rect 116824 79566 116830 79630
rect 116894 79566 117036 79630
rect 116824 79494 117036 79566
rect 116824 79430 116966 79494
rect 117030 79430 117036 79494
rect 116824 79424 117036 79430
rect 136816 79494 137572 79500
rect 136816 79430 137502 79494
rect 137566 79430 137572 79494
rect 136816 79424 137572 79430
rect 136816 79368 137028 79424
rect 136816 79312 136944 79368
rect 137000 79312 137028 79368
rect 136816 79288 137028 79312
rect 115192 79222 115404 79228
rect 115192 79158 115198 79222
rect 115262 79158 115404 79222
rect 115192 79086 115404 79158
rect 115192 79022 115198 79086
rect 115262 79022 115404 79086
rect 115192 79016 115404 79022
rect 115600 79222 115812 79228
rect 115600 79158 115606 79222
rect 115670 79158 115812 79222
rect 115600 79086 115812 79158
rect 115600 79022 115742 79086
rect 115806 79022 115812 79086
rect 115600 79016 115812 79022
rect 116008 79092 116220 79228
rect 116416 79222 116628 79228
rect 116416 79158 116558 79222
rect 116622 79158 116628 79222
rect 116416 79092 116628 79158
rect 116008 79086 116628 79092
rect 116008 79022 116014 79086
rect 116078 79022 116628 79086
rect 116008 79016 116628 79022
rect 116824 79222 117036 79228
rect 116824 79158 116966 79222
rect 117030 79158 117036 79222
rect 116824 79086 117036 79158
rect 116824 79022 116966 79086
rect 117030 79022 117036 79086
rect 116824 79016 117036 79022
rect 22304 78956 22380 79016
rect 28288 78956 28364 79016
rect 110296 78956 110372 79016
rect 116144 78956 116220 79016
rect 22304 78880 22652 78956
rect 22576 78820 22652 78880
rect 28288 78950 28636 78956
rect 28288 78886 28294 78950
rect 28358 78886 28636 78950
rect 21760 78814 21972 78820
rect 21760 78750 21766 78814
rect 21830 78750 21972 78814
rect 21760 78678 21972 78750
rect 21760 78614 21902 78678
rect 21966 78614 21972 78678
rect 21760 78608 21972 78614
rect 22168 78678 22380 78820
rect 22168 78614 22310 78678
rect 22374 78614 22380 78678
rect 22168 78608 22380 78614
rect 22576 78678 22788 78820
rect 22576 78614 22582 78678
rect 22646 78614 22788 78678
rect 22576 78608 22788 78614
rect 22984 78814 23196 78820
rect 22984 78750 23126 78814
rect 23190 78750 23196 78814
rect 22984 78678 23196 78750
rect 22984 78614 22990 78678
rect 23054 78614 23196 78678
rect 22984 78608 23196 78614
rect 23392 78814 23604 78820
rect 23392 78750 23398 78814
rect 23462 78750 23604 78814
rect 23392 78678 23604 78750
rect 28288 78744 28636 78886
rect 110160 78744 110508 78956
rect 116144 78880 116492 78956
rect 116416 78820 116492 78880
rect 115192 78814 115404 78820
rect 115192 78750 115198 78814
rect 115262 78750 115404 78814
rect 28424 78684 28500 78744
rect 110296 78684 110372 78744
rect 23392 78614 23398 78678
rect 23462 78614 23604 78678
rect 23392 78608 23604 78614
rect 28288 78472 28636 78684
rect 110160 78472 110508 78684
rect 115192 78678 115404 78750
rect 115192 78614 115334 78678
rect 115398 78614 115404 78678
rect 115192 78608 115404 78614
rect 115600 78814 115812 78820
rect 115600 78750 115742 78814
rect 115806 78750 115812 78814
rect 115600 78678 115812 78750
rect 115600 78614 115742 78678
rect 115806 78614 115812 78678
rect 115600 78608 115812 78614
rect 116008 78814 116220 78820
rect 116008 78750 116014 78814
rect 116078 78750 116220 78814
rect 116008 78678 116220 78750
rect 116008 78614 116014 78678
rect 116078 78614 116220 78678
rect 116008 78608 116220 78614
rect 116416 78608 116628 78820
rect 116824 78814 117036 78820
rect 116824 78750 116966 78814
rect 117030 78750 117036 78814
rect 116824 78678 117036 78750
rect 116824 78614 116966 78678
rect 117030 78614 117036 78678
rect 116824 78608 117036 78614
rect 28424 78412 28500 78472
rect 110160 78412 110236 78472
rect 21760 78406 21972 78412
rect 21760 78342 21902 78406
rect 21966 78342 21972 78406
rect 21760 78270 21972 78342
rect 21760 78206 21902 78270
rect 21966 78206 21972 78270
rect 21760 78200 21972 78206
rect 22168 78406 22380 78412
rect 22168 78342 22310 78406
rect 22374 78342 22380 78406
rect 22168 78276 22380 78342
rect 22576 78406 22788 78412
rect 22576 78342 22582 78406
rect 22646 78342 22788 78406
rect 22576 78276 22788 78342
rect 22168 78270 22788 78276
rect 22168 78206 22310 78270
rect 22374 78206 22788 78270
rect 22168 78200 22788 78206
rect 22984 78406 23196 78412
rect 22984 78342 22990 78406
rect 23054 78342 23196 78406
rect 22984 78270 23196 78342
rect 22984 78206 22990 78270
rect 23054 78206 23196 78270
rect 22984 78200 23196 78206
rect 23392 78406 23604 78412
rect 23392 78342 23398 78406
rect 23462 78342 23604 78406
rect 23392 78270 23604 78342
rect 23392 78206 23398 78270
rect 23462 78206 23604 78270
rect 23392 78200 23604 78206
rect 28288 78200 28636 78412
rect 110160 78200 110508 78412
rect 115192 78406 115404 78412
rect 115192 78342 115334 78406
rect 115398 78342 115404 78406
rect 115192 78270 115404 78342
rect 115192 78206 115334 78270
rect 115398 78206 115404 78270
rect 115192 78200 115404 78206
rect 115600 78406 115812 78412
rect 115600 78342 115742 78406
rect 115806 78342 115812 78406
rect 115600 78270 115812 78342
rect 115600 78206 115606 78270
rect 115670 78206 115812 78270
rect 115600 78200 115812 78206
rect 116008 78406 116220 78412
rect 116008 78342 116014 78406
rect 116078 78342 116220 78406
rect 116008 78276 116220 78342
rect 116416 78276 116628 78412
rect 116008 78270 116628 78276
rect 116008 78206 116014 78270
rect 116078 78206 116628 78270
rect 116008 78200 116628 78206
rect 116824 78406 117036 78412
rect 116824 78342 116966 78406
rect 117030 78342 117036 78406
rect 116824 78270 117036 78342
rect 116824 78206 116966 78270
rect 117030 78206 117036 78270
rect 116824 78200 117036 78206
rect 22304 78140 22380 78200
rect 28288 78140 28364 78200
rect 110432 78140 110508 78200
rect 22304 78064 22652 78140
rect 22576 78004 22652 78064
rect 21760 77998 21972 78004
rect 21760 77934 21902 77998
rect 21966 77934 21972 77998
rect 21760 77792 21972 77934
rect 22168 77998 22380 78004
rect 22168 77934 22310 77998
rect 22374 77934 22380 77998
rect 22168 77868 22380 77934
rect 22168 77862 22516 77868
rect 22168 77798 22446 77862
rect 22510 77798 22516 77862
rect 22168 77792 22516 77798
rect 22576 77792 22788 78004
rect 22984 77998 23196 78004
rect 22984 77934 22990 77998
rect 23054 77934 23196 77998
rect 22984 77862 23196 77934
rect 22984 77798 23126 77862
rect 23190 77798 23196 77862
rect 22984 77792 23196 77798
rect 23392 77998 23604 78004
rect 23392 77934 23398 77998
rect 23462 77934 23604 77998
rect 23392 77862 23604 77934
rect 23392 77798 23534 77862
rect 23598 77798 23604 77862
rect 23392 77792 23604 77798
rect 28288 77928 28636 78140
rect 110160 77928 110508 78140
rect 115192 77998 115404 78004
rect 115192 77934 115334 77998
rect 115398 77934 115404 77998
rect 28288 77868 28364 77928
rect 110296 77868 110372 77928
rect 21760 77732 21836 77792
rect 1224 77726 1980 77732
rect 1224 77662 1230 77726
rect 1294 77688 1980 77726
rect 1294 77662 1798 77688
rect 1224 77656 1798 77662
rect 1768 77632 1798 77656
rect 1854 77632 1980 77688
rect 1768 77520 1980 77632
rect 21760 77384 21972 77732
rect 28288 77726 28636 77868
rect 28288 77662 28294 77726
rect 28358 77662 28636 77726
rect 28288 77656 28636 77662
rect 110160 77726 110508 77868
rect 115192 77862 115404 77934
rect 115192 77798 115334 77862
rect 115398 77798 115404 77862
rect 115192 77792 115404 77798
rect 115600 77998 115812 78004
rect 115600 77934 115606 77998
rect 115670 77934 115812 77998
rect 115600 77862 115812 77934
rect 115600 77798 115742 77862
rect 115806 77798 115812 77862
rect 115600 77792 115812 77798
rect 116008 77998 116628 78004
rect 116008 77934 116014 77998
rect 116078 77934 116628 77998
rect 116008 77928 116628 77934
rect 116008 77868 116220 77928
rect 116008 77862 116356 77868
rect 116008 77798 116286 77862
rect 116350 77798 116356 77862
rect 116008 77792 116356 77798
rect 116416 77792 116628 77928
rect 116824 77998 117036 78004
rect 116824 77934 116966 77998
rect 117030 77934 117036 77998
rect 116824 77792 117036 77934
rect 110160 77662 110438 77726
rect 110502 77662 110508 77726
rect 110160 77656 110508 77662
rect 116824 77732 116900 77792
rect 28560 77596 28636 77656
rect 110296 77596 110372 77656
rect 21896 77324 21972 77384
rect 21760 76976 21972 77324
rect 22168 77384 22380 77596
rect 22478 77590 22788 77596
rect 22440 77526 22446 77590
rect 22510 77526 22788 77590
rect 22478 77520 22788 77526
rect 22576 77384 22788 77520
rect 22984 77590 23196 77596
rect 22984 77526 23126 77590
rect 23190 77526 23196 77590
rect 22984 77454 23196 77526
rect 22984 77390 22990 77454
rect 23054 77390 23196 77454
rect 22984 77384 23196 77390
rect 23392 77590 23604 77596
rect 23392 77526 23534 77590
rect 23598 77526 23604 77590
rect 23392 77454 23604 77526
rect 23392 77390 23398 77454
rect 23462 77390 23604 77454
rect 23392 77384 23604 77390
rect 28288 77454 28636 77596
rect 28288 77390 28294 77454
rect 28358 77390 28636 77454
rect 22168 77324 22244 77384
rect 22576 77324 22652 77384
rect 22168 77188 22380 77324
rect 22576 77188 22788 77324
rect 22168 77112 22788 77188
rect 22168 76976 22380 77112
rect 22576 77046 22788 77112
rect 22576 76982 22582 77046
rect 22646 76982 22788 77046
rect 22576 76976 22788 76982
rect 22984 77182 23196 77188
rect 22984 77118 22990 77182
rect 23054 77118 23196 77182
rect 22984 77046 23196 77118
rect 22984 76982 22990 77046
rect 23054 76982 23196 77046
rect 22984 76976 23196 76982
rect 23392 77182 23604 77188
rect 23392 77118 23398 77182
rect 23462 77118 23604 77182
rect 23392 77046 23604 77118
rect 28288 77112 28636 77390
rect 110160 77454 110508 77596
rect 110160 77390 110438 77454
rect 110502 77390 110508 77454
rect 110160 77112 110508 77390
rect 115192 77590 115404 77596
rect 115192 77526 115334 77590
rect 115398 77526 115404 77590
rect 115192 77454 115404 77526
rect 115192 77390 115334 77454
rect 115398 77390 115404 77454
rect 115192 77384 115404 77390
rect 115600 77590 115812 77596
rect 115600 77526 115742 77590
rect 115806 77526 115812 77590
rect 115600 77454 115812 77526
rect 115600 77390 115606 77454
rect 115670 77390 115812 77454
rect 115600 77384 115812 77390
rect 116008 77460 116220 77596
rect 116318 77590 116628 77596
rect 116280 77526 116286 77590
rect 116350 77526 116628 77590
rect 116318 77520 116628 77526
rect 116416 77460 116628 77520
rect 116008 77384 116628 77460
rect 116824 77384 117036 77732
rect 136816 77688 137028 77732
rect 136816 77632 136944 77688
rect 137000 77632 137028 77688
rect 136816 77596 137028 77632
rect 136816 77590 137572 77596
rect 136816 77526 137502 77590
rect 137566 77526 137572 77590
rect 136816 77520 137572 77526
rect 116008 77324 116084 77384
rect 116552 77324 116628 77384
rect 116960 77324 117036 77384
rect 115192 77182 115404 77188
rect 115192 77118 115334 77182
rect 115398 77118 115404 77182
rect 28560 77052 28636 77112
rect 110296 77052 110372 77112
rect 23392 76982 23534 77046
rect 23598 76982 23604 77046
rect 23392 76976 23604 76982
rect 21760 76916 21836 76976
rect 21760 76774 21972 76916
rect 28288 76840 28636 77052
rect 110160 76910 110508 77052
rect 115192 77046 115404 77118
rect 115192 76982 115334 77046
rect 115398 76982 115404 77046
rect 115192 76976 115404 76982
rect 115600 77182 115812 77188
rect 115600 77118 115606 77182
rect 115670 77118 115812 77182
rect 115600 77046 115812 77118
rect 115600 76982 115742 77046
rect 115806 76982 115812 77046
rect 115600 76976 115812 76982
rect 116008 77046 116220 77324
rect 116008 76982 116014 77046
rect 116078 76982 116220 77046
rect 116008 76976 116220 76982
rect 116416 76976 116628 77324
rect 116824 76976 117036 77324
rect 110160 76846 110438 76910
rect 110502 76846 110508 76910
rect 110160 76840 110508 76846
rect 28424 76780 28500 76840
rect 110432 76780 110508 76840
rect 116824 76916 116900 76976
rect 21760 76710 21766 76774
rect 21830 76710 21972 76774
rect 21760 76704 21972 76710
rect 22168 76568 22380 76780
rect 22576 76774 22788 76780
rect 22576 76710 22582 76774
rect 22646 76710 22788 76774
rect 22576 76568 22788 76710
rect 22984 76774 23196 76780
rect 22984 76710 22990 76774
rect 23054 76710 23196 76774
rect 22984 76568 23196 76710
rect 23392 76774 23604 76780
rect 23392 76710 23534 76774
rect 23598 76710 23604 76774
rect 23392 76568 23604 76710
rect 22168 76508 22244 76568
rect 22576 76508 22652 76568
rect 22984 76508 23060 76568
rect 23528 76508 23604 76568
rect 21760 76502 21972 76508
rect 21760 76438 21766 76502
rect 21830 76438 21972 76502
rect 21760 76366 21972 76438
rect 21760 76302 21902 76366
rect 21966 76302 21972 76366
rect 21760 76296 21972 76302
rect 22168 76372 22380 76508
rect 22576 76372 22788 76508
rect 22168 76366 22788 76372
rect 22168 76302 22582 76366
rect 22646 76302 22788 76366
rect 22168 76296 22788 76302
rect 22984 76160 23196 76508
rect 23392 76160 23604 76508
rect 28288 76502 28636 76780
rect 28288 76438 28294 76502
rect 28358 76438 28636 76502
rect 28288 76432 28636 76438
rect 110160 76638 110508 76780
rect 110160 76574 110438 76638
rect 110502 76574 110508 76638
rect 110160 76502 110508 76574
rect 115192 76774 115404 76780
rect 115192 76710 115334 76774
rect 115398 76710 115404 76774
rect 115192 76568 115404 76710
rect 115328 76508 115404 76568
rect 110160 76438 110302 76502
rect 110366 76438 110508 76502
rect 110160 76432 110508 76438
rect 28288 76230 28636 76236
rect 28288 76166 28294 76230
rect 28358 76166 28636 76230
rect 22984 76100 23060 76160
rect 23392 76100 23468 76160
rect 1768 76008 1980 76100
rect 1768 75964 1798 76008
rect 1224 75958 1798 75964
rect 1224 75894 1230 75958
rect 1294 75952 1798 75958
rect 1854 75952 1980 76008
rect 1294 75894 1980 75952
rect 1224 75888 1980 75894
rect 21760 76094 21972 76100
rect 21760 76030 21902 76094
rect 21966 76030 21972 76094
rect 21760 75958 21972 76030
rect 21760 75894 21766 75958
rect 21830 75894 21972 75958
rect 21760 75888 21972 75894
rect 22168 76094 22788 76100
rect 22168 76030 22582 76094
rect 22646 76030 22788 76094
rect 22168 76024 22788 76030
rect 22168 75828 22380 76024
rect 22168 75752 22516 75828
rect 22576 75752 22788 76024
rect 22984 75752 23196 76100
rect 23392 75752 23604 76100
rect 22168 75692 22244 75752
rect 22440 75692 22516 75752
rect 22984 75692 23060 75752
rect 23528 75692 23604 75752
rect 21760 75686 21972 75692
rect 21760 75622 21766 75686
rect 21830 75622 21972 75686
rect 21760 75550 21972 75622
rect 21760 75486 21766 75550
rect 21830 75486 21972 75550
rect 21760 75480 21972 75486
rect 22168 75480 22380 75692
rect 22440 75616 22788 75692
rect 22576 75556 22788 75616
rect 22478 75550 22788 75556
rect 22440 75486 22446 75550
rect 22510 75486 22788 75550
rect 22478 75480 22788 75486
rect 22984 75550 23196 75692
rect 22984 75486 22990 75550
rect 23054 75486 23196 75550
rect 22984 75480 23196 75486
rect 23392 75550 23604 75692
rect 28288 76094 28636 76166
rect 28288 76030 28566 76094
rect 28630 76030 28636 76094
rect 28288 75822 28636 76030
rect 28288 75758 28566 75822
rect 28630 75758 28636 75822
rect 28288 75616 28636 75758
rect 110160 76230 110508 76236
rect 110160 76166 110302 76230
rect 110366 76166 110508 76230
rect 110160 75616 110508 76166
rect 115192 76160 115404 76508
rect 115600 76774 115812 76780
rect 115600 76710 115742 76774
rect 115806 76710 115812 76774
rect 115600 76568 115812 76710
rect 116008 76774 116220 76780
rect 116008 76710 116014 76774
rect 116078 76710 116220 76774
rect 116008 76568 116220 76710
rect 115600 76508 115676 76568
rect 116144 76508 116220 76568
rect 115600 76160 115812 76508
rect 116008 76366 116220 76508
rect 116008 76302 116150 76366
rect 116214 76302 116220 76366
rect 116008 76296 116220 76302
rect 116416 76568 116628 76780
rect 116824 76774 117036 76916
rect 116824 76710 116830 76774
rect 116894 76710 117036 76774
rect 116824 76704 117036 76710
rect 116416 76508 116492 76568
rect 116416 76366 116628 76508
rect 116416 76302 116558 76366
rect 116622 76302 116628 76366
rect 116416 76296 116628 76302
rect 116824 76502 117036 76508
rect 116824 76438 116830 76502
rect 116894 76438 117036 76502
rect 116824 76366 117036 76438
rect 116824 76302 116966 76366
rect 117030 76302 117036 76366
rect 116824 76296 117036 76302
rect 115192 76100 115268 76160
rect 115600 76100 115676 76160
rect 115192 75752 115404 76100
rect 115600 75752 115812 76100
rect 116008 76094 116628 76100
rect 116008 76030 116150 76094
rect 116214 76030 116558 76094
rect 116622 76030 116628 76094
rect 116008 76024 116628 76030
rect 116008 75828 116220 76024
rect 116008 75752 116356 75828
rect 116416 75752 116628 76024
rect 116824 76094 117036 76100
rect 116824 76030 116966 76094
rect 117030 76030 117036 76094
rect 116824 75958 117036 76030
rect 116824 75894 116830 75958
rect 116894 75894 117036 75958
rect 116824 75888 117036 75894
rect 136816 76008 137028 76100
rect 136816 75952 136944 76008
rect 137000 75964 137028 76008
rect 137000 75958 137572 75964
rect 137000 75952 137502 75958
rect 136816 75894 137502 75952
rect 137566 75894 137572 75958
rect 136816 75888 137572 75894
rect 115328 75692 115404 75752
rect 115736 75692 115812 75752
rect 116144 75692 116220 75752
rect 28424 75556 28500 75616
rect 110432 75556 110508 75616
rect 23392 75486 23534 75550
rect 23598 75486 23604 75550
rect 23392 75480 23604 75486
rect 21760 75278 21972 75284
rect 21760 75214 21766 75278
rect 21830 75214 21972 75278
rect 21760 75142 21972 75214
rect 21760 75078 21902 75142
rect 21966 75078 21972 75142
rect 21760 75072 21972 75078
rect 22168 75278 22516 75284
rect 22168 75214 22446 75278
rect 22510 75214 22516 75278
rect 22168 75208 22516 75214
rect 22168 75148 22380 75208
rect 22576 75148 22788 75284
rect 22168 75142 22788 75148
rect 22168 75078 22718 75142
rect 22782 75078 22788 75142
rect 22168 75072 22788 75078
rect 22984 75278 23196 75284
rect 22984 75214 22990 75278
rect 23054 75214 23196 75278
rect 22984 75142 23196 75214
rect 22984 75078 23126 75142
rect 23190 75078 23196 75142
rect 22984 75072 23196 75078
rect 23392 75278 23604 75284
rect 23392 75214 23534 75278
rect 23598 75214 23604 75278
rect 23392 75142 23604 75214
rect 23392 75078 23398 75142
rect 23462 75078 23604 75142
rect 23392 75072 23604 75078
rect 28288 75278 28636 75556
rect 28288 75214 28430 75278
rect 28494 75214 28636 75278
rect 28288 75072 28636 75214
rect 110160 75072 110508 75556
rect 115192 75550 115404 75692
rect 115192 75486 115334 75550
rect 115398 75486 115404 75550
rect 115192 75480 115404 75486
rect 115600 75550 115812 75692
rect 115600 75486 115742 75550
rect 115806 75486 115812 75550
rect 115600 75480 115812 75486
rect 116008 75550 116220 75692
rect 116280 75692 116356 75752
rect 116280 75616 116628 75692
rect 116008 75486 116150 75550
rect 116214 75486 116220 75550
rect 116008 75480 116220 75486
rect 116416 75550 116628 75616
rect 116416 75486 116422 75550
rect 116486 75486 116628 75550
rect 116416 75480 116628 75486
rect 116824 75686 117036 75692
rect 116824 75622 116830 75686
rect 116894 75622 117036 75686
rect 116824 75550 117036 75622
rect 116824 75486 116830 75550
rect 116894 75486 117036 75550
rect 116824 75480 117036 75486
rect 115192 75278 115404 75284
rect 115192 75214 115334 75278
rect 115398 75214 115404 75278
rect 115192 75142 115404 75214
rect 115192 75078 115198 75142
rect 115262 75078 115404 75142
rect 115192 75072 115404 75078
rect 115600 75278 115812 75284
rect 115600 75214 115742 75278
rect 115806 75214 115812 75278
rect 115600 75142 115812 75214
rect 115600 75078 115606 75142
rect 115670 75078 115812 75142
rect 115600 75072 115812 75078
rect 116008 75278 116220 75284
rect 116008 75214 116150 75278
rect 116214 75214 116220 75278
rect 116008 75072 116220 75214
rect 116416 75278 116628 75284
rect 116416 75214 116422 75278
rect 116486 75214 116628 75278
rect 116416 75142 116628 75214
rect 116416 75078 116558 75142
rect 116622 75078 116628 75142
rect 116416 75072 116628 75078
rect 116824 75278 117036 75284
rect 116824 75214 116830 75278
rect 116894 75214 117036 75278
rect 116824 75142 117036 75214
rect 116824 75078 116966 75142
rect 117030 75078 117036 75142
rect 116824 75072 117036 75078
rect 28424 75012 28500 75072
rect 110432 75012 110508 75072
rect 28288 75006 28636 75012
rect 28288 74942 28430 75006
rect 28494 74942 28636 75006
rect 21760 74870 21972 74876
rect 21760 74806 21902 74870
rect 21966 74806 21972 74870
rect 21760 74734 21972 74806
rect 21760 74670 21766 74734
rect 21830 74670 21972 74734
rect 21760 74664 21972 74670
rect 22168 74870 22788 74876
rect 22168 74806 22718 74870
rect 22782 74806 22788 74870
rect 22168 74800 22788 74806
rect 22168 74740 22380 74800
rect 22168 74734 22516 74740
rect 22168 74670 22174 74734
rect 22238 74670 22446 74734
rect 22510 74670 22516 74734
rect 22168 74664 22516 74670
rect 22576 74664 22788 74800
rect 22984 74870 23196 74876
rect 22984 74806 23126 74870
rect 23190 74806 23196 74870
rect 22984 74734 23196 74806
rect 22984 74670 23126 74734
rect 23190 74670 23196 74734
rect 22984 74664 23196 74670
rect 23392 74870 23604 74876
rect 23392 74806 23398 74870
rect 23462 74806 23604 74870
rect 23392 74734 23604 74806
rect 28288 74800 28636 74942
rect 28560 74740 28636 74800
rect 23392 74670 23398 74734
rect 23462 74670 23604 74734
rect 23392 74664 23604 74670
rect 28288 74528 28636 74740
rect 110160 74800 110508 75012
rect 115192 74870 115404 74876
rect 115192 74806 115198 74870
rect 115262 74806 115404 74870
rect 110160 74740 110236 74800
rect 110160 74528 110508 74740
rect 115192 74734 115404 74806
rect 115192 74670 115198 74734
rect 115262 74670 115404 74734
rect 115192 74664 115404 74670
rect 115600 74870 115812 74876
rect 115600 74806 115606 74870
rect 115670 74806 115812 74870
rect 115600 74734 115812 74806
rect 115600 74670 115606 74734
rect 115670 74670 115812 74734
rect 115600 74664 115812 74670
rect 116008 74740 116220 74876
rect 116416 74870 116628 74876
rect 116416 74806 116558 74870
rect 116622 74806 116628 74870
rect 116416 74740 116628 74806
rect 116008 74734 116628 74740
rect 116008 74670 116014 74734
rect 116078 74670 116628 74734
rect 116008 74664 116628 74670
rect 116824 74870 117036 74876
rect 116824 74806 116966 74870
rect 117030 74806 117036 74870
rect 116824 74734 117036 74806
rect 116824 74670 116966 74734
rect 117030 74670 117036 74734
rect 116824 74664 117036 74670
rect 116144 74604 116220 74664
rect 116144 74528 116492 74604
rect 28288 74468 28364 74528
rect 110296 74468 110372 74528
rect 116416 74468 116492 74528
rect 1768 74328 1980 74468
rect 1768 74272 1798 74328
rect 1854 74272 1980 74328
rect 1768 74196 1980 74272
rect 21760 74462 21972 74468
rect 21760 74398 21766 74462
rect 21830 74398 21972 74462
rect 21760 74326 21972 74398
rect 21760 74262 21766 74326
rect 21830 74262 21972 74326
rect 21760 74256 21972 74262
rect 22168 74462 22380 74468
rect 22478 74462 22788 74468
rect 22168 74398 22174 74462
rect 22238 74398 22380 74462
rect 22440 74398 22446 74462
rect 22510 74398 22788 74462
rect 22168 74256 22380 74398
rect 22478 74392 22788 74398
rect 22576 74326 22788 74392
rect 22576 74262 22582 74326
rect 22646 74262 22788 74326
rect 22576 74256 22788 74262
rect 22984 74462 23196 74468
rect 22984 74398 23126 74462
rect 23190 74398 23196 74462
rect 22984 74326 23196 74398
rect 22984 74262 22990 74326
rect 23054 74262 23196 74326
rect 22984 74256 23196 74262
rect 23392 74462 23604 74468
rect 23392 74398 23398 74462
rect 23462 74398 23604 74462
rect 23392 74326 23604 74398
rect 23392 74262 23398 74326
rect 23462 74262 23604 74326
rect 23392 74256 23604 74262
rect 28288 74256 28636 74468
rect 110160 74256 110508 74468
rect 115192 74462 115404 74468
rect 115192 74398 115198 74462
rect 115262 74398 115404 74462
rect 115192 74326 115404 74398
rect 115192 74262 115198 74326
rect 115262 74262 115404 74326
rect 115192 74256 115404 74262
rect 115600 74462 115812 74468
rect 115600 74398 115606 74462
rect 115670 74398 115812 74462
rect 115600 74326 115812 74398
rect 115600 74262 115606 74326
rect 115670 74262 115812 74326
rect 115600 74256 115812 74262
rect 116008 74462 116220 74468
rect 116008 74398 116014 74462
rect 116078 74398 116220 74462
rect 116008 74326 116220 74398
rect 116008 74262 116014 74326
rect 116078 74262 116220 74326
rect 116008 74256 116220 74262
rect 116416 74256 116628 74468
rect 116824 74462 117036 74468
rect 116824 74398 116966 74462
rect 117030 74398 117036 74462
rect 116824 74326 117036 74398
rect 116824 74262 116966 74326
rect 117030 74262 117036 74326
rect 116824 74256 117036 74262
rect 136816 74332 137028 74468
rect 136816 74328 137572 74332
rect 136816 74272 136944 74328
rect 137000 74326 137572 74328
rect 137000 74272 137502 74326
rect 136816 74262 137502 74272
rect 137566 74262 137572 74326
rect 136816 74256 137572 74262
rect 28424 74196 28500 74256
rect 110432 74196 110508 74256
rect 1224 74190 1980 74196
rect 1224 74126 1230 74190
rect 1294 74126 1980 74190
rect 1224 74120 1980 74126
rect 21760 74054 21972 74060
rect 21760 73990 21766 74054
rect 21830 73990 21972 74054
rect 21760 73848 21972 73990
rect 22168 73924 22380 74060
rect 22576 74054 22788 74060
rect 22576 73990 22582 74054
rect 22646 73990 22788 74054
rect 22576 73924 22788 73990
rect 22168 73918 22788 73924
rect 22168 73854 22718 73918
rect 22782 73854 22788 73918
rect 22168 73848 22788 73854
rect 22984 74054 23196 74060
rect 22984 73990 22990 74054
rect 23054 73990 23196 74054
rect 22984 73918 23196 73990
rect 22984 73854 22990 73918
rect 23054 73854 23196 73918
rect 22984 73848 23196 73854
rect 23392 74054 23604 74060
rect 23392 73990 23398 74054
rect 23462 73990 23604 74054
rect 23392 73918 23604 73990
rect 28288 73984 28636 74196
rect 110160 73984 110508 74196
rect 136816 74120 137028 74256
rect 28424 73924 28500 73984
rect 110432 73924 110508 73984
rect 23392 73854 23398 73918
rect 23462 73854 23604 73918
rect 23392 73848 23604 73854
rect 21896 73788 21972 73848
rect 21760 73510 21972 73788
rect 28288 73712 28636 73924
rect 110160 73712 110508 73924
rect 115192 74054 115404 74060
rect 115192 73990 115198 74054
rect 115262 73990 115404 74054
rect 115192 73918 115404 73990
rect 115192 73854 115198 73918
rect 115262 73854 115404 73918
rect 115192 73848 115404 73854
rect 115600 74054 115812 74060
rect 115600 73990 115606 74054
rect 115670 73990 115812 74054
rect 115600 73918 115812 73990
rect 115600 73854 115606 73918
rect 115670 73854 115812 73918
rect 115600 73848 115812 73854
rect 116008 74054 116220 74060
rect 116008 73990 116014 74054
rect 116078 73990 116220 74054
rect 116008 73924 116220 73990
rect 116416 73924 116628 74060
rect 116008 73918 116628 73924
rect 116008 73854 116150 73918
rect 116214 73854 116628 73918
rect 116008 73848 116628 73854
rect 116824 74054 117036 74060
rect 116824 73990 116966 74054
rect 117030 73990 117036 74054
rect 116824 73848 117036 73990
rect 28560 73652 28636 73712
rect 110432 73652 110508 73712
rect 116824 73788 116900 73848
rect 21760 73446 21902 73510
rect 21966 73446 21972 73510
rect 21760 73440 21972 73446
rect 22168 73516 22380 73652
rect 22576 73646 22788 73652
rect 22576 73582 22718 73646
rect 22782 73582 22788 73646
rect 22576 73516 22788 73582
rect 22168 73510 22788 73516
rect 22168 73446 22174 73510
rect 22238 73446 22788 73510
rect 22168 73440 22788 73446
rect 22984 73646 23196 73652
rect 22984 73582 22990 73646
rect 23054 73582 23196 73646
rect 22984 73510 23196 73582
rect 22984 73446 22990 73510
rect 23054 73446 23196 73510
rect 22984 73440 23196 73446
rect 23392 73646 23604 73652
rect 23392 73582 23398 73646
rect 23462 73582 23604 73646
rect 23392 73510 23604 73582
rect 23392 73446 23534 73510
rect 23598 73446 23604 73510
rect 23392 73440 23604 73446
rect 28288 73440 28636 73652
rect 110160 73440 110508 73652
rect 115192 73646 115404 73652
rect 115192 73582 115198 73646
rect 115262 73582 115404 73646
rect 115192 73510 115404 73582
rect 115192 73446 115334 73510
rect 115398 73446 115404 73510
rect 115192 73440 115404 73446
rect 115600 73646 115812 73652
rect 115600 73582 115606 73646
rect 115670 73582 115812 73646
rect 115600 73510 115812 73582
rect 115600 73446 115742 73510
rect 115806 73446 115812 73510
rect 115600 73440 115812 73446
rect 116008 73646 116220 73652
rect 116008 73582 116150 73646
rect 116214 73582 116220 73646
rect 116008 73516 116220 73582
rect 116416 73516 116628 73652
rect 116008 73510 116628 73516
rect 116008 73446 116014 73510
rect 116078 73446 116628 73510
rect 116008 73440 116628 73446
rect 116824 73510 117036 73788
rect 116824 73446 116830 73510
rect 116894 73446 117036 73510
rect 116824 73440 117036 73446
rect 22304 73380 22380 73440
rect 28560 73380 28636 73440
rect 110296 73380 110372 73440
rect 22304 73304 22652 73380
rect 22576 73244 22652 73304
rect 21760 73238 21972 73244
rect 21760 73174 21902 73238
rect 21966 73174 21972 73238
rect 21760 73032 21972 73174
rect 22168 73238 22380 73244
rect 22168 73174 22174 73238
rect 22238 73174 22380 73238
rect 22168 73032 22380 73174
rect 22576 73108 22788 73244
rect 22478 73102 22788 73108
rect 22440 73038 22446 73102
rect 22510 73038 22788 73102
rect 22478 73032 22788 73038
rect 22984 73238 23196 73244
rect 22984 73174 22990 73238
rect 23054 73174 23196 73238
rect 22984 73102 23196 73174
rect 22984 73038 22990 73102
rect 23054 73038 23196 73102
rect 22984 73032 23196 73038
rect 23392 73238 23604 73244
rect 23392 73174 23534 73238
rect 23598 73174 23604 73238
rect 23392 73102 23604 73174
rect 28288 73168 28636 73380
rect 110160 73168 110508 73380
rect 28424 73108 28500 73168
rect 110432 73108 110508 73168
rect 23392 73038 23398 73102
rect 23462 73038 23604 73102
rect 23392 73032 23604 73038
rect 21896 72972 21972 73032
rect 21760 72830 21972 72972
rect 28288 72966 28636 73108
rect 28288 72902 28430 72966
rect 28494 72902 28636 72966
rect 28288 72896 28636 72902
rect 28560 72836 28636 72896
rect 21760 72766 21902 72830
rect 21966 72766 21972 72830
rect 21760 72760 21972 72766
rect 22168 72830 22516 72836
rect 22168 72766 22446 72830
rect 22510 72766 22516 72830
rect 22168 72760 22516 72766
rect 22168 72700 22380 72760
rect 1224 72694 1980 72700
rect 1224 72630 1230 72694
rect 1294 72648 1980 72694
rect 1294 72630 1798 72648
rect 1224 72624 1798 72630
rect 1768 72592 1798 72624
rect 1854 72592 1980 72648
rect 22168 72624 22516 72700
rect 22576 72624 22788 72836
rect 1768 72488 1980 72592
rect 22304 72564 22380 72624
rect 21760 72558 21972 72564
rect 21760 72494 21902 72558
rect 21966 72494 21972 72558
rect 21760 72422 21972 72494
rect 21760 72358 21766 72422
rect 21830 72358 21972 72422
rect 21760 72352 21972 72358
rect 22168 72422 22380 72564
rect 22440 72564 22516 72624
rect 22712 72564 22788 72624
rect 22440 72488 22788 72564
rect 22168 72358 22174 72422
rect 22238 72358 22380 72422
rect 22168 72352 22380 72358
rect 22576 72422 22788 72488
rect 22576 72358 22582 72422
rect 22646 72358 22788 72422
rect 22576 72352 22788 72358
rect 22984 72830 23196 72836
rect 22984 72766 22990 72830
rect 23054 72766 23196 72830
rect 22984 72624 23196 72766
rect 23392 72830 23604 72836
rect 23392 72766 23398 72830
rect 23462 72766 23604 72830
rect 23392 72624 23604 72766
rect 28288 72694 28636 72836
rect 28288 72630 28430 72694
rect 28494 72630 28636 72694
rect 22984 72564 23060 72624
rect 23392 72564 23468 72624
rect 22984 72216 23196 72564
rect 23392 72216 23604 72564
rect 28288 72558 28636 72630
rect 28288 72494 28430 72558
rect 28494 72494 28636 72558
rect 28288 72488 28636 72494
rect 110160 72896 110508 73108
rect 115192 73238 115404 73244
rect 115192 73174 115334 73238
rect 115398 73174 115404 73238
rect 115192 73102 115404 73174
rect 115192 73038 115334 73102
rect 115398 73038 115404 73102
rect 115192 73032 115404 73038
rect 115600 73238 115812 73244
rect 115600 73174 115742 73238
rect 115806 73174 115812 73238
rect 115600 73102 115812 73174
rect 115600 73038 115742 73102
rect 115806 73038 115812 73102
rect 115600 73032 115812 73038
rect 116008 73238 116220 73244
rect 116008 73174 116014 73238
rect 116078 73174 116220 73238
rect 116008 73108 116220 73174
rect 116416 73108 116628 73244
rect 116008 73102 116628 73108
rect 116008 73038 116014 73102
rect 116078 73038 116422 73102
rect 116486 73038 116628 73102
rect 116008 73032 116628 73038
rect 116824 73238 117036 73244
rect 116824 73174 116830 73238
rect 116894 73174 117036 73238
rect 116824 73032 117036 73174
rect 116960 72972 117036 73032
rect 110160 72836 110236 72896
rect 110160 72558 110508 72836
rect 110160 72494 110438 72558
rect 110502 72494 110508 72558
rect 110160 72488 110508 72494
rect 115192 72830 115404 72836
rect 115192 72766 115334 72830
rect 115398 72766 115404 72830
rect 115192 72624 115404 72766
rect 115600 72830 115812 72836
rect 115600 72766 115742 72830
rect 115806 72766 115812 72830
rect 115600 72624 115812 72766
rect 116008 72830 116220 72836
rect 116008 72766 116014 72830
rect 116078 72766 116220 72830
rect 116008 72624 116220 72766
rect 116416 72830 116628 72836
rect 116416 72766 116422 72830
rect 116486 72766 116628 72830
rect 116416 72624 116628 72766
rect 116824 72830 117036 72972
rect 116824 72766 116966 72830
rect 117030 72766 117036 72830
rect 116824 72760 117036 72766
rect 136816 72694 137572 72700
rect 136816 72648 137502 72694
rect 115192 72564 115268 72624
rect 115600 72564 115676 72624
rect 116144 72564 116220 72624
rect 136816 72592 136944 72648
rect 137000 72630 137502 72648
rect 137566 72630 137572 72694
rect 137000 72624 137572 72630
rect 137000 72592 137028 72624
rect 23120 72156 23196 72216
rect 23528 72156 23604 72216
rect 21760 72150 21972 72156
rect 21760 72086 21766 72150
rect 21830 72086 21972 72150
rect 21760 72014 21972 72086
rect 21760 71950 21902 72014
rect 21966 71950 21972 72014
rect 21760 71944 21972 71950
rect 22168 72150 22380 72156
rect 22168 72086 22174 72150
rect 22238 72086 22380 72150
rect 22168 71808 22380 72086
rect 22576 72150 22788 72156
rect 22576 72086 22582 72150
rect 22646 72086 22788 72150
rect 22576 71808 22788 72086
rect 22984 71808 23196 72156
rect 22304 71748 22380 71808
rect 23120 71748 23196 71808
rect 21760 71742 21972 71748
rect 21760 71678 21902 71742
rect 21966 71678 21972 71742
rect 21760 71606 21972 71678
rect 21760 71542 21902 71606
rect 21966 71542 21972 71606
rect 21760 71536 21972 71542
rect 22168 71672 22788 71748
rect 22168 71536 22380 71672
rect 22576 71612 22788 71672
rect 22478 71606 22788 71612
rect 22440 71542 22446 71606
rect 22510 71542 22718 71606
rect 22782 71542 22788 71606
rect 22478 71536 22788 71542
rect 22984 71606 23196 71748
rect 22984 71542 22990 71606
rect 23054 71542 23196 71606
rect 22984 71536 23196 71542
rect 23392 71808 23604 72156
rect 28288 72286 28636 72292
rect 28288 72222 28430 72286
rect 28494 72222 28636 72286
rect 28288 72150 28636 72222
rect 28288 72086 28294 72150
rect 28358 72086 28636 72150
rect 28288 71878 28636 72086
rect 28288 71814 28294 71878
rect 28358 71814 28636 71878
rect 23392 71748 23468 71808
rect 23392 71606 23604 71748
rect 28288 71672 28636 71814
rect 28560 71612 28636 71672
rect 23392 71542 23534 71606
rect 23598 71542 23604 71606
rect 23392 71536 23604 71542
rect 21760 71334 21972 71340
rect 21760 71270 21902 71334
rect 21966 71270 21972 71334
rect 21760 71198 21972 71270
rect 21760 71134 21766 71198
rect 21830 71134 21972 71198
rect 21760 71128 21972 71134
rect 22168 71334 22516 71340
rect 22168 71270 22446 71334
rect 22510 71270 22516 71334
rect 22168 71264 22516 71270
rect 22576 71334 22788 71340
rect 22576 71270 22718 71334
rect 22782 71270 22788 71334
rect 22168 71198 22380 71264
rect 22168 71134 22174 71198
rect 22238 71134 22380 71198
rect 22168 71128 22380 71134
rect 22576 71198 22788 71270
rect 22576 71134 22582 71198
rect 22646 71134 22788 71198
rect 22576 71128 22788 71134
rect 22984 71334 23196 71340
rect 22984 71270 22990 71334
rect 23054 71270 23196 71334
rect 22984 71198 23196 71270
rect 22984 71134 22990 71198
rect 23054 71134 23196 71198
rect 22984 71128 23196 71134
rect 23392 71334 23604 71340
rect 23392 71270 23534 71334
rect 23598 71270 23604 71334
rect 23392 71198 23604 71270
rect 23392 71134 23534 71198
rect 23598 71134 23604 71198
rect 23392 71128 23604 71134
rect 28288 71128 28636 71612
rect 110160 72286 110508 72292
rect 110160 72222 110438 72286
rect 110502 72222 110508 72286
rect 110160 71672 110508 72222
rect 115192 72216 115404 72564
rect 115600 72216 115812 72564
rect 116008 72422 116220 72564
rect 116008 72358 116014 72422
rect 116078 72358 116220 72422
rect 116008 72352 116220 72358
rect 116416 72352 116628 72564
rect 116824 72558 117036 72564
rect 116824 72494 116966 72558
rect 117030 72494 117036 72558
rect 116824 72422 117036 72494
rect 136816 72488 137028 72592
rect 116824 72358 116830 72422
rect 116894 72358 117036 72422
rect 116824 72352 117036 72358
rect 116416 72292 116492 72352
rect 115328 72156 115404 72216
rect 115736 72156 115812 72216
rect 116144 72216 116492 72292
rect 116144 72156 116220 72216
rect 115192 71808 115404 72156
rect 115600 71808 115812 72156
rect 116008 72150 116628 72156
rect 116008 72086 116014 72150
rect 116078 72086 116628 72150
rect 116008 72080 116628 72086
rect 116008 71808 116220 72080
rect 116416 71808 116628 72080
rect 116824 72150 117036 72156
rect 116824 72086 116830 72150
rect 116894 72086 117036 72150
rect 116824 72014 117036 72086
rect 116824 71950 116830 72014
rect 116894 71950 117036 72014
rect 116824 71944 117036 71950
rect 115192 71748 115268 71808
rect 115600 71748 115676 71808
rect 116416 71748 116492 71808
rect 110160 71612 110236 71672
rect 110160 71128 110508 71612
rect 115192 71606 115404 71748
rect 115192 71542 115198 71606
rect 115262 71542 115404 71606
rect 115192 71536 115404 71542
rect 115600 71606 115812 71748
rect 115600 71542 115742 71606
rect 115806 71542 115812 71606
rect 115600 71536 115812 71542
rect 116008 71672 116628 71748
rect 116008 71612 116220 71672
rect 116008 71606 116356 71612
rect 116008 71542 116014 71606
rect 116078 71542 116286 71606
rect 116350 71542 116356 71606
rect 116008 71536 116356 71542
rect 116416 71536 116628 71672
rect 116824 71742 117036 71748
rect 116824 71678 116830 71742
rect 116894 71678 117036 71742
rect 116824 71606 117036 71678
rect 116824 71542 116830 71606
rect 116894 71542 117036 71606
rect 116824 71536 117036 71542
rect 115192 71334 115404 71340
rect 115192 71270 115198 71334
rect 115262 71270 115404 71334
rect 115192 71198 115404 71270
rect 115192 71134 115334 71198
rect 115398 71134 115404 71198
rect 115192 71128 115404 71134
rect 115600 71334 115812 71340
rect 115600 71270 115742 71334
rect 115806 71270 115812 71334
rect 115600 71198 115812 71270
rect 115600 71134 115742 71198
rect 115806 71134 115812 71198
rect 115600 71128 115812 71134
rect 116008 71334 116220 71340
rect 116318 71334 116628 71340
rect 116008 71270 116014 71334
rect 116078 71270 116220 71334
rect 116280 71270 116286 71334
rect 116350 71270 116628 71334
rect 116008 71128 116220 71270
rect 116318 71264 116628 71270
rect 116416 71204 116628 71264
rect 116318 71198 116628 71204
rect 116280 71134 116286 71198
rect 116350 71134 116628 71198
rect 116318 71128 116628 71134
rect 116824 71334 117036 71340
rect 116824 71270 116830 71334
rect 116894 71270 117036 71334
rect 116824 71198 117036 71270
rect 116824 71134 116830 71198
rect 116894 71134 117036 71198
rect 116824 71128 117036 71134
rect 28288 71068 28364 71128
rect 110432 71068 110508 71128
rect 1224 71062 1980 71068
rect 1224 70998 1230 71062
rect 1294 70998 1980 71062
rect 1224 70992 1980 70998
rect 1768 70968 1980 70992
rect 1768 70912 1798 70968
rect 1854 70912 1980 70968
rect 1768 70856 1980 70912
rect 21760 70926 21972 70932
rect 21760 70862 21766 70926
rect 21830 70862 21972 70926
rect 21760 70790 21972 70862
rect 21760 70726 21902 70790
rect 21966 70726 21972 70790
rect 21760 70720 21972 70726
rect 22168 70926 22380 70932
rect 22168 70862 22174 70926
rect 22238 70862 22380 70926
rect 22168 70720 22380 70862
rect 22576 70926 22788 70932
rect 22576 70862 22582 70926
rect 22646 70862 22788 70926
rect 22576 70790 22788 70862
rect 22576 70726 22718 70790
rect 22782 70726 22788 70790
rect 22576 70720 22788 70726
rect 22984 70926 23196 70932
rect 22984 70862 22990 70926
rect 23054 70862 23196 70926
rect 22984 70790 23196 70862
rect 22984 70726 23126 70790
rect 23190 70726 23196 70790
rect 22984 70720 23196 70726
rect 23392 70926 23604 70932
rect 23392 70862 23534 70926
rect 23598 70862 23604 70926
rect 23392 70790 23604 70862
rect 28288 70856 28636 71068
rect 110160 70856 110508 71068
rect 136816 71062 137572 71068
rect 136816 70998 137502 71062
rect 137566 70998 137572 71062
rect 136816 70992 137572 70998
rect 136816 70968 137028 70992
rect 28560 70796 28636 70856
rect 110432 70796 110508 70856
rect 23392 70726 23398 70790
rect 23462 70726 23604 70790
rect 23392 70720 23604 70726
rect 25160 70584 27004 70660
rect 28288 70584 28636 70796
rect 25160 70524 25236 70584
rect 26928 70524 27004 70584
rect 28560 70524 28636 70584
rect 21760 70518 21972 70524
rect 21760 70454 21902 70518
rect 21966 70454 21972 70518
rect 21760 70382 21972 70454
rect 21760 70318 21902 70382
rect 21966 70318 21972 70382
rect 21760 70312 21972 70318
rect 22168 70518 22788 70524
rect 22168 70454 22718 70518
rect 22782 70454 22788 70518
rect 22168 70448 22788 70454
rect 22168 70388 22380 70448
rect 22168 70382 22516 70388
rect 22168 70318 22446 70382
rect 22510 70318 22516 70382
rect 22168 70312 22516 70318
rect 22576 70312 22788 70448
rect 22984 70518 23196 70524
rect 22984 70454 23126 70518
rect 23190 70454 23196 70518
rect 22984 70382 23196 70454
rect 22984 70318 23126 70382
rect 23190 70318 23196 70382
rect 22984 70312 23196 70318
rect 23392 70518 23604 70524
rect 23392 70454 23398 70518
rect 23462 70454 23604 70518
rect 23392 70382 23604 70454
rect 23392 70318 23534 70382
rect 23598 70318 23604 70382
rect 23392 70312 23604 70318
rect 23800 70388 24012 70524
rect 24208 70448 25236 70524
rect 23800 70312 24148 70388
rect 24208 70382 24556 70448
rect 24208 70318 24214 70382
rect 24278 70318 24556 70382
rect 24208 70312 24556 70318
rect 25296 70388 25508 70524
rect 25296 70312 26868 70388
rect 26928 70312 27140 70524
rect 28288 70388 28636 70524
rect 28152 70312 28636 70388
rect 110160 70584 110508 70796
rect 115192 70926 115404 70932
rect 115192 70862 115334 70926
rect 115398 70862 115404 70926
rect 115192 70790 115404 70862
rect 115192 70726 115198 70790
rect 115262 70726 115404 70790
rect 115192 70720 115404 70726
rect 115600 70926 115812 70932
rect 115600 70862 115742 70926
rect 115806 70862 115812 70926
rect 115600 70790 115812 70862
rect 115600 70726 115606 70790
rect 115670 70726 115812 70790
rect 115600 70720 115812 70726
rect 116008 70926 116356 70932
rect 116008 70862 116286 70926
rect 116350 70862 116356 70926
rect 116008 70856 116356 70862
rect 116008 70796 116220 70856
rect 116416 70796 116628 70932
rect 116008 70790 116628 70796
rect 116008 70726 116558 70790
rect 116622 70726 116628 70790
rect 116008 70720 116628 70726
rect 116824 70926 117036 70932
rect 116824 70862 116830 70926
rect 116894 70862 117036 70926
rect 116824 70790 117036 70862
rect 136816 70912 136944 70968
rect 137000 70912 137028 70968
rect 136816 70856 137028 70912
rect 116824 70726 116966 70790
rect 117030 70726 117036 70790
rect 116824 70720 117036 70726
rect 114240 70584 114860 70660
rect 110160 70524 110236 70584
rect 114240 70524 114316 70584
rect 114784 70524 114860 70584
rect 115056 70584 115676 70660
rect 115056 70524 115132 70584
rect 115600 70524 115676 70584
rect 110160 70312 110508 70524
rect 111656 70388 111868 70524
rect 113288 70448 114316 70524
rect 111656 70312 113228 70388
rect 113288 70382 113500 70448
rect 113288 70318 113294 70382
rect 113358 70318 113500 70382
rect 113288 70312 113500 70318
rect 114376 70388 114588 70524
rect 114784 70448 115132 70524
rect 115192 70518 115404 70524
rect 115192 70454 115198 70518
rect 115262 70454 115404 70518
rect 114376 70312 114724 70388
rect 114784 70312 114996 70448
rect 115192 70382 115404 70454
rect 115192 70318 115198 70382
rect 115262 70318 115404 70382
rect 115192 70312 115404 70318
rect 115600 70518 115812 70524
rect 115600 70454 115606 70518
rect 115670 70454 115812 70518
rect 115600 70382 115812 70454
rect 115600 70318 115742 70382
rect 115806 70318 115812 70382
rect 115600 70312 115812 70318
rect 116008 70388 116220 70524
rect 116416 70518 116628 70524
rect 116416 70454 116558 70518
rect 116622 70454 116628 70518
rect 116416 70388 116628 70454
rect 116008 70382 116628 70388
rect 116008 70318 116150 70382
rect 116214 70318 116628 70382
rect 116008 70312 116628 70318
rect 116824 70518 117036 70524
rect 116824 70454 116966 70518
rect 117030 70454 117036 70518
rect 116824 70382 117036 70454
rect 116824 70318 116966 70382
rect 117030 70318 117036 70382
rect 116824 70312 117036 70318
rect 23800 70252 23876 70312
rect 23256 70176 23876 70252
rect 24072 70252 24148 70312
rect 25296 70252 25372 70312
rect 24072 70176 25372 70252
rect 26792 70252 26868 70312
rect 28152 70252 28228 70312
rect 28560 70252 28636 70312
rect 110296 70252 110372 70312
rect 113152 70252 113228 70312
rect 114376 70252 114452 70312
rect 26792 70176 28228 70252
rect 23256 70116 23332 70176
rect 21760 70110 21972 70116
rect 21760 70046 21902 70110
rect 21966 70046 21972 70110
rect 21760 69904 21972 70046
rect 22168 69974 22380 70116
rect 22478 70110 22788 70116
rect 22440 70046 22446 70110
rect 22510 70046 22788 70110
rect 22478 70040 22788 70046
rect 22168 69910 22174 69974
rect 22238 69910 22380 69974
rect 22168 69904 22380 69910
rect 22576 69974 22788 70040
rect 22576 69910 22582 69974
rect 22646 69910 22788 69974
rect 22576 69904 22788 69910
rect 22984 70110 23332 70116
rect 22984 70046 23126 70110
rect 23190 70046 23332 70110
rect 22984 70040 23332 70046
rect 23392 70110 24284 70116
rect 23392 70046 23534 70110
rect 23598 70046 24214 70110
rect 24278 70046 24284 70110
rect 23392 70040 24284 70046
rect 28288 70040 28636 70252
rect 110160 70040 110508 70252
rect 113152 70176 114452 70252
rect 114648 70252 114724 70312
rect 115192 70252 115268 70312
rect 116144 70252 116220 70312
rect 114648 70176 115268 70252
rect 115464 70176 116084 70252
rect 116144 70176 116492 70252
rect 115464 70116 115540 70176
rect 116008 70116 116084 70176
rect 116416 70116 116492 70176
rect 115192 70110 115540 70116
rect 115192 70046 115198 70110
rect 115262 70046 115540 70110
rect 115192 70040 115540 70046
rect 115600 70110 115812 70116
rect 115600 70046 115742 70110
rect 115806 70046 115812 70110
rect 22984 69974 23196 70040
rect 22984 69910 22990 69974
rect 23054 69910 23196 69974
rect 22984 69904 23196 69910
rect 23392 69974 23604 70040
rect 28424 69980 28500 70040
rect 110296 69980 110372 70040
rect 23392 69910 23398 69974
rect 23462 69910 23604 69974
rect 23392 69904 23604 69910
rect 21760 69844 21836 69904
rect 21760 69566 21972 69844
rect 28288 69768 28636 69980
rect 110160 69768 110508 69980
rect 115192 69974 115404 70040
rect 115192 69910 115198 69974
rect 115262 69910 115404 69974
rect 115192 69904 115404 69910
rect 115600 69974 115812 70046
rect 115600 69910 115606 69974
rect 115670 69910 115812 69974
rect 115600 69904 115812 69910
rect 116008 70110 116220 70116
rect 116008 70046 116150 70110
rect 116214 70046 116220 70110
rect 116008 69974 116220 70046
rect 116008 69910 116014 69974
rect 116078 69910 116220 69974
rect 116008 69904 116220 69910
rect 116416 69974 116628 70116
rect 116416 69910 116558 69974
rect 116622 69910 116628 69974
rect 116416 69904 116628 69910
rect 116824 70110 117036 70116
rect 116824 70046 116966 70110
rect 117030 70046 117036 70110
rect 116824 69904 117036 70046
rect 116824 69844 116900 69904
rect 28424 69708 28500 69768
rect 110160 69708 110236 69768
rect 21760 69502 21902 69566
rect 21966 69502 21972 69566
rect 21760 69496 21972 69502
rect 22168 69702 22788 69708
rect 22168 69638 22174 69702
rect 22238 69638 22582 69702
rect 22646 69638 22788 69702
rect 22168 69632 22788 69638
rect 22168 69496 22380 69632
rect 22576 69572 22788 69632
rect 22478 69566 22788 69572
rect 22440 69502 22446 69566
rect 22510 69502 22788 69566
rect 22478 69496 22788 69502
rect 22984 69702 23196 69708
rect 22984 69638 22990 69702
rect 23054 69638 23196 69702
rect 22984 69566 23196 69638
rect 22984 69502 22990 69566
rect 23054 69502 23196 69566
rect 22984 69496 23196 69502
rect 23392 69702 23604 69708
rect 23392 69638 23398 69702
rect 23462 69638 23604 69702
rect 23392 69566 23604 69638
rect 23392 69502 23398 69566
rect 23462 69502 23604 69566
rect 23392 69496 23604 69502
rect 28288 69496 28636 69708
rect 110160 69702 113364 69708
rect 110160 69638 113294 69702
rect 113358 69638 113364 69702
rect 110160 69632 113364 69638
rect 115192 69702 115404 69708
rect 115192 69638 115198 69702
rect 115262 69638 115404 69702
rect 110160 69496 110508 69632
rect 115192 69566 115404 69638
rect 115192 69502 115198 69566
rect 115262 69502 115404 69566
rect 115192 69496 115404 69502
rect 115600 69702 115812 69708
rect 115600 69638 115606 69702
rect 115670 69638 115812 69702
rect 115600 69566 115812 69638
rect 115600 69502 115606 69566
rect 115670 69502 115812 69566
rect 115600 69496 115812 69502
rect 116008 69702 116220 69708
rect 116008 69638 116014 69702
rect 116078 69638 116220 69702
rect 116008 69566 116220 69638
rect 116008 69502 116150 69566
rect 116214 69502 116220 69566
rect 116008 69496 116220 69502
rect 116416 69702 116628 69708
rect 116416 69638 116558 69702
rect 116622 69638 116628 69702
rect 116416 69496 116628 69638
rect 116824 69566 117036 69844
rect 116824 69502 116830 69566
rect 116894 69502 117036 69566
rect 116824 69496 117036 69502
rect 22304 69436 22380 69496
rect 28288 69436 28364 69496
rect 110432 69436 110508 69496
rect 1768 69300 1980 69436
rect 22304 69360 22652 69436
rect 22576 69300 22652 69360
rect 1224 69294 1980 69300
rect 1224 69230 1230 69294
rect 1294 69288 1980 69294
rect 1294 69232 1798 69288
rect 1854 69232 1980 69288
rect 1294 69230 1980 69232
rect 1224 69224 1980 69230
rect 1768 69088 1980 69224
rect 21760 69294 21972 69300
rect 21760 69230 21902 69294
rect 21966 69230 21972 69294
rect 21760 69088 21972 69230
rect 22168 69294 22516 69300
rect 22168 69230 22446 69294
rect 22510 69230 22516 69294
rect 22168 69224 22516 69230
rect 22168 69088 22380 69224
rect 22576 69158 22788 69300
rect 22576 69094 22582 69158
rect 22646 69094 22788 69158
rect 22576 69088 22788 69094
rect 22984 69294 23196 69300
rect 22984 69230 22990 69294
rect 23054 69230 23196 69294
rect 22984 69158 23196 69230
rect 22984 69094 23126 69158
rect 23190 69094 23196 69158
rect 22984 69088 23196 69094
rect 23392 69294 23604 69300
rect 23392 69230 23398 69294
rect 23462 69230 23604 69294
rect 23392 69158 23604 69230
rect 23392 69094 23534 69158
rect 23598 69094 23604 69158
rect 23392 69088 23604 69094
rect 28288 69224 28636 69436
rect 110160 69224 110508 69436
rect 136816 69300 137028 69436
rect 115192 69294 115404 69300
rect 115192 69230 115198 69294
rect 115262 69230 115404 69294
rect 28288 69164 28364 69224
rect 110296 69164 110372 69224
rect 21760 69028 21836 69088
rect 21760 68886 21972 69028
rect 28288 69022 28636 69164
rect 28288 68958 28294 69022
rect 28358 68958 28636 69022
rect 28288 68952 28636 68958
rect 110160 69022 110508 69164
rect 115192 69158 115404 69230
rect 115192 69094 115334 69158
rect 115398 69094 115404 69158
rect 115192 69088 115404 69094
rect 115600 69294 115812 69300
rect 115600 69230 115606 69294
rect 115670 69230 115812 69294
rect 115600 69158 115812 69230
rect 115600 69094 115742 69158
rect 115806 69094 115812 69158
rect 115600 69088 115812 69094
rect 116008 69294 116628 69300
rect 116008 69230 116150 69294
rect 116214 69230 116628 69294
rect 116008 69224 116628 69230
rect 116008 69164 116220 69224
rect 116008 69158 116356 69164
rect 116008 69094 116286 69158
rect 116350 69094 116356 69158
rect 116008 69088 116356 69094
rect 116416 69088 116628 69224
rect 116824 69294 117036 69300
rect 116824 69230 116830 69294
rect 116894 69230 117036 69294
rect 116824 69088 117036 69230
rect 136816 69294 137572 69300
rect 136816 69288 137502 69294
rect 136816 69232 136944 69288
rect 137000 69232 137502 69288
rect 136816 69230 137502 69232
rect 137566 69230 137572 69294
rect 136816 69224 137572 69230
rect 136816 69088 137028 69224
rect 110160 68958 110438 69022
rect 110502 68958 110508 69022
rect 110160 68952 110508 68958
rect 116824 69028 116900 69088
rect 28560 68892 28636 68952
rect 110296 68892 110372 68952
rect 21760 68822 21902 68886
rect 21966 68822 21972 68886
rect 21760 68816 21972 68822
rect 22168 68680 22380 68892
rect 22576 68886 22788 68892
rect 22576 68822 22582 68886
rect 22646 68822 22788 68886
rect 22576 68680 22788 68822
rect 22984 68886 23196 68892
rect 22984 68822 23126 68886
rect 23190 68822 23196 68886
rect 22984 68750 23196 68822
rect 22984 68686 23126 68750
rect 23190 68686 23196 68750
rect 22984 68680 23196 68686
rect 23392 68886 23604 68892
rect 23392 68822 23534 68886
rect 23598 68822 23604 68886
rect 23392 68750 23604 68822
rect 23392 68686 23398 68750
rect 23462 68686 23604 68750
rect 23392 68680 23604 68686
rect 28288 68750 28636 68892
rect 28288 68686 28294 68750
rect 28358 68686 28430 68750
rect 28494 68686 28636 68750
rect 22168 68620 22244 68680
rect 22576 68620 22652 68680
rect 21760 68614 21972 68620
rect 21760 68550 21902 68614
rect 21966 68550 21972 68614
rect 21760 68272 21972 68550
rect 22168 68484 22380 68620
rect 22576 68484 22788 68620
rect 22168 68408 22788 68484
rect 22168 68342 22380 68408
rect 22168 68278 22174 68342
rect 22238 68278 22380 68342
rect 22168 68272 22380 68278
rect 22576 68342 22788 68408
rect 22576 68278 22582 68342
rect 22646 68278 22788 68342
rect 22576 68272 22788 68278
rect 22984 68478 23196 68484
rect 22984 68414 23126 68478
rect 23190 68414 23196 68478
rect 22984 68272 23196 68414
rect 21760 68212 21836 68272
rect 23120 68212 23196 68272
rect 21760 68070 21972 68212
rect 21760 68006 21766 68070
rect 21830 68006 21972 68070
rect 21760 68000 21972 68006
rect 22168 68070 22380 68076
rect 22168 68006 22174 68070
rect 22238 68006 22380 68070
rect 22168 67864 22380 68006
rect 22576 68070 22788 68076
rect 22576 68006 22582 68070
rect 22646 68006 22788 68070
rect 22576 67864 22788 68006
rect 22984 67864 23196 68212
rect 23392 68478 23604 68484
rect 23392 68414 23398 68478
rect 23462 68414 23604 68478
rect 23392 68272 23604 68414
rect 28288 68408 28636 68686
rect 110160 68750 110508 68892
rect 110160 68686 110438 68750
rect 110502 68686 110508 68750
rect 110160 68408 110508 68686
rect 115192 68886 115404 68892
rect 115192 68822 115334 68886
rect 115398 68822 115404 68886
rect 115192 68750 115404 68822
rect 115192 68686 115334 68750
rect 115398 68686 115404 68750
rect 115192 68680 115404 68686
rect 115600 68886 115812 68892
rect 115600 68822 115742 68886
rect 115806 68822 115812 68886
rect 115600 68750 115812 68822
rect 115600 68686 115742 68750
rect 115806 68686 115812 68750
rect 115600 68680 115812 68686
rect 116008 68756 116220 68892
rect 116318 68886 116628 68892
rect 116280 68822 116286 68886
rect 116350 68822 116628 68886
rect 116318 68816 116628 68822
rect 116824 68886 117036 69028
rect 116824 68822 116966 68886
rect 117030 68822 117036 68886
rect 116824 68816 117036 68822
rect 116008 68680 116356 68756
rect 116416 68680 116628 68816
rect 116144 68620 116220 68680
rect 110432 68348 110508 68408
rect 28288 68342 28636 68348
rect 28288 68278 28430 68342
rect 28494 68278 28636 68342
rect 23392 68212 23468 68272
rect 23392 67864 23604 68212
rect 22168 67804 22244 67864
rect 22576 67804 22652 67864
rect 23120 67804 23196 67864
rect 23528 67804 23604 67864
rect 21760 67798 21972 67804
rect 21760 67734 21766 67798
rect 21830 67734 21972 67798
rect 1224 67662 1980 67668
rect 1224 67598 1230 67662
rect 1294 67608 1980 67662
rect 1294 67598 1798 67608
rect 1224 67592 1798 67598
rect 1768 67552 1798 67592
rect 1854 67552 1980 67608
rect 21760 67662 21972 67734
rect 21760 67598 21766 67662
rect 21830 67598 21972 67662
rect 21760 67592 21972 67598
rect 22168 67592 22380 67804
rect 22576 67662 22788 67804
rect 22576 67598 22582 67662
rect 22646 67598 22788 67662
rect 22576 67592 22788 67598
rect 1768 67456 1980 67552
rect 22984 67456 23196 67804
rect 23392 67456 23604 67804
rect 28288 67728 28636 68278
rect 110160 68206 110508 68348
rect 110160 68142 110438 68206
rect 110502 68142 110508 68206
rect 110160 67934 110508 68142
rect 110160 67870 110438 67934
rect 110502 67870 110508 67934
rect 110160 67728 110508 67870
rect 115192 68478 115404 68484
rect 115192 68414 115334 68478
rect 115398 68414 115404 68478
rect 115192 68272 115404 68414
rect 115600 68478 115812 68484
rect 115600 68414 115742 68478
rect 115806 68414 115812 68478
rect 115600 68272 115812 68414
rect 116008 68342 116220 68620
rect 116280 68620 116356 68680
rect 116552 68620 116628 68680
rect 116280 68544 116628 68620
rect 116008 68278 116014 68342
rect 116078 68278 116220 68342
rect 116008 68272 116220 68278
rect 116416 68272 116628 68544
rect 116824 68614 117036 68620
rect 116824 68550 116966 68614
rect 117030 68550 117036 68614
rect 116824 68272 117036 68550
rect 115192 68212 115268 68272
rect 115600 68212 115676 68272
rect 116824 68212 116900 68272
rect 115192 67864 115404 68212
rect 115328 67804 115404 67864
rect 28424 67668 28500 67728
rect 110296 67668 110372 67728
rect 28288 67592 28636 67668
rect 110160 67592 110508 67668
rect 22984 67396 23060 67456
rect 23392 67396 23468 67456
rect 28406 67396 28504 67592
rect 110294 67396 110392 67592
rect 115192 67456 115404 67804
rect 115600 67864 115812 68212
rect 116008 68070 116220 68076
rect 116008 68006 116014 68070
rect 116078 68006 116220 68070
rect 116008 67864 116220 68006
rect 116416 67864 116628 68076
rect 116824 68070 117036 68212
rect 116824 68006 116830 68070
rect 116894 68006 117036 68070
rect 116824 68000 117036 68006
rect 115600 67804 115676 67864
rect 116008 67804 116084 67864
rect 116416 67804 116492 67864
rect 115600 67456 115812 67804
rect 116008 67668 116220 67804
rect 116416 67668 116628 67804
rect 116008 67662 116628 67668
rect 116008 67598 116558 67662
rect 116622 67598 116628 67662
rect 116008 67592 116628 67598
rect 116824 67798 117036 67804
rect 116824 67734 116830 67798
rect 116894 67734 117036 67798
rect 116824 67662 117036 67734
rect 116824 67598 116830 67662
rect 116894 67598 117036 67662
rect 116824 67592 117036 67598
rect 136816 67608 137028 67668
rect 136816 67552 136944 67608
rect 137000 67552 137028 67608
rect 136816 67532 137028 67552
rect 136816 67526 137572 67532
rect 136816 67462 137502 67526
rect 137566 67462 137572 67526
rect 136816 67456 137572 67462
rect 115192 67396 115268 67456
rect 115600 67396 115676 67456
rect 21760 67390 21972 67396
rect 21760 67326 21766 67390
rect 21830 67326 21972 67390
rect 21760 67254 21972 67326
rect 21760 67190 21902 67254
rect 21966 67190 21972 67254
rect 21760 67184 21972 67190
rect 22168 67390 22788 67396
rect 22168 67326 22582 67390
rect 22646 67326 22788 67390
rect 22168 67320 22788 67326
rect 22168 67048 22380 67320
rect 22576 67048 22788 67320
rect 22984 67254 23196 67396
rect 22984 67190 22990 67254
rect 23054 67190 23196 67254
rect 22984 67184 23196 67190
rect 23392 67254 23604 67396
rect 23392 67190 23534 67254
rect 23598 67190 23604 67254
rect 23392 67184 23604 67190
rect 28288 67184 28636 67396
rect 110160 67390 110508 67396
rect 110160 67326 110302 67390
rect 110366 67326 110508 67390
rect 110160 67184 110508 67326
rect 115192 67254 115404 67396
rect 115192 67190 115198 67254
rect 115262 67190 115404 67254
rect 115192 67184 115404 67190
rect 115600 67254 115812 67396
rect 115600 67190 115606 67254
rect 115670 67190 115812 67254
rect 115600 67184 115812 67190
rect 116008 67390 116628 67396
rect 116008 67326 116558 67390
rect 116622 67326 116628 67390
rect 116008 67320 116628 67326
rect 28424 67124 28500 67184
rect 110160 67124 110236 67184
rect 116008 67124 116220 67320
rect 22168 66988 22244 67048
rect 22576 66988 22652 67048
rect 21760 66982 21972 66988
rect 21760 66918 21902 66982
rect 21966 66918 21972 66982
rect 21760 66846 21972 66918
rect 21760 66782 21766 66846
rect 21830 66782 21972 66846
rect 21760 66776 21972 66782
rect 22168 66776 22380 66988
rect 22576 66846 22788 66988
rect 22576 66782 22582 66846
rect 22646 66782 22788 66846
rect 22576 66776 22788 66782
rect 22984 66982 23196 66988
rect 22984 66918 22990 66982
rect 23054 66918 23196 66982
rect 22984 66846 23196 66918
rect 22984 66782 22990 66846
rect 23054 66782 23196 66846
rect 22984 66776 23196 66782
rect 23392 66982 23604 66988
rect 23392 66918 23534 66982
rect 23598 66918 23604 66982
rect 23392 66846 23604 66918
rect 28288 66912 28636 67124
rect 110160 67118 110508 67124
rect 110160 67054 110302 67118
rect 110366 67054 110508 67118
rect 110160 66912 110508 67054
rect 116008 67048 116356 67124
rect 116416 67048 116628 67320
rect 116824 67390 117036 67396
rect 116824 67326 116830 67390
rect 116894 67326 117036 67390
rect 116824 67254 117036 67326
rect 116824 67190 116966 67254
rect 117030 67190 117036 67254
rect 116824 67184 117036 67190
rect 116008 66988 116084 67048
rect 116280 66988 116356 67048
rect 28424 66852 28500 66912
rect 110432 66852 110508 66912
rect 23392 66782 23534 66846
rect 23598 66782 23604 66846
rect 23392 66776 23604 66782
rect 28288 66640 28636 66852
rect 110160 66640 110508 66852
rect 115192 66982 115404 66988
rect 115192 66918 115198 66982
rect 115262 66918 115404 66982
rect 115192 66846 115404 66918
rect 115192 66782 115334 66846
rect 115398 66782 115404 66846
rect 115192 66776 115404 66782
rect 115600 66982 115812 66988
rect 115600 66918 115606 66982
rect 115670 66918 115812 66982
rect 115600 66846 115812 66918
rect 115600 66782 115742 66846
rect 115806 66782 115812 66846
rect 115600 66776 115812 66782
rect 116008 66776 116220 66988
rect 116280 66912 116628 66988
rect 116416 66852 116628 66912
rect 116318 66846 116628 66852
rect 116280 66782 116286 66846
rect 116350 66782 116628 66846
rect 116318 66776 116628 66782
rect 116824 66982 117036 66988
rect 116824 66918 116966 66982
rect 117030 66918 117036 66982
rect 116824 66846 117036 66918
rect 116824 66782 116830 66846
rect 116894 66782 117036 66846
rect 116824 66776 117036 66782
rect 28288 66580 28364 66640
rect 110160 66580 110236 66640
rect 21760 66574 21972 66580
rect 21760 66510 21766 66574
rect 21830 66510 21972 66574
rect 21760 66438 21972 66510
rect 21760 66374 21902 66438
rect 21966 66374 21972 66438
rect 21760 66368 21972 66374
rect 22168 66574 22788 66580
rect 22168 66510 22582 66574
rect 22646 66510 22788 66574
rect 22168 66504 22788 66510
rect 22168 66444 22380 66504
rect 22168 66438 22516 66444
rect 22168 66374 22446 66438
rect 22510 66374 22516 66438
rect 22168 66368 22516 66374
rect 22576 66368 22788 66504
rect 22984 66574 23196 66580
rect 22984 66510 22990 66574
rect 23054 66510 23196 66574
rect 22984 66438 23196 66510
rect 22984 66374 23126 66438
rect 23190 66374 23196 66438
rect 22984 66368 23196 66374
rect 23392 66574 23604 66580
rect 23392 66510 23534 66574
rect 23598 66510 23604 66574
rect 23392 66438 23604 66510
rect 23392 66374 23398 66438
rect 23462 66374 23604 66438
rect 23392 66368 23604 66374
rect 28288 66368 28636 66580
rect 110160 66368 110508 66580
rect 115192 66574 115404 66580
rect 115192 66510 115334 66574
rect 115398 66510 115404 66574
rect 115192 66438 115404 66510
rect 115192 66374 115198 66438
rect 115262 66374 115404 66438
rect 115192 66368 115404 66374
rect 115600 66574 115812 66580
rect 115600 66510 115742 66574
rect 115806 66510 115812 66574
rect 115600 66438 115812 66510
rect 115600 66374 115606 66438
rect 115670 66374 115812 66438
rect 115600 66368 115812 66374
rect 116008 66574 116356 66580
rect 116008 66510 116286 66574
rect 116350 66510 116356 66574
rect 116008 66504 116356 66510
rect 116008 66444 116220 66504
rect 116416 66444 116628 66580
rect 116008 66438 116628 66444
rect 116008 66374 116558 66438
rect 116622 66374 116628 66438
rect 116008 66368 116628 66374
rect 116824 66574 117036 66580
rect 116824 66510 116830 66574
rect 116894 66510 117036 66574
rect 116824 66438 117036 66510
rect 116824 66374 116966 66438
rect 117030 66374 117036 66438
rect 116824 66368 117036 66374
rect 28424 66308 28500 66368
rect 110432 66308 110508 66368
rect 21760 66166 21972 66172
rect 21760 66102 21902 66166
rect 21966 66102 21972 66166
rect 1768 65928 1980 66036
rect 21760 66030 21972 66102
rect 21760 65966 21766 66030
rect 21830 65966 21972 66030
rect 21760 65960 21972 65966
rect 22168 66036 22380 66172
rect 22478 66166 22788 66172
rect 22440 66102 22446 66166
rect 22510 66102 22788 66166
rect 22478 66096 22788 66102
rect 22576 66036 22788 66096
rect 22168 66030 22788 66036
rect 22168 65966 22310 66030
rect 22374 65966 22788 66030
rect 22168 65960 22788 65966
rect 22984 66166 23196 66172
rect 22984 66102 23126 66166
rect 23190 66102 23196 66166
rect 22984 66030 23196 66102
rect 22984 65966 23126 66030
rect 23190 65966 23196 66030
rect 22984 65960 23196 65966
rect 23392 66166 23604 66172
rect 23392 66102 23398 66166
rect 23462 66102 23604 66166
rect 23392 66030 23604 66102
rect 28288 66096 28636 66308
rect 110160 66096 110508 66308
rect 115192 66166 115404 66172
rect 115192 66102 115198 66166
rect 115262 66102 115404 66166
rect 28424 66036 28500 66096
rect 110296 66036 110372 66096
rect 23392 65966 23534 66030
rect 23598 65966 23604 66030
rect 23392 65960 23604 65966
rect 1768 65900 1798 65928
rect 1224 65894 1798 65900
rect 1224 65830 1230 65894
rect 1294 65872 1798 65894
rect 1854 65872 1980 65928
rect 1294 65830 1980 65872
rect 1224 65824 1980 65830
rect 22304 65900 22380 65960
rect 22304 65824 22652 65900
rect 22576 65764 22652 65824
rect 28288 65824 28636 66036
rect 110160 65824 110508 66036
rect 115192 66030 115404 66102
rect 115192 65966 115198 66030
rect 115262 65966 115404 66030
rect 115192 65960 115404 65966
rect 115600 66166 115812 66172
rect 115600 66102 115606 66166
rect 115670 66102 115812 66166
rect 115600 66030 115812 66102
rect 115600 65966 115606 66030
rect 115670 65966 115812 66030
rect 115600 65960 115812 65966
rect 116008 66036 116220 66172
rect 116416 66166 116628 66172
rect 116416 66102 116558 66166
rect 116622 66102 116628 66166
rect 116416 66036 116628 66102
rect 116008 66030 116628 66036
rect 116008 65966 116150 66030
rect 116214 65966 116422 66030
rect 116486 65966 116628 66030
rect 116008 65960 116628 65966
rect 116824 66166 117036 66172
rect 116824 66102 116966 66166
rect 117030 66102 117036 66166
rect 116824 66030 117036 66102
rect 116824 65966 116830 66030
rect 116894 65966 117036 66030
rect 116824 65960 117036 65966
rect 136816 66030 137572 66036
rect 136816 65966 137502 66030
rect 137566 65966 137572 66030
rect 136816 65960 137572 65966
rect 136816 65928 137028 65960
rect 136816 65872 136944 65928
rect 137000 65872 137028 65928
rect 136816 65824 137028 65872
rect 28288 65764 28364 65824
rect 110296 65764 110372 65824
rect 21760 65758 21972 65764
rect 21760 65694 21766 65758
rect 21830 65694 21972 65758
rect 21760 65622 21972 65694
rect 21760 65558 21902 65622
rect 21966 65558 21972 65622
rect 21760 65552 21972 65558
rect 22168 65758 22380 65764
rect 22168 65694 22310 65758
rect 22374 65694 22380 65758
rect 22168 65552 22380 65694
rect 22576 65622 22788 65764
rect 22576 65558 22582 65622
rect 22646 65558 22788 65622
rect 22576 65552 22788 65558
rect 22984 65758 23196 65764
rect 22984 65694 23126 65758
rect 23190 65694 23196 65758
rect 22984 65622 23196 65694
rect 22984 65558 22990 65622
rect 23054 65558 23196 65622
rect 22984 65552 23196 65558
rect 23392 65758 23604 65764
rect 23392 65694 23534 65758
rect 23598 65694 23604 65758
rect 23392 65622 23604 65694
rect 23392 65558 23534 65622
rect 23598 65558 23604 65622
rect 23392 65552 23604 65558
rect 28288 65552 28636 65764
rect 110160 65552 110508 65764
rect 115192 65758 115404 65764
rect 115192 65694 115198 65758
rect 115262 65694 115404 65758
rect 115192 65622 115404 65694
rect 115192 65558 115198 65622
rect 115262 65558 115404 65622
rect 115192 65552 115404 65558
rect 115600 65758 115812 65764
rect 115600 65694 115606 65758
rect 115670 65694 115812 65758
rect 115600 65622 115812 65694
rect 115600 65558 115606 65622
rect 115670 65558 115812 65622
rect 115600 65552 115812 65558
rect 116008 65758 116220 65764
rect 116008 65694 116150 65758
rect 116214 65694 116220 65758
rect 116008 65622 116220 65694
rect 116008 65558 116014 65622
rect 116078 65558 116220 65622
rect 116008 65552 116220 65558
rect 116416 65758 116628 65764
rect 116416 65694 116422 65758
rect 116486 65694 116628 65758
rect 116416 65552 116628 65694
rect 116824 65758 117036 65764
rect 116824 65694 116830 65758
rect 116894 65694 117036 65758
rect 116824 65622 117036 65694
rect 116824 65558 116830 65622
rect 116894 65558 117036 65622
rect 116824 65552 117036 65558
rect 28424 65492 28500 65552
rect 110432 65492 110508 65552
rect 21760 65350 21972 65356
rect 21760 65286 21902 65350
rect 21966 65286 21972 65350
rect 21760 65144 21972 65286
rect 22168 65350 22788 65356
rect 22168 65286 22582 65350
rect 22646 65286 22788 65350
rect 22168 65280 22788 65286
rect 22168 65220 22380 65280
rect 22168 65214 22516 65220
rect 22168 65150 22310 65214
rect 22374 65150 22446 65214
rect 22510 65150 22516 65214
rect 22168 65144 22516 65150
rect 22576 65144 22788 65280
rect 22984 65350 23196 65356
rect 22984 65286 22990 65350
rect 23054 65286 23196 65350
rect 22984 65214 23196 65286
rect 22984 65150 23126 65214
rect 23190 65150 23196 65214
rect 22984 65144 23196 65150
rect 23392 65350 23604 65356
rect 23392 65286 23534 65350
rect 23598 65286 23604 65350
rect 23392 65214 23604 65286
rect 28288 65280 28636 65492
rect 110160 65280 110508 65492
rect 115192 65350 115404 65356
rect 115192 65286 115198 65350
rect 115262 65286 115404 65350
rect 28424 65220 28500 65280
rect 110160 65220 110236 65280
rect 23392 65150 23398 65214
rect 23462 65150 23604 65214
rect 23392 65144 23604 65150
rect 21896 65084 21972 65144
rect 21760 64736 21972 65084
rect 28288 65008 28636 65220
rect 110160 65008 110508 65220
rect 115192 65214 115404 65286
rect 115192 65150 115198 65214
rect 115262 65150 115404 65214
rect 115192 65144 115404 65150
rect 115600 65350 115812 65356
rect 115600 65286 115606 65350
rect 115670 65286 115812 65350
rect 115600 65214 115812 65286
rect 115600 65150 115606 65214
rect 115670 65150 115812 65214
rect 115600 65144 115812 65150
rect 116008 65350 116220 65356
rect 116008 65286 116014 65350
rect 116078 65286 116220 65350
rect 116008 65220 116220 65286
rect 116416 65220 116628 65356
rect 116008 65214 116628 65220
rect 116008 65150 116150 65214
rect 116214 65150 116628 65214
rect 116008 65144 116628 65150
rect 116824 65350 117036 65356
rect 116824 65286 116830 65350
rect 116894 65286 117036 65350
rect 116824 65144 117036 65286
rect 116960 65084 117036 65144
rect 28560 64948 28636 65008
rect 110432 64948 110508 65008
rect 22168 64942 22380 64948
rect 22478 64942 22788 64948
rect 22168 64878 22310 64942
rect 22374 64878 22380 64942
rect 22440 64878 22446 64942
rect 22510 64878 22788 64942
rect 22168 64736 22380 64878
rect 22478 64872 22788 64878
rect 22576 64736 22788 64872
rect 22984 64942 23196 64948
rect 22984 64878 23126 64942
rect 23190 64878 23196 64942
rect 22984 64806 23196 64878
rect 22984 64742 22990 64806
rect 23054 64742 23196 64806
rect 22984 64736 23196 64742
rect 23392 64942 23604 64948
rect 23392 64878 23398 64942
rect 23462 64878 23604 64942
rect 23392 64806 23604 64878
rect 23392 64742 23534 64806
rect 23598 64742 23604 64806
rect 23392 64736 23604 64742
rect 21760 64676 21836 64736
rect 22576 64676 22652 64736
rect 1224 64398 1980 64404
rect 1224 64334 1230 64398
rect 1294 64334 1980 64398
rect 1224 64328 1980 64334
rect 21760 64328 21972 64676
rect 22168 64398 22380 64676
rect 22168 64334 22174 64398
rect 22238 64334 22380 64398
rect 22168 64328 22380 64334
rect 22576 64398 22788 64676
rect 22576 64334 22582 64398
rect 22646 64334 22788 64398
rect 22576 64328 22788 64334
rect 22984 64534 23196 64540
rect 22984 64470 22990 64534
rect 23054 64470 23196 64534
rect 22984 64328 23196 64470
rect 23392 64534 23604 64540
rect 23392 64470 23534 64534
rect 23598 64470 23604 64534
rect 23392 64328 23604 64470
rect 28288 64464 28636 64948
rect 110160 64464 110508 64948
rect 115192 64942 115404 64948
rect 115192 64878 115198 64942
rect 115262 64878 115404 64942
rect 115192 64806 115404 64878
rect 115192 64742 115334 64806
rect 115398 64742 115404 64806
rect 115192 64736 115404 64742
rect 115600 64942 115812 64948
rect 115600 64878 115606 64942
rect 115670 64878 115812 64942
rect 115600 64806 115812 64878
rect 115600 64742 115742 64806
rect 115806 64742 115812 64806
rect 115600 64736 115812 64742
rect 116008 64942 116220 64948
rect 116008 64878 116150 64942
rect 116214 64878 116220 64942
rect 116008 64736 116220 64878
rect 116416 64736 116628 64948
rect 116824 64736 117036 65084
rect 116008 64676 116084 64736
rect 116552 64676 116628 64736
rect 116960 64676 117036 64736
rect 28288 64404 28364 64464
rect 110432 64404 110508 64464
rect 1768 64248 1980 64328
rect 21896 64268 21972 64328
rect 1768 64192 1798 64248
rect 1854 64192 1980 64248
rect 1768 64056 1980 64192
rect 21760 64126 21972 64268
rect 22984 64268 23060 64328
rect 23392 64268 23468 64328
rect 21760 64062 21902 64126
rect 21966 64062 21972 64126
rect 21760 64056 21972 64062
rect 22168 64126 22380 64132
rect 22168 64062 22174 64126
rect 22238 64062 22380 64126
rect 22168 63920 22380 64062
rect 22576 64126 22788 64132
rect 22576 64062 22582 64126
rect 22646 64062 22788 64126
rect 22576 63996 22788 64062
rect 22304 63860 22380 63920
rect 22440 63920 22788 63996
rect 22440 63860 22516 63920
rect 22712 63860 22788 63920
rect 21760 63854 21972 63860
rect 21760 63790 21902 63854
rect 21966 63790 21972 63854
rect 21760 63718 21972 63790
rect 21760 63654 21766 63718
rect 21830 63654 21972 63718
rect 21760 63648 21972 63654
rect 22168 63784 22516 63860
rect 22168 63718 22380 63784
rect 22168 63654 22310 63718
rect 22374 63654 22380 63718
rect 22168 63648 22380 63654
rect 22576 63648 22788 63860
rect 22984 63920 23196 64268
rect 23392 63920 23604 64268
rect 22984 63860 23060 63920
rect 23392 63860 23468 63920
rect 22984 63512 23196 63860
rect 23392 63512 23604 63860
rect 28288 63854 28636 64404
rect 28288 63790 28566 63854
rect 28630 63790 28636 63854
rect 28288 63784 28636 63790
rect 110160 64262 110508 64404
rect 115192 64534 115404 64540
rect 115192 64470 115334 64534
rect 115398 64470 115404 64534
rect 115192 64328 115404 64470
rect 115600 64534 115812 64540
rect 115600 64470 115742 64534
rect 115806 64470 115812 64534
rect 115600 64328 115812 64470
rect 116008 64398 116220 64676
rect 116008 64334 116014 64398
rect 116078 64334 116220 64398
rect 116008 64328 116220 64334
rect 116416 64398 116628 64676
rect 116416 64334 116558 64398
rect 116622 64334 116628 64398
rect 116416 64328 116628 64334
rect 116824 64328 117036 64676
rect 115328 64268 115404 64328
rect 115736 64268 115812 64328
rect 110160 64198 110166 64262
rect 110230 64198 110508 64262
rect 110160 63990 110508 64198
rect 110160 63926 110166 63990
rect 110230 63926 110508 63990
rect 110160 63854 110508 63926
rect 110160 63790 110438 63854
rect 110502 63790 110508 63854
rect 110160 63784 110508 63790
rect 115192 63920 115404 64268
rect 115600 63920 115812 64268
rect 116824 64268 116900 64328
rect 136816 64268 137028 64404
rect 116008 64126 116220 64132
rect 116008 64062 116014 64126
rect 116078 64062 116220 64126
rect 116008 63996 116220 64062
rect 116416 64126 116628 64132
rect 116416 64062 116558 64126
rect 116622 64062 116628 64126
rect 116008 63920 116356 63996
rect 116416 63920 116628 64062
rect 116824 64126 117036 64268
rect 116824 64062 116830 64126
rect 116894 64062 117036 64126
rect 116824 64056 117036 64062
rect 136816 64262 137572 64268
rect 136816 64248 137502 64262
rect 136816 64192 136944 64248
rect 137000 64198 137502 64248
rect 137566 64198 137572 64262
rect 137000 64192 137572 64198
rect 136816 64056 137028 64192
rect 115192 63860 115268 63920
rect 115736 63860 115812 63920
rect 116144 63860 116220 63920
rect 23120 63452 23196 63512
rect 23528 63452 23604 63512
rect 21760 63446 21972 63452
rect 21760 63382 21766 63446
rect 21830 63382 21972 63446
rect 21760 63310 21972 63382
rect 21760 63246 21902 63310
rect 21966 63246 21972 63310
rect 21760 63240 21972 63246
rect 22168 63446 22380 63452
rect 22168 63382 22310 63446
rect 22374 63382 22380 63446
rect 22168 63104 22380 63382
rect 22576 63180 22788 63452
rect 22984 63310 23196 63452
rect 22984 63246 23126 63310
rect 23190 63246 23196 63310
rect 22984 63240 23196 63246
rect 23392 63310 23604 63452
rect 23392 63246 23398 63310
rect 23462 63246 23604 63310
rect 23392 63240 23604 63246
rect 28288 63582 28636 63588
rect 28288 63518 28566 63582
rect 28630 63518 28636 63582
rect 28288 63446 28636 63518
rect 28288 63382 28294 63446
rect 28358 63382 28636 63446
rect 28288 63240 28636 63382
rect 110160 63582 110508 63588
rect 110160 63518 110438 63582
rect 110502 63518 110508 63582
rect 110160 63240 110508 63518
rect 115192 63512 115404 63860
rect 115600 63512 115812 63860
rect 116008 63648 116220 63860
rect 116280 63860 116356 63920
rect 116552 63860 116628 63920
rect 116280 63784 116628 63860
rect 116416 63724 116628 63784
rect 116318 63718 116628 63724
rect 116280 63654 116286 63718
rect 116350 63654 116628 63718
rect 116318 63648 116628 63654
rect 116824 63854 117036 63860
rect 116824 63790 116830 63854
rect 116894 63790 117036 63854
rect 116824 63718 117036 63790
rect 116824 63654 116830 63718
rect 116894 63654 117036 63718
rect 116824 63648 117036 63654
rect 115328 63452 115404 63512
rect 115736 63452 115812 63512
rect 115192 63310 115404 63452
rect 115192 63246 115198 63310
rect 115262 63246 115404 63310
rect 115192 63240 115404 63246
rect 115600 63310 115812 63452
rect 115600 63246 115606 63310
rect 115670 63246 115812 63310
rect 115600 63240 115812 63246
rect 116008 63446 116356 63452
rect 116008 63382 116286 63446
rect 116350 63382 116356 63446
rect 116008 63376 116356 63382
rect 116008 63316 116220 63376
rect 116416 63316 116628 63452
rect 116008 63240 116628 63316
rect 116824 63446 117036 63452
rect 116824 63382 116830 63446
rect 116894 63382 117036 63446
rect 116824 63310 117036 63382
rect 116824 63246 116966 63310
rect 117030 63246 117036 63310
rect 116824 63240 117036 63246
rect 22304 63044 22380 63104
rect 22440 63104 22788 63180
rect 28288 63180 28364 63240
rect 110432 63180 110508 63240
rect 28288 63174 28636 63180
rect 28288 63110 28294 63174
rect 28358 63110 28636 63174
rect 22440 63044 22516 63104
rect 21760 63038 21972 63044
rect 21760 62974 21902 63038
rect 21966 62974 21972 63038
rect 21760 62902 21972 62974
rect 21760 62838 21766 62902
rect 21830 62838 21972 62902
rect 21760 62832 21972 62838
rect 22168 62968 22516 63044
rect 22168 62908 22380 62968
rect 22576 62908 22788 63044
rect 22984 63038 23196 63044
rect 22984 62974 23126 63038
rect 23190 62974 23196 63038
rect 22168 62902 22924 62908
rect 22168 62838 22582 62902
rect 22646 62838 22924 62902
rect 22168 62832 22924 62838
rect 22984 62902 23196 62974
rect 22984 62838 22990 62902
rect 23054 62838 23196 62902
rect 22984 62832 23196 62838
rect 23392 63038 23604 63044
rect 23392 62974 23398 63038
rect 23462 62974 23604 63038
rect 23392 62902 23604 62974
rect 28288 62968 28636 63110
rect 110160 62968 110508 63180
rect 116008 63104 116220 63240
rect 116416 63180 116628 63240
rect 116280 63104 116628 63180
rect 116280 63044 116356 63104
rect 116552 63044 116628 63104
rect 115192 63038 115404 63044
rect 115192 62974 115198 63038
rect 115262 62974 115404 63038
rect 28424 62908 28500 62968
rect 110296 62908 110372 62968
rect 23392 62838 23398 62902
rect 23462 62838 23604 62902
rect 23392 62832 23604 62838
rect 22848 62772 22924 62832
rect 22848 62696 23468 62772
rect 23392 62636 23468 62696
rect 1224 62630 1980 62636
rect 1224 62566 1230 62630
rect 1294 62568 1980 62630
rect 1294 62566 1798 62568
rect 1224 62560 1798 62566
rect 1768 62512 1798 62560
rect 1854 62512 1980 62568
rect 1768 62424 1980 62512
rect 21760 62630 21972 62636
rect 21760 62566 21766 62630
rect 21830 62566 21972 62630
rect 21760 62494 21972 62566
rect 21760 62430 21766 62494
rect 21830 62430 21972 62494
rect 21760 62424 21972 62430
rect 22168 62494 22380 62636
rect 22168 62430 22174 62494
rect 22238 62430 22380 62494
rect 22168 62424 22380 62430
rect 22576 62630 22788 62636
rect 22576 62566 22582 62630
rect 22646 62566 22788 62630
rect 22576 62424 22788 62566
rect 22984 62630 23196 62636
rect 22984 62566 22990 62630
rect 23054 62566 23196 62630
rect 22984 62494 23196 62566
rect 22984 62430 22990 62494
rect 23054 62430 23196 62494
rect 22984 62424 23196 62430
rect 23392 62630 23604 62636
rect 23392 62566 23398 62630
rect 23462 62566 23604 62630
rect 23392 62494 23604 62566
rect 23392 62430 23534 62494
rect 23598 62430 23604 62494
rect 23392 62424 23604 62430
rect 28288 62424 28636 62908
rect 110160 62630 110508 62908
rect 115192 62902 115404 62974
rect 115192 62838 115198 62902
rect 115262 62838 115404 62902
rect 115192 62832 115404 62838
rect 115600 63038 115812 63044
rect 115600 62974 115606 63038
rect 115670 62974 115812 63038
rect 115600 62902 115812 62974
rect 115600 62838 115606 62902
rect 115670 62838 115812 62902
rect 115600 62832 115812 62838
rect 116008 62968 116356 63044
rect 116008 62908 116220 62968
rect 116008 62902 116356 62908
rect 116008 62838 116150 62902
rect 116214 62838 116286 62902
rect 116350 62838 116356 62902
rect 116008 62832 116356 62838
rect 116416 62832 116628 63044
rect 116824 63038 117036 63044
rect 116824 62974 116966 63038
rect 117030 62974 117036 63038
rect 116824 62902 117036 62974
rect 116824 62838 116966 62902
rect 117030 62838 117036 62902
rect 116824 62832 117036 62838
rect 110160 62566 110166 62630
rect 110230 62566 110508 62630
rect 110160 62424 110508 62566
rect 115192 62630 115404 62636
rect 115192 62566 115198 62630
rect 115262 62566 115404 62630
rect 115192 62494 115404 62566
rect 115192 62430 115334 62494
rect 115398 62430 115404 62494
rect 115192 62424 115404 62430
rect 115600 62630 115812 62636
rect 115600 62566 115606 62630
rect 115670 62566 115812 62630
rect 115600 62494 115812 62566
rect 115600 62430 115742 62494
rect 115806 62430 115812 62494
rect 115600 62424 115812 62430
rect 116008 62630 116220 62636
rect 116318 62630 116628 62636
rect 116008 62566 116150 62630
rect 116214 62566 116220 62630
rect 116280 62566 116286 62630
rect 116350 62566 116628 62630
rect 116008 62424 116220 62566
rect 116318 62560 116628 62566
rect 116416 62494 116628 62560
rect 116416 62430 116422 62494
rect 116486 62430 116628 62494
rect 116416 62424 116628 62430
rect 116824 62630 117036 62636
rect 116824 62566 116966 62630
rect 117030 62566 117036 62630
rect 116824 62494 117036 62566
rect 116824 62430 116830 62494
rect 116894 62430 117036 62494
rect 116824 62424 117036 62430
rect 136816 62630 137572 62636
rect 136816 62568 137502 62630
rect 136816 62512 136944 62568
rect 137000 62566 137502 62568
rect 137566 62566 137572 62630
rect 137000 62560 137572 62566
rect 137000 62512 137028 62560
rect 136816 62424 137028 62512
rect 22576 62364 22652 62424
rect 22304 62288 22652 62364
rect 28288 62364 28364 62424
rect 110432 62364 110508 62424
rect 22304 62228 22380 62288
rect 21760 62222 21972 62228
rect 21760 62158 21766 62222
rect 21830 62158 21972 62222
rect 21760 62086 21972 62158
rect 21760 62022 21902 62086
rect 21966 62022 21972 62086
rect 21760 62016 21972 62022
rect 22168 62222 22788 62228
rect 22168 62158 22174 62222
rect 22238 62158 22788 62222
rect 22168 62152 22788 62158
rect 22168 62092 22380 62152
rect 22168 62086 22516 62092
rect 22168 62022 22446 62086
rect 22510 62022 22516 62086
rect 22168 62016 22516 62022
rect 22576 62016 22788 62152
rect 22984 62222 23196 62228
rect 22984 62158 22990 62222
rect 23054 62158 23196 62222
rect 22984 62086 23196 62158
rect 22984 62022 22990 62086
rect 23054 62022 23196 62086
rect 22984 62016 23196 62022
rect 23392 62222 23604 62228
rect 23392 62158 23534 62222
rect 23598 62158 23604 62222
rect 23392 62086 23604 62158
rect 28288 62152 28636 62364
rect 110160 62358 110508 62364
rect 110160 62294 110166 62358
rect 110230 62294 110508 62358
rect 110160 62152 110508 62294
rect 28560 62092 28636 62152
rect 110432 62092 110508 62152
rect 23392 62022 23398 62086
rect 23462 62022 23604 62086
rect 23392 62016 23604 62022
rect 28288 61880 28636 62092
rect 28560 61820 28636 61880
rect 21760 61814 21972 61820
rect 21760 61750 21902 61814
rect 21966 61750 21972 61814
rect 21760 61678 21972 61750
rect 21760 61614 21902 61678
rect 21966 61614 21972 61678
rect 21760 61608 21972 61614
rect 22168 61684 22380 61820
rect 22478 61814 22788 61820
rect 22440 61750 22446 61814
rect 22510 61750 22788 61814
rect 22478 61744 22788 61750
rect 22168 61678 22516 61684
rect 22168 61614 22310 61678
rect 22374 61614 22446 61678
rect 22510 61614 22516 61678
rect 22168 61608 22516 61614
rect 22576 61608 22788 61744
rect 22984 61814 23196 61820
rect 22984 61750 22990 61814
rect 23054 61750 23196 61814
rect 22984 61678 23196 61750
rect 22984 61614 22990 61678
rect 23054 61614 23196 61678
rect 22984 61608 23196 61614
rect 23392 61814 23604 61820
rect 23392 61750 23398 61814
rect 23462 61750 23604 61814
rect 23392 61678 23604 61750
rect 23392 61614 23534 61678
rect 23598 61614 23604 61678
rect 23392 61608 23604 61614
rect 28288 61608 28636 61820
rect 110160 61880 110508 62092
rect 115192 62222 115404 62228
rect 115192 62158 115334 62222
rect 115398 62158 115404 62222
rect 115192 62086 115404 62158
rect 115192 62022 115198 62086
rect 115262 62022 115404 62086
rect 115192 62016 115404 62022
rect 115600 62222 115812 62228
rect 115600 62158 115742 62222
rect 115806 62158 115812 62222
rect 115600 62086 115812 62158
rect 115600 62022 115606 62086
rect 115670 62022 115812 62086
rect 115600 62016 115812 62022
rect 116008 62222 116628 62228
rect 116008 62158 116422 62222
rect 116486 62158 116628 62222
rect 116008 62152 116628 62158
rect 116008 62016 116220 62152
rect 116416 62086 116628 62152
rect 116416 62022 116558 62086
rect 116622 62022 116628 62086
rect 116416 62016 116628 62022
rect 116824 62222 117036 62228
rect 116824 62158 116830 62222
rect 116894 62158 117036 62222
rect 116824 62086 117036 62158
rect 116824 62022 116966 62086
rect 117030 62022 117036 62086
rect 116824 62016 117036 62022
rect 110160 61820 110236 61880
rect 110160 61608 110508 61820
rect 115192 61814 115404 61820
rect 115192 61750 115198 61814
rect 115262 61750 115404 61814
rect 115192 61678 115404 61750
rect 115192 61614 115334 61678
rect 115398 61614 115404 61678
rect 115192 61608 115404 61614
rect 115600 61814 115812 61820
rect 115600 61750 115606 61814
rect 115670 61750 115812 61814
rect 115600 61678 115812 61750
rect 115600 61614 115742 61678
rect 115806 61614 115812 61678
rect 115600 61608 115812 61614
rect 116008 61684 116220 61820
rect 116416 61814 116628 61820
rect 116416 61750 116558 61814
rect 116622 61750 116628 61814
rect 116416 61684 116628 61750
rect 116008 61678 116628 61684
rect 116008 61614 116150 61678
rect 116214 61614 116628 61678
rect 116008 61608 116628 61614
rect 116824 61814 117036 61820
rect 116824 61750 116966 61814
rect 117030 61750 117036 61814
rect 116824 61678 117036 61750
rect 116824 61614 116830 61678
rect 116894 61614 117036 61678
rect 116824 61608 117036 61614
rect 22304 61548 22380 61608
rect 22576 61548 22652 61608
rect 28560 61548 28636 61608
rect 110296 61548 110372 61608
rect 116144 61548 116220 61608
rect 22304 61472 22652 61548
rect 21760 61406 21972 61412
rect 21760 61342 21902 61406
rect 21966 61342 21972 61406
rect 21760 61200 21972 61342
rect 22168 61406 22380 61412
rect 22478 61406 22788 61412
rect 22168 61342 22310 61406
rect 22374 61342 22380 61406
rect 22440 61342 22446 61406
rect 22510 61342 22788 61406
rect 22168 61200 22380 61342
rect 22478 61336 22788 61342
rect 22576 61270 22788 61336
rect 22576 61206 22718 61270
rect 22782 61206 22788 61270
rect 22576 61200 22788 61206
rect 22984 61406 23196 61412
rect 22984 61342 22990 61406
rect 23054 61342 23196 61406
rect 22984 61270 23196 61342
rect 22984 61206 22990 61270
rect 23054 61206 23196 61270
rect 22984 61200 23196 61206
rect 23392 61406 23604 61412
rect 23392 61342 23534 61406
rect 23598 61342 23604 61406
rect 23392 61270 23604 61342
rect 28288 61336 28636 61548
rect 110160 61336 110508 61548
rect 116144 61472 116492 61548
rect 116416 61412 116492 61472
rect 28424 61276 28500 61336
rect 110432 61276 110508 61336
rect 23392 61206 23534 61270
rect 23598 61206 23604 61270
rect 23392 61200 23604 61206
rect 21760 61140 21836 61200
rect 1224 60998 1980 61004
rect 1224 60934 1230 60998
rect 1294 60934 1980 60998
rect 1224 60928 1980 60934
rect 1768 60888 1980 60928
rect 1768 60832 1798 60888
rect 1854 60832 1980 60888
rect 1768 60792 1980 60832
rect 21760 60792 21972 61140
rect 28288 61064 28636 61276
rect 110160 61134 110508 61276
rect 115192 61406 115404 61412
rect 115192 61342 115334 61406
rect 115398 61342 115404 61406
rect 115192 61270 115404 61342
rect 115192 61206 115198 61270
rect 115262 61206 115404 61270
rect 115192 61200 115404 61206
rect 115600 61406 115812 61412
rect 115600 61342 115742 61406
rect 115806 61342 115812 61406
rect 115600 61270 115812 61342
rect 115600 61206 115742 61270
rect 115806 61206 115812 61270
rect 115600 61200 115812 61206
rect 116008 61406 116220 61412
rect 116008 61342 116150 61406
rect 116214 61342 116220 61406
rect 116008 61270 116220 61342
rect 116008 61206 116014 61270
rect 116078 61206 116220 61270
rect 116008 61200 116220 61206
rect 116416 61270 116628 61412
rect 116416 61206 116558 61270
rect 116622 61206 116628 61270
rect 116416 61200 116628 61206
rect 116824 61406 117036 61412
rect 116824 61342 116830 61406
rect 116894 61342 117036 61406
rect 116824 61200 117036 61342
rect 110160 61070 110438 61134
rect 110502 61070 110508 61134
rect 110160 61064 110508 61070
rect 116824 61140 116900 61200
rect 28424 61004 28500 61064
rect 110160 61004 110236 61064
rect 22168 60998 22516 61004
rect 22168 60934 22446 60998
rect 22510 60934 22516 60998
rect 22168 60928 22516 60934
rect 22576 60998 22788 61004
rect 22576 60934 22718 60998
rect 22782 60934 22788 60998
rect 22168 60868 22380 60928
rect 22576 60868 22788 60934
rect 22168 60792 22788 60868
rect 22984 60998 23196 61004
rect 22984 60934 22990 60998
rect 23054 60934 23196 60998
rect 22984 60862 23196 60934
rect 22984 60798 23126 60862
rect 23190 60798 23196 60862
rect 22984 60792 23196 60798
rect 23392 60998 23604 61004
rect 23392 60934 23534 60998
rect 23598 60934 23604 60998
rect 23392 60862 23604 60934
rect 23392 60798 23398 60862
rect 23462 60798 23604 60862
rect 23392 60792 23604 60798
rect 21896 60732 21972 60792
rect 22304 60732 22380 60792
rect 21760 60384 21972 60732
rect 22168 60454 22380 60732
rect 22478 60726 22788 60732
rect 22440 60662 22446 60726
rect 22510 60662 22788 60726
rect 22478 60656 22788 60662
rect 22168 60390 22174 60454
rect 22238 60390 22380 60454
rect 22168 60384 22380 60390
rect 22576 60384 22788 60656
rect 22984 60590 23196 60596
rect 22984 60526 23126 60590
rect 23190 60526 23196 60590
rect 22984 60454 23196 60526
rect 22984 60390 23126 60454
rect 23190 60390 23196 60454
rect 22984 60384 23196 60390
rect 23392 60590 23604 60596
rect 23392 60526 23398 60590
rect 23462 60526 23604 60590
rect 23392 60454 23604 60526
rect 23392 60390 23534 60454
rect 23598 60390 23604 60454
rect 23392 60384 23604 60390
rect 28288 60520 28636 61004
rect 110160 60862 110508 61004
rect 110160 60798 110438 60862
rect 110502 60798 110508 60862
rect 110160 60520 110508 60798
rect 115192 60998 115404 61004
rect 115192 60934 115198 60998
rect 115262 60934 115404 60998
rect 115192 60862 115404 60934
rect 115192 60798 115198 60862
rect 115262 60798 115404 60862
rect 115192 60792 115404 60798
rect 115600 60998 115812 61004
rect 115600 60934 115742 60998
rect 115806 60934 115812 60998
rect 115600 60862 115812 60934
rect 115600 60798 115606 60862
rect 115670 60798 115812 60862
rect 115600 60792 115812 60798
rect 116008 60998 116220 61004
rect 116008 60934 116014 60998
rect 116078 60934 116220 60998
rect 116008 60792 116220 60934
rect 116416 60998 116628 61004
rect 116416 60934 116558 60998
rect 116622 60934 116628 60998
rect 116416 60792 116628 60934
rect 116824 60792 117036 61140
rect 136816 60998 137572 61004
rect 136816 60934 137502 60998
rect 137566 60934 137572 60998
rect 136816 60928 137572 60934
rect 136816 60888 137028 60928
rect 136816 60832 136944 60888
rect 137000 60832 137028 60888
rect 136816 60792 137028 60832
rect 116008 60732 116084 60792
rect 116824 60732 116900 60792
rect 115192 60590 115404 60596
rect 115192 60526 115198 60590
rect 115262 60526 115404 60590
rect 28288 60460 28364 60520
rect 110160 60460 110236 60520
rect 21896 60324 21972 60384
rect 21760 60182 21972 60324
rect 28288 60318 28636 60460
rect 28288 60254 28566 60318
rect 28630 60254 28636 60318
rect 28288 60248 28636 60254
rect 110160 60248 110508 60460
rect 115192 60454 115404 60526
rect 115192 60390 115334 60454
rect 115398 60390 115404 60454
rect 115192 60384 115404 60390
rect 115600 60590 115812 60596
rect 115600 60526 115606 60590
rect 115670 60526 115812 60590
rect 115600 60454 115812 60526
rect 115600 60390 115742 60454
rect 115806 60390 115812 60454
rect 115600 60384 115812 60390
rect 116008 60454 116220 60732
rect 116008 60390 116014 60454
rect 116078 60390 116220 60454
rect 116008 60384 116220 60390
rect 116416 60454 116628 60732
rect 116416 60390 116422 60454
rect 116486 60390 116628 60454
rect 116416 60384 116628 60390
rect 116824 60384 117036 60732
rect 116824 60324 116900 60384
rect 28424 60188 28500 60248
rect 110296 60188 110372 60248
rect 21760 60118 21902 60182
rect 21966 60118 21972 60182
rect 21760 60112 21972 60118
rect 22168 60182 22380 60188
rect 22168 60118 22174 60182
rect 22238 60118 22380 60182
rect 22168 59976 22380 60118
rect 22576 59976 22788 60188
rect 22984 60182 23196 60188
rect 22984 60118 23126 60182
rect 23190 60118 23196 60182
rect 22984 59976 23196 60118
rect 23392 60182 23604 60188
rect 23392 60118 23534 60182
rect 23598 60118 23604 60182
rect 23392 59976 23604 60118
rect 22168 59916 22244 59976
rect 22712 59916 22788 59976
rect 23120 59916 23196 59976
rect 23528 59916 23604 59976
rect 21760 59910 21972 59916
rect 21760 59846 21902 59910
rect 21966 59846 21972 59910
rect 21760 59774 21972 59846
rect 21760 59710 21902 59774
rect 21966 59710 21972 59774
rect 21760 59704 21972 59710
rect 22168 59780 22380 59916
rect 22576 59780 22788 59916
rect 22168 59774 22788 59780
rect 22168 59710 22310 59774
rect 22374 59710 22788 59774
rect 22168 59704 22788 59710
rect 22304 59644 22380 59704
rect 22304 59568 22652 59644
rect 22576 59508 22652 59568
rect 22984 59568 23196 59916
rect 23392 59568 23604 59916
rect 28288 60046 28636 60188
rect 28288 59982 28294 60046
rect 28358 59982 28566 60046
rect 28630 59982 28636 60046
rect 28288 59840 28636 59982
rect 110160 59910 110508 60188
rect 115192 60182 115404 60188
rect 115192 60118 115334 60182
rect 115398 60118 115404 60182
rect 115192 59976 115404 60118
rect 115600 60182 115812 60188
rect 115600 60118 115742 60182
rect 115806 60118 115812 60182
rect 115600 59976 115812 60118
rect 115328 59916 115404 59976
rect 115736 59916 115812 59976
rect 110160 59846 110166 59910
rect 110230 59846 110508 59910
rect 110160 59840 110508 59846
rect 28288 59638 28636 59644
rect 28288 59574 28294 59638
rect 28358 59574 28636 59638
rect 22984 59508 23060 59568
rect 23392 59508 23468 59568
rect 21760 59502 21972 59508
rect 21760 59438 21902 59502
rect 21966 59438 21972 59502
rect 21760 59366 21972 59438
rect 21760 59302 21766 59366
rect 21830 59302 21972 59366
rect 21760 59296 21972 59302
rect 22168 59502 22380 59508
rect 22168 59438 22310 59502
rect 22374 59438 22380 59502
rect 1224 59230 1980 59236
rect 1224 59166 1230 59230
rect 1294 59208 1980 59230
rect 1294 59166 1798 59208
rect 1224 59160 1798 59166
rect 1768 59152 1798 59160
rect 1854 59152 1980 59208
rect 22168 59160 22380 59438
rect 22576 59160 22788 59508
rect 22984 59366 23196 59508
rect 22984 59302 22990 59366
rect 23054 59302 23196 59366
rect 22984 59296 23196 59302
rect 23392 59366 23604 59508
rect 23392 59302 23534 59366
rect 23598 59302 23604 59366
rect 23392 59296 23604 59302
rect 28288 59296 28636 59574
rect 110160 59638 110508 59644
rect 110160 59574 110166 59638
rect 110230 59574 110508 59638
rect 110160 59502 110508 59574
rect 110160 59438 110438 59502
rect 110502 59438 110508 59502
rect 110160 59296 110508 59438
rect 115192 59568 115404 59916
rect 115600 59568 115812 59916
rect 116008 60182 116220 60188
rect 116008 60118 116014 60182
rect 116078 60118 116220 60182
rect 116008 60052 116220 60118
rect 116416 60182 116628 60188
rect 116416 60118 116422 60182
rect 116486 60118 116628 60182
rect 116416 60052 116628 60118
rect 116824 60182 117036 60324
rect 116824 60118 116830 60182
rect 116894 60118 117036 60182
rect 116824 60112 117036 60118
rect 116008 59976 116628 60052
rect 116008 59916 116084 59976
rect 116552 59916 116628 59976
rect 116008 59704 116220 59916
rect 116416 59774 116628 59916
rect 116416 59710 116558 59774
rect 116622 59710 116628 59774
rect 116416 59704 116628 59710
rect 116824 59910 117036 59916
rect 116824 59846 116830 59910
rect 116894 59846 117036 59910
rect 116824 59774 117036 59846
rect 116824 59710 116966 59774
rect 117030 59710 117036 59774
rect 116824 59704 117036 59710
rect 115192 59508 115268 59568
rect 115600 59508 115676 59568
rect 115192 59366 115404 59508
rect 115192 59302 115334 59366
rect 115398 59302 115404 59366
rect 115192 59296 115404 59302
rect 115600 59366 115812 59508
rect 115600 59302 115742 59366
rect 115806 59302 115812 59366
rect 115600 59296 115812 59302
rect 28424 59236 28500 59296
rect 110432 59236 110508 59296
rect 1768 59024 1980 59152
rect 22304 59100 22380 59160
rect 21760 59094 21972 59100
rect 21760 59030 21766 59094
rect 21830 59030 21972 59094
rect 21760 58958 21972 59030
rect 21760 58894 21902 58958
rect 21966 58894 21972 58958
rect 21760 58888 21972 58894
rect 22168 58958 22380 59100
rect 22168 58894 22310 58958
rect 22374 58894 22380 58958
rect 22168 58888 22380 58894
rect 22576 58888 22788 59100
rect 22984 59094 23196 59100
rect 22984 59030 22990 59094
rect 23054 59030 23196 59094
rect 22984 58958 23196 59030
rect 22984 58894 22990 58958
rect 23054 58894 23196 58958
rect 22984 58888 23196 58894
rect 23392 59094 23604 59100
rect 23392 59030 23534 59094
rect 23598 59030 23604 59094
rect 23392 58958 23604 59030
rect 23392 58894 23398 58958
rect 23462 58894 23604 58958
rect 23392 58888 23604 58894
rect 28288 59024 28636 59236
rect 110160 59230 110508 59236
rect 110160 59166 110438 59230
rect 110502 59166 110508 59230
rect 110160 59024 110508 59166
rect 116008 59160 116220 59508
rect 116144 59100 116220 59160
rect 115192 59094 115404 59100
rect 115192 59030 115334 59094
rect 115398 59030 115404 59094
rect 28288 58964 28364 59024
rect 110296 58964 110372 59024
rect 22576 58828 22652 58888
rect 22304 58752 22652 58828
rect 22304 58692 22380 58752
rect 21760 58686 21972 58692
rect 21760 58622 21902 58686
rect 21966 58622 21972 58686
rect 21760 58550 21972 58622
rect 21760 58486 21902 58550
rect 21966 58486 21972 58550
rect 21760 58480 21972 58486
rect 22168 58686 22788 58692
rect 22168 58622 22310 58686
rect 22374 58622 22788 58686
rect 22168 58616 22788 58622
rect 22168 58550 22380 58616
rect 22168 58486 22174 58550
rect 22238 58486 22380 58550
rect 22168 58480 22380 58486
rect 22576 58550 22788 58616
rect 22576 58486 22718 58550
rect 22782 58486 22788 58550
rect 22576 58480 22788 58486
rect 22984 58686 23196 58692
rect 22984 58622 22990 58686
rect 23054 58622 23196 58686
rect 22984 58550 23196 58622
rect 22984 58486 22990 58550
rect 23054 58486 23196 58550
rect 22984 58480 23196 58486
rect 23392 58686 23604 58692
rect 23392 58622 23398 58686
rect 23462 58622 23604 58686
rect 23392 58550 23604 58622
rect 23392 58486 23398 58550
rect 23462 58486 23604 58550
rect 23392 58480 23604 58486
rect 28288 58686 28636 58964
rect 28288 58622 28566 58686
rect 28630 58622 28636 58686
rect 28288 58480 28636 58622
rect 110160 58686 110508 58964
rect 115192 58958 115404 59030
rect 115192 58894 115198 58958
rect 115262 58894 115404 58958
rect 115192 58888 115404 58894
rect 115600 59094 115812 59100
rect 115600 59030 115742 59094
rect 115806 59030 115812 59094
rect 115600 58958 115812 59030
rect 115600 58894 115742 58958
rect 115806 58894 115812 58958
rect 115600 58888 115812 58894
rect 116008 58958 116220 59100
rect 116008 58894 116150 58958
rect 116214 58894 116220 58958
rect 116008 58888 116220 58894
rect 116416 59502 116628 59508
rect 116416 59438 116558 59502
rect 116622 59438 116628 59502
rect 116416 59160 116628 59438
rect 116824 59502 117036 59508
rect 116824 59438 116966 59502
rect 117030 59438 117036 59502
rect 116824 59366 117036 59438
rect 116824 59302 116830 59366
rect 116894 59302 117036 59366
rect 116824 59296 117036 59302
rect 136816 59208 137028 59236
rect 116416 59100 116492 59160
rect 136816 59152 136944 59208
rect 137000 59152 137028 59208
rect 136816 59100 137028 59152
rect 116416 58958 116628 59100
rect 116416 58894 116558 58958
rect 116622 58894 116628 58958
rect 116416 58888 116628 58894
rect 116824 59094 117036 59100
rect 116824 59030 116830 59094
rect 116894 59030 117036 59094
rect 116824 58958 117036 59030
rect 136816 59094 137572 59100
rect 136816 59030 137502 59094
rect 137566 59030 137572 59094
rect 136816 59024 137572 59030
rect 116824 58894 116830 58958
rect 116894 58894 117036 58958
rect 116824 58888 117036 58894
rect 110160 58622 110438 58686
rect 110502 58622 110508 58686
rect 110160 58480 110508 58622
rect 115192 58686 115404 58692
rect 115192 58622 115198 58686
rect 115262 58622 115404 58686
rect 115192 58550 115404 58622
rect 115192 58486 115198 58550
rect 115262 58486 115404 58550
rect 115192 58480 115404 58486
rect 115600 58686 115812 58692
rect 115600 58622 115742 58686
rect 115806 58622 115812 58686
rect 115600 58550 115812 58622
rect 115600 58486 115742 58550
rect 115806 58486 115812 58550
rect 115600 58480 115812 58486
rect 116008 58686 116220 58692
rect 116008 58622 116150 58686
rect 116214 58622 116220 58686
rect 116008 58556 116220 58622
rect 116416 58686 116628 58692
rect 116416 58622 116558 58686
rect 116622 58622 116628 58686
rect 116416 58556 116628 58622
rect 116008 58550 116628 58556
rect 116008 58486 116014 58550
rect 116078 58486 116628 58550
rect 116008 58480 116628 58486
rect 116824 58686 117036 58692
rect 116824 58622 116830 58686
rect 116894 58622 117036 58686
rect 116824 58550 117036 58622
rect 116824 58486 116830 58550
rect 116894 58486 117036 58550
rect 116824 58480 117036 58486
rect 28288 58420 28364 58480
rect 110432 58420 110508 58480
rect 28288 58414 28636 58420
rect 28288 58350 28566 58414
rect 28630 58350 28636 58414
rect 21760 58278 21972 58284
rect 21760 58214 21902 58278
rect 21966 58214 21972 58278
rect 21760 58142 21972 58214
rect 21760 58078 21766 58142
rect 21830 58078 21972 58142
rect 21760 58072 21972 58078
rect 22168 58278 22380 58284
rect 22168 58214 22174 58278
rect 22238 58214 22380 58278
rect 22168 58072 22380 58214
rect 22576 58278 22788 58284
rect 22576 58214 22718 58278
rect 22782 58214 22788 58278
rect 22576 58148 22788 58214
rect 22478 58142 22788 58148
rect 22440 58078 22446 58142
rect 22510 58078 22788 58142
rect 22478 58072 22788 58078
rect 22984 58278 23196 58284
rect 22984 58214 22990 58278
rect 23054 58214 23196 58278
rect 22984 58142 23196 58214
rect 22984 58078 22990 58142
rect 23054 58078 23196 58142
rect 22984 58072 23196 58078
rect 23392 58278 23604 58284
rect 23392 58214 23398 58278
rect 23462 58214 23604 58278
rect 23392 58142 23604 58214
rect 23392 58078 23534 58142
rect 23598 58078 23604 58142
rect 23392 58072 23604 58078
rect 28288 58208 28636 58350
rect 110160 58414 110508 58420
rect 110160 58350 110438 58414
rect 110502 58350 110508 58414
rect 110160 58208 110508 58350
rect 116144 58420 116220 58480
rect 116144 58344 116492 58420
rect 116416 58284 116492 58344
rect 115192 58278 115404 58284
rect 115192 58214 115198 58278
rect 115262 58214 115404 58278
rect 28288 58148 28364 58208
rect 110296 58148 110372 58208
rect 28288 57936 28636 58148
rect 110160 57936 110508 58148
rect 115192 58142 115404 58214
rect 115192 58078 115198 58142
rect 115262 58078 115404 58142
rect 115192 58072 115404 58078
rect 115600 58278 115812 58284
rect 115600 58214 115742 58278
rect 115806 58214 115812 58278
rect 115600 58142 115812 58214
rect 115600 58078 115742 58142
rect 115806 58078 115812 58142
rect 115600 58072 115812 58078
rect 116008 58278 116220 58284
rect 116008 58214 116014 58278
rect 116078 58214 116220 58278
rect 116008 58072 116220 58214
rect 116416 58072 116628 58284
rect 116824 58278 117036 58284
rect 116824 58214 116830 58278
rect 116894 58214 117036 58278
rect 116824 58142 117036 58214
rect 116824 58078 116830 58142
rect 116894 58078 117036 58142
rect 116824 58072 117036 58078
rect 116416 58012 116492 58072
rect 116144 57936 116492 58012
rect 28288 57876 28364 57936
rect 110296 57876 110372 57936
rect 116144 57876 116220 57936
rect 21760 57870 21972 57876
rect 21760 57806 21766 57870
rect 21830 57806 21972 57870
rect 21760 57734 21972 57806
rect 21760 57670 21902 57734
rect 21966 57670 21972 57734
rect 21760 57664 21972 57670
rect 22168 57870 22516 57876
rect 22168 57806 22446 57870
rect 22510 57806 22516 57870
rect 22168 57800 22516 57806
rect 22168 57740 22380 57800
rect 22576 57740 22788 57876
rect 22168 57734 22788 57740
rect 22168 57670 22718 57734
rect 22782 57670 22788 57734
rect 22168 57664 22788 57670
rect 22984 57870 23196 57876
rect 22984 57806 22990 57870
rect 23054 57806 23196 57870
rect 22984 57734 23196 57806
rect 22984 57670 23126 57734
rect 23190 57670 23196 57734
rect 22984 57664 23196 57670
rect 23392 57870 23604 57876
rect 23392 57806 23534 57870
rect 23598 57806 23604 57870
rect 23392 57734 23604 57806
rect 23392 57670 23398 57734
rect 23462 57670 23604 57734
rect 23392 57664 23604 57670
rect 28288 57664 28636 57876
rect 110160 57664 110508 57876
rect 115192 57870 115404 57876
rect 115192 57806 115198 57870
rect 115262 57806 115404 57870
rect 115192 57734 115404 57806
rect 115192 57670 115198 57734
rect 115262 57670 115404 57734
rect 115192 57664 115404 57670
rect 115600 57870 115812 57876
rect 115600 57806 115742 57870
rect 115806 57806 115812 57870
rect 115600 57734 115812 57806
rect 115600 57670 115606 57734
rect 115670 57670 115812 57734
rect 115600 57664 115812 57670
rect 116008 57800 116628 57876
rect 116008 57664 116220 57800
rect 116416 57734 116628 57800
rect 116416 57670 116558 57734
rect 116622 57670 116628 57734
rect 116416 57664 116628 57670
rect 116824 57870 117036 57876
rect 116824 57806 116830 57870
rect 116894 57806 117036 57870
rect 116824 57734 117036 57806
rect 116824 57670 116966 57734
rect 117030 57670 117036 57734
rect 116824 57664 117036 57670
rect 28424 57604 28500 57664
rect 110432 57604 110508 57664
rect 1768 57528 1980 57604
rect 1768 57472 1798 57528
rect 1854 57472 1980 57528
rect 1768 57468 1980 57472
rect 1224 57462 1980 57468
rect 1224 57398 1230 57462
rect 1294 57398 1980 57462
rect 1224 57392 1980 57398
rect 21760 57462 21972 57468
rect 21760 57398 21902 57462
rect 21966 57398 21972 57462
rect 21760 57256 21972 57398
rect 22168 57332 22380 57468
rect 22576 57462 22788 57468
rect 22576 57398 22718 57462
rect 22782 57398 22788 57462
rect 22576 57332 22788 57398
rect 22168 57256 22788 57332
rect 22984 57462 23196 57468
rect 22984 57398 23126 57462
rect 23190 57398 23196 57462
rect 22984 57326 23196 57398
rect 22984 57262 23126 57326
rect 23190 57262 23196 57326
rect 22984 57256 23196 57262
rect 23392 57462 23604 57468
rect 23392 57398 23398 57462
rect 23462 57398 23604 57462
rect 23392 57326 23604 57398
rect 28288 57392 28636 57604
rect 110160 57392 110508 57604
rect 136816 57528 137028 57604
rect 136816 57472 136944 57528
rect 137000 57472 137028 57528
rect 136816 57468 137028 57472
rect 115192 57462 115404 57468
rect 115192 57398 115198 57462
rect 115262 57398 115404 57462
rect 28560 57332 28636 57392
rect 110296 57332 110372 57392
rect 23392 57262 23534 57326
rect 23598 57262 23604 57326
rect 23392 57256 23604 57262
rect 21896 57196 21972 57256
rect 21760 56848 21972 57196
rect 22304 57196 22380 57256
rect 22304 57120 22652 57196
rect 22576 57060 22652 57120
rect 28288 57120 28636 57332
rect 110160 57120 110508 57332
rect 115192 57326 115404 57398
rect 115192 57262 115334 57326
rect 115398 57262 115404 57326
rect 115192 57256 115404 57262
rect 115600 57462 115812 57468
rect 115600 57398 115606 57462
rect 115670 57398 115812 57462
rect 115600 57326 115812 57398
rect 115600 57262 115742 57326
rect 115806 57262 115812 57326
rect 115600 57256 115812 57262
rect 116008 57462 116628 57468
rect 116008 57398 116558 57462
rect 116622 57398 116628 57462
rect 116008 57392 116628 57398
rect 116008 57332 116220 57392
rect 116008 57326 116356 57332
rect 116008 57262 116150 57326
rect 116214 57262 116286 57326
rect 116350 57262 116356 57326
rect 116008 57256 116356 57262
rect 116416 57256 116628 57392
rect 116824 57462 117036 57468
rect 116824 57398 116966 57462
rect 117030 57398 117036 57462
rect 116824 57256 117036 57398
rect 136816 57462 137572 57468
rect 136816 57398 137502 57462
rect 137566 57398 137572 57462
rect 136816 57392 137572 57398
rect 116960 57196 117036 57256
rect 28288 57060 28364 57120
rect 110296 57060 110372 57120
rect 22168 56848 22380 57060
rect 22576 56924 22788 57060
rect 22478 56918 22788 56924
rect 22440 56854 22446 56918
rect 22510 56854 22788 56918
rect 22478 56848 22788 56854
rect 22984 57054 23196 57060
rect 22984 56990 23126 57054
rect 23190 56990 23196 57054
rect 22984 56918 23196 56990
rect 22984 56854 22990 56918
rect 23054 56854 23196 56918
rect 22984 56848 23196 56854
rect 23392 57054 23604 57060
rect 23392 56990 23534 57054
rect 23598 56990 23604 57054
rect 23392 56918 23604 56990
rect 23392 56854 23534 56918
rect 23598 56854 23604 56918
rect 23392 56848 23604 56854
rect 28288 56848 28636 57060
rect 110160 56848 110508 57060
rect 115192 57054 115404 57060
rect 115192 56990 115334 57054
rect 115398 56990 115404 57054
rect 115192 56918 115404 56990
rect 115192 56854 115198 56918
rect 115262 56854 115404 56918
rect 115192 56848 115404 56854
rect 115600 57054 115812 57060
rect 115600 56990 115742 57054
rect 115806 56990 115812 57054
rect 115600 56918 115812 56990
rect 115600 56854 115606 56918
rect 115670 56854 115812 56918
rect 115600 56848 115812 56854
rect 116008 57054 116220 57060
rect 116318 57054 116628 57060
rect 116008 56990 116150 57054
rect 116214 56990 116220 57054
rect 116280 56990 116286 57054
rect 116350 56990 116628 57054
rect 116008 56848 116220 56990
rect 116318 56984 116628 56990
rect 21760 56788 21836 56848
rect 22168 56788 22244 56848
rect 21760 56440 21972 56788
rect 22168 56712 22788 56788
rect 22168 56652 22380 56712
rect 22168 56646 22516 56652
rect 22168 56582 22446 56646
rect 22510 56582 22516 56646
rect 22168 56576 22516 56582
rect 22168 56440 22380 56576
rect 22576 56516 22788 56712
rect 28406 56652 28504 56848
rect 110294 56652 110392 56848
rect 116144 56788 116220 56848
rect 22478 56510 22788 56516
rect 22440 56446 22446 56510
rect 22510 56446 22718 56510
rect 22782 56446 22788 56510
rect 22478 56440 22788 56446
rect 22984 56646 23196 56652
rect 22984 56582 22990 56646
rect 23054 56582 23196 56646
rect 22984 56510 23196 56582
rect 22984 56446 22990 56510
rect 23054 56446 23196 56510
rect 22984 56440 23196 56446
rect 23392 56646 23604 56652
rect 23392 56582 23534 56646
rect 23598 56582 23604 56646
rect 23392 56510 23604 56582
rect 28288 56576 28636 56652
rect 110160 56576 110508 56652
rect 28424 56516 28500 56576
rect 110432 56516 110508 56576
rect 23392 56446 23398 56510
rect 23462 56446 23604 56510
rect 23392 56440 23604 56446
rect 21896 56380 21972 56440
rect 21760 56238 21972 56380
rect 28288 56304 28636 56516
rect 110160 56374 110508 56516
rect 115192 56646 115404 56652
rect 115192 56582 115198 56646
rect 115262 56582 115404 56646
rect 115192 56510 115404 56582
rect 115192 56446 115198 56510
rect 115262 56446 115404 56510
rect 115192 56440 115404 56446
rect 115600 56646 115812 56652
rect 115600 56582 115606 56646
rect 115670 56582 115812 56646
rect 115600 56510 115812 56582
rect 115600 56446 115606 56510
rect 115670 56446 115812 56510
rect 115600 56440 115812 56446
rect 116008 56440 116220 56788
rect 116416 56848 116628 56984
rect 116824 56848 117036 57196
rect 116416 56788 116492 56848
rect 116824 56788 116900 56848
rect 116416 56510 116628 56788
rect 116416 56446 116558 56510
rect 116622 56446 116628 56510
rect 116416 56440 116628 56446
rect 116824 56440 117036 56788
rect 110160 56310 110438 56374
rect 110502 56310 110508 56374
rect 110160 56304 110508 56310
rect 116824 56380 116900 56440
rect 28288 56244 28364 56304
rect 110296 56244 110372 56304
rect 21760 56174 21902 56238
rect 21966 56174 21972 56238
rect 21760 56168 21972 56174
rect 22168 56238 22516 56244
rect 22168 56174 22446 56238
rect 22510 56174 22516 56238
rect 22168 56168 22516 56174
rect 22576 56238 22788 56244
rect 22576 56174 22718 56238
rect 22782 56174 22788 56238
rect 22168 56032 22380 56168
rect 22576 56032 22788 56174
rect 22984 56238 23196 56244
rect 22984 56174 22990 56238
rect 23054 56174 23196 56238
rect 22984 56032 23196 56174
rect 23392 56238 23604 56244
rect 23392 56174 23398 56238
rect 23462 56174 23604 56238
rect 23392 56032 23604 56174
rect 22168 55972 22244 56032
rect 22576 55972 22652 56032
rect 23120 55972 23196 56032
rect 23528 55972 23604 56032
rect 1768 55848 1980 55972
rect 1768 55836 1798 55848
rect 1224 55830 1798 55836
rect 1224 55766 1230 55830
rect 1294 55792 1798 55830
rect 1854 55792 1980 55848
rect 1294 55766 1980 55792
rect 1224 55760 1980 55766
rect 21760 55966 21972 55972
rect 21760 55902 21902 55966
rect 21966 55902 21972 55966
rect 21760 55830 21972 55902
rect 21760 55766 21766 55830
rect 21830 55766 21972 55830
rect 21760 55760 21972 55766
rect 22168 55760 22380 55972
rect 22576 55830 22788 55972
rect 22576 55766 22582 55830
rect 22646 55766 22788 55830
rect 22576 55760 22788 55766
rect 22984 55624 23196 55972
rect 23392 55624 23604 55972
rect 28288 55966 28636 56244
rect 28288 55902 28566 55966
rect 28630 55902 28636 55966
rect 28288 55896 28636 55902
rect 110160 56102 110508 56244
rect 110160 56038 110438 56102
rect 110502 56038 110508 56102
rect 110160 55966 110508 56038
rect 115192 56238 115404 56244
rect 115192 56174 115198 56238
rect 115262 56174 115404 56238
rect 115192 56032 115404 56174
rect 115600 56238 115812 56244
rect 115600 56174 115606 56238
rect 115670 56174 115812 56238
rect 115600 56032 115812 56174
rect 115328 55972 115404 56032
rect 115736 55972 115812 56032
rect 110160 55902 110438 55966
rect 110502 55902 110508 55966
rect 110160 55896 110508 55902
rect 22984 55564 23060 55624
rect 23528 55564 23604 55624
rect 21760 55558 21972 55564
rect 21760 55494 21766 55558
rect 21830 55494 21972 55558
rect 21760 55422 21972 55494
rect 21760 55358 21902 55422
rect 21966 55358 21972 55422
rect 21760 55352 21972 55358
rect 22168 55428 22380 55564
rect 22576 55558 22788 55564
rect 22576 55494 22582 55558
rect 22646 55494 22788 55558
rect 22576 55428 22788 55494
rect 22168 55352 22788 55428
rect 22168 55216 22380 55352
rect 22576 55216 22788 55352
rect 22984 55216 23196 55564
rect 22304 55156 22380 55216
rect 22712 55156 22788 55216
rect 23120 55156 23196 55216
rect 21760 55150 21972 55156
rect 21760 55086 21902 55150
rect 21966 55086 21972 55150
rect 21760 55014 21972 55086
rect 21760 54950 21766 55014
rect 21830 54950 21972 55014
rect 21760 54944 21972 54950
rect 22168 55014 22380 55156
rect 22168 54950 22174 55014
rect 22238 54950 22380 55014
rect 22168 54944 22380 54950
rect 22576 54944 22788 55156
rect 22984 55014 23196 55156
rect 22984 54950 22990 55014
rect 23054 54950 23196 55014
rect 22984 54944 23196 54950
rect 23392 55216 23604 55564
rect 28288 55694 28636 55700
rect 28288 55630 28566 55694
rect 28630 55630 28636 55694
rect 28288 55558 28636 55630
rect 28288 55494 28566 55558
rect 28630 55494 28636 55558
rect 28288 55286 28636 55494
rect 28288 55222 28566 55286
rect 28630 55222 28636 55286
rect 23392 55156 23468 55216
rect 23392 55014 23604 55156
rect 28288 55080 28636 55222
rect 110160 55694 110508 55700
rect 110160 55630 110438 55694
rect 110502 55630 110508 55694
rect 110160 55558 110508 55630
rect 110160 55494 110438 55558
rect 110502 55494 110508 55558
rect 110160 55286 110508 55494
rect 110160 55222 110438 55286
rect 110502 55222 110508 55286
rect 110160 55080 110508 55222
rect 28424 55020 28500 55080
rect 110432 55020 110508 55080
rect 23392 54950 23534 55014
rect 23598 54950 23604 55014
rect 23392 54944 23604 54950
rect 21760 54742 21972 54748
rect 21760 54678 21766 54742
rect 21830 54678 21972 54742
rect 21760 54606 21972 54678
rect 21760 54542 21902 54606
rect 21966 54542 21972 54606
rect 21760 54536 21972 54542
rect 22168 54742 22380 54748
rect 22168 54678 22174 54742
rect 22238 54678 22380 54742
rect 22168 54606 22380 54678
rect 22576 54612 22788 54748
rect 22478 54606 22788 54612
rect 22168 54542 22310 54606
rect 22374 54542 22380 54606
rect 22440 54542 22446 54606
rect 22510 54542 22788 54606
rect 22168 54536 22380 54542
rect 22478 54536 22788 54542
rect 22984 54742 23196 54748
rect 22984 54678 22990 54742
rect 23054 54678 23196 54742
rect 22984 54606 23196 54678
rect 22984 54542 22990 54606
rect 23054 54542 23196 54606
rect 22984 54536 23196 54542
rect 23392 54742 23604 54748
rect 23392 54678 23534 54742
rect 23598 54678 23604 54742
rect 23392 54606 23604 54678
rect 23392 54542 23534 54606
rect 23598 54542 23604 54606
rect 23392 54536 23604 54542
rect 28288 54742 28636 55020
rect 28288 54678 28294 54742
rect 28358 54678 28636 54742
rect 28288 54536 28636 54678
rect 110160 54536 110508 55020
rect 115192 55624 115404 55972
rect 115600 55624 115812 55972
rect 116008 56108 116220 56244
rect 116416 56238 116628 56244
rect 116416 56174 116558 56238
rect 116622 56174 116628 56238
rect 116416 56108 116628 56174
rect 116824 56238 117036 56380
rect 116824 56174 116966 56238
rect 117030 56174 117036 56238
rect 116824 56168 117036 56174
rect 116008 56032 116628 56108
rect 116008 55972 116084 56032
rect 116416 55972 116492 56032
rect 116008 55760 116220 55972
rect 116416 55830 116628 55972
rect 116416 55766 116558 55830
rect 116622 55766 116628 55830
rect 116416 55760 116628 55766
rect 116824 55966 117036 55972
rect 116824 55902 116966 55966
rect 117030 55902 117036 55966
rect 116824 55830 117036 55902
rect 116824 55766 116966 55830
rect 117030 55766 117036 55830
rect 116824 55760 117036 55766
rect 136816 55848 137028 55972
rect 136816 55792 136944 55848
rect 137000 55836 137028 55848
rect 137000 55830 137572 55836
rect 137000 55792 137502 55830
rect 136816 55766 137502 55792
rect 137566 55766 137572 55830
rect 136816 55760 137572 55766
rect 115192 55564 115268 55624
rect 115736 55564 115812 55624
rect 115192 55216 115404 55564
rect 115600 55216 115812 55564
rect 116008 55292 116220 55564
rect 116416 55558 116628 55564
rect 116416 55494 116558 55558
rect 116622 55494 116628 55558
rect 116416 55292 116628 55494
rect 116824 55558 117036 55564
rect 116824 55494 116966 55558
rect 117030 55494 117036 55558
rect 116824 55422 117036 55494
rect 116824 55358 116966 55422
rect 117030 55358 117036 55422
rect 116824 55352 117036 55358
rect 116008 55216 116628 55292
rect 115192 55156 115268 55216
rect 115600 55156 115676 55216
rect 116144 55156 116220 55216
rect 116552 55156 116628 55216
rect 115192 55014 115404 55156
rect 115192 54950 115198 55014
rect 115262 54950 115404 55014
rect 115192 54944 115404 54950
rect 115600 55014 115812 55156
rect 115600 54950 115742 55014
rect 115806 54950 115812 55014
rect 115600 54944 115812 54950
rect 116008 55020 116220 55156
rect 116008 55014 116356 55020
rect 116008 54950 116286 55014
rect 116350 54950 116356 55014
rect 116008 54944 116356 54950
rect 116416 54944 116628 55156
rect 116824 55150 117036 55156
rect 116824 55086 116966 55150
rect 117030 55086 117036 55150
rect 116824 55014 117036 55086
rect 116824 54950 116830 55014
rect 116894 54950 117036 55014
rect 116824 54944 117036 54950
rect 115192 54742 115404 54748
rect 115192 54678 115198 54742
rect 115262 54678 115404 54742
rect 115192 54606 115404 54678
rect 115192 54542 115334 54606
rect 115398 54542 115404 54606
rect 115192 54536 115404 54542
rect 115600 54742 115812 54748
rect 115600 54678 115742 54742
rect 115806 54678 115812 54742
rect 115600 54606 115812 54678
rect 115600 54542 115742 54606
rect 115806 54542 115812 54606
rect 115600 54536 115812 54542
rect 116008 54606 116220 54748
rect 116318 54742 116628 54748
rect 116280 54678 116286 54742
rect 116350 54678 116628 54742
rect 116318 54672 116628 54678
rect 116416 54612 116628 54672
rect 116318 54606 116628 54612
rect 116008 54542 116150 54606
rect 116214 54542 116220 54606
rect 116280 54542 116286 54606
rect 116350 54542 116628 54606
rect 116008 54536 116220 54542
rect 116318 54536 116628 54542
rect 116824 54742 117036 54748
rect 116824 54678 116830 54742
rect 116894 54678 117036 54742
rect 116824 54606 117036 54678
rect 116824 54542 116830 54606
rect 116894 54542 117036 54606
rect 116824 54536 117036 54542
rect 28288 54476 28364 54536
rect 110296 54476 110372 54536
rect 28288 54470 28636 54476
rect 28288 54406 28294 54470
rect 28358 54406 28636 54470
rect 21760 54334 21972 54340
rect 21760 54270 21902 54334
rect 21966 54270 21972 54334
rect 1224 54198 1980 54204
rect 1224 54134 1230 54198
rect 1294 54168 1980 54198
rect 1294 54134 1798 54168
rect 1224 54128 1798 54134
rect 1768 54112 1798 54128
rect 1854 54112 1980 54168
rect 21760 54198 21972 54270
rect 21760 54134 21902 54198
rect 21966 54134 21972 54198
rect 21760 54128 21972 54134
rect 22168 54334 22516 54340
rect 22168 54270 22310 54334
rect 22374 54270 22446 54334
rect 22510 54270 22516 54334
rect 22168 54264 22516 54270
rect 22168 54204 22380 54264
rect 22576 54204 22788 54340
rect 22168 54198 22788 54204
rect 22168 54134 22174 54198
rect 22238 54134 22788 54198
rect 22168 54128 22788 54134
rect 22984 54334 23196 54340
rect 22984 54270 22990 54334
rect 23054 54270 23196 54334
rect 22984 54198 23196 54270
rect 22984 54134 22990 54198
rect 23054 54134 23196 54198
rect 22984 54128 23196 54134
rect 23392 54334 23604 54340
rect 23392 54270 23534 54334
rect 23598 54270 23604 54334
rect 23392 54198 23604 54270
rect 28288 54264 28636 54406
rect 110160 54264 110508 54476
rect 115192 54334 115404 54340
rect 115192 54270 115334 54334
rect 115398 54270 115404 54334
rect 28424 54204 28500 54264
rect 110296 54204 110372 54264
rect 23392 54134 23398 54198
rect 23462 54134 23604 54198
rect 23392 54128 23604 54134
rect 1768 53992 1980 54112
rect 28288 53992 28636 54204
rect 110160 53992 110508 54204
rect 115192 54198 115404 54270
rect 115192 54134 115334 54198
rect 115398 54134 115404 54198
rect 115192 54128 115404 54134
rect 115600 54334 115812 54340
rect 115600 54270 115742 54334
rect 115806 54270 115812 54334
rect 115600 54198 115812 54270
rect 115600 54134 115606 54198
rect 115670 54134 115812 54198
rect 115600 54128 115812 54134
rect 116008 54334 116356 54340
rect 116008 54270 116150 54334
rect 116214 54270 116286 54334
rect 116350 54270 116356 54334
rect 116008 54264 116356 54270
rect 116008 54204 116220 54264
rect 116416 54204 116628 54340
rect 116008 54198 116628 54204
rect 116008 54134 116014 54198
rect 116078 54134 116422 54198
rect 116486 54134 116628 54198
rect 116008 54128 116628 54134
rect 116824 54334 117036 54340
rect 116824 54270 116830 54334
rect 116894 54270 117036 54334
rect 116824 54198 117036 54270
rect 116824 54134 116830 54198
rect 116894 54134 117036 54198
rect 116824 54128 117036 54134
rect 136816 54198 137572 54204
rect 136816 54168 137502 54198
rect 136816 54112 136944 54168
rect 137000 54134 137502 54168
rect 137566 54134 137572 54198
rect 137000 54128 137572 54134
rect 137000 54112 137028 54128
rect 136816 53992 137028 54112
rect 28288 53932 28364 53992
rect 110432 53932 110508 53992
rect 21760 53926 21972 53932
rect 21760 53862 21902 53926
rect 21966 53862 21972 53926
rect 21760 53790 21972 53862
rect 21760 53726 21766 53790
rect 21830 53726 21972 53790
rect 21760 53720 21972 53726
rect 22168 53926 22380 53932
rect 22168 53862 22174 53926
rect 22238 53862 22380 53926
rect 22168 53796 22380 53862
rect 22576 53796 22788 53932
rect 22168 53790 22788 53796
rect 22168 53726 22174 53790
rect 22238 53726 22582 53790
rect 22646 53726 22788 53790
rect 22168 53720 22788 53726
rect 22984 53926 23196 53932
rect 22984 53862 22990 53926
rect 23054 53862 23196 53926
rect 22984 53790 23196 53862
rect 22984 53726 23126 53790
rect 23190 53726 23196 53790
rect 22984 53720 23196 53726
rect 23392 53926 23604 53932
rect 23392 53862 23398 53926
rect 23462 53862 23604 53926
rect 23392 53790 23604 53862
rect 23392 53726 23534 53790
rect 23598 53726 23604 53790
rect 23392 53720 23604 53726
rect 28288 53720 28636 53932
rect 110160 53720 110508 53932
rect 115192 53926 115404 53932
rect 115192 53862 115334 53926
rect 115398 53862 115404 53926
rect 115192 53790 115404 53862
rect 115192 53726 115334 53790
rect 115398 53726 115404 53790
rect 115192 53720 115404 53726
rect 115600 53926 115812 53932
rect 115600 53862 115606 53926
rect 115670 53862 115812 53926
rect 115600 53790 115812 53862
rect 115600 53726 115742 53790
rect 115806 53726 115812 53790
rect 115600 53720 115812 53726
rect 116008 53926 116220 53932
rect 116008 53862 116014 53926
rect 116078 53862 116220 53926
rect 116008 53720 116220 53862
rect 116416 53926 116628 53932
rect 116416 53862 116422 53926
rect 116486 53862 116628 53926
rect 116416 53796 116628 53862
rect 116318 53790 116628 53796
rect 116280 53726 116286 53790
rect 116350 53726 116628 53790
rect 116318 53720 116628 53726
rect 116824 53926 117036 53932
rect 116824 53862 116830 53926
rect 116894 53862 117036 53926
rect 116824 53790 117036 53862
rect 116824 53726 116830 53790
rect 116894 53726 117036 53790
rect 116824 53720 117036 53726
rect 28288 53660 28364 53720
rect 110160 53660 110236 53720
rect 21760 53518 21972 53524
rect 21760 53454 21766 53518
rect 21830 53454 21972 53518
rect 21760 53312 21972 53454
rect 22168 53518 22380 53524
rect 22168 53454 22174 53518
rect 22238 53454 22380 53518
rect 22168 53312 22380 53454
rect 22576 53518 22788 53524
rect 22576 53454 22582 53518
rect 22646 53454 22788 53518
rect 22576 53382 22788 53454
rect 22576 53318 22718 53382
rect 22782 53318 22788 53382
rect 22576 53312 22788 53318
rect 22984 53518 23196 53524
rect 22984 53454 23126 53518
rect 23190 53454 23196 53518
rect 22984 53382 23196 53454
rect 22984 53318 22990 53382
rect 23054 53318 23196 53382
rect 22984 53312 23196 53318
rect 23392 53518 23604 53524
rect 23392 53454 23534 53518
rect 23598 53454 23604 53518
rect 23392 53382 23604 53454
rect 28288 53448 28636 53660
rect 110160 53448 110508 53660
rect 28424 53388 28500 53448
rect 110432 53388 110508 53448
rect 23392 53318 23398 53382
rect 23462 53318 23604 53382
rect 23392 53312 23604 53318
rect 21760 53252 21836 53312
rect 21760 52974 21972 53252
rect 28288 53176 28636 53388
rect 28560 53116 28636 53176
rect 21760 52910 21766 52974
rect 21830 52910 21972 52974
rect 21760 52904 21972 52910
rect 22168 53110 22788 53116
rect 22168 53046 22718 53110
rect 22782 53046 22788 53110
rect 22168 53040 22788 53046
rect 22168 52980 22380 53040
rect 22168 52974 22516 52980
rect 22168 52910 22446 52974
rect 22510 52910 22516 52974
rect 22168 52904 22516 52910
rect 22576 52904 22788 53040
rect 22984 53110 23196 53116
rect 22984 53046 22990 53110
rect 23054 53046 23196 53110
rect 22984 52974 23196 53046
rect 22984 52910 23126 52974
rect 23190 52910 23196 52974
rect 22984 52904 23196 52910
rect 23392 53110 23604 53116
rect 23392 53046 23398 53110
rect 23462 53046 23604 53110
rect 23392 52974 23604 53046
rect 23392 52910 23534 52974
rect 23598 52910 23604 52974
rect 23392 52904 23604 52910
rect 28288 52904 28636 53116
rect 110160 53176 110508 53388
rect 115192 53518 115404 53524
rect 115192 53454 115334 53518
rect 115398 53454 115404 53518
rect 115192 53382 115404 53454
rect 115192 53318 115198 53382
rect 115262 53318 115404 53382
rect 115192 53312 115404 53318
rect 115600 53518 115812 53524
rect 115600 53454 115742 53518
rect 115806 53454 115812 53518
rect 115600 53382 115812 53454
rect 115600 53318 115606 53382
rect 115670 53318 115812 53382
rect 115600 53312 115812 53318
rect 116008 53518 116356 53524
rect 116008 53454 116286 53518
rect 116350 53454 116356 53518
rect 116008 53448 116356 53454
rect 116008 53388 116220 53448
rect 116416 53388 116628 53524
rect 116008 53382 116628 53388
rect 116008 53318 116558 53382
rect 116622 53318 116628 53382
rect 116008 53312 116628 53318
rect 116824 53518 117036 53524
rect 116824 53454 116830 53518
rect 116894 53454 117036 53518
rect 116824 53312 117036 53454
rect 116824 53252 116900 53312
rect 110160 53116 110236 53176
rect 110160 52904 110508 53116
rect 115192 53110 115404 53116
rect 115192 53046 115198 53110
rect 115262 53046 115404 53110
rect 115192 52974 115404 53046
rect 115192 52910 115334 52974
rect 115398 52910 115404 52974
rect 115192 52904 115404 52910
rect 115600 53110 115812 53116
rect 115600 53046 115606 53110
rect 115670 53046 115812 53110
rect 115600 52974 115812 53046
rect 115600 52910 115742 52974
rect 115806 52910 115812 52974
rect 115600 52904 115812 52910
rect 116008 52980 116220 53116
rect 116416 53110 116628 53116
rect 116416 53046 116558 53110
rect 116622 53046 116628 53110
rect 116008 52974 116356 52980
rect 116008 52910 116150 52974
rect 116214 52910 116286 52974
rect 116350 52910 116356 52974
rect 116008 52904 116356 52910
rect 116416 52974 116628 53046
rect 116416 52910 116422 52974
rect 116486 52910 116628 52974
rect 116416 52904 116628 52910
rect 116824 52974 117036 53252
rect 116824 52910 116830 52974
rect 116894 52910 117036 52974
rect 116824 52904 117036 52910
rect 28288 52844 28364 52904
rect 110296 52844 110372 52904
rect 21760 52702 21972 52708
rect 21760 52638 21766 52702
rect 21830 52638 21972 52702
rect 1224 52566 1980 52572
rect 1224 52502 1230 52566
rect 1294 52502 1980 52566
rect 1224 52496 1980 52502
rect 1768 52488 1980 52496
rect 1768 52432 1798 52488
rect 1854 52432 1980 52488
rect 1768 52360 1980 52432
rect 21760 52496 21972 52638
rect 22168 52566 22380 52708
rect 22478 52702 22788 52708
rect 22440 52638 22446 52702
rect 22510 52638 22788 52702
rect 22478 52632 22788 52638
rect 22168 52502 22174 52566
rect 22238 52502 22380 52566
rect 22168 52496 22380 52502
rect 22576 52566 22788 52632
rect 22576 52502 22718 52566
rect 22782 52502 22788 52566
rect 22576 52496 22788 52502
rect 22984 52702 23196 52708
rect 22984 52638 23126 52702
rect 23190 52638 23196 52702
rect 22984 52566 23196 52638
rect 22984 52502 22990 52566
rect 23054 52502 23196 52566
rect 22984 52496 23196 52502
rect 23392 52702 23604 52708
rect 23392 52638 23534 52702
rect 23598 52638 23604 52702
rect 23392 52566 23604 52638
rect 23392 52502 23398 52566
rect 23462 52502 23604 52566
rect 23392 52496 23604 52502
rect 28288 52632 28636 52844
rect 110160 52632 110508 52844
rect 28288 52572 28364 52632
rect 110432 52572 110508 52632
rect 21760 52436 21836 52496
rect 21760 52294 21972 52436
rect 28288 52360 28636 52572
rect 110160 52430 110508 52572
rect 115192 52702 115404 52708
rect 115192 52638 115334 52702
rect 115398 52638 115404 52702
rect 115192 52566 115404 52638
rect 115192 52502 115334 52566
rect 115398 52502 115404 52566
rect 115192 52496 115404 52502
rect 115600 52702 115812 52708
rect 115600 52638 115742 52702
rect 115806 52638 115812 52702
rect 115600 52566 115812 52638
rect 115600 52502 115742 52566
rect 115806 52502 115812 52566
rect 115600 52496 115812 52502
rect 116008 52702 116220 52708
rect 116318 52702 116628 52708
rect 116008 52638 116150 52702
rect 116214 52638 116220 52702
rect 116280 52638 116286 52702
rect 116350 52638 116422 52702
rect 116486 52638 116628 52702
rect 116008 52572 116220 52638
rect 116318 52632 116628 52638
rect 116008 52566 116356 52572
rect 116008 52502 116014 52566
rect 116078 52502 116286 52566
rect 116350 52502 116356 52566
rect 116008 52496 116356 52502
rect 116416 52496 116628 52632
rect 116824 52702 117036 52708
rect 116824 52638 116830 52702
rect 116894 52638 117036 52702
rect 116824 52496 117036 52638
rect 136816 52566 137572 52572
rect 136816 52502 137502 52566
rect 137566 52502 137572 52566
rect 136816 52496 137572 52502
rect 110160 52366 110438 52430
rect 110502 52366 110508 52430
rect 110160 52360 110508 52366
rect 116824 52436 116900 52496
rect 136816 52488 137028 52496
rect 28424 52300 28500 52360
rect 110160 52300 110236 52360
rect 21760 52230 21902 52294
rect 21966 52230 21972 52294
rect 21760 52224 21972 52230
rect 22168 52294 22380 52300
rect 22168 52230 22174 52294
rect 22238 52230 22380 52294
rect 22168 52088 22380 52230
rect 22576 52294 22788 52300
rect 22576 52230 22718 52294
rect 22782 52230 22788 52294
rect 22576 52164 22788 52230
rect 22304 52028 22380 52088
rect 22440 52088 22788 52164
rect 22984 52294 23196 52300
rect 22984 52230 22990 52294
rect 23054 52230 23196 52294
rect 22984 52158 23196 52230
rect 22984 52094 22990 52158
rect 23054 52094 23196 52158
rect 22984 52088 23196 52094
rect 23392 52294 23604 52300
rect 23392 52230 23398 52294
rect 23462 52230 23604 52294
rect 23392 52158 23604 52230
rect 23392 52094 23398 52158
rect 23462 52094 23604 52158
rect 23392 52088 23604 52094
rect 22440 52028 22516 52088
rect 21760 52022 21972 52028
rect 21760 51958 21902 52022
rect 21966 51958 21972 52022
rect 21760 51680 21972 51958
rect 22168 51952 22516 52028
rect 22168 51892 22380 51952
rect 22576 51892 22788 52028
rect 22168 51816 22788 51892
rect 22168 51750 22380 51816
rect 22168 51686 22174 51750
rect 22238 51686 22380 51750
rect 22168 51680 22380 51686
rect 22576 51680 22788 51816
rect 22984 51886 23196 51892
rect 22984 51822 22990 51886
rect 23054 51822 23196 51886
rect 22984 51680 23196 51822
rect 23392 51886 23604 51892
rect 23392 51822 23398 51886
rect 23462 51822 23604 51886
rect 23392 51680 23604 51822
rect 21896 51620 21972 51680
rect 23120 51620 23196 51680
rect 23528 51620 23604 51680
rect 21760 51478 21972 51620
rect 21760 51414 21766 51478
rect 21830 51414 21972 51478
rect 21760 51408 21972 51414
rect 22168 51478 22380 51484
rect 22168 51414 22174 51478
rect 22238 51414 22380 51478
rect 22168 51272 22380 51414
rect 22576 51348 22788 51484
rect 22440 51272 22788 51348
rect 22984 51272 23196 51620
rect 23392 51272 23604 51620
rect 28288 51886 28636 52300
rect 28288 51822 28430 51886
rect 28494 51822 28636 51886
rect 28288 51816 28636 51822
rect 110160 52158 110508 52300
rect 110160 52094 110438 52158
rect 110502 52094 110508 52158
rect 110160 51816 110508 52094
rect 115192 52294 115404 52300
rect 115192 52230 115334 52294
rect 115398 52230 115404 52294
rect 115192 52158 115404 52230
rect 115192 52094 115198 52158
rect 115262 52094 115404 52158
rect 115192 52088 115404 52094
rect 115600 52294 115812 52300
rect 115600 52230 115742 52294
rect 115806 52230 115812 52294
rect 115600 52158 115812 52230
rect 115600 52094 115606 52158
rect 115670 52094 115812 52158
rect 115600 52088 115812 52094
rect 116008 52294 116220 52300
rect 116318 52294 116628 52300
rect 116008 52230 116014 52294
rect 116078 52230 116220 52294
rect 116280 52230 116286 52294
rect 116350 52230 116628 52294
rect 116008 52088 116220 52230
rect 116318 52224 116628 52230
rect 116824 52294 117036 52436
rect 136816 52432 136944 52488
rect 137000 52432 137028 52488
rect 136816 52360 137028 52432
rect 116824 52230 116966 52294
rect 117030 52230 117036 52294
rect 116824 52224 117036 52230
rect 116416 52088 116628 52224
rect 116008 52028 116084 52088
rect 115192 51886 115404 51892
rect 115192 51822 115198 51886
rect 115262 51822 115404 51886
rect 28288 51756 28364 51816
rect 110296 51756 110372 51816
rect 28288 51614 28636 51756
rect 28288 51550 28430 51614
rect 28494 51550 28566 51614
rect 28630 51550 28636 51614
rect 28288 51342 28636 51550
rect 28288 51278 28566 51342
rect 28630 51278 28636 51342
rect 22168 51212 22244 51272
rect 22440 51212 22516 51272
rect 21760 51206 21972 51212
rect 21760 51142 21766 51206
rect 21830 51142 21972 51206
rect 21760 51070 21972 51142
rect 21760 51006 21902 51070
rect 21966 51006 21972 51070
rect 21760 51000 21972 51006
rect 22168 51136 22516 51212
rect 22576 51212 22652 51272
rect 22984 51212 23060 51272
rect 23392 51212 23468 51272
rect 22168 51076 22380 51136
rect 22168 51070 22516 51076
rect 22168 51006 22310 51070
rect 22374 51006 22446 51070
rect 22510 51006 22516 51070
rect 22168 51000 22516 51006
rect 22576 51000 22788 51212
rect 22984 51070 23196 51212
rect 22984 51006 22990 51070
rect 23054 51006 23196 51070
rect 22984 51000 23196 51006
rect 23392 51070 23604 51212
rect 28288 51136 28636 51278
rect 28560 51076 28636 51136
rect 23392 51006 23398 51070
rect 23462 51006 23604 51070
rect 23392 51000 23604 51006
rect 1224 50934 1980 50940
rect 1224 50870 1230 50934
rect 1294 50870 1980 50934
rect 1224 50864 1980 50870
rect 1768 50808 1980 50864
rect 1768 50752 1798 50808
rect 1854 50752 1980 50808
rect 1768 50728 1980 50752
rect 21760 50798 21972 50804
rect 21760 50734 21902 50798
rect 21966 50734 21972 50798
rect 21760 50662 21972 50734
rect 21760 50598 21766 50662
rect 21830 50598 21972 50662
rect 21760 50592 21972 50598
rect 22168 50798 22380 50804
rect 22478 50798 22788 50804
rect 22168 50734 22310 50798
rect 22374 50734 22380 50798
rect 22440 50734 22446 50798
rect 22510 50734 22788 50798
rect 22168 50662 22380 50734
rect 22478 50728 22788 50734
rect 22168 50598 22174 50662
rect 22238 50598 22380 50662
rect 22168 50592 22380 50598
rect 22576 50662 22788 50728
rect 22576 50598 22582 50662
rect 22646 50598 22788 50662
rect 22576 50592 22788 50598
rect 22984 50798 23196 50804
rect 22984 50734 22990 50798
rect 23054 50734 23196 50798
rect 22984 50662 23196 50734
rect 22984 50598 22990 50662
rect 23054 50598 23196 50662
rect 22984 50592 23196 50598
rect 23392 50798 23604 50804
rect 23392 50734 23398 50798
rect 23462 50734 23604 50798
rect 23392 50662 23604 50734
rect 23392 50598 23534 50662
rect 23598 50598 23604 50662
rect 23392 50592 23604 50598
rect 28288 50592 28636 51076
rect 110160 51136 110508 51756
rect 115192 51680 115404 51822
rect 115600 51886 115812 51892
rect 115600 51822 115606 51886
rect 115670 51822 115812 51886
rect 115600 51680 115812 51822
rect 116008 51750 116220 52028
rect 116008 51686 116014 51750
rect 116078 51686 116220 51750
rect 116008 51680 116220 51686
rect 116416 51750 116628 52028
rect 116416 51686 116422 51750
rect 116486 51686 116628 51750
rect 116416 51680 116628 51686
rect 116824 52022 117036 52028
rect 116824 51958 116966 52022
rect 117030 51958 117036 52022
rect 116824 51680 117036 51958
rect 115328 51620 115404 51680
rect 115736 51620 115812 51680
rect 115192 51272 115404 51620
rect 115328 51212 115404 51272
rect 110160 51076 110236 51136
rect 110160 50798 110508 51076
rect 115192 51070 115404 51212
rect 115192 51006 115198 51070
rect 115262 51006 115404 51070
rect 115192 51000 115404 51006
rect 115600 51272 115812 51620
rect 116824 51620 116900 51680
rect 116008 51478 116220 51484
rect 116008 51414 116014 51478
rect 116078 51414 116220 51478
rect 116008 51348 116220 51414
rect 116416 51478 116628 51484
rect 116416 51414 116422 51478
rect 116486 51414 116628 51478
rect 116008 51272 116356 51348
rect 115600 51212 115676 51272
rect 116144 51212 116220 51272
rect 115600 51070 115812 51212
rect 115600 51006 115606 51070
rect 115670 51006 115812 51070
rect 115600 51000 115812 51006
rect 116008 51000 116220 51212
rect 116280 51212 116356 51272
rect 116416 51272 116628 51414
rect 116824 51478 117036 51620
rect 116824 51414 116830 51478
rect 116894 51414 117036 51478
rect 116824 51408 117036 51414
rect 116416 51212 116492 51272
rect 116280 51136 116628 51212
rect 116416 51070 116628 51136
rect 116416 51006 116558 51070
rect 116622 51006 116628 51070
rect 116416 51000 116628 51006
rect 116824 51206 117036 51212
rect 116824 51142 116830 51206
rect 116894 51142 117036 51206
rect 116824 51070 117036 51142
rect 116824 51006 116830 51070
rect 116894 51006 117036 51070
rect 116824 51000 117036 51006
rect 136816 50934 137572 50940
rect 136816 50870 137502 50934
rect 137566 50870 137572 50934
rect 136816 50864 137572 50870
rect 136816 50808 137028 50864
rect 110160 50734 110438 50798
rect 110502 50734 110508 50798
rect 110160 50592 110508 50734
rect 115192 50798 115404 50804
rect 115192 50734 115198 50798
rect 115262 50734 115404 50798
rect 115192 50662 115404 50734
rect 115192 50598 115334 50662
rect 115398 50598 115404 50662
rect 115192 50592 115404 50598
rect 115600 50798 115812 50804
rect 115600 50734 115606 50798
rect 115670 50734 115812 50798
rect 115600 50662 115812 50734
rect 115600 50598 115742 50662
rect 115806 50598 115812 50662
rect 115600 50592 115812 50598
rect 116008 50662 116220 50804
rect 116008 50598 116014 50662
rect 116078 50598 116220 50662
rect 116008 50592 116220 50598
rect 116416 50798 116628 50804
rect 116416 50734 116558 50798
rect 116622 50734 116628 50798
rect 116416 50662 116628 50734
rect 116416 50598 116422 50662
rect 116486 50598 116628 50662
rect 116416 50592 116628 50598
rect 116824 50798 117036 50804
rect 116824 50734 116830 50798
rect 116894 50734 117036 50798
rect 116824 50662 117036 50734
rect 136816 50752 136944 50808
rect 137000 50752 137028 50808
rect 136816 50728 137028 50752
rect 116824 50598 116830 50662
rect 116894 50598 117036 50662
rect 116824 50592 117036 50598
rect 28424 50532 28500 50592
rect 110432 50532 110508 50592
rect 21760 50390 21972 50396
rect 21760 50326 21766 50390
rect 21830 50326 21972 50390
rect 21760 50254 21972 50326
rect 21760 50190 21902 50254
rect 21966 50190 21972 50254
rect 21760 50184 21972 50190
rect 22168 50390 22380 50396
rect 22168 50326 22174 50390
rect 22238 50326 22380 50390
rect 22168 50184 22380 50326
rect 22576 50390 22788 50396
rect 22576 50326 22582 50390
rect 22646 50326 22788 50390
rect 22576 50260 22788 50326
rect 22478 50254 22788 50260
rect 22440 50190 22446 50254
rect 22510 50190 22788 50254
rect 22478 50184 22788 50190
rect 22984 50390 23196 50396
rect 22984 50326 22990 50390
rect 23054 50326 23196 50390
rect 22984 50254 23196 50326
rect 22984 50190 23126 50254
rect 23190 50190 23196 50254
rect 22984 50184 23196 50190
rect 23392 50390 23604 50396
rect 23392 50326 23534 50390
rect 23598 50326 23604 50390
rect 23392 50254 23604 50326
rect 23392 50190 23534 50254
rect 23598 50190 23604 50254
rect 23392 50184 23604 50190
rect 28288 50320 28636 50532
rect 110160 50526 110508 50532
rect 110160 50462 110438 50526
rect 110502 50462 110508 50526
rect 110160 50320 110508 50462
rect 115192 50390 115404 50396
rect 115192 50326 115334 50390
rect 115398 50326 115404 50390
rect 28288 50260 28364 50320
rect 110296 50260 110372 50320
rect 28288 50048 28636 50260
rect 110160 50048 110508 50260
rect 115192 50254 115404 50326
rect 115192 50190 115334 50254
rect 115398 50190 115404 50254
rect 115192 50184 115404 50190
rect 115600 50390 115812 50396
rect 115600 50326 115742 50390
rect 115806 50326 115812 50390
rect 115600 50254 115812 50326
rect 115600 50190 115606 50254
rect 115670 50190 115812 50254
rect 115600 50184 115812 50190
rect 116008 50390 116220 50396
rect 116008 50326 116014 50390
rect 116078 50326 116220 50390
rect 116008 50254 116220 50326
rect 116416 50390 116628 50396
rect 116416 50326 116422 50390
rect 116486 50326 116628 50390
rect 116416 50260 116628 50326
rect 116318 50254 116628 50260
rect 116008 50190 116150 50254
rect 116214 50190 116220 50254
rect 116280 50190 116286 50254
rect 116350 50190 116628 50254
rect 116008 50184 116220 50190
rect 116318 50184 116628 50190
rect 116824 50390 117036 50396
rect 116824 50326 116830 50390
rect 116894 50326 117036 50390
rect 116824 50254 117036 50326
rect 116824 50190 116966 50254
rect 117030 50190 117036 50254
rect 116824 50184 117036 50190
rect 28288 49988 28364 50048
rect 110432 49988 110508 50048
rect 21760 49982 21972 49988
rect 21760 49918 21902 49982
rect 21966 49918 21972 49982
rect 21760 49846 21972 49918
rect 21760 49782 21902 49846
rect 21966 49782 21972 49846
rect 21760 49776 21972 49782
rect 22168 49982 22516 49988
rect 22168 49918 22446 49982
rect 22510 49918 22516 49982
rect 22168 49912 22516 49918
rect 22168 49852 22380 49912
rect 22576 49852 22788 49988
rect 22168 49846 22788 49852
rect 22168 49782 22174 49846
rect 22238 49782 22582 49846
rect 22646 49782 22788 49846
rect 22168 49776 22788 49782
rect 22984 49982 23196 49988
rect 22984 49918 23126 49982
rect 23190 49918 23196 49982
rect 22984 49846 23196 49918
rect 22984 49782 22990 49846
rect 23054 49782 23196 49846
rect 22984 49776 23196 49782
rect 23392 49982 23604 49988
rect 23392 49918 23534 49982
rect 23598 49918 23604 49982
rect 23392 49846 23604 49918
rect 23392 49782 23534 49846
rect 23598 49782 23604 49846
rect 23392 49776 23604 49782
rect 28288 49776 28636 49988
rect 110160 49776 110508 49988
rect 115192 49982 115404 49988
rect 115192 49918 115334 49982
rect 115398 49918 115404 49982
rect 115192 49846 115404 49918
rect 115192 49782 115334 49846
rect 115398 49782 115404 49846
rect 115192 49776 115404 49782
rect 115600 49982 115812 49988
rect 115600 49918 115606 49982
rect 115670 49918 115812 49982
rect 115600 49846 115812 49918
rect 115600 49782 115742 49846
rect 115806 49782 115812 49846
rect 115600 49776 115812 49782
rect 116008 49982 116356 49988
rect 116008 49918 116150 49982
rect 116214 49918 116286 49982
rect 116350 49918 116356 49982
rect 116008 49912 116356 49918
rect 116008 49852 116220 49912
rect 116416 49852 116628 49988
rect 116008 49846 116628 49852
rect 116008 49782 116014 49846
rect 116078 49782 116628 49846
rect 116008 49776 116628 49782
rect 116824 49982 117036 49988
rect 116824 49918 116966 49982
rect 117030 49918 117036 49982
rect 116824 49846 117036 49918
rect 116824 49782 116966 49846
rect 117030 49782 117036 49846
rect 116824 49776 117036 49782
rect 28424 49716 28500 49776
rect 110160 49716 110236 49776
rect 116144 49716 116220 49776
rect 21760 49574 21972 49580
rect 21760 49510 21902 49574
rect 21966 49510 21972 49574
rect 21760 49438 21972 49510
rect 21760 49374 21766 49438
rect 21830 49374 21972 49438
rect 21760 49368 21972 49374
rect 22168 49574 22380 49580
rect 22168 49510 22174 49574
rect 22238 49510 22380 49574
rect 22168 49368 22380 49510
rect 22576 49574 22788 49580
rect 22576 49510 22582 49574
rect 22646 49510 22788 49574
rect 22576 49438 22788 49510
rect 22576 49374 22582 49438
rect 22646 49374 22788 49438
rect 22576 49368 22788 49374
rect 22984 49574 23196 49580
rect 22984 49510 22990 49574
rect 23054 49510 23196 49574
rect 22984 49438 23196 49510
rect 22984 49374 22990 49438
rect 23054 49374 23196 49438
rect 22984 49368 23196 49374
rect 23392 49574 23604 49580
rect 23392 49510 23534 49574
rect 23598 49510 23604 49574
rect 23392 49438 23604 49510
rect 23392 49374 23534 49438
rect 23598 49374 23604 49438
rect 23392 49368 23604 49374
rect 28288 49504 28636 49716
rect 110160 49504 110508 49716
rect 116144 49640 116492 49716
rect 116416 49580 116492 49640
rect 115192 49574 115404 49580
rect 115192 49510 115334 49574
rect 115398 49510 115404 49574
rect 28288 49444 28364 49504
rect 110296 49444 110372 49504
rect 28288 49232 28636 49444
rect 110160 49232 110508 49444
rect 115192 49438 115404 49510
rect 115192 49374 115334 49438
rect 115398 49374 115404 49438
rect 115192 49368 115404 49374
rect 115600 49574 115812 49580
rect 115600 49510 115742 49574
rect 115806 49510 115812 49574
rect 115600 49438 115812 49510
rect 115600 49374 115742 49438
rect 115806 49374 115812 49438
rect 115600 49368 115812 49374
rect 116008 49574 116220 49580
rect 116008 49510 116014 49574
rect 116078 49510 116220 49574
rect 116008 49368 116220 49510
rect 116416 49438 116628 49580
rect 116416 49374 116422 49438
rect 116486 49374 116628 49438
rect 116416 49368 116628 49374
rect 116824 49574 117036 49580
rect 116824 49510 116966 49574
rect 117030 49510 117036 49574
rect 116824 49438 117036 49510
rect 116824 49374 116830 49438
rect 116894 49374 117036 49438
rect 116824 49368 117036 49374
rect 28288 49172 28364 49232
rect 110296 49172 110372 49232
rect 1224 49166 1980 49172
rect 1224 49102 1230 49166
rect 1294 49128 1980 49166
rect 1294 49102 1798 49128
rect 1224 49096 1798 49102
rect 1768 49072 1798 49096
rect 1854 49072 1980 49128
rect 1768 48960 1980 49072
rect 21760 49166 21972 49172
rect 21760 49102 21766 49166
rect 21830 49102 21972 49166
rect 21760 49030 21972 49102
rect 21760 48966 21902 49030
rect 21966 48966 21972 49030
rect 21760 48960 21972 48966
rect 22168 49036 22380 49172
rect 22576 49166 22788 49172
rect 22576 49102 22582 49166
rect 22646 49102 22788 49166
rect 22576 49036 22788 49102
rect 22168 49030 22788 49036
rect 22168 48966 22718 49030
rect 22782 48966 22788 49030
rect 22168 48960 22788 48966
rect 22984 49166 23196 49172
rect 22984 49102 22990 49166
rect 23054 49102 23196 49166
rect 22984 49030 23196 49102
rect 22984 48966 23126 49030
rect 23190 48966 23196 49030
rect 22984 48960 23196 48966
rect 23392 49166 23604 49172
rect 23392 49102 23534 49166
rect 23598 49102 23604 49166
rect 23392 49030 23604 49102
rect 23392 48966 23398 49030
rect 23462 48966 23604 49030
rect 23392 48960 23604 48966
rect 28288 48960 28636 49172
rect 110160 48960 110508 49172
rect 115192 49166 115404 49172
rect 115192 49102 115334 49166
rect 115398 49102 115404 49166
rect 115192 49030 115404 49102
rect 115192 48966 115198 49030
rect 115262 48966 115404 49030
rect 115192 48960 115404 48966
rect 115600 49166 115812 49172
rect 115600 49102 115742 49166
rect 115806 49102 115812 49166
rect 115600 49030 115812 49102
rect 115600 48966 115606 49030
rect 115670 48966 115812 49030
rect 115600 48960 115812 48966
rect 116008 49166 116628 49172
rect 116008 49102 116422 49166
rect 116486 49102 116628 49166
rect 116008 49096 116628 49102
rect 116008 48960 116220 49096
rect 116416 49030 116628 49096
rect 116416 48966 116558 49030
rect 116622 48966 116628 49030
rect 116416 48960 116628 48966
rect 116824 49166 117036 49172
rect 116824 49102 116830 49166
rect 116894 49102 117036 49166
rect 116824 49030 117036 49102
rect 116824 48966 116966 49030
rect 117030 48966 117036 49030
rect 116824 48960 117036 48966
rect 136816 49128 137028 49172
rect 136816 49072 136944 49128
rect 137000 49072 137028 49128
rect 136816 49036 137028 49072
rect 136816 49030 137572 49036
rect 136816 48966 137502 49030
rect 137566 48966 137572 49030
rect 136816 48960 137572 48966
rect 28424 48900 28500 48960
rect 110160 48900 110236 48960
rect 21760 48758 21972 48764
rect 21760 48694 21902 48758
rect 21966 48694 21972 48758
rect 21760 48552 21972 48694
rect 22168 48628 22380 48764
rect 22576 48758 22788 48764
rect 22576 48694 22718 48758
rect 22782 48694 22788 48758
rect 22576 48628 22788 48694
rect 22168 48622 22788 48628
rect 22168 48558 22310 48622
rect 22374 48558 22788 48622
rect 22168 48552 22788 48558
rect 22984 48758 23196 48764
rect 22984 48694 23126 48758
rect 23190 48694 23196 48758
rect 22984 48622 23196 48694
rect 22984 48558 23126 48622
rect 23190 48558 23196 48622
rect 22984 48552 23196 48558
rect 23392 48758 23604 48764
rect 23392 48694 23398 48758
rect 23462 48694 23604 48758
rect 23392 48622 23604 48694
rect 28288 48688 28636 48900
rect 28560 48628 28636 48688
rect 23392 48558 23398 48622
rect 23462 48558 23604 48622
rect 23392 48552 23604 48558
rect 21760 48492 21836 48552
rect 22304 48492 22380 48552
rect 21760 48350 21972 48492
rect 22304 48416 22652 48492
rect 22576 48356 22652 48416
rect 28288 48416 28636 48628
rect 110160 48688 110508 48900
rect 115192 48758 115404 48764
rect 115192 48694 115198 48758
rect 115262 48694 115404 48758
rect 110160 48628 110236 48688
rect 110160 48416 110508 48628
rect 115192 48622 115404 48694
rect 115192 48558 115334 48622
rect 115398 48558 115404 48622
rect 115192 48552 115404 48558
rect 115600 48758 115812 48764
rect 115600 48694 115606 48758
rect 115670 48694 115812 48758
rect 115600 48622 115812 48694
rect 115600 48558 115742 48622
rect 115806 48558 115812 48622
rect 115600 48552 115812 48558
rect 116008 48622 116220 48764
rect 116416 48758 116628 48764
rect 116416 48694 116558 48758
rect 116622 48694 116628 48758
rect 116416 48628 116628 48694
rect 116318 48622 116628 48628
rect 116008 48558 116150 48622
rect 116214 48558 116220 48622
rect 116280 48558 116286 48622
rect 116350 48558 116628 48622
rect 116008 48552 116220 48558
rect 116318 48552 116628 48558
rect 116824 48758 117036 48764
rect 116824 48694 116966 48758
rect 117030 48694 117036 48758
rect 116824 48552 117036 48694
rect 116824 48492 116900 48552
rect 28288 48356 28364 48416
rect 110296 48356 110372 48416
rect 21760 48286 21766 48350
rect 21830 48286 21972 48350
rect 21760 48280 21972 48286
rect 22168 48350 22380 48356
rect 22168 48286 22310 48350
rect 22374 48286 22380 48350
rect 22168 48144 22380 48286
rect 22304 48084 22380 48144
rect 21760 48078 21972 48084
rect 21760 48014 21766 48078
rect 21830 48014 21972 48078
rect 21760 47736 21972 48014
rect 22168 47736 22380 48084
rect 22576 48144 22788 48356
rect 22984 48350 23196 48356
rect 22984 48286 23126 48350
rect 23190 48286 23196 48350
rect 22984 48214 23196 48286
rect 22984 48150 22990 48214
rect 23054 48150 23196 48214
rect 22984 48144 23196 48150
rect 23392 48350 23604 48356
rect 23392 48286 23398 48350
rect 23462 48286 23604 48350
rect 23392 48214 23604 48286
rect 23392 48150 23398 48214
rect 23462 48150 23604 48214
rect 23392 48144 23604 48150
rect 22576 48084 22652 48144
rect 22576 47806 22788 48084
rect 22576 47742 22718 47806
rect 22782 47742 22788 47806
rect 22576 47736 22788 47742
rect 22984 47942 23196 47948
rect 22984 47878 22990 47942
rect 23054 47878 23196 47942
rect 22984 47736 23196 47878
rect 23392 47942 23604 47948
rect 23392 47878 23398 47942
rect 23462 47878 23604 47942
rect 23392 47736 23604 47878
rect 28288 47872 28636 48356
rect 110160 47872 110508 48356
rect 115192 48350 115404 48356
rect 115192 48286 115334 48350
rect 115398 48286 115404 48350
rect 115192 48214 115404 48286
rect 115192 48150 115198 48214
rect 115262 48150 115404 48214
rect 115192 48144 115404 48150
rect 115600 48350 115812 48356
rect 115600 48286 115742 48350
rect 115806 48286 115812 48350
rect 115600 48214 115812 48286
rect 115600 48150 115742 48214
rect 115806 48150 115812 48214
rect 115600 48144 115812 48150
rect 116008 48350 116356 48356
rect 116008 48286 116150 48350
rect 116214 48286 116286 48350
rect 116350 48286 116356 48350
rect 116008 48280 116356 48286
rect 116008 48220 116220 48280
rect 116416 48220 116628 48356
rect 116824 48350 117036 48492
rect 116824 48286 116830 48350
rect 116894 48286 117036 48350
rect 116824 48280 117036 48286
rect 116008 48214 116628 48220
rect 116008 48150 116150 48214
rect 116214 48150 116628 48214
rect 116008 48144 116628 48150
rect 116144 48084 116220 48144
rect 115192 47942 115404 47948
rect 115192 47878 115198 47942
rect 115262 47878 115404 47942
rect 28288 47812 28364 47872
rect 110160 47812 110236 47872
rect 21896 47676 21972 47736
rect 1768 47448 1980 47540
rect 21760 47534 21972 47676
rect 22984 47676 23060 47736
rect 23392 47676 23468 47736
rect 21760 47470 21766 47534
rect 21830 47470 21972 47534
rect 21760 47464 21972 47470
rect 1768 47404 1798 47448
rect 1224 47398 1798 47404
rect 1224 47334 1230 47398
rect 1294 47392 1798 47398
rect 1854 47392 1980 47448
rect 1294 47334 1980 47392
rect 1224 47328 1980 47334
rect 22168 47404 22380 47540
rect 22576 47534 22788 47540
rect 22576 47470 22718 47534
rect 22782 47470 22788 47534
rect 22168 47328 22516 47404
rect 22168 47268 22244 47328
rect 22440 47268 22516 47328
rect 22576 47328 22788 47470
rect 22984 47328 23196 47676
rect 23392 47328 23604 47676
rect 22576 47268 22652 47328
rect 23120 47268 23196 47328
rect 23528 47268 23604 47328
rect 21760 47262 21972 47268
rect 21760 47198 21766 47262
rect 21830 47198 21972 47262
rect 21760 47126 21972 47198
rect 21760 47062 21766 47126
rect 21830 47062 21972 47126
rect 21760 47056 21972 47062
rect 22168 47132 22380 47268
rect 22440 47192 22788 47268
rect 22168 47126 22516 47132
rect 22168 47062 22446 47126
rect 22510 47062 22516 47126
rect 22168 47056 22516 47062
rect 22576 47056 22788 47192
rect 22984 46920 23196 47268
rect 23392 46920 23604 47268
rect 28288 47262 28636 47812
rect 28288 47198 28294 47262
rect 28358 47198 28636 47262
rect 28288 47192 28636 47198
rect 110160 47670 110508 47812
rect 110160 47606 110166 47670
rect 110230 47606 110508 47670
rect 110160 47398 110508 47606
rect 110160 47334 110166 47398
rect 110230 47334 110508 47398
rect 110160 47262 110508 47334
rect 115192 47736 115404 47878
rect 115600 47942 115812 47948
rect 115600 47878 115742 47942
rect 115806 47878 115812 47942
rect 115600 47736 115812 47878
rect 116008 47736 116220 48084
rect 116318 48078 116628 48084
rect 116280 48014 116286 48078
rect 116350 48014 116628 48078
rect 116318 48008 116628 48014
rect 116416 47806 116628 48008
rect 116416 47742 116558 47806
rect 116622 47742 116628 47806
rect 116416 47736 116628 47742
rect 116824 48078 117036 48084
rect 116824 48014 116830 48078
rect 116894 48014 117036 48078
rect 116824 47736 117036 48014
rect 115192 47676 115268 47736
rect 115600 47676 115676 47736
rect 116824 47676 116900 47736
rect 115192 47328 115404 47676
rect 115600 47328 115812 47676
rect 115328 47268 115404 47328
rect 115736 47268 115812 47328
rect 110160 47198 110302 47262
rect 110366 47198 110508 47262
rect 110160 47192 110508 47198
rect 22984 46860 23060 46920
rect 23528 46860 23604 46920
rect 21760 46854 21972 46860
rect 21760 46790 21766 46854
rect 21830 46790 21972 46854
rect 21760 46718 21972 46790
rect 21760 46654 21902 46718
rect 21966 46654 21972 46718
rect 21760 46648 21972 46654
rect 22168 46724 22380 46860
rect 22478 46854 22788 46860
rect 22440 46790 22446 46854
rect 22510 46790 22788 46854
rect 22478 46784 22788 46790
rect 22576 46724 22788 46784
rect 22168 46648 22788 46724
rect 22984 46718 23196 46860
rect 22984 46654 22990 46718
rect 23054 46654 23196 46718
rect 22984 46648 23196 46654
rect 23392 46718 23604 46860
rect 23392 46654 23398 46718
rect 23462 46654 23604 46718
rect 23392 46648 23604 46654
rect 28288 46990 28636 46996
rect 28288 46926 28294 46990
rect 28358 46926 28636 46990
rect 28288 46648 28636 46926
rect 110160 46990 110508 46996
rect 110160 46926 110302 46990
rect 110366 46926 110508 46990
rect 110160 46854 110508 46926
rect 110160 46790 110438 46854
rect 110502 46790 110508 46854
rect 110160 46648 110508 46790
rect 115192 46920 115404 47268
rect 115600 46920 115812 47268
rect 116008 47328 116220 47540
rect 116416 47534 116628 47540
rect 116416 47470 116558 47534
rect 116622 47470 116628 47534
rect 116416 47328 116628 47470
rect 116824 47534 117036 47676
rect 116824 47470 116966 47534
rect 117030 47470 117036 47534
rect 116824 47464 117036 47470
rect 136816 47534 137572 47540
rect 136816 47470 137502 47534
rect 137566 47470 137572 47534
rect 136816 47464 137572 47470
rect 136816 47448 137028 47464
rect 136816 47392 136944 47448
rect 137000 47392 137028 47448
rect 136816 47328 137028 47392
rect 116008 47268 116084 47328
rect 116416 47268 116492 47328
rect 116008 47192 116628 47268
rect 116008 47132 116220 47192
rect 116008 47126 116356 47132
rect 116008 47062 116150 47126
rect 116214 47062 116286 47126
rect 116350 47062 116356 47126
rect 116008 47056 116356 47062
rect 116416 47056 116628 47192
rect 116824 47262 117036 47268
rect 116824 47198 116966 47262
rect 117030 47198 117036 47262
rect 116824 47126 117036 47198
rect 116824 47062 116830 47126
rect 116894 47062 117036 47126
rect 116824 47056 117036 47062
rect 115192 46860 115268 46920
rect 115600 46860 115676 46920
rect 115192 46718 115404 46860
rect 115192 46654 115198 46718
rect 115262 46654 115404 46718
rect 115192 46648 115404 46654
rect 115600 46718 115812 46860
rect 115600 46654 115606 46718
rect 115670 46654 115812 46718
rect 115600 46648 115812 46654
rect 116008 46854 116220 46860
rect 116318 46854 116628 46860
rect 116008 46790 116150 46854
rect 116214 46790 116220 46854
rect 116280 46790 116286 46854
rect 116350 46790 116628 46854
rect 22168 46512 22380 46648
rect 22576 46512 22788 46648
rect 28560 46588 28636 46648
rect 110432 46588 110508 46648
rect 22168 46452 22244 46512
rect 22712 46452 22788 46512
rect 21760 46446 21972 46452
rect 21760 46382 21902 46446
rect 21966 46382 21972 46446
rect 21760 46310 21972 46382
rect 21760 46246 21766 46310
rect 21830 46246 21972 46310
rect 21760 46240 21972 46246
rect 22168 46310 22380 46452
rect 22168 46246 22174 46310
rect 22238 46246 22380 46310
rect 22168 46240 22380 46246
rect 22576 46240 22788 46452
rect 22984 46446 23196 46452
rect 22984 46382 22990 46446
rect 23054 46382 23196 46446
rect 22984 46310 23196 46382
rect 22984 46246 23126 46310
rect 23190 46246 23196 46310
rect 22984 46240 23196 46246
rect 23392 46446 23604 46452
rect 23392 46382 23398 46446
rect 23462 46382 23604 46446
rect 23392 46310 23604 46382
rect 28288 46446 28636 46588
rect 28288 46382 28294 46446
rect 28358 46382 28636 46446
rect 28288 46376 28636 46382
rect 110160 46582 110508 46588
rect 110160 46518 110438 46582
rect 110502 46518 110508 46582
rect 110160 46376 110508 46518
rect 116008 46588 116220 46790
rect 116318 46784 116628 46790
rect 116008 46512 116356 46588
rect 116416 46512 116628 46784
rect 116824 46854 117036 46860
rect 116824 46790 116830 46854
rect 116894 46790 117036 46854
rect 116824 46718 117036 46790
rect 116824 46654 116830 46718
rect 116894 46654 117036 46718
rect 116824 46648 117036 46654
rect 116144 46452 116220 46512
rect 115192 46446 115404 46452
rect 115192 46382 115198 46446
rect 115262 46382 115404 46446
rect 28424 46316 28500 46376
rect 110160 46316 110236 46376
rect 23392 46246 23534 46310
rect 23598 46246 23604 46310
rect 23392 46240 23604 46246
rect 28288 46240 28636 46316
rect 110160 46240 110508 46316
rect 115192 46310 115404 46382
rect 115192 46246 115334 46310
rect 115398 46246 115404 46310
rect 115192 46240 115404 46246
rect 115600 46446 115812 46452
rect 115600 46382 115606 46446
rect 115670 46382 115812 46446
rect 115600 46310 115812 46382
rect 115600 46246 115742 46310
rect 115806 46246 115812 46310
rect 115600 46240 115812 46246
rect 116008 46310 116220 46452
rect 116280 46452 116356 46512
rect 116280 46376 116628 46452
rect 116008 46246 116014 46310
rect 116078 46246 116220 46310
rect 116008 46240 116220 46246
rect 116416 46240 116628 46376
rect 116824 46446 117036 46452
rect 116824 46382 116830 46446
rect 116894 46382 117036 46446
rect 116824 46310 117036 46382
rect 116824 46246 116830 46310
rect 116894 46246 117036 46310
rect 116824 46240 117036 46246
rect 28406 46044 28504 46240
rect 110294 46044 110392 46240
rect 21760 46038 21972 46044
rect 21760 45974 21766 46038
rect 21830 45974 21972 46038
rect 1768 45768 1980 45908
rect 21760 45902 21972 45974
rect 21760 45838 21902 45902
rect 21966 45838 21972 45902
rect 21760 45832 21972 45838
rect 22168 46038 22380 46044
rect 22168 45974 22174 46038
rect 22238 45974 22380 46038
rect 22168 45902 22380 45974
rect 22168 45838 22310 45902
rect 22374 45838 22380 45902
rect 22168 45832 22380 45838
rect 22576 45832 22788 46044
rect 22984 46038 23196 46044
rect 22984 45974 23126 46038
rect 23190 45974 23196 46038
rect 22984 45902 23196 45974
rect 22984 45838 23126 45902
rect 23190 45838 23196 45902
rect 22984 45832 23196 45838
rect 23392 46038 23604 46044
rect 23392 45974 23534 46038
rect 23598 45974 23604 46038
rect 23392 45902 23604 45974
rect 23392 45838 23398 45902
rect 23462 45838 23604 45902
rect 23392 45832 23604 45838
rect 28288 46038 28636 46044
rect 28288 45974 28294 46038
rect 28358 45974 28636 46038
rect 28288 45832 28636 45974
rect 110160 45832 110508 46044
rect 115192 46038 115404 46044
rect 115192 45974 115334 46038
rect 115398 45974 115404 46038
rect 115192 45902 115404 45974
rect 115192 45838 115198 45902
rect 115262 45838 115404 45902
rect 115192 45832 115404 45838
rect 115600 46038 115812 46044
rect 115600 45974 115742 46038
rect 115806 45974 115812 46038
rect 115600 45902 115812 45974
rect 115600 45838 115606 45902
rect 115670 45838 115812 45902
rect 115600 45832 115812 45838
rect 116008 46038 116220 46044
rect 116008 45974 116014 46038
rect 116078 45974 116220 46038
rect 116008 45908 116220 45974
rect 116008 45832 116356 45908
rect 116416 45902 116628 46044
rect 116416 45838 116422 45902
rect 116486 45838 116628 45902
rect 116416 45832 116628 45838
rect 116824 46038 117036 46044
rect 116824 45974 116830 46038
rect 116894 45974 117036 46038
rect 116824 45902 117036 45974
rect 116824 45838 116966 45902
rect 117030 45838 117036 45902
rect 116824 45832 117036 45838
rect 22576 45772 22652 45832
rect 1768 45712 1798 45768
rect 1854 45712 1980 45768
rect 1768 45636 1980 45712
rect 22304 45696 22652 45772
rect 28288 45772 28364 45832
rect 110296 45772 110372 45832
rect 116280 45772 116356 45832
rect 22304 45636 22380 45696
rect 1224 45630 1980 45636
rect 1224 45566 1230 45630
rect 1294 45566 1980 45630
rect 1224 45560 1980 45566
rect 21760 45630 21972 45636
rect 21760 45566 21902 45630
rect 21966 45566 21972 45630
rect 21760 45494 21972 45566
rect 21760 45430 21902 45494
rect 21966 45430 21972 45494
rect 21760 45424 21972 45430
rect 22168 45630 22788 45636
rect 22168 45566 22310 45630
rect 22374 45566 22788 45630
rect 22168 45560 22788 45566
rect 22168 45424 22380 45560
rect 22576 45494 22788 45560
rect 22576 45430 22582 45494
rect 22646 45430 22788 45494
rect 22576 45424 22788 45430
rect 22984 45630 23196 45636
rect 22984 45566 23126 45630
rect 23190 45566 23196 45630
rect 22984 45494 23196 45566
rect 22984 45430 22990 45494
rect 23054 45430 23196 45494
rect 22984 45424 23196 45430
rect 23392 45630 23604 45636
rect 23392 45566 23398 45630
rect 23462 45566 23604 45630
rect 23392 45494 23604 45566
rect 28288 45560 28636 45772
rect 110160 45560 110508 45772
rect 116280 45696 116492 45772
rect 116416 45636 116492 45696
rect 136816 45768 137028 45908
rect 136816 45712 136944 45768
rect 137000 45712 137028 45768
rect 136816 45636 137028 45712
rect 115192 45630 115404 45636
rect 115192 45566 115198 45630
rect 115262 45566 115404 45630
rect 28424 45500 28500 45560
rect 110160 45500 110236 45560
rect 23392 45430 23398 45494
rect 23462 45430 23604 45494
rect 23392 45424 23604 45430
rect 28288 45288 28636 45500
rect 110160 45288 110508 45500
rect 115192 45494 115404 45566
rect 115192 45430 115334 45494
rect 115398 45430 115404 45494
rect 115192 45424 115404 45430
rect 115600 45630 115812 45636
rect 115600 45566 115606 45630
rect 115670 45566 115812 45630
rect 115600 45494 115812 45566
rect 115600 45430 115742 45494
rect 115806 45430 115812 45494
rect 115600 45424 115812 45430
rect 116008 45630 116628 45636
rect 116008 45566 116422 45630
rect 116486 45566 116628 45630
rect 116008 45560 116628 45566
rect 116008 45500 116220 45560
rect 116008 45494 116356 45500
rect 116008 45430 116150 45494
rect 116214 45430 116286 45494
rect 116350 45430 116356 45494
rect 116008 45424 116356 45430
rect 116416 45424 116628 45560
rect 116824 45630 117036 45636
rect 116824 45566 116966 45630
rect 117030 45566 117036 45630
rect 116824 45494 117036 45566
rect 136816 45630 137572 45636
rect 136816 45566 137502 45630
rect 137566 45566 137572 45630
rect 136816 45560 137572 45566
rect 116824 45430 116966 45494
rect 117030 45430 117036 45494
rect 116824 45424 117036 45430
rect 28288 45228 28364 45288
rect 110432 45228 110508 45288
rect 21760 45222 21972 45228
rect 21760 45158 21902 45222
rect 21966 45158 21972 45222
rect 21760 45086 21972 45158
rect 21760 45022 21766 45086
rect 21830 45022 21972 45086
rect 21760 45016 21972 45022
rect 22168 45086 22380 45228
rect 22168 45022 22174 45086
rect 22238 45022 22380 45086
rect 22168 45016 22380 45022
rect 22576 45222 22788 45228
rect 22576 45158 22582 45222
rect 22646 45158 22788 45222
rect 22576 45086 22788 45158
rect 22576 45022 22582 45086
rect 22646 45022 22788 45086
rect 22576 45016 22788 45022
rect 22984 45222 23196 45228
rect 22984 45158 22990 45222
rect 23054 45158 23196 45222
rect 22984 45086 23196 45158
rect 22984 45022 22990 45086
rect 23054 45022 23196 45086
rect 22984 45016 23196 45022
rect 23392 45222 23604 45228
rect 23392 45158 23398 45222
rect 23462 45158 23604 45222
rect 23392 45086 23604 45158
rect 23392 45022 23534 45086
rect 23598 45022 23604 45086
rect 23392 45016 23604 45022
rect 28288 45016 28636 45228
rect 110160 45016 110508 45228
rect 115192 45222 115404 45228
rect 115192 45158 115334 45222
rect 115398 45158 115404 45222
rect 115192 45086 115404 45158
rect 115192 45022 115334 45086
rect 115398 45022 115404 45086
rect 115192 45016 115404 45022
rect 115600 45222 115812 45228
rect 115600 45158 115742 45222
rect 115806 45158 115812 45222
rect 115600 45086 115812 45158
rect 115600 45022 115742 45086
rect 115806 45022 115812 45086
rect 115600 45016 115812 45022
rect 116008 45222 116220 45228
rect 116318 45222 116628 45228
rect 116008 45158 116150 45222
rect 116214 45158 116220 45222
rect 116280 45158 116286 45222
rect 116350 45158 116628 45222
rect 116008 45016 116220 45158
rect 116318 45152 116628 45158
rect 116416 45086 116628 45152
rect 116416 45022 116422 45086
rect 116486 45022 116628 45086
rect 116416 45016 116628 45022
rect 116824 45222 117036 45228
rect 116824 45158 116966 45222
rect 117030 45158 117036 45222
rect 116824 45086 117036 45158
rect 116824 45022 116830 45086
rect 116894 45022 117036 45086
rect 116824 45016 117036 45022
rect 28288 44956 28364 45016
rect 110432 44956 110508 45016
rect 21760 44814 21972 44820
rect 21760 44750 21766 44814
rect 21830 44750 21972 44814
rect 21760 44608 21972 44750
rect 22168 44814 22380 44820
rect 22168 44750 22174 44814
rect 22238 44750 22380 44814
rect 22168 44678 22380 44750
rect 22168 44614 22310 44678
rect 22374 44614 22380 44678
rect 22168 44608 22380 44614
rect 22576 44814 22788 44820
rect 22576 44750 22582 44814
rect 22646 44750 22788 44814
rect 22576 44678 22788 44750
rect 22576 44614 22718 44678
rect 22782 44614 22788 44678
rect 22576 44608 22788 44614
rect 22984 44814 23196 44820
rect 22984 44750 22990 44814
rect 23054 44750 23196 44814
rect 22984 44678 23196 44750
rect 22984 44614 23126 44678
rect 23190 44614 23196 44678
rect 22984 44608 23196 44614
rect 23392 44814 23604 44820
rect 23392 44750 23534 44814
rect 23598 44750 23604 44814
rect 23392 44678 23604 44750
rect 28288 44744 28636 44956
rect 110160 44744 110508 44956
rect 28424 44684 28500 44744
rect 110432 44684 110508 44744
rect 23392 44614 23398 44678
rect 23462 44614 23604 44678
rect 23392 44608 23604 44614
rect 21760 44548 21836 44608
rect 21760 44200 21972 44548
rect 28288 44472 28636 44684
rect 28560 44412 28636 44472
rect 22168 44406 22788 44412
rect 22168 44342 22310 44406
rect 22374 44342 22718 44406
rect 22782 44342 22788 44406
rect 22168 44336 22788 44342
rect 22168 44276 22380 44336
rect 22168 44200 22516 44276
rect 22576 44200 22788 44336
rect 22984 44406 23196 44412
rect 22984 44342 23126 44406
rect 23190 44342 23196 44406
rect 22984 44270 23196 44342
rect 22984 44206 22990 44270
rect 23054 44206 23196 44270
rect 22984 44200 23196 44206
rect 23392 44406 23604 44412
rect 23392 44342 23398 44406
rect 23462 44342 23604 44406
rect 23392 44270 23604 44342
rect 23392 44206 23398 44270
rect 23462 44206 23604 44270
rect 23392 44200 23604 44206
rect 21896 44140 21972 44200
rect 22440 44140 22516 44200
rect 1224 44134 1980 44140
rect 1224 44070 1230 44134
rect 1294 44088 1980 44134
rect 1294 44070 1798 44088
rect 1224 44064 1798 44070
rect 1768 44032 1798 44064
rect 1854 44032 1980 44088
rect 1768 43928 1980 44032
rect 21760 43792 21972 44140
rect 22168 43862 22380 44140
rect 22440 44064 22788 44140
rect 22168 43798 22174 43862
rect 22238 43798 22380 43862
rect 22168 43792 22380 43798
rect 22576 43862 22788 44064
rect 22576 43798 22582 43862
rect 22646 43798 22788 43862
rect 22576 43792 22788 43798
rect 22984 43998 23196 44004
rect 22984 43934 22990 43998
rect 23054 43934 23196 43998
rect 22984 43862 23196 43934
rect 22984 43798 22990 43862
rect 23054 43798 23196 43862
rect 22984 43792 23196 43798
rect 23392 43998 23604 44004
rect 23392 43934 23398 43998
rect 23462 43934 23604 43998
rect 23392 43862 23604 43934
rect 23392 43798 23398 43862
rect 23462 43798 23604 43862
rect 23392 43792 23604 43798
rect 28288 43928 28636 44412
rect 110160 44542 110508 44684
rect 115192 44814 115404 44820
rect 115192 44750 115334 44814
rect 115398 44750 115404 44814
rect 115192 44678 115404 44750
rect 115192 44614 115198 44678
rect 115262 44614 115404 44678
rect 115192 44608 115404 44614
rect 115600 44814 115812 44820
rect 115600 44750 115742 44814
rect 115806 44750 115812 44814
rect 115600 44678 115812 44750
rect 115600 44614 115606 44678
rect 115670 44614 115812 44678
rect 115600 44608 115812 44614
rect 116008 44814 116628 44820
rect 116008 44750 116422 44814
rect 116486 44750 116628 44814
rect 116008 44744 116628 44750
rect 116008 44608 116220 44744
rect 116416 44678 116628 44744
rect 116416 44614 116558 44678
rect 116622 44614 116628 44678
rect 116416 44608 116628 44614
rect 116824 44814 117036 44820
rect 116824 44750 116830 44814
rect 116894 44750 117036 44814
rect 116824 44608 117036 44750
rect 110160 44478 110166 44542
rect 110230 44478 110508 44542
rect 110160 44472 110508 44478
rect 116824 44548 116900 44608
rect 110160 44412 110236 44472
rect 110160 44270 110508 44412
rect 110160 44206 110166 44270
rect 110230 44206 110508 44270
rect 110160 43928 110508 44206
rect 115192 44406 115404 44412
rect 115192 44342 115198 44406
rect 115262 44342 115404 44406
rect 115192 44270 115404 44342
rect 115192 44206 115198 44270
rect 115262 44206 115404 44270
rect 115192 44200 115404 44206
rect 115600 44406 115812 44412
rect 115600 44342 115606 44406
rect 115670 44342 115812 44406
rect 115600 44270 115812 44342
rect 115600 44206 115606 44270
rect 115670 44206 115812 44270
rect 115600 44200 115812 44206
rect 116008 44406 116356 44412
rect 116008 44342 116286 44406
rect 116350 44342 116356 44406
rect 116008 44336 116356 44342
rect 116416 44406 116628 44412
rect 116416 44342 116558 44406
rect 116622 44342 116628 44406
rect 116008 44276 116220 44336
rect 116416 44276 116628 44342
rect 116008 44200 116628 44276
rect 116824 44200 117036 44548
rect 116144 44140 116220 44200
rect 116960 44140 117036 44200
rect 28288 43868 28364 43928
rect 110432 43868 110508 43928
rect 21760 43732 21836 43792
rect 21760 43590 21972 43732
rect 28288 43656 28636 43868
rect 110160 43726 110508 43868
rect 115192 43998 115404 44004
rect 115192 43934 115198 43998
rect 115262 43934 115404 43998
rect 115192 43862 115404 43934
rect 115192 43798 115198 43862
rect 115262 43798 115404 43862
rect 115192 43792 115404 43798
rect 115600 43998 115812 44004
rect 115600 43934 115606 43998
rect 115670 43934 115812 43998
rect 115600 43862 115812 43934
rect 115600 43798 115606 43862
rect 115670 43798 115812 43862
rect 115600 43792 115812 43798
rect 116008 43862 116220 44140
rect 116318 44134 116628 44140
rect 116280 44070 116286 44134
rect 116350 44070 116628 44134
rect 116318 44064 116628 44070
rect 116008 43798 116014 43862
rect 116078 43798 116220 43862
rect 116008 43792 116220 43798
rect 116416 43862 116628 44064
rect 116416 43798 116558 43862
rect 116622 43798 116628 43862
rect 116416 43792 116628 43798
rect 116824 43792 117036 44140
rect 136816 44134 137572 44140
rect 136816 44088 137502 44134
rect 136816 44032 136944 44088
rect 137000 44070 137502 44088
rect 137566 44070 137572 44134
rect 137000 44064 137572 44070
rect 137000 44032 137028 44064
rect 136816 43928 137028 44032
rect 110160 43662 110438 43726
rect 110502 43662 110508 43726
rect 110160 43656 110508 43662
rect 116824 43732 116900 43792
rect 28424 43596 28500 43656
rect 110160 43596 110236 43656
rect 21760 43526 21902 43590
rect 21966 43526 21972 43590
rect 21760 43520 21972 43526
rect 22168 43590 22516 43596
rect 22168 43526 22174 43590
rect 22238 43526 22446 43590
rect 22510 43526 22516 43590
rect 22168 43520 22516 43526
rect 22576 43590 22788 43596
rect 22576 43526 22582 43590
rect 22646 43526 22788 43590
rect 22168 43384 22380 43520
rect 22576 43460 22788 43526
rect 22440 43384 22788 43460
rect 22440 43324 22516 43384
rect 22712 43324 22788 43384
rect 21760 43318 21972 43324
rect 21760 43254 21902 43318
rect 21966 43254 21972 43318
rect 21760 43182 21972 43254
rect 21760 43118 21766 43182
rect 21830 43118 21972 43182
rect 21760 43112 21972 43118
rect 22168 43248 22516 43324
rect 22576 43318 22788 43324
rect 22576 43254 22582 43318
rect 22646 43254 22788 43318
rect 22168 43188 22380 43248
rect 22168 43182 22516 43188
rect 22168 43118 22446 43182
rect 22510 43118 22516 43182
rect 22168 43112 22516 43118
rect 22576 43112 22788 43254
rect 22984 43590 23196 43596
rect 22984 43526 22990 43590
rect 23054 43526 23196 43590
rect 22984 43384 23196 43526
rect 23392 43590 23604 43596
rect 23392 43526 23398 43590
rect 23462 43526 23604 43590
rect 23392 43384 23604 43526
rect 22984 43324 23060 43384
rect 23392 43324 23468 43384
rect 22984 42976 23196 43324
rect 23392 42976 23604 43324
rect 28288 43318 28636 43596
rect 28288 43254 28294 43318
rect 28358 43254 28636 43318
rect 28288 43248 28636 43254
rect 110160 43454 110508 43596
rect 110160 43390 110438 43454
rect 110502 43390 110508 43454
rect 110160 43318 110508 43390
rect 110160 43254 110166 43318
rect 110230 43254 110508 43318
rect 110160 43248 110508 43254
rect 115192 43590 115404 43596
rect 115192 43526 115198 43590
rect 115262 43526 115404 43590
rect 115192 43384 115404 43526
rect 115600 43590 115812 43596
rect 115600 43526 115606 43590
rect 115670 43526 115812 43590
rect 115600 43384 115812 43526
rect 116008 43590 116220 43596
rect 116008 43526 116014 43590
rect 116078 43526 116220 43590
rect 116008 43384 116220 43526
rect 116416 43590 116628 43596
rect 116416 43526 116558 43590
rect 116622 43526 116628 43590
rect 116416 43384 116628 43526
rect 116824 43590 117036 43732
rect 116824 43526 116966 43590
rect 117030 43526 117036 43590
rect 116824 43520 117036 43526
rect 115192 43324 115268 43384
rect 115600 43324 115676 43384
rect 116144 43324 116220 43384
rect 116552 43324 116628 43384
rect 23120 42916 23196 42976
rect 23528 42916 23604 42976
rect 21760 42910 21972 42916
rect 21760 42846 21766 42910
rect 21830 42846 21972 42910
rect 21760 42774 21972 42846
rect 21760 42710 21766 42774
rect 21830 42710 21972 42774
rect 21760 42704 21972 42710
rect 22168 42568 22380 42916
rect 22478 42910 22788 42916
rect 22440 42846 22446 42910
rect 22510 42846 22788 42910
rect 22478 42840 22788 42846
rect 22576 42568 22788 42840
rect 22984 42774 23196 42916
rect 22984 42710 23126 42774
rect 23190 42710 23196 42774
rect 22984 42704 23196 42710
rect 23392 42774 23604 42916
rect 23392 42710 23398 42774
rect 23462 42710 23604 42774
rect 23392 42704 23604 42710
rect 28288 43046 28636 43052
rect 28288 42982 28294 43046
rect 28358 42982 28636 43046
rect 28288 42910 28636 42982
rect 28288 42846 28294 42910
rect 28358 42846 28636 42910
rect 28288 42704 28636 42846
rect 110160 43046 110508 43052
rect 110160 42982 110166 43046
rect 110230 42982 110508 43046
rect 110160 42704 110508 42982
rect 115192 42976 115404 43324
rect 115600 42976 115812 43324
rect 116008 43188 116220 43324
rect 116008 43112 116356 43188
rect 116416 43112 116628 43324
rect 116824 43318 117036 43324
rect 116824 43254 116966 43318
rect 117030 43254 117036 43318
rect 116824 43182 117036 43254
rect 116824 43118 116966 43182
rect 117030 43118 117036 43182
rect 116824 43112 117036 43118
rect 116280 43052 116356 43112
rect 116280 42976 116492 43052
rect 115328 42916 115404 42976
rect 115736 42916 115812 42976
rect 116416 42916 116492 42976
rect 115192 42774 115404 42916
rect 115192 42710 115334 42774
rect 115398 42710 115404 42774
rect 115192 42704 115404 42710
rect 115600 42774 115812 42916
rect 115600 42710 115606 42774
rect 115670 42710 115812 42774
rect 115600 42704 115812 42710
rect 116008 42840 116628 42916
rect 28424 42644 28500 42704
rect 110296 42644 110372 42704
rect 22304 42508 22380 42568
rect 22712 42508 22788 42568
rect 28288 42638 28636 42644
rect 28288 42574 28294 42638
rect 28358 42574 28636 42638
rect 1224 42502 1980 42508
rect 1224 42438 1230 42502
rect 1294 42438 1980 42502
rect 1224 42432 1980 42438
rect 1768 42408 1980 42432
rect 1768 42352 1798 42408
rect 1854 42352 1980 42408
rect 1768 42296 1980 42352
rect 21760 42502 21972 42508
rect 21760 42438 21766 42502
rect 21830 42438 21972 42502
rect 21760 42366 21972 42438
rect 21760 42302 21902 42366
rect 21966 42302 21972 42366
rect 21760 42296 21972 42302
rect 22168 42372 22380 42508
rect 22576 42372 22788 42508
rect 22168 42296 22788 42372
rect 22984 42502 23196 42508
rect 22984 42438 23126 42502
rect 23190 42438 23196 42502
rect 22984 42366 23196 42438
rect 22984 42302 23126 42366
rect 23190 42302 23196 42366
rect 22984 42296 23196 42302
rect 23392 42502 23604 42508
rect 23392 42438 23398 42502
rect 23462 42438 23604 42502
rect 23392 42366 23604 42438
rect 28288 42432 28636 42574
rect 110160 42432 110508 42644
rect 116008 42568 116220 42840
rect 116416 42568 116628 42840
rect 116824 42910 117036 42916
rect 116824 42846 116966 42910
rect 117030 42846 117036 42910
rect 116824 42774 117036 42846
rect 116824 42710 116966 42774
rect 117030 42710 117036 42774
rect 116824 42704 117036 42710
rect 116144 42508 116220 42568
rect 116552 42508 116628 42568
rect 115192 42502 115404 42508
rect 115192 42438 115334 42502
rect 115398 42438 115404 42502
rect 28560 42372 28636 42432
rect 110296 42372 110372 42432
rect 23392 42302 23398 42366
rect 23462 42302 23604 42366
rect 23392 42296 23604 42302
rect 22304 42236 22380 42296
rect 22304 42160 22652 42236
rect 22576 42100 22652 42160
rect 21760 42094 21972 42100
rect 21760 42030 21902 42094
rect 21966 42030 21972 42094
rect 21760 41958 21972 42030
rect 21760 41894 21766 41958
rect 21830 41894 21972 41958
rect 21760 41888 21972 41894
rect 22168 42024 22788 42100
rect 22168 41964 22380 42024
rect 22168 41958 22516 41964
rect 22168 41894 22174 41958
rect 22238 41894 22446 41958
rect 22510 41894 22516 41958
rect 22168 41888 22516 41894
rect 22576 41888 22788 42024
rect 22984 42094 23196 42100
rect 22984 42030 23126 42094
rect 23190 42030 23196 42094
rect 22984 41958 23196 42030
rect 22984 41894 23126 41958
rect 23190 41894 23196 41958
rect 22984 41888 23196 41894
rect 23392 42094 23604 42100
rect 23392 42030 23398 42094
rect 23462 42030 23604 42094
rect 23392 41958 23604 42030
rect 23392 41894 23534 41958
rect 23598 41894 23604 41958
rect 23392 41888 23604 41894
rect 28288 41888 28636 42372
rect 110160 42094 110508 42372
rect 115192 42366 115404 42438
rect 115192 42302 115198 42366
rect 115262 42302 115404 42366
rect 115192 42296 115404 42302
rect 115600 42502 115812 42508
rect 115600 42438 115606 42502
rect 115670 42438 115812 42502
rect 115600 42366 115812 42438
rect 115600 42302 115606 42366
rect 115670 42302 115812 42366
rect 115600 42296 115812 42302
rect 116008 42366 116220 42508
rect 116008 42302 116150 42366
rect 116214 42302 116220 42366
rect 116008 42296 116220 42302
rect 116416 42296 116628 42508
rect 116824 42502 117036 42508
rect 116824 42438 116966 42502
rect 117030 42438 117036 42502
rect 116824 42366 117036 42438
rect 116824 42302 116966 42366
rect 117030 42302 117036 42366
rect 116824 42296 117036 42302
rect 136816 42502 137572 42508
rect 136816 42438 137502 42502
rect 137566 42438 137572 42502
rect 136816 42432 137572 42438
rect 136816 42408 137028 42432
rect 136816 42352 136944 42408
rect 137000 42352 137028 42408
rect 136816 42296 137028 42352
rect 110160 42030 110438 42094
rect 110502 42030 110508 42094
rect 110160 41888 110508 42030
rect 115192 42094 115404 42100
rect 115192 42030 115198 42094
rect 115262 42030 115404 42094
rect 115192 41958 115404 42030
rect 115192 41894 115334 41958
rect 115398 41894 115404 41958
rect 115192 41888 115404 41894
rect 115600 42094 115812 42100
rect 115600 42030 115606 42094
rect 115670 42030 115812 42094
rect 115600 41958 115812 42030
rect 115600 41894 115742 41958
rect 115806 41894 115812 41958
rect 115600 41888 115812 41894
rect 116008 42094 116220 42100
rect 116008 42030 116150 42094
rect 116214 42030 116220 42094
rect 116008 41958 116220 42030
rect 116008 41894 116014 41958
rect 116078 41894 116220 41958
rect 116008 41888 116220 41894
rect 116416 41958 116628 42100
rect 116416 41894 116422 41958
rect 116486 41894 116628 41958
rect 116416 41888 116628 41894
rect 116824 42094 117036 42100
rect 116824 42030 116966 42094
rect 117030 42030 117036 42094
rect 116824 41958 117036 42030
rect 116824 41894 116830 41958
rect 116894 41894 117036 41958
rect 116824 41888 117036 41894
rect 28424 41828 28500 41888
rect 110432 41828 110508 41888
rect 21760 41686 21972 41692
rect 21760 41622 21766 41686
rect 21830 41622 21972 41686
rect 21760 41550 21972 41622
rect 21760 41486 21766 41550
rect 21830 41486 21972 41550
rect 21760 41480 21972 41486
rect 22168 41686 22380 41692
rect 22478 41686 22788 41692
rect 22168 41622 22174 41686
rect 22238 41622 22380 41686
rect 22440 41622 22446 41686
rect 22510 41622 22788 41686
rect 22168 41480 22380 41622
rect 22478 41616 22788 41622
rect 22576 41480 22788 41616
rect 22984 41686 23196 41692
rect 22984 41622 23126 41686
rect 23190 41622 23196 41686
rect 22984 41550 23196 41622
rect 22984 41486 23126 41550
rect 23190 41486 23196 41550
rect 22984 41480 23196 41486
rect 23392 41686 23604 41692
rect 23392 41622 23534 41686
rect 23598 41622 23604 41686
rect 23392 41550 23604 41622
rect 23392 41486 23398 41550
rect 23462 41486 23604 41550
rect 23392 41480 23604 41486
rect 28288 41616 28636 41828
rect 110160 41822 110508 41828
rect 110160 41758 110438 41822
rect 110502 41758 110508 41822
rect 110160 41616 110508 41758
rect 115192 41686 115404 41692
rect 115192 41622 115334 41686
rect 115398 41622 115404 41686
rect 28288 41556 28364 41616
rect 110296 41556 110372 41616
rect 22576 41420 22652 41480
rect 22304 41344 22652 41420
rect 28288 41344 28636 41556
rect 110160 41344 110508 41556
rect 115192 41550 115404 41622
rect 115192 41486 115198 41550
rect 115262 41486 115404 41550
rect 115192 41480 115404 41486
rect 115600 41686 115812 41692
rect 115600 41622 115742 41686
rect 115806 41622 115812 41686
rect 115600 41550 115812 41622
rect 115600 41486 115606 41550
rect 115670 41486 115812 41550
rect 115600 41480 115812 41486
rect 116008 41686 116220 41692
rect 116008 41622 116014 41686
rect 116078 41622 116220 41686
rect 116008 41550 116220 41622
rect 116416 41686 116628 41692
rect 116416 41622 116422 41686
rect 116486 41622 116628 41686
rect 116416 41556 116628 41622
rect 116318 41550 116628 41556
rect 116008 41486 116014 41550
rect 116078 41486 116220 41550
rect 116280 41486 116286 41550
rect 116350 41486 116558 41550
rect 116622 41486 116628 41550
rect 116008 41480 116220 41486
rect 116318 41480 116628 41486
rect 116824 41686 117036 41692
rect 116824 41622 116830 41686
rect 116894 41622 117036 41686
rect 116824 41550 117036 41622
rect 116824 41486 116966 41550
rect 117030 41486 117036 41550
rect 116824 41480 117036 41486
rect 22304 41284 22380 41344
rect 28560 41284 28636 41344
rect 110432 41284 110508 41344
rect 21760 41278 21972 41284
rect 21760 41214 21766 41278
rect 21830 41214 21972 41278
rect 21760 41142 21972 41214
rect 21760 41078 21766 41142
rect 21830 41078 21972 41142
rect 21760 41072 21972 41078
rect 22168 41208 22788 41284
rect 22168 41142 22380 41208
rect 22168 41078 22174 41142
rect 22238 41078 22380 41142
rect 22168 41072 22380 41078
rect 22576 41142 22788 41208
rect 22576 41078 22718 41142
rect 22782 41078 22788 41142
rect 22576 41072 22788 41078
rect 22984 41278 23196 41284
rect 22984 41214 23126 41278
rect 23190 41214 23196 41278
rect 22984 41142 23196 41214
rect 22984 41078 22990 41142
rect 23054 41078 23196 41142
rect 22984 41072 23196 41078
rect 23392 41278 23604 41284
rect 23392 41214 23398 41278
rect 23462 41214 23604 41278
rect 23392 41142 23604 41214
rect 23392 41078 23534 41142
rect 23598 41078 23604 41142
rect 23392 41072 23604 41078
rect 28288 41072 28636 41284
rect 110160 41072 110508 41284
rect 115192 41278 115404 41284
rect 115192 41214 115198 41278
rect 115262 41214 115404 41278
rect 115192 41142 115404 41214
rect 115192 41078 115198 41142
rect 115262 41078 115404 41142
rect 115192 41072 115404 41078
rect 115600 41278 115812 41284
rect 115600 41214 115606 41278
rect 115670 41214 115812 41278
rect 115600 41142 115812 41214
rect 115600 41078 115742 41142
rect 115806 41078 115812 41142
rect 115600 41072 115812 41078
rect 116008 41278 116356 41284
rect 116008 41214 116014 41278
rect 116078 41214 116286 41278
rect 116350 41214 116356 41278
rect 116008 41208 116356 41214
rect 116416 41278 116628 41284
rect 116416 41214 116558 41278
rect 116622 41214 116628 41278
rect 116008 41142 116220 41208
rect 116008 41078 116014 41142
rect 116078 41078 116220 41142
rect 116008 41072 116220 41078
rect 116416 41072 116628 41214
rect 116824 41278 117036 41284
rect 116824 41214 116966 41278
rect 117030 41214 117036 41278
rect 116824 41142 117036 41214
rect 116824 41078 116966 41142
rect 117030 41078 117036 41142
rect 116824 41072 117036 41078
rect 28424 41012 28500 41072
rect 110432 41012 110508 41072
rect 1768 40740 1980 40876
rect 21760 40870 21972 40876
rect 21760 40806 21766 40870
rect 21830 40806 21972 40870
rect 1224 40734 1980 40740
rect 1224 40670 1230 40734
rect 1294 40728 1980 40734
rect 1294 40672 1798 40728
rect 1854 40672 1980 40728
rect 1294 40670 1980 40672
rect 1224 40664 1980 40670
rect 1768 40528 1980 40664
rect 14552 40598 14764 40740
rect 21760 40664 21972 40806
rect 22168 40870 22380 40876
rect 22168 40806 22174 40870
rect 22238 40806 22380 40870
rect 22168 40664 22380 40806
rect 22576 40870 22788 40876
rect 22576 40806 22718 40870
rect 22782 40806 22788 40870
rect 22576 40734 22788 40806
rect 22576 40670 22582 40734
rect 22646 40670 22788 40734
rect 22576 40664 22788 40670
rect 22984 40870 23196 40876
rect 22984 40806 22990 40870
rect 23054 40806 23196 40870
rect 22984 40734 23196 40806
rect 22984 40670 23126 40734
rect 23190 40670 23196 40734
rect 22984 40664 23196 40670
rect 23392 40870 23604 40876
rect 23392 40806 23534 40870
rect 23598 40806 23604 40870
rect 23392 40734 23604 40806
rect 28288 40800 28636 41012
rect 110160 40800 110508 41012
rect 28424 40740 28500 40800
rect 110432 40740 110508 40800
rect 23392 40670 23534 40734
rect 23598 40670 23604 40734
rect 23392 40664 23604 40670
rect 21896 40604 21972 40664
rect 14552 40534 14694 40598
rect 14758 40534 14764 40598
rect 14552 40528 14764 40534
rect 21760 40256 21972 40604
rect 28288 40528 28636 40740
rect 28560 40468 28636 40528
rect 22168 40256 22380 40468
rect 22576 40462 22788 40468
rect 22576 40398 22582 40462
rect 22646 40398 22788 40462
rect 22576 40332 22788 40398
rect 21760 40196 21836 40256
rect 22304 40196 22380 40256
rect 22440 40256 22788 40332
rect 22984 40462 23196 40468
rect 22984 40398 23126 40462
rect 23190 40398 23196 40462
rect 22984 40326 23196 40398
rect 22984 40262 22990 40326
rect 23054 40262 23196 40326
rect 22984 40256 23196 40262
rect 23392 40462 23604 40468
rect 23392 40398 23534 40462
rect 23598 40398 23604 40462
rect 23392 40326 23604 40398
rect 23392 40262 23398 40326
rect 23462 40262 23604 40326
rect 23392 40256 23604 40262
rect 22440 40196 22516 40256
rect 0 40120 14356 40196
rect 14144 40102 14356 40120
rect 14144 40046 14212 40102
rect 14268 40046 14356 40102
rect 14144 39984 14356 40046
rect 15152 40033 15218 40036
rect 15966 40033 16032 40036
rect 15152 40031 16032 40033
rect 15152 39975 15157 40031
rect 15213 39975 15971 40031
rect 16027 39975 16032 40031
rect 15152 39973 16032 39975
rect 15152 39970 15218 39973
rect 15966 39970 16032 39973
rect 21760 39848 21972 40196
rect 22168 40120 22516 40196
rect 22168 39924 22380 40120
rect 22576 39924 22788 40196
rect 22168 39918 22788 39924
rect 22168 39854 22582 39918
rect 22646 39854 22788 39918
rect 22168 39848 22788 39854
rect 22984 40054 23196 40060
rect 22984 39990 22990 40054
rect 23054 39990 23196 40054
rect 22984 39918 23196 39990
rect 22984 39854 23126 39918
rect 23190 39854 23196 39918
rect 22984 39848 23196 39854
rect 23392 40054 23604 40060
rect 23392 39990 23398 40054
rect 23462 39990 23604 40054
rect 23392 39918 23604 39990
rect 28288 39984 28636 40468
rect 110160 40598 110508 40740
rect 115192 40870 115404 40876
rect 115192 40806 115198 40870
rect 115262 40806 115404 40870
rect 115192 40734 115404 40806
rect 115192 40670 115198 40734
rect 115262 40670 115404 40734
rect 115192 40664 115404 40670
rect 115600 40870 115812 40876
rect 115600 40806 115742 40870
rect 115806 40806 115812 40870
rect 115600 40734 115812 40806
rect 115600 40670 115742 40734
rect 115806 40670 115812 40734
rect 115600 40664 115812 40670
rect 116008 40870 116220 40876
rect 116008 40806 116014 40870
rect 116078 40806 116220 40870
rect 116008 40734 116220 40806
rect 116008 40670 116014 40734
rect 116078 40670 116220 40734
rect 116008 40664 116220 40670
rect 116416 40664 116628 40876
rect 116824 40870 117036 40876
rect 116824 40806 116966 40870
rect 117030 40806 117036 40870
rect 116824 40664 117036 40806
rect 136816 40740 137028 40876
rect 136816 40734 137572 40740
rect 136816 40728 137502 40734
rect 136816 40672 136944 40728
rect 137000 40672 137502 40728
rect 136816 40670 137502 40672
rect 137566 40670 137572 40734
rect 136816 40664 137572 40670
rect 116416 40604 116492 40664
rect 110160 40534 110166 40598
rect 110230 40534 110508 40598
rect 110160 40528 110508 40534
rect 116144 40528 116492 40604
rect 116824 40604 116900 40664
rect 110160 40468 110236 40528
rect 116144 40468 116220 40528
rect 110160 40326 110508 40468
rect 110160 40262 110166 40326
rect 110230 40262 110508 40326
rect 110160 39984 110508 40262
rect 115192 40462 115404 40468
rect 115192 40398 115198 40462
rect 115262 40398 115404 40462
rect 115192 40326 115404 40398
rect 115192 40262 115198 40326
rect 115262 40262 115404 40326
rect 115192 40256 115404 40262
rect 115600 40462 115812 40468
rect 115600 40398 115742 40462
rect 115806 40398 115812 40462
rect 115600 40326 115812 40398
rect 115600 40262 115606 40326
rect 115670 40262 115812 40326
rect 115600 40256 115812 40262
rect 116008 40462 116628 40468
rect 116008 40398 116014 40462
rect 116078 40398 116628 40462
rect 116008 40392 116628 40398
rect 116008 40332 116220 40392
rect 116008 40256 116356 40332
rect 116416 40256 116628 40392
rect 116824 40256 117036 40604
rect 136816 40528 137028 40664
rect 116144 40196 116220 40256
rect 115192 40054 115404 40060
rect 115192 39990 115198 40054
rect 115262 39990 115404 40054
rect 28560 39924 28636 39984
rect 110296 39924 110372 39984
rect 23392 39854 23534 39918
rect 23598 39854 23604 39918
rect 23392 39848 23604 39854
rect 21760 39788 21836 39848
rect 21760 39646 21972 39788
rect 28288 39782 28636 39924
rect 28288 39718 28430 39782
rect 28494 39718 28636 39782
rect 28288 39712 28636 39718
rect 110160 39712 110508 39924
rect 115192 39918 115404 39990
rect 115192 39854 115198 39918
rect 115262 39854 115404 39918
rect 115192 39848 115404 39854
rect 115600 40054 115812 40060
rect 115600 39990 115606 40054
rect 115670 39990 115812 40054
rect 115600 39918 115812 39990
rect 115600 39854 115606 39918
rect 115670 39854 115812 39918
rect 115600 39848 115812 39854
rect 116008 39848 116220 40196
rect 116280 40196 116356 40256
rect 116824 40196 116900 40256
rect 116280 40120 116628 40196
rect 116416 39918 116628 40120
rect 116416 39854 116422 39918
rect 116486 39854 116628 39918
rect 116416 39848 116628 39854
rect 116824 39848 117036 40196
rect 116960 39788 117036 39848
rect 28288 39652 28364 39712
rect 110296 39652 110372 39712
rect 21760 39582 21766 39646
rect 21830 39582 21972 39646
rect 21760 39576 21972 39582
rect 22168 39440 22380 39652
rect 22576 39646 22788 39652
rect 22576 39582 22582 39646
rect 22646 39582 22788 39646
rect 22576 39516 22788 39582
rect 22440 39440 22788 39516
rect 22984 39646 23196 39652
rect 22984 39582 23126 39646
rect 23190 39582 23196 39646
rect 22984 39440 23196 39582
rect 23392 39646 23604 39652
rect 23392 39582 23534 39646
rect 23598 39582 23604 39646
rect 23392 39440 23604 39582
rect 22168 39380 22244 39440
rect 22440 39380 22516 39440
rect 14552 39238 14764 39380
rect 14552 39174 14558 39238
rect 14622 39174 14764 39238
rect 14552 39168 14764 39174
rect 21760 39374 21972 39380
rect 21760 39310 21766 39374
rect 21830 39310 21972 39374
rect 21760 39238 21972 39310
rect 21760 39174 21902 39238
rect 21966 39174 21972 39238
rect 21760 39168 21972 39174
rect 22168 39304 22516 39380
rect 22576 39380 22652 39440
rect 23120 39380 23196 39440
rect 23528 39380 23604 39440
rect 22168 39244 22380 39304
rect 22168 39238 22516 39244
rect 22168 39174 22310 39238
rect 22374 39174 22446 39238
rect 22510 39174 22516 39238
rect 22168 39168 22516 39174
rect 22576 39168 22788 39380
rect 1224 39102 1980 39108
rect 1224 39038 1230 39102
rect 1294 39048 1980 39102
rect 1294 39038 1798 39048
rect 1224 39032 1798 39038
rect 1768 38992 1798 39032
rect 1854 38992 1980 39048
rect 1768 38896 1980 38992
rect 22984 39032 23196 39380
rect 23392 39032 23604 39380
rect 28288 39510 28636 39652
rect 28288 39446 28430 39510
rect 28494 39446 28636 39510
rect 28288 39374 28636 39446
rect 28288 39310 28294 39374
rect 28358 39310 28636 39374
rect 28288 39304 28636 39310
rect 110160 39374 110508 39652
rect 115192 39646 115404 39652
rect 115192 39582 115198 39646
rect 115262 39582 115404 39646
rect 115192 39440 115404 39582
rect 115600 39646 115812 39652
rect 115600 39582 115606 39646
rect 115670 39582 115812 39646
rect 115600 39440 115812 39582
rect 116008 39440 116220 39652
rect 115328 39380 115404 39440
rect 115736 39380 115812 39440
rect 116144 39380 116220 39440
rect 116416 39646 116628 39652
rect 116416 39582 116422 39646
rect 116486 39582 116628 39646
rect 116416 39440 116628 39582
rect 116824 39646 117036 39788
rect 116824 39582 116830 39646
rect 116894 39582 117036 39646
rect 116824 39576 117036 39582
rect 116416 39380 116492 39440
rect 110160 39310 110438 39374
rect 110502 39310 110508 39374
rect 110160 39304 110508 39310
rect 28288 39102 28636 39108
rect 28288 39038 28294 39102
rect 28358 39038 28636 39102
rect 22984 38972 23060 39032
rect 23392 38972 23468 39032
rect 21760 38966 21972 38972
rect 21760 38902 21902 38966
rect 21966 38902 21972 38966
rect 21760 38830 21972 38902
rect 21760 38766 21902 38830
rect 21966 38766 21972 38830
rect 21760 38760 21972 38766
rect 22168 38966 22380 38972
rect 22478 38966 22788 38972
rect 22168 38902 22310 38966
rect 22374 38902 22380 38966
rect 22440 38902 22446 38966
rect 22510 38902 22788 38966
rect 22168 38624 22380 38902
rect 22478 38896 22788 38902
rect 22576 38624 22788 38896
rect 22984 38624 23196 38972
rect 23392 38624 23604 38972
rect 22168 38564 22244 38624
rect 23120 38564 23196 38624
rect 23528 38564 23604 38624
rect 21760 38558 21972 38564
rect 21760 38494 21902 38558
rect 21966 38494 21972 38558
rect 15152 38475 15218 38478
rect 15886 38475 15952 38478
rect 15152 38473 15952 38475
rect 14144 38402 14356 38428
rect 15152 38417 15157 38473
rect 15213 38417 15891 38473
rect 15947 38417 15952 38473
rect 15152 38415 15952 38417
rect 15152 38412 15218 38415
rect 15886 38412 15952 38415
rect 21760 38422 21972 38494
rect 14144 38346 14212 38402
rect 14268 38346 14356 38402
rect 21760 38358 21902 38422
rect 21966 38358 21972 38422
rect 21760 38352 21972 38358
rect 22168 38422 22380 38564
rect 22168 38358 22174 38422
rect 22238 38358 22380 38422
rect 22168 38352 22380 38358
rect 22576 38422 22788 38564
rect 22576 38358 22718 38422
rect 22782 38358 22788 38422
rect 22576 38352 22788 38358
rect 22984 38422 23196 38564
rect 22984 38358 22990 38422
rect 23054 38358 23196 38422
rect 22984 38352 23196 38358
rect 23392 38422 23604 38564
rect 28288 38966 28636 39038
rect 28288 38902 28294 38966
rect 28358 38902 28636 38966
rect 28288 38694 28636 38902
rect 28288 38630 28294 38694
rect 28358 38630 28636 38694
rect 28288 38488 28636 38630
rect 110160 39102 110508 39108
rect 110160 39038 110438 39102
rect 110502 39038 110508 39102
rect 110160 38694 110508 39038
rect 110160 38630 110166 38694
rect 110230 38630 110508 38694
rect 110160 38488 110508 38630
rect 115192 39032 115404 39380
rect 115600 39032 115812 39380
rect 116008 39304 116628 39380
rect 116008 39168 116220 39304
rect 116416 39238 116628 39304
rect 116416 39174 116558 39238
rect 116622 39174 116628 39238
rect 116416 39168 116628 39174
rect 116824 39374 117036 39380
rect 116824 39310 116830 39374
rect 116894 39310 117036 39374
rect 116824 39238 117036 39310
rect 116824 39174 116966 39238
rect 117030 39174 117036 39238
rect 116824 39168 117036 39174
rect 136816 39048 137028 39108
rect 115192 38972 115268 39032
rect 115600 38972 115676 39032
rect 136816 38992 136944 39048
rect 137000 38992 137028 39048
rect 136816 38972 137028 38992
rect 115192 38624 115404 38972
rect 115600 38624 115812 38972
rect 115328 38564 115404 38624
rect 115736 38564 115812 38624
rect 28560 38428 28636 38488
rect 110296 38428 110372 38488
rect 23392 38358 23398 38422
rect 23462 38358 23604 38422
rect 23392 38352 23604 38358
rect 14144 38292 14356 38346
rect 0 38216 14356 38292
rect 21760 38150 21972 38156
rect 21760 38086 21902 38150
rect 21966 38086 21972 38150
rect 21760 38014 21972 38086
rect 21760 37950 21902 38014
rect 21966 37950 21972 38014
rect 21760 37944 21972 37950
rect 22168 38150 22380 38156
rect 22168 38086 22174 38150
rect 22238 38086 22380 38150
rect 22168 38020 22380 38086
rect 22576 38150 22788 38156
rect 22576 38086 22718 38150
rect 22782 38086 22788 38150
rect 22576 38020 22788 38086
rect 22168 37944 22788 38020
rect 22984 38150 23196 38156
rect 22984 38086 22990 38150
rect 23054 38086 23196 38150
rect 22984 38014 23196 38086
rect 22984 37950 22990 38014
rect 23054 37950 23196 38014
rect 22984 37944 23196 37950
rect 23392 38150 23604 38156
rect 23392 38086 23398 38150
rect 23462 38086 23604 38150
rect 23392 38014 23604 38086
rect 23392 37950 23398 38014
rect 23462 37950 23604 38014
rect 23392 37944 23604 37950
rect 28288 37944 28636 38428
rect 110160 38422 110508 38428
rect 110160 38358 110166 38422
rect 110230 38358 110508 38422
rect 110160 37944 110508 38358
rect 115192 38422 115404 38564
rect 115192 38358 115334 38422
rect 115398 38358 115404 38422
rect 115192 38352 115404 38358
rect 115600 38422 115812 38564
rect 115600 38358 115742 38422
rect 115806 38358 115812 38422
rect 115600 38352 115812 38358
rect 116008 38836 116220 38972
rect 116416 38966 116628 38972
rect 116416 38902 116558 38966
rect 116622 38902 116628 38966
rect 116416 38836 116628 38902
rect 116008 38760 116628 38836
rect 116824 38966 117036 38972
rect 116824 38902 116966 38966
rect 117030 38902 117036 38966
rect 116824 38830 117036 38902
rect 136816 38966 137572 38972
rect 136816 38902 137502 38966
rect 137566 38902 137572 38966
rect 136816 38896 137572 38902
rect 116824 38766 116966 38830
rect 117030 38766 117036 38830
rect 116824 38760 117036 38766
rect 116008 38624 116220 38760
rect 116416 38624 116628 38760
rect 116008 38564 116084 38624
rect 116416 38564 116492 38624
rect 116008 38422 116220 38564
rect 116008 38358 116014 38422
rect 116078 38358 116220 38422
rect 116008 38352 116220 38358
rect 116416 38352 116628 38564
rect 116824 38558 117036 38564
rect 116824 38494 116966 38558
rect 117030 38494 117036 38558
rect 116824 38422 117036 38494
rect 116824 38358 116830 38422
rect 116894 38358 117036 38422
rect 116824 38352 117036 38358
rect 115192 38150 115404 38156
rect 115192 38086 115334 38150
rect 115398 38086 115404 38150
rect 115192 38014 115404 38086
rect 115192 37950 115198 38014
rect 115262 37950 115404 38014
rect 115192 37944 115404 37950
rect 115600 38150 115812 38156
rect 115600 38086 115742 38150
rect 115806 38086 115812 38150
rect 115600 38014 115812 38086
rect 115600 37950 115606 38014
rect 115670 37950 115812 38014
rect 115600 37944 115812 37950
rect 116008 38150 116220 38156
rect 116008 38086 116014 38150
rect 116078 38086 116220 38150
rect 116008 38020 116220 38086
rect 116416 38020 116628 38156
rect 116008 38014 116628 38020
rect 116008 37950 116014 38014
rect 116078 37950 116628 38014
rect 116008 37944 116628 37950
rect 116824 38150 117036 38156
rect 116824 38086 116830 38150
rect 116894 38086 117036 38150
rect 116824 38014 117036 38086
rect 116824 37950 116966 38014
rect 117030 37950 117036 38014
rect 116824 37944 117036 37950
rect 22304 37884 22380 37944
rect 28424 37884 28500 37944
rect 110432 37884 110508 37944
rect 14552 37878 14764 37884
rect 14552 37814 14694 37878
rect 14758 37814 14764 37878
rect 14552 37748 14764 37814
rect 22304 37808 22652 37884
rect 22576 37748 22652 37808
rect 14552 37742 14900 37748
rect 14552 37678 14830 37742
rect 14894 37678 14900 37742
rect 14552 37672 14900 37678
rect 21760 37742 21972 37748
rect 21760 37678 21902 37742
rect 21966 37678 21972 37742
rect 21760 37606 21972 37678
rect 21760 37542 21766 37606
rect 21830 37542 21972 37606
rect 21760 37536 21972 37542
rect 22168 37672 22788 37748
rect 22168 37612 22380 37672
rect 22168 37606 22516 37612
rect 22168 37542 22174 37606
rect 22238 37542 22446 37606
rect 22510 37542 22516 37606
rect 22168 37536 22516 37542
rect 22576 37536 22788 37672
rect 22984 37742 23196 37748
rect 22984 37678 22990 37742
rect 23054 37678 23196 37742
rect 22984 37606 23196 37678
rect 22984 37542 23126 37606
rect 23190 37542 23196 37606
rect 22984 37536 23196 37542
rect 23392 37742 23604 37748
rect 23392 37678 23398 37742
rect 23462 37678 23604 37742
rect 23392 37606 23604 37678
rect 28288 37672 28636 37884
rect 110160 37672 110508 37884
rect 115192 37742 115404 37748
rect 115192 37678 115198 37742
rect 115262 37678 115404 37742
rect 28424 37612 28500 37672
rect 110160 37612 110236 37672
rect 23392 37542 23534 37606
rect 23598 37542 23604 37606
rect 23392 37536 23604 37542
rect 1224 37470 1980 37476
rect 1224 37406 1230 37470
rect 1294 37406 1980 37470
rect 1224 37400 1980 37406
rect 28288 37400 28636 37612
rect 110160 37400 110508 37612
rect 115192 37606 115404 37678
rect 115192 37542 115334 37606
rect 115398 37542 115404 37606
rect 115192 37536 115404 37542
rect 115600 37742 115812 37748
rect 115600 37678 115606 37742
rect 115670 37678 115812 37742
rect 115600 37606 115812 37678
rect 115600 37542 115742 37606
rect 115806 37542 115812 37606
rect 115600 37536 115812 37542
rect 116008 37742 116220 37748
rect 116008 37678 116014 37742
rect 116078 37678 116220 37742
rect 116008 37606 116220 37678
rect 116416 37612 116628 37748
rect 116318 37606 116628 37612
rect 116008 37542 116150 37606
rect 116214 37542 116220 37606
rect 116280 37542 116286 37606
rect 116350 37542 116628 37606
rect 116008 37536 116220 37542
rect 116318 37536 116628 37542
rect 116824 37742 117036 37748
rect 116824 37678 116966 37742
rect 117030 37678 117036 37742
rect 116824 37606 117036 37678
rect 116824 37542 116830 37606
rect 116894 37542 117036 37606
rect 116824 37536 117036 37542
rect 1777 37368 1875 37400
rect 1777 37312 1798 37368
rect 1854 37312 1875 37368
rect 28288 37340 28364 37400
rect 110296 37340 110372 37400
rect 136816 37368 137028 37476
rect 1777 37291 1875 37312
rect 14144 37274 14356 37340
rect 14144 37218 14212 37274
rect 14268 37218 14356 37274
rect 14144 37204 14356 37218
rect 21760 37334 21972 37340
rect 21760 37270 21766 37334
rect 21830 37270 21972 37334
rect 0 37128 14356 37204
rect 15152 37205 15218 37208
rect 15806 37205 15872 37208
rect 15152 37203 15872 37205
rect 15152 37147 15157 37203
rect 15213 37147 15811 37203
rect 15867 37147 15872 37203
rect 15152 37145 15872 37147
rect 15152 37142 15218 37145
rect 15806 37142 15872 37145
rect 21760 37198 21972 37270
rect 21760 37134 21902 37198
rect 21966 37134 21972 37198
rect 21760 37128 21972 37134
rect 22168 37334 22380 37340
rect 22478 37334 22788 37340
rect 22168 37270 22174 37334
rect 22238 37270 22380 37334
rect 22440 37270 22446 37334
rect 22510 37270 22788 37334
rect 22168 37128 22380 37270
rect 22478 37264 22788 37270
rect 22576 37128 22788 37264
rect 22984 37334 23196 37340
rect 22984 37270 23126 37334
rect 23190 37270 23196 37334
rect 22984 37198 23196 37270
rect 22984 37134 22990 37198
rect 23054 37134 23196 37198
rect 22984 37128 23196 37134
rect 23392 37334 23604 37340
rect 23392 37270 23534 37334
rect 23598 37270 23604 37334
rect 23392 37198 23604 37270
rect 23392 37134 23398 37198
rect 23462 37134 23604 37198
rect 23392 37128 23604 37134
rect 28288 37128 28636 37340
rect 110160 37128 110508 37340
rect 115192 37334 115404 37340
rect 115192 37270 115334 37334
rect 115398 37270 115404 37334
rect 115192 37198 115404 37270
rect 115192 37134 115334 37198
rect 115398 37134 115404 37198
rect 115192 37128 115404 37134
rect 115600 37334 115812 37340
rect 115600 37270 115742 37334
rect 115806 37270 115812 37334
rect 115600 37198 115812 37270
rect 115600 37134 115606 37198
rect 115670 37134 115812 37198
rect 115600 37128 115812 37134
rect 116008 37334 116356 37340
rect 116008 37270 116150 37334
rect 116214 37270 116286 37334
rect 116350 37270 116356 37334
rect 116008 37264 116356 37270
rect 116008 37204 116220 37264
rect 116008 37198 116356 37204
rect 116008 37134 116150 37198
rect 116214 37134 116286 37198
rect 116350 37134 116356 37198
rect 116008 37128 116356 37134
rect 116416 37198 116628 37340
rect 116416 37134 116558 37198
rect 116622 37134 116628 37198
rect 116416 37128 116628 37134
rect 116824 37334 117036 37340
rect 116824 37270 116830 37334
rect 116894 37270 117036 37334
rect 116824 37198 117036 37270
rect 136816 37312 136944 37368
rect 137000 37340 137028 37368
rect 137000 37334 137572 37340
rect 137000 37312 137502 37334
rect 136816 37270 137502 37312
rect 137566 37270 137572 37334
rect 136816 37264 137572 37270
rect 116824 37134 116830 37198
rect 116894 37134 117036 37198
rect 116824 37128 117036 37134
rect 22576 37068 22652 37128
rect 22304 36992 22652 37068
rect 28288 37068 28364 37128
rect 110296 37068 110372 37128
rect 22304 36932 22380 36992
rect 21760 36926 21972 36932
rect 21760 36862 21902 36926
rect 21966 36862 21972 36926
rect 21760 36720 21972 36862
rect 22168 36856 22788 36932
rect 22168 36790 22380 36856
rect 22168 36726 22174 36790
rect 22238 36726 22380 36790
rect 22168 36720 22380 36726
rect 22576 36790 22788 36856
rect 22576 36726 22718 36790
rect 22782 36726 22788 36790
rect 22576 36720 22788 36726
rect 22984 36926 23196 36932
rect 22984 36862 22990 36926
rect 23054 36862 23196 36926
rect 22984 36790 23196 36862
rect 22984 36726 22990 36790
rect 23054 36726 23196 36790
rect 22984 36720 23196 36726
rect 23392 36926 23604 36932
rect 23392 36862 23398 36926
rect 23462 36862 23604 36926
rect 23392 36790 23604 36862
rect 28288 36856 28636 37068
rect 28560 36796 28636 36856
rect 23392 36726 23398 36790
rect 23462 36726 23604 36790
rect 23392 36720 23604 36726
rect 21896 36660 21972 36720
rect 14552 36518 14764 36524
rect 14552 36454 14558 36518
rect 14622 36454 14764 36518
rect 14552 36382 14764 36454
rect 14552 36318 14694 36382
rect 14758 36318 14764 36382
rect 14552 36312 14764 36318
rect 21760 36382 21972 36660
rect 28288 36584 28636 36796
rect 110160 36856 110508 37068
rect 115192 36926 115404 36932
rect 115192 36862 115334 36926
rect 115398 36862 115404 36926
rect 110160 36796 110236 36856
rect 110160 36584 110508 36796
rect 115192 36790 115404 36862
rect 115192 36726 115198 36790
rect 115262 36726 115404 36790
rect 115192 36720 115404 36726
rect 115600 36926 115812 36932
rect 115600 36862 115606 36926
rect 115670 36862 115812 36926
rect 115600 36790 115812 36862
rect 115600 36726 115606 36790
rect 115670 36726 115812 36790
rect 115600 36720 115812 36726
rect 116008 36926 116220 36932
rect 116318 36926 116628 36932
rect 116008 36862 116150 36926
rect 116214 36862 116220 36926
rect 116280 36862 116286 36926
rect 116350 36862 116558 36926
rect 116622 36862 116628 36926
rect 116008 36796 116220 36862
rect 116318 36856 116628 36862
rect 116008 36790 116356 36796
rect 116008 36726 116014 36790
rect 116078 36726 116286 36790
rect 116350 36726 116356 36790
rect 116008 36720 116356 36726
rect 116416 36720 116628 36856
rect 116824 36926 117036 36932
rect 116824 36862 116830 36926
rect 116894 36862 117036 36926
rect 116824 36720 117036 36862
rect 116960 36660 117036 36720
rect 28288 36524 28364 36584
rect 110296 36524 110372 36584
rect 21760 36318 21902 36382
rect 21966 36318 21972 36382
rect 21760 36312 21972 36318
rect 22168 36518 22380 36524
rect 22168 36454 22174 36518
rect 22238 36454 22380 36518
rect 22168 36382 22380 36454
rect 22168 36318 22174 36382
rect 22238 36318 22380 36382
rect 22168 36312 22380 36318
rect 22576 36518 22788 36524
rect 22576 36454 22718 36518
rect 22782 36454 22788 36518
rect 22576 36382 22788 36454
rect 22576 36318 22582 36382
rect 22646 36318 22788 36382
rect 22576 36312 22788 36318
rect 22984 36518 23196 36524
rect 22984 36454 22990 36518
rect 23054 36454 23196 36518
rect 22984 36382 23196 36454
rect 22984 36318 22990 36382
rect 23054 36318 23196 36382
rect 22984 36312 23196 36318
rect 23392 36518 23604 36524
rect 23392 36454 23398 36518
rect 23462 36454 23604 36518
rect 23392 36382 23604 36454
rect 23392 36318 23534 36382
rect 23598 36318 23604 36382
rect 23392 36312 23604 36318
rect 28288 36312 28636 36524
rect 110160 36312 110508 36524
rect 115192 36518 115404 36524
rect 115192 36454 115198 36518
rect 115262 36454 115404 36518
rect 115192 36382 115404 36454
rect 115192 36318 115334 36382
rect 115398 36318 115404 36382
rect 115192 36312 115404 36318
rect 115600 36518 115812 36524
rect 115600 36454 115606 36518
rect 115670 36454 115812 36518
rect 115600 36382 115812 36454
rect 115600 36318 115742 36382
rect 115806 36318 115812 36382
rect 115600 36312 115812 36318
rect 116008 36518 116220 36524
rect 116318 36518 116628 36524
rect 116008 36454 116014 36518
rect 116078 36454 116220 36518
rect 116280 36454 116286 36518
rect 116350 36454 116628 36518
rect 116008 36312 116220 36454
rect 116318 36448 116628 36454
rect 116416 36388 116628 36448
rect 116318 36382 116628 36388
rect 116280 36318 116286 36382
rect 116350 36318 116628 36382
rect 116318 36312 116628 36318
rect 116824 36382 117036 36660
rect 116824 36318 116966 36382
rect 117030 36318 117036 36382
rect 116824 36312 117036 36318
rect 28288 36252 28364 36312
rect 110160 36252 110236 36312
rect 21760 36110 21972 36116
rect 21760 36046 21902 36110
rect 21966 36046 21972 36110
rect 21760 35904 21972 36046
rect 22168 36110 22380 36116
rect 22168 36046 22174 36110
rect 22238 36046 22380 36110
rect 22168 35904 22380 36046
rect 22576 36110 22788 36116
rect 22576 36046 22582 36110
rect 22646 36046 22788 36110
rect 22576 35974 22788 36046
rect 22576 35910 22718 35974
rect 22782 35910 22788 35974
rect 22576 35904 22788 35910
rect 22984 36110 23196 36116
rect 22984 36046 22990 36110
rect 23054 36046 23196 36110
rect 22984 35974 23196 36046
rect 22984 35910 23126 35974
rect 23190 35910 23196 35974
rect 22984 35904 23196 35910
rect 23392 36110 23604 36116
rect 23392 36046 23534 36110
rect 23598 36046 23604 36110
rect 23392 35974 23604 36046
rect 28288 36040 28636 36252
rect 110160 36040 110508 36252
rect 115192 36110 115404 36116
rect 115192 36046 115334 36110
rect 115398 36046 115404 36110
rect 28424 35980 28500 36040
rect 110296 35980 110372 36040
rect 23392 35910 23398 35974
rect 23462 35910 23604 35974
rect 23392 35904 23604 35910
rect 21896 35844 21972 35904
rect 1224 35838 1980 35844
rect 1224 35774 1230 35838
rect 1294 35774 1980 35838
rect 1224 35768 1980 35774
rect 1768 35688 1875 35768
rect 1768 35632 1798 35688
rect 1854 35632 1875 35688
rect 1777 35611 1875 35632
rect 14144 35574 14356 35708
rect 21760 35702 21972 35844
rect 28288 35838 28636 35980
rect 28288 35774 28566 35838
rect 28630 35774 28636 35838
rect 28288 35768 28636 35774
rect 28560 35708 28636 35768
rect 15152 35647 15218 35650
rect 15726 35647 15792 35650
rect 15152 35645 15792 35647
rect 15152 35589 15157 35645
rect 15213 35589 15731 35645
rect 15787 35589 15792 35645
rect 21760 35638 21902 35702
rect 21966 35638 21972 35702
rect 21760 35632 21972 35638
rect 22168 35702 22788 35708
rect 22168 35638 22718 35702
rect 22782 35638 22788 35702
rect 22168 35632 22788 35638
rect 15152 35587 15792 35589
rect 15152 35584 15218 35587
rect 15726 35584 15792 35587
rect 14144 35572 14212 35574
rect 2040 35518 14212 35572
rect 14268 35518 14356 35574
rect 2040 35496 14356 35518
rect 22168 35572 22380 35632
rect 22168 35496 22516 35572
rect 22576 35496 22788 35632
rect 22984 35702 23196 35708
rect 22984 35638 23126 35702
rect 23190 35638 23196 35702
rect 22984 35496 23196 35638
rect 2040 35436 2116 35496
rect 22168 35436 22244 35496
rect 22440 35436 22516 35496
rect 23120 35436 23196 35496
rect 0 35360 2116 35436
rect 21760 35430 21972 35436
rect 21760 35366 21902 35430
rect 21966 35366 21972 35430
rect 21760 35294 21972 35366
rect 21760 35230 21766 35294
rect 21830 35230 21972 35294
rect 21760 35224 21972 35230
rect 22168 35224 22380 35436
rect 22440 35360 22788 35436
rect 22576 35294 22788 35360
rect 22576 35230 22582 35294
rect 22646 35230 22788 35294
rect 22576 35224 22788 35230
rect 14552 35158 14862 35164
rect 14552 35094 14830 35158
rect 14894 35094 14900 35158
rect 14552 35088 14862 35094
rect 22984 35088 23196 35436
rect 14552 34886 14764 35088
rect 23120 35028 23196 35088
rect 14552 34822 14558 34886
rect 14622 34822 14764 34886
rect 14552 34816 14764 34822
rect 21760 35022 21972 35028
rect 21760 34958 21766 35022
rect 21830 34958 21972 35022
rect 21760 34886 21972 34958
rect 21760 34822 21902 34886
rect 21966 34822 21972 34886
rect 21760 34816 21972 34822
rect 22168 34886 22788 34892
rect 22168 34822 22582 34886
rect 22646 34822 22788 34886
rect 22168 34816 22788 34822
rect 22168 34680 22380 34816
rect 22576 34756 22788 34816
rect 22440 34680 22788 34756
rect 22984 34680 23196 35028
rect 22440 34620 22516 34680
rect 22712 34620 22788 34680
rect 23120 34620 23196 34680
rect 21760 34614 21972 34620
rect 21760 34550 21902 34614
rect 21966 34550 21972 34614
rect 14144 34446 14356 34484
rect 14144 34390 14212 34446
rect 14268 34390 14356 34446
rect 21760 34478 21972 34550
rect 21760 34414 21902 34478
rect 21966 34414 21972 34478
rect 21760 34408 21972 34414
rect 22168 34544 22516 34620
rect 22168 34484 22380 34544
rect 22168 34478 22516 34484
rect 22168 34414 22446 34478
rect 22510 34414 22516 34478
rect 22168 34408 22516 34414
rect 22576 34408 22788 34620
rect 22984 34478 23196 34620
rect 22984 34414 23126 34478
rect 23190 34414 23196 34478
rect 22984 34408 23196 34414
rect 23392 35702 23604 35708
rect 23392 35638 23398 35702
rect 23462 35638 23604 35702
rect 23392 35496 23604 35638
rect 28288 35566 28636 35708
rect 28288 35502 28566 35566
rect 28630 35502 28636 35566
rect 28288 35496 28636 35502
rect 110160 35838 110508 35980
rect 115192 35974 115404 36046
rect 115192 35910 115334 35974
rect 115398 35910 115404 35974
rect 115192 35904 115404 35910
rect 115600 36110 115812 36116
rect 115600 36046 115742 36110
rect 115806 36046 115812 36110
rect 115600 35974 115812 36046
rect 115600 35910 115606 35974
rect 115670 35910 115812 35974
rect 115600 35904 115812 35910
rect 116008 36110 116356 36116
rect 116008 36046 116286 36110
rect 116350 36046 116356 36110
rect 116008 36040 116356 36046
rect 116008 35980 116220 36040
rect 116416 35980 116628 36116
rect 116008 35974 116628 35980
rect 116008 35910 116558 35974
rect 116622 35910 116628 35974
rect 116008 35904 116628 35910
rect 116824 36110 117036 36116
rect 116824 36046 116966 36110
rect 117030 36046 117036 36110
rect 116824 35904 117036 36046
rect 116960 35844 117036 35904
rect 110160 35774 110302 35838
rect 110366 35774 110508 35838
rect 110160 35768 110508 35774
rect 110160 35708 110236 35768
rect 110160 35566 110508 35708
rect 110160 35502 110302 35566
rect 110366 35502 110508 35566
rect 110160 35496 110508 35502
rect 115192 35702 115404 35708
rect 115192 35638 115334 35702
rect 115398 35638 115404 35702
rect 115192 35496 115404 35638
rect 23392 35436 23468 35496
rect 23392 35088 23604 35436
rect 28406 35300 28504 35496
rect 110294 35300 110392 35496
rect 115328 35436 115404 35496
rect 28288 35224 28636 35300
rect 110160 35224 110508 35300
rect 28288 35164 28364 35224
rect 110432 35164 110508 35224
rect 23392 35028 23468 35088
rect 23392 34680 23604 35028
rect 23392 34620 23468 34680
rect 23392 34478 23604 34620
rect 23392 34414 23398 34478
rect 23462 34414 23604 34478
rect 23392 34408 23604 34414
rect 28288 34544 28636 35164
rect 110160 35022 110508 35164
rect 115192 35088 115404 35436
rect 115600 35702 115812 35708
rect 115600 35638 115606 35702
rect 115670 35638 115812 35702
rect 115600 35496 115812 35638
rect 116008 35702 116356 35708
rect 116008 35638 116286 35702
rect 116350 35638 116356 35702
rect 116008 35632 116356 35638
rect 116416 35702 116628 35708
rect 116416 35638 116558 35702
rect 116622 35638 116628 35702
rect 116008 35572 116220 35632
rect 116416 35572 116628 35638
rect 116824 35702 117036 35844
rect 116824 35638 116966 35702
rect 117030 35638 117036 35702
rect 116824 35632 117036 35638
rect 136816 35708 137028 35844
rect 136816 35702 137572 35708
rect 136816 35688 137502 35702
rect 136816 35632 136944 35688
rect 137000 35638 137502 35688
rect 137566 35638 137572 35702
rect 137000 35632 137572 35638
rect 116008 35496 116628 35572
rect 136816 35496 137028 35632
rect 115600 35436 115676 35496
rect 116008 35436 116084 35496
rect 115600 35088 115812 35436
rect 116008 35224 116220 35436
rect 116318 35430 116628 35436
rect 116280 35366 116286 35430
rect 116350 35366 116628 35430
rect 116318 35360 116628 35366
rect 116416 35294 116628 35360
rect 116416 35230 116558 35294
rect 116622 35230 116628 35294
rect 116416 35224 116628 35230
rect 116824 35430 117036 35436
rect 116824 35366 116966 35430
rect 117030 35366 117036 35430
rect 116824 35294 117036 35366
rect 116824 35230 116830 35294
rect 116894 35230 117036 35294
rect 116824 35224 117036 35230
rect 115328 35028 115404 35088
rect 115736 35028 115812 35088
rect 110160 34958 110438 35022
rect 110502 34958 110508 35022
rect 110160 34750 110508 34958
rect 110160 34686 110166 34750
rect 110230 34686 110438 34750
rect 110502 34686 110508 34750
rect 110160 34544 110508 34686
rect 115192 34680 115404 35028
rect 115328 34620 115404 34680
rect 28288 34484 28364 34544
rect 110432 34484 110508 34544
rect 14144 34348 14356 34390
rect 0 34272 14356 34348
rect 15152 34377 15218 34380
rect 15646 34377 15712 34380
rect 15152 34375 15712 34377
rect 15152 34319 15157 34375
rect 15213 34319 15651 34375
rect 15707 34319 15712 34375
rect 15152 34317 15712 34319
rect 15152 34314 15218 34317
rect 15646 34314 15712 34317
rect 21760 34206 21972 34212
rect 21760 34142 21902 34206
rect 21966 34142 21972 34206
rect 1224 34070 1980 34076
rect 1224 34006 1230 34070
rect 1294 34008 1980 34070
rect 1294 34006 1798 34008
rect 1224 34000 1798 34006
rect 1768 33952 1798 34000
rect 1854 33952 1980 34008
rect 21760 34070 21972 34142
rect 21760 34006 21766 34070
rect 21830 34006 21972 34070
rect 21760 34000 21972 34006
rect 22168 34070 22380 34212
rect 22478 34206 22788 34212
rect 22440 34142 22446 34206
rect 22510 34142 22788 34206
rect 22478 34136 22788 34142
rect 22168 34006 22174 34070
rect 22238 34006 22380 34070
rect 22168 34000 22380 34006
rect 22576 34070 22788 34136
rect 22576 34006 22718 34070
rect 22782 34006 22788 34070
rect 22576 34000 22788 34006
rect 22984 34206 23196 34212
rect 22984 34142 23126 34206
rect 23190 34142 23196 34206
rect 22984 34070 23196 34142
rect 22984 34006 22990 34070
rect 23054 34006 23196 34070
rect 22984 34000 23196 34006
rect 23392 34206 23604 34212
rect 23392 34142 23398 34206
rect 23462 34142 23604 34206
rect 23392 34070 23604 34142
rect 23392 34006 23534 34070
rect 23598 34006 23604 34070
rect 23392 34000 23604 34006
rect 28288 34206 28636 34484
rect 28288 34142 28294 34206
rect 28358 34142 28636 34206
rect 28288 34000 28636 34142
rect 110160 34478 110508 34484
rect 110160 34414 110166 34478
rect 110230 34414 110508 34478
rect 110160 34000 110508 34414
rect 115192 34478 115404 34620
rect 115192 34414 115334 34478
rect 115398 34414 115404 34478
rect 115192 34408 115404 34414
rect 115600 34680 115812 35028
rect 116824 35022 117036 35028
rect 116824 34958 116830 35022
rect 116894 34958 117036 35022
rect 116008 34680 116220 34892
rect 116416 34886 116628 34892
rect 116416 34822 116558 34886
rect 116622 34822 116628 34886
rect 116416 34756 116628 34822
rect 116824 34886 117036 34958
rect 116824 34822 116966 34886
rect 117030 34822 117036 34886
rect 116824 34816 117036 34822
rect 115600 34620 115676 34680
rect 116144 34620 116220 34680
rect 116280 34680 116628 34756
rect 116280 34620 116356 34680
rect 115600 34478 115812 34620
rect 115600 34414 115606 34478
rect 115670 34414 115812 34478
rect 115600 34408 115812 34414
rect 116008 34544 116356 34620
rect 116008 34484 116220 34544
rect 116416 34484 116628 34620
rect 116008 34478 116628 34484
rect 116008 34414 116014 34478
rect 116078 34414 116628 34478
rect 116008 34408 116628 34414
rect 116824 34614 117036 34620
rect 116824 34550 116966 34614
rect 117030 34550 117036 34614
rect 116824 34478 117036 34550
rect 116824 34414 116966 34478
rect 117030 34414 117036 34478
rect 116824 34408 117036 34414
rect 116144 34348 116220 34408
rect 116144 34272 116492 34348
rect 116416 34212 116492 34272
rect 115192 34206 115404 34212
rect 115192 34142 115334 34206
rect 115398 34142 115404 34206
rect 115192 34070 115404 34142
rect 115192 34006 115334 34070
rect 115398 34006 115404 34070
rect 115192 34000 115404 34006
rect 115600 34206 115812 34212
rect 115600 34142 115606 34206
rect 115670 34142 115812 34206
rect 115600 34070 115812 34142
rect 115600 34006 115606 34070
rect 115670 34006 115812 34070
rect 115600 34000 115812 34006
rect 116008 34206 116220 34212
rect 116008 34142 116014 34206
rect 116078 34142 116220 34206
rect 116008 34000 116220 34142
rect 116416 34076 116628 34212
rect 116318 34070 116628 34076
rect 116280 34006 116286 34070
rect 116350 34006 116558 34070
rect 116622 34006 116628 34070
rect 116318 34000 116628 34006
rect 116824 34206 117036 34212
rect 116824 34142 116966 34206
rect 117030 34142 117036 34206
rect 116824 34070 117036 34142
rect 116824 34006 116830 34070
rect 116894 34006 117036 34070
rect 116824 34000 117036 34006
rect 136816 34070 137572 34076
rect 136816 34008 137502 34070
rect 1768 33864 1980 33952
rect 28424 33940 28500 34000
rect 110432 33940 110508 34000
rect 28288 33934 28636 33940
rect 28288 33870 28294 33934
rect 28358 33870 28636 33934
rect 21760 33798 21972 33804
rect 21760 33734 21766 33798
rect 21830 33734 21972 33798
rect 14552 33662 14764 33668
rect 14552 33598 14694 33662
rect 14758 33598 14764 33662
rect 14552 33526 14764 33598
rect 21760 33662 21972 33734
rect 21760 33598 21902 33662
rect 21966 33598 21972 33662
rect 21760 33592 21972 33598
rect 22168 33798 22380 33804
rect 22168 33734 22174 33798
rect 22238 33734 22380 33798
rect 22168 33668 22380 33734
rect 22576 33798 22788 33804
rect 22576 33734 22718 33798
rect 22782 33734 22788 33798
rect 22576 33668 22788 33734
rect 22168 33592 22788 33668
rect 22984 33798 23196 33804
rect 22984 33734 22990 33798
rect 23054 33734 23196 33798
rect 22984 33662 23196 33734
rect 22984 33598 23126 33662
rect 23190 33598 23196 33662
rect 22984 33592 23196 33598
rect 23392 33798 23604 33804
rect 23392 33734 23534 33798
rect 23598 33734 23604 33798
rect 23392 33662 23604 33734
rect 28288 33728 28636 33870
rect 28560 33668 28636 33728
rect 23392 33598 23398 33662
rect 23462 33598 23604 33662
rect 23392 33592 23604 33598
rect 14552 33462 14694 33526
rect 14758 33462 14764 33526
rect 14552 33456 14764 33462
rect 22304 33532 22380 33592
rect 22304 33456 22652 33532
rect 28288 33456 28636 33668
rect 110160 33728 110508 33940
rect 136816 33952 136944 34008
rect 137000 34006 137502 34008
rect 137566 34006 137572 34070
rect 137000 34000 137572 34006
rect 137000 33952 137028 34000
rect 136816 33864 137028 33952
rect 115192 33798 115404 33804
rect 115192 33734 115334 33798
rect 115398 33734 115404 33798
rect 110160 33668 110236 33728
rect 110160 33456 110508 33668
rect 115192 33662 115404 33734
rect 115192 33598 115198 33662
rect 115262 33598 115404 33662
rect 115192 33592 115404 33598
rect 115600 33798 115812 33804
rect 115600 33734 115606 33798
rect 115670 33734 115812 33798
rect 115600 33662 115812 33734
rect 115600 33598 115606 33662
rect 115670 33598 115812 33662
rect 115600 33592 115812 33598
rect 116008 33798 116356 33804
rect 116008 33734 116286 33798
rect 116350 33734 116356 33798
rect 116008 33728 116356 33734
rect 116416 33798 116628 33804
rect 116416 33734 116558 33798
rect 116622 33734 116628 33798
rect 116008 33662 116220 33728
rect 116008 33598 116150 33662
rect 116214 33598 116220 33662
rect 116008 33592 116220 33598
rect 116416 33592 116628 33734
rect 116824 33798 117036 33804
rect 116824 33734 116830 33798
rect 116894 33734 117036 33798
rect 116824 33662 117036 33734
rect 116824 33598 116966 33662
rect 117030 33598 117036 33662
rect 116824 33592 117036 33598
rect 22576 33396 22652 33456
rect 28424 33396 28500 33456
rect 110160 33396 110236 33456
rect 21760 33390 21972 33396
rect 21760 33326 21902 33390
rect 21966 33326 21972 33390
rect 21760 33254 21972 33326
rect 21760 33190 21766 33254
rect 21830 33190 21972 33254
rect 21760 33184 21972 33190
rect 22168 33254 22380 33396
rect 22168 33190 22174 33254
rect 22238 33190 22380 33254
rect 22168 33184 22380 33190
rect 22576 33254 22788 33396
rect 22576 33190 22582 33254
rect 22646 33190 22788 33254
rect 22576 33184 22788 33190
rect 22984 33390 23196 33396
rect 22984 33326 23126 33390
rect 23190 33326 23196 33390
rect 22984 33254 23196 33326
rect 22984 33190 22990 33254
rect 23054 33190 23196 33254
rect 22984 33184 23196 33190
rect 23392 33390 23604 33396
rect 23392 33326 23398 33390
rect 23462 33326 23604 33390
rect 23392 33254 23604 33326
rect 23392 33190 23534 33254
rect 23598 33190 23604 33254
rect 23392 33184 23604 33190
rect 28288 33184 28636 33396
rect 110160 33184 110508 33396
rect 115192 33390 115404 33396
rect 115192 33326 115198 33390
rect 115262 33326 115404 33390
rect 115192 33254 115404 33326
rect 115192 33190 115334 33254
rect 115398 33190 115404 33254
rect 115192 33184 115404 33190
rect 115600 33390 115812 33396
rect 115600 33326 115606 33390
rect 115670 33326 115812 33390
rect 115600 33254 115812 33326
rect 115600 33190 115742 33254
rect 115806 33190 115812 33254
rect 115600 33184 115812 33190
rect 116008 33390 116220 33396
rect 116008 33326 116150 33390
rect 116214 33326 116220 33390
rect 116008 33254 116220 33326
rect 116008 33190 116150 33254
rect 116214 33190 116220 33254
rect 116008 33184 116220 33190
rect 116416 33254 116628 33396
rect 116416 33190 116422 33254
rect 116486 33190 116628 33254
rect 116416 33184 116628 33190
rect 116824 33390 117036 33396
rect 116824 33326 116966 33390
rect 117030 33326 117036 33390
rect 116824 33254 117036 33326
rect 116824 33190 116830 33254
rect 116894 33190 117036 33254
rect 116824 33184 117036 33190
rect 28424 33124 28500 33184
rect 110432 33124 110508 33184
rect 21760 32982 21972 32988
rect 21760 32918 21766 32982
rect 21830 32918 21972 32982
rect 0 32776 14356 32852
rect 21760 32846 21972 32918
rect 14144 32746 14356 32776
rect 15152 32819 15218 32822
rect 15566 32819 15632 32822
rect 15152 32817 15632 32819
rect 15152 32761 15157 32817
rect 15213 32761 15571 32817
rect 15627 32761 15632 32817
rect 21760 32782 21902 32846
rect 21966 32782 21972 32846
rect 21760 32776 21972 32782
rect 22168 32982 22380 32988
rect 22168 32918 22174 32982
rect 22238 32918 22380 32982
rect 22168 32846 22380 32918
rect 22576 32982 22788 32988
rect 22576 32918 22582 32982
rect 22646 32918 22788 32982
rect 22576 32852 22788 32918
rect 22478 32846 22788 32852
rect 22168 32782 22310 32846
rect 22374 32782 22380 32846
rect 22440 32782 22446 32846
rect 22510 32782 22788 32846
rect 22168 32776 22380 32782
rect 22478 32776 22788 32782
rect 22984 32982 23196 32988
rect 22984 32918 22990 32982
rect 23054 32918 23196 32982
rect 22984 32846 23196 32918
rect 22984 32782 22990 32846
rect 23054 32782 23196 32846
rect 22984 32776 23196 32782
rect 23392 32982 23604 32988
rect 23392 32918 23534 32982
rect 23598 32918 23604 32982
rect 23392 32846 23604 32918
rect 23392 32782 23534 32846
rect 23598 32782 23604 32846
rect 23392 32776 23604 32782
rect 28288 32912 28636 33124
rect 110160 32912 110508 33124
rect 115192 32982 115404 32988
rect 115192 32918 115334 32982
rect 115398 32918 115404 32982
rect 28288 32852 28364 32912
rect 110296 32852 110372 32912
rect 15152 32759 15632 32761
rect 15152 32756 15218 32759
rect 15566 32756 15632 32759
rect 14144 32690 14212 32746
rect 14268 32690 14356 32746
rect 14144 32640 14356 32690
rect 28288 32640 28636 32852
rect 110160 32640 110508 32852
rect 115192 32846 115404 32918
rect 115192 32782 115334 32846
rect 115398 32782 115404 32846
rect 115192 32776 115404 32782
rect 115600 32982 115812 32988
rect 115600 32918 115742 32982
rect 115806 32918 115812 32982
rect 115600 32846 115812 32918
rect 115600 32782 115606 32846
rect 115670 32782 115812 32846
rect 115600 32776 115812 32782
rect 116008 32982 116628 32988
rect 116008 32918 116150 32982
rect 116214 32918 116422 32982
rect 116486 32918 116628 32982
rect 116008 32912 116628 32918
rect 116008 32852 116220 32912
rect 116008 32846 116356 32852
rect 116008 32782 116014 32846
rect 116078 32782 116286 32846
rect 116350 32782 116356 32846
rect 116008 32776 116356 32782
rect 116416 32776 116628 32912
rect 116824 32982 117036 32988
rect 116824 32918 116830 32982
rect 116894 32918 117036 32982
rect 116824 32846 117036 32918
rect 116824 32782 116830 32846
rect 116894 32782 117036 32846
rect 116824 32776 117036 32782
rect 28288 32580 28364 32640
rect 110296 32580 110372 32640
rect 21760 32574 21972 32580
rect 21760 32510 21902 32574
rect 21966 32510 21972 32574
rect 1224 32438 1980 32444
rect 1224 32374 1230 32438
rect 1294 32374 1980 32438
rect 1224 32368 1980 32374
rect 21760 32438 21972 32510
rect 21760 32374 21902 32438
rect 21966 32374 21972 32438
rect 21760 32368 21972 32374
rect 22168 32574 22516 32580
rect 22168 32510 22310 32574
rect 22374 32510 22446 32574
rect 22510 32510 22516 32574
rect 22168 32504 22516 32510
rect 22168 32444 22380 32504
rect 22576 32444 22788 32580
rect 22168 32368 22788 32444
rect 22984 32574 23196 32580
rect 22984 32510 22990 32574
rect 23054 32510 23196 32574
rect 22984 32438 23196 32510
rect 22984 32374 22990 32438
rect 23054 32374 23196 32438
rect 22984 32368 23196 32374
rect 23392 32574 23604 32580
rect 23392 32510 23534 32574
rect 23598 32510 23604 32574
rect 23392 32438 23604 32510
rect 23392 32374 23398 32438
rect 23462 32374 23604 32438
rect 23392 32368 23604 32374
rect 28288 32368 28636 32580
rect 110160 32368 110508 32580
rect 115192 32574 115404 32580
rect 115192 32510 115334 32574
rect 115398 32510 115404 32574
rect 115192 32438 115404 32510
rect 115192 32374 115198 32438
rect 115262 32374 115404 32438
rect 115192 32368 115404 32374
rect 115600 32574 115812 32580
rect 115600 32510 115606 32574
rect 115670 32510 115812 32574
rect 115600 32438 115812 32510
rect 115600 32374 115606 32438
rect 115670 32374 115812 32438
rect 115600 32368 115812 32374
rect 116008 32574 116220 32580
rect 116318 32574 116628 32580
rect 116008 32510 116014 32574
rect 116078 32510 116220 32574
rect 116280 32510 116286 32574
rect 116350 32510 116628 32574
rect 116008 32444 116220 32510
rect 116318 32504 116628 32510
rect 116008 32438 116356 32444
rect 116008 32374 116014 32438
rect 116078 32374 116286 32438
rect 116350 32374 116356 32438
rect 116008 32368 116356 32374
rect 116416 32368 116628 32504
rect 116824 32574 117036 32580
rect 116824 32510 116830 32574
rect 116894 32510 117036 32574
rect 116824 32438 117036 32510
rect 116824 32374 116966 32438
rect 117030 32374 117036 32438
rect 116824 32368 117036 32374
rect 136816 32438 137572 32444
rect 136816 32374 137502 32438
rect 137566 32374 137572 32438
rect 136816 32368 137572 32374
rect 1768 32328 1980 32368
rect 1768 32272 1798 32328
rect 1854 32272 1980 32328
rect 22576 32308 22652 32368
rect 1768 32232 1980 32272
rect 14552 32302 14764 32308
rect 14552 32238 14558 32302
rect 14622 32238 14764 32302
rect 14552 32166 14764 32238
rect 22440 32232 22652 32308
rect 28288 32308 28364 32368
rect 110160 32308 110236 32368
rect 136816 32328 137028 32368
rect 22440 32172 22516 32232
rect 14552 32102 14558 32166
rect 14622 32102 14764 32166
rect 14552 32096 14764 32102
rect 21760 32166 21972 32172
rect 21760 32102 21902 32166
rect 21966 32102 21972 32166
rect 21760 31960 21972 32102
rect 22168 32096 22516 32172
rect 22168 32036 22380 32096
rect 22576 32036 22788 32172
rect 22168 32030 22788 32036
rect 22168 31966 22582 32030
rect 22646 31966 22788 32030
rect 22168 31960 22788 31966
rect 22984 32166 23196 32172
rect 22984 32102 22990 32166
rect 23054 32102 23196 32166
rect 22984 32030 23196 32102
rect 22984 31966 23126 32030
rect 23190 31966 23196 32030
rect 22984 31960 23196 31966
rect 23392 32166 23604 32172
rect 23392 32102 23398 32166
rect 23462 32102 23604 32166
rect 23392 32030 23604 32102
rect 28288 32096 28636 32308
rect 110160 32096 110508 32308
rect 136816 32272 136944 32328
rect 137000 32272 137028 32328
rect 136816 32232 137028 32272
rect 115192 32166 115404 32172
rect 115192 32102 115198 32166
rect 115262 32102 115404 32166
rect 28424 32036 28500 32096
rect 110296 32036 110372 32096
rect 23392 31966 23534 32030
rect 23598 31966 23604 32030
rect 23392 31960 23604 31966
rect 21760 31900 21836 31960
rect 14144 31618 14356 31764
rect 21760 31758 21972 31900
rect 28288 31824 28636 32036
rect 110160 31894 110508 32036
rect 115192 32030 115404 32102
rect 115192 31966 115334 32030
rect 115398 31966 115404 32030
rect 115192 31960 115404 31966
rect 115600 32166 115812 32172
rect 115600 32102 115606 32166
rect 115670 32102 115812 32166
rect 115600 32030 115812 32102
rect 115600 31966 115742 32030
rect 115806 31966 115812 32030
rect 115600 31960 115812 31966
rect 116008 32166 116220 32172
rect 116318 32166 116628 32172
rect 116008 32102 116014 32166
rect 116078 32102 116220 32166
rect 116280 32102 116286 32166
rect 116350 32102 116628 32166
rect 116008 31960 116220 32102
rect 116318 32096 116628 32102
rect 116416 31960 116628 32096
rect 116824 32166 117036 32172
rect 116824 32102 116966 32166
rect 117030 32102 117036 32166
rect 116824 31960 117036 32102
rect 116416 31900 116492 31960
rect 110160 31830 110166 31894
rect 110230 31830 110508 31894
rect 110160 31824 110508 31830
rect 116144 31824 116492 31900
rect 116824 31900 116900 31960
rect 28288 31764 28364 31824
rect 110160 31764 110236 31824
rect 116144 31764 116220 31824
rect 21760 31694 21766 31758
rect 21830 31694 21972 31758
rect 21760 31688 21972 31694
rect 22168 31758 22788 31764
rect 22168 31694 22582 31758
rect 22646 31694 22788 31758
rect 22168 31688 22788 31694
rect 14144 31562 14212 31618
rect 14268 31562 14356 31618
rect 14144 31492 14356 31562
rect 22168 31628 22380 31688
rect 22168 31552 22516 31628
rect 22576 31552 22788 31688
rect 22984 31758 23196 31764
rect 22984 31694 23126 31758
rect 23190 31694 23196 31758
rect 22984 31622 23196 31694
rect 22984 31558 22990 31622
rect 23054 31558 23196 31622
rect 22984 31552 23196 31558
rect 23392 31758 23604 31764
rect 23392 31694 23534 31758
rect 23598 31694 23604 31758
rect 23392 31622 23604 31694
rect 23392 31558 23398 31622
rect 23462 31558 23604 31622
rect 23392 31552 23604 31558
rect 0 31416 14356 31492
rect 15152 31549 15218 31552
rect 15486 31549 15552 31552
rect 15152 31547 15552 31549
rect 15152 31491 15157 31547
rect 15213 31491 15491 31547
rect 15547 31491 15552 31547
rect 22304 31492 22380 31552
rect 15152 31489 15552 31491
rect 15152 31486 15218 31489
rect 15486 31486 15552 31489
rect 21760 31486 21972 31492
rect 21760 31422 21766 31486
rect 21830 31422 21972 31486
rect 21760 31144 21972 31422
rect 22168 31144 22380 31492
rect 22440 31492 22516 31552
rect 22440 31416 22788 31492
rect 22576 31214 22788 31416
rect 22576 31150 22582 31214
rect 22646 31150 22788 31214
rect 22576 31144 22788 31150
rect 22984 31350 23196 31356
rect 22984 31286 22990 31350
rect 23054 31286 23196 31350
rect 22984 31144 23196 31286
rect 21896 31084 21972 31144
rect 23120 31084 23196 31144
rect 21760 30942 21972 31084
rect 21760 30878 21766 30942
rect 21830 30878 21972 30942
rect 21760 30872 21972 30878
rect 14552 30806 14764 30812
rect 14552 30742 14694 30806
rect 14758 30742 14764 30806
rect 14552 30676 14764 30742
rect 22168 30736 22380 30948
rect 22576 30942 22788 30948
rect 22576 30878 22582 30942
rect 22646 30878 22788 30942
rect 22576 30812 22788 30878
rect 22440 30736 22788 30812
rect 22984 30736 23196 31084
rect 23392 31350 23604 31356
rect 23392 31286 23398 31350
rect 23462 31286 23604 31350
rect 23392 31144 23604 31286
rect 28288 31280 28636 31764
rect 110160 31622 110508 31764
rect 110160 31558 110166 31622
rect 110230 31558 110508 31622
rect 110160 31280 110508 31558
rect 115192 31758 115404 31764
rect 115192 31694 115334 31758
rect 115398 31694 115404 31758
rect 115192 31622 115404 31694
rect 115192 31558 115198 31622
rect 115262 31558 115404 31622
rect 115192 31552 115404 31558
rect 115600 31758 115812 31764
rect 115600 31694 115742 31758
rect 115806 31694 115812 31758
rect 115600 31622 115812 31694
rect 115600 31558 115606 31622
rect 115670 31558 115812 31622
rect 115600 31552 115812 31558
rect 116008 31758 116356 31764
rect 116008 31694 116150 31758
rect 116214 31694 116286 31758
rect 116350 31694 116356 31758
rect 116008 31688 116356 31694
rect 116416 31758 116628 31764
rect 116416 31694 116422 31758
rect 116486 31694 116628 31758
rect 116008 31552 116220 31688
rect 116416 31628 116628 31694
rect 116824 31758 117036 31900
rect 116824 31694 116830 31758
rect 116894 31694 117036 31758
rect 116824 31688 117036 31694
rect 116280 31552 116628 31628
rect 116280 31492 116356 31552
rect 116008 31416 116356 31492
rect 116416 31486 116628 31492
rect 116416 31422 116422 31486
rect 116486 31422 116628 31486
rect 115192 31350 115404 31356
rect 115192 31286 115198 31350
rect 115262 31286 115404 31350
rect 28560 31220 28636 31280
rect 110296 31220 110372 31280
rect 23392 31084 23468 31144
rect 23392 30736 23604 31084
rect 22168 30676 22244 30736
rect 22440 30676 22516 30736
rect 1224 30670 1980 30676
rect 1224 30606 1230 30670
rect 1294 30648 1980 30670
rect 1294 30606 1798 30648
rect 1224 30600 1798 30606
rect 1768 30592 1798 30600
rect 1854 30592 1980 30648
rect 14552 30670 18572 30676
rect 14552 30606 18502 30670
rect 18566 30606 18572 30670
rect 14552 30600 18572 30606
rect 21760 30670 21972 30676
rect 21760 30606 21766 30670
rect 21830 30606 21972 30670
rect 1768 30464 1980 30592
rect 21760 30534 21972 30606
rect 21760 30470 21902 30534
rect 21966 30470 21972 30534
rect 21760 30464 21972 30470
rect 22168 30600 22516 30676
rect 22576 30676 22652 30736
rect 23120 30676 23196 30736
rect 23528 30676 23604 30736
rect 22168 30464 22380 30600
rect 22576 30540 22788 30676
rect 22478 30534 22788 30540
rect 22440 30470 22446 30534
rect 22510 30470 22718 30534
rect 22782 30470 22788 30534
rect 22478 30464 22788 30470
rect 22984 30328 23196 30676
rect 23120 30268 23196 30328
rect 21760 30262 21972 30268
rect 21760 30198 21902 30262
rect 21966 30198 21972 30262
rect 21760 30126 21972 30198
rect 21760 30062 21766 30126
rect 21830 30062 21972 30126
rect 21760 30056 21972 30062
rect 22168 30262 22516 30268
rect 22168 30198 22446 30262
rect 22510 30198 22516 30262
rect 22168 30192 22516 30198
rect 22576 30262 22788 30268
rect 22576 30198 22718 30262
rect 22782 30198 22788 30262
rect 14144 29918 14356 29996
rect 15152 29991 15218 29994
rect 15406 29991 15472 29994
rect 15152 29989 15472 29991
rect 15152 29933 15157 29989
rect 15213 29933 15411 29989
rect 15467 29933 15472 29989
rect 15152 29931 15472 29933
rect 15152 29928 15218 29931
rect 15406 29928 15472 29931
rect 14144 29862 14212 29918
rect 14268 29862 14356 29918
rect 14144 29860 14356 29862
rect 22168 29920 22380 30192
rect 22576 29920 22788 30198
rect 22984 30126 23196 30268
rect 22984 30062 23126 30126
rect 23190 30062 23196 30126
rect 22984 30056 23196 30062
rect 23392 30328 23604 30676
rect 28288 31078 28636 31220
rect 28288 31014 28294 31078
rect 28358 31014 28636 31078
rect 28288 30806 28636 31014
rect 28288 30742 28294 30806
rect 28358 30742 28636 30806
rect 28288 30670 28636 30742
rect 28288 30606 28294 30670
rect 28358 30606 28636 30670
rect 28288 30600 28636 30606
rect 110160 30670 110508 31220
rect 115192 31144 115404 31286
rect 115328 31084 115404 31144
rect 110160 30606 110438 30670
rect 110502 30606 110508 30670
rect 110160 30600 110508 30606
rect 115192 30736 115404 31084
rect 115600 31350 115812 31356
rect 115600 31286 115606 31350
rect 115670 31286 115812 31350
rect 115600 31144 115812 31286
rect 116008 31214 116220 31416
rect 116008 31150 116014 31214
rect 116078 31150 116220 31214
rect 116008 31144 116220 31150
rect 116416 31144 116628 31422
rect 116824 31486 117036 31492
rect 116824 31422 116830 31486
rect 116894 31422 117036 31486
rect 116824 31144 117036 31422
rect 115600 31084 115676 31144
rect 116824 31084 116900 31144
rect 115600 30736 115812 31084
rect 115192 30676 115268 30736
rect 115736 30676 115812 30736
rect 28288 30398 28636 30404
rect 28288 30334 28294 30398
rect 28358 30334 28636 30398
rect 23392 30268 23468 30328
rect 23392 30126 23604 30268
rect 23392 30062 23398 30126
rect 23462 30062 23604 30126
rect 23392 30056 23604 30062
rect 28288 30262 28636 30334
rect 28288 30198 28294 30262
rect 28358 30198 28636 30262
rect 28288 30056 28636 30198
rect 110160 30398 110508 30404
rect 110160 30334 110438 30398
rect 110502 30334 110508 30398
rect 110160 30262 110508 30334
rect 110160 30198 110166 30262
rect 110230 30198 110508 30262
rect 110160 30056 110508 30198
rect 115192 30328 115404 30676
rect 115600 30328 115812 30676
rect 116008 30942 116220 30948
rect 116008 30878 116014 30942
rect 116078 30878 116220 30942
rect 116008 30736 116220 30878
rect 116416 30736 116628 30948
rect 116824 30942 117036 31084
rect 116824 30878 116830 30942
rect 116894 30878 117036 30942
rect 116824 30872 117036 30878
rect 116008 30676 116084 30736
rect 116416 30676 116492 30736
rect 116008 30600 116628 30676
rect 116008 30540 116220 30600
rect 116008 30534 116356 30540
rect 116008 30470 116286 30534
rect 116350 30470 116356 30534
rect 116008 30464 116356 30470
rect 116416 30464 116628 30600
rect 116824 30670 117036 30676
rect 116824 30606 116830 30670
rect 116894 30606 117036 30670
rect 116824 30534 117036 30606
rect 116824 30470 116966 30534
rect 117030 30470 117036 30534
rect 116824 30464 117036 30470
rect 136816 30648 137028 30676
rect 136816 30592 136944 30648
rect 137000 30592 137028 30648
rect 136816 30540 137028 30592
rect 136816 30534 137572 30540
rect 136816 30470 137502 30534
rect 137566 30470 137572 30534
rect 136816 30464 137572 30470
rect 115192 30268 115268 30328
rect 115736 30268 115812 30328
rect 115192 30126 115404 30268
rect 115192 30062 115334 30126
rect 115398 30062 115404 30126
rect 115192 30056 115404 30062
rect 115600 30126 115812 30268
rect 115600 30062 115742 30126
rect 115806 30062 115812 30126
rect 115600 30056 115812 30062
rect 28288 29996 28364 30056
rect 110160 29996 110236 30056
rect 28288 29990 28636 29996
rect 28288 29926 28294 29990
rect 28358 29926 28636 29990
rect 22168 29860 22244 29920
rect 22576 29860 22652 29920
rect 0 29784 14356 29860
rect 21760 29854 21972 29860
rect 21760 29790 21766 29854
rect 21830 29790 21972 29854
rect 21760 29718 21972 29790
rect 15238 29667 15322 29671
rect 15238 29662 15355 29667
rect 15238 29606 15294 29662
rect 15350 29606 15355 29662
rect 21760 29654 21766 29718
rect 21830 29654 21972 29718
rect 21760 29648 21972 29654
rect 22168 29648 22380 29860
rect 22576 29718 22788 29860
rect 22576 29654 22582 29718
rect 22646 29654 22788 29718
rect 22576 29648 22788 29654
rect 22984 29854 23196 29860
rect 22984 29790 23126 29854
rect 23190 29790 23196 29854
rect 22984 29718 23196 29790
rect 22984 29654 22990 29718
rect 23054 29654 23196 29718
rect 22984 29648 23196 29654
rect 23392 29854 23604 29860
rect 23392 29790 23398 29854
rect 23462 29790 23604 29854
rect 23392 29718 23604 29790
rect 28288 29784 28636 29926
rect 110160 29990 110508 29996
rect 110160 29926 110166 29990
rect 110230 29926 110508 29990
rect 110160 29784 110508 29926
rect 116008 29920 116220 30268
rect 116318 30262 116628 30268
rect 116280 30198 116286 30262
rect 116350 30198 116628 30262
rect 116318 30192 116628 30198
rect 116416 29920 116628 30192
rect 116824 30262 117036 30268
rect 116824 30198 116966 30262
rect 117030 30198 117036 30262
rect 116824 30126 117036 30198
rect 116824 30062 116966 30126
rect 117030 30062 117036 30126
rect 116824 30056 117036 30062
rect 116008 29860 116084 29920
rect 116416 29860 116492 29920
rect 115192 29854 115404 29860
rect 115192 29790 115334 29854
rect 115398 29790 115404 29854
rect 28560 29724 28636 29784
rect 110296 29724 110372 29784
rect 23392 29654 23398 29718
rect 23462 29654 23604 29718
rect 23392 29648 23604 29654
rect 15238 29601 15355 29606
rect 15238 29597 15322 29601
rect 28288 29512 28636 29724
rect 110160 29512 110508 29724
rect 115192 29718 115404 29790
rect 115192 29654 115198 29718
rect 115262 29654 115404 29718
rect 115192 29648 115404 29654
rect 115600 29854 115812 29860
rect 115600 29790 115742 29854
rect 115806 29790 115812 29854
rect 115600 29718 115812 29790
rect 115600 29654 115606 29718
rect 115670 29654 115812 29718
rect 115600 29648 115812 29654
rect 116008 29724 116220 29860
rect 116416 29724 116628 29860
rect 116008 29718 116628 29724
rect 116008 29654 116014 29718
rect 116078 29654 116628 29718
rect 116008 29648 116628 29654
rect 116824 29854 117036 29860
rect 116824 29790 116966 29854
rect 117030 29790 117036 29854
rect 116824 29718 117036 29790
rect 116824 29654 116966 29718
rect 117030 29654 117036 29718
rect 116824 29648 117036 29654
rect 28288 29452 28364 29512
rect 110160 29452 110236 29512
rect 14552 29446 14764 29452
rect 14552 29382 14558 29446
rect 14622 29382 14764 29446
rect 14552 29316 14764 29382
rect 21760 29446 21972 29452
rect 21760 29382 21766 29446
rect 21830 29382 21972 29446
rect 14552 29310 16668 29316
rect 14552 29246 16598 29310
rect 16662 29246 16668 29310
rect 14552 29240 16668 29246
rect 21760 29310 21972 29382
rect 21760 29246 21902 29310
rect 21966 29246 21972 29310
rect 21760 29240 21972 29246
rect 22168 29316 22380 29452
rect 22576 29446 22788 29452
rect 22576 29382 22582 29446
rect 22646 29382 22788 29446
rect 22576 29316 22788 29382
rect 22168 29310 22788 29316
rect 22168 29246 22718 29310
rect 22782 29246 22788 29310
rect 22168 29240 22788 29246
rect 22984 29446 23196 29452
rect 22984 29382 22990 29446
rect 23054 29382 23196 29446
rect 22984 29310 23196 29382
rect 22984 29246 22990 29310
rect 23054 29246 23196 29310
rect 22984 29240 23196 29246
rect 23392 29446 23604 29452
rect 23392 29382 23398 29446
rect 23462 29382 23604 29446
rect 23392 29310 23604 29382
rect 23392 29246 23398 29310
rect 23462 29246 23604 29310
rect 23392 29240 23604 29246
rect 28288 29240 28636 29452
rect 110160 29240 110508 29452
rect 115192 29446 115404 29452
rect 115192 29382 115198 29446
rect 115262 29382 115404 29446
rect 115192 29310 115404 29382
rect 115192 29246 115198 29310
rect 115262 29246 115404 29310
rect 115192 29240 115404 29246
rect 115600 29446 115812 29452
rect 115600 29382 115606 29446
rect 115670 29382 115812 29446
rect 115600 29310 115812 29382
rect 115600 29246 115606 29310
rect 115670 29246 115812 29310
rect 115600 29240 115812 29246
rect 116008 29446 116220 29452
rect 116008 29382 116014 29446
rect 116078 29382 116220 29446
rect 116008 29316 116220 29382
rect 116416 29316 116628 29452
rect 116008 29310 116628 29316
rect 116008 29246 116150 29310
rect 116214 29246 116628 29310
rect 116008 29240 116628 29246
rect 116824 29446 117036 29452
rect 116824 29382 116966 29446
rect 117030 29382 117036 29446
rect 116824 29310 117036 29382
rect 116824 29246 116966 29310
rect 117030 29246 117036 29310
rect 116824 29240 117036 29246
rect 22168 29180 22244 29240
rect 28560 29180 28636 29240
rect 110296 29180 110372 29240
rect 19176 29104 19796 29180
rect 19176 29044 19252 29104
rect 19720 29044 19796 29104
rect 21624 29104 22244 29180
rect 21624 29044 21700 29104
rect 1768 28968 1980 29044
rect 1768 28912 1798 28968
rect 1854 28912 1980 28968
rect 1768 28908 1980 28912
rect 1224 28902 1980 28908
rect 1224 28838 1230 28902
rect 1294 28838 1980 28902
rect 1224 28832 1980 28838
rect 18088 28902 18300 29044
rect 18088 28838 18094 28902
rect 18158 28838 18300 28902
rect 18088 28832 18300 28838
rect 18496 29038 19252 29044
rect 18496 28974 18502 29038
rect 18566 28974 19252 29038
rect 18496 28968 19252 28974
rect 18496 28832 18708 28968
rect 18904 28902 19116 28968
rect 18904 28838 18910 28902
rect 18974 28838 19116 28902
rect 18904 28832 19116 28838
rect 19312 28902 19524 29044
rect 19312 28838 19454 28902
rect 19518 28838 19524 28902
rect 19312 28832 19524 28838
rect 19720 28968 21700 29044
rect 21760 29038 21972 29044
rect 21760 28974 21902 29038
rect 21966 28974 21972 29038
rect 19720 28832 19932 28968
rect 21760 28902 21972 28974
rect 21760 28838 21766 28902
rect 21830 28838 21972 28902
rect 21760 28832 21972 28838
rect 22168 29038 22788 29044
rect 22168 28974 22718 29038
rect 22782 28974 22788 29038
rect 22168 28968 22788 28974
rect 22168 28908 22380 28968
rect 22168 28902 22516 28908
rect 22168 28838 22174 28902
rect 22238 28838 22446 28902
rect 22510 28838 22516 28902
rect 22168 28832 22516 28838
rect 22576 28832 22788 28968
rect 22984 29038 23196 29044
rect 22984 28974 22990 29038
rect 23054 28974 23196 29038
rect 22984 28902 23196 28974
rect 22984 28838 22990 28902
rect 23054 28838 23196 28902
rect 22984 28832 23196 28838
rect 23392 29038 23604 29044
rect 23392 28974 23398 29038
rect 23462 28974 23604 29038
rect 23392 28902 23604 28974
rect 28288 28968 28636 29180
rect 110160 28968 110508 29180
rect 115192 29038 115404 29044
rect 115192 28974 115198 29038
rect 115262 28974 115404 29038
rect 28424 28908 28500 28968
rect 110160 28908 110236 28968
rect 23392 28838 23534 28902
rect 23598 28838 23604 28902
rect 23392 28832 23604 28838
rect 28288 28696 28636 28908
rect 110160 28696 110508 28908
rect 115192 28902 115404 28974
rect 115192 28838 115334 28902
rect 115398 28838 115404 28902
rect 115192 28832 115404 28838
rect 115600 29038 115812 29044
rect 115600 28974 115606 29038
rect 115670 28974 115812 29038
rect 115600 28902 115812 28974
rect 115600 28838 115742 28902
rect 115806 28838 115812 28902
rect 115600 28832 115812 28838
rect 116008 29038 116220 29044
rect 116008 28974 116150 29038
rect 116214 28974 116220 29038
rect 116008 28908 116220 28974
rect 116416 28908 116628 29044
rect 116008 28902 116628 28908
rect 116008 28838 116014 28902
rect 116078 28838 116628 28902
rect 116008 28832 116628 28838
rect 116824 29038 117036 29044
rect 116824 28974 116966 29038
rect 117030 28974 117036 29038
rect 116824 28902 117036 28974
rect 116824 28838 116830 28902
rect 116894 28838 117036 28902
rect 116824 28832 117036 28838
rect 118864 28902 119076 29044
rect 118864 28838 119006 28902
rect 119070 28838 119076 28902
rect 118864 28832 119076 28838
rect 119272 28902 119484 29044
rect 119272 28838 119278 28902
rect 119342 28838 119484 28902
rect 119272 28832 119484 28838
rect 119680 28968 120300 29044
rect 119680 28832 119892 28968
rect 120088 28908 120300 28968
rect 119990 28902 120300 28908
rect 119952 28838 119958 28902
rect 120022 28838 120300 28902
rect 119990 28832 120300 28838
rect 120496 28902 120708 29044
rect 120496 28838 120502 28902
rect 120566 28838 120708 28902
rect 120496 28832 120708 28838
rect 136816 29038 137572 29044
rect 136816 28974 137502 29038
rect 137566 28974 137572 29038
rect 136816 28968 137572 28974
rect 136816 28912 136944 28968
rect 137000 28912 137028 28968
rect 136816 28832 137028 28912
rect 28424 28636 28500 28696
rect 110296 28636 110372 28696
rect 21760 28630 21972 28636
rect 21760 28566 21766 28630
rect 21830 28566 21972 28630
rect 21760 28494 21972 28566
rect 21760 28430 21766 28494
rect 21830 28430 21972 28494
rect 21760 28424 21972 28430
rect 22168 28630 22380 28636
rect 22478 28630 22788 28636
rect 22168 28566 22174 28630
rect 22238 28566 22380 28630
rect 22440 28566 22446 28630
rect 22510 28566 22788 28630
rect 22168 28424 22380 28566
rect 22478 28560 22788 28566
rect 22576 28424 22788 28560
rect 22984 28630 23196 28636
rect 22984 28566 22990 28630
rect 23054 28566 23196 28630
rect 22984 28494 23196 28566
rect 22984 28430 22990 28494
rect 23054 28430 23196 28494
rect 22984 28424 23196 28430
rect 23392 28630 23604 28636
rect 23392 28566 23534 28630
rect 23598 28566 23604 28630
rect 23392 28494 23604 28566
rect 23392 28430 23398 28494
rect 23462 28430 23604 28494
rect 23392 28424 23604 28430
rect 28288 28424 28636 28636
rect 110160 28424 110508 28636
rect 115192 28630 115404 28636
rect 115192 28566 115334 28630
rect 115398 28566 115404 28630
rect 115192 28494 115404 28566
rect 115192 28430 115334 28494
rect 115398 28430 115404 28494
rect 115192 28424 115404 28430
rect 115600 28630 115812 28636
rect 115600 28566 115742 28630
rect 115806 28566 115812 28630
rect 115600 28494 115812 28566
rect 115600 28430 115742 28494
rect 115806 28430 115812 28494
rect 115600 28424 115812 28430
rect 116008 28630 116220 28636
rect 116008 28566 116014 28630
rect 116078 28566 116220 28630
rect 116008 28500 116220 28566
rect 116416 28500 116628 28636
rect 116008 28424 116628 28500
rect 116824 28630 117036 28636
rect 116824 28566 116830 28630
rect 116894 28566 117036 28630
rect 116824 28494 117036 28566
rect 116824 28430 116966 28494
rect 117030 28430 117036 28494
rect 116824 28424 117036 28430
rect 22576 28364 22652 28424
rect 19176 28288 19796 28364
rect 19176 28228 19252 28288
rect 19720 28228 19796 28288
rect 22304 28288 22652 28364
rect 28288 28364 28364 28424
rect 110296 28364 110372 28424
rect 116144 28364 116220 28424
rect 22304 28228 22380 28288
rect 18088 28222 18300 28228
rect 18088 28158 18094 28222
rect 18158 28158 18300 28222
rect 18088 28086 18300 28158
rect 18088 28022 18094 28086
rect 18158 28022 18300 28086
rect 18088 28016 18300 28022
rect 18496 28222 19252 28228
rect 18496 28158 18910 28222
rect 18974 28158 19252 28222
rect 18496 28152 19252 28158
rect 19312 28222 19524 28228
rect 19312 28158 19454 28222
rect 19518 28158 19524 28222
rect 18496 28016 18708 28152
rect 18904 28086 19116 28152
rect 18904 28022 19046 28086
rect 19110 28022 19116 28086
rect 18904 28016 19116 28022
rect 19312 28086 19524 28158
rect 19312 28022 19454 28086
rect 19518 28022 19524 28086
rect 19312 28016 19524 28022
rect 19720 28086 19932 28228
rect 19720 28022 19726 28086
rect 19790 28022 19932 28086
rect 19720 28016 19932 28022
rect 21760 28222 21972 28228
rect 21760 28158 21766 28222
rect 21830 28158 21972 28222
rect 21760 28016 21972 28158
rect 22168 28152 22788 28228
rect 22168 28086 22380 28152
rect 22168 28022 22310 28086
rect 22374 28022 22380 28086
rect 22168 28016 22380 28022
rect 22576 28086 22788 28152
rect 22576 28022 22718 28086
rect 22782 28022 22788 28086
rect 22576 28016 22788 28022
rect 22984 28222 23196 28228
rect 22984 28158 22990 28222
rect 23054 28158 23196 28222
rect 22984 28086 23196 28158
rect 22984 28022 22990 28086
rect 23054 28022 23196 28086
rect 22984 28016 23196 28022
rect 23392 28222 23604 28228
rect 23392 28158 23398 28222
rect 23462 28158 23604 28222
rect 23392 28086 23604 28158
rect 28288 28152 28636 28364
rect 28560 28092 28636 28152
rect 23392 28022 23398 28086
rect 23462 28022 23604 28086
rect 23392 28016 23604 28022
rect 21896 27956 21972 28016
rect 18360 27678 19388 27684
rect 18360 27614 19318 27678
rect 19382 27614 19388 27678
rect 18360 27608 19388 27614
rect 21760 27608 21972 27956
rect 28288 27950 28636 28092
rect 28288 27886 28294 27950
rect 28358 27886 28636 27950
rect 28288 27880 28636 27886
rect 110160 28152 110508 28364
rect 116144 28288 116492 28364
rect 116416 28228 116492 28288
rect 119816 28288 120164 28364
rect 119816 28228 119892 28288
rect 120088 28228 120164 28288
rect 115192 28222 115404 28228
rect 115192 28158 115334 28222
rect 115398 28158 115404 28222
rect 110160 28092 110236 28152
rect 110160 27880 110508 28092
rect 115192 28086 115404 28158
rect 115192 28022 115334 28086
rect 115398 28022 115404 28086
rect 115192 28016 115404 28022
rect 115600 28222 115812 28228
rect 115600 28158 115742 28222
rect 115806 28158 115812 28222
rect 115600 28086 115812 28158
rect 115600 28022 115742 28086
rect 115806 28022 115812 28086
rect 115600 28016 115812 28022
rect 116008 28092 116220 28228
rect 116416 28092 116628 28228
rect 116008 28086 116628 28092
rect 116008 28022 116014 28086
rect 116078 28022 116628 28086
rect 116008 28016 116628 28022
rect 116824 28222 117036 28228
rect 116824 28158 116966 28222
rect 117030 28158 117036 28222
rect 116824 28016 117036 28158
rect 118864 28222 119076 28228
rect 118864 28158 119006 28222
rect 119070 28158 119076 28222
rect 118864 28086 119076 28158
rect 118864 28022 119006 28086
rect 119070 28022 119076 28086
rect 118864 28016 119076 28022
rect 119272 28222 119484 28228
rect 119272 28158 119278 28222
rect 119342 28158 119484 28222
rect 119272 28092 119484 28158
rect 119680 28222 120028 28228
rect 119680 28158 119958 28222
rect 120022 28158 120028 28222
rect 119680 28152 120028 28158
rect 119680 28092 119892 28152
rect 119272 28086 119620 28092
rect 119272 28022 119414 28086
rect 119478 28022 119620 28086
rect 119272 28016 119620 28022
rect 119680 28086 120028 28092
rect 119680 28022 119958 28086
rect 120022 28022 120028 28086
rect 119680 28016 120028 28022
rect 120088 28016 120300 28228
rect 120496 28222 120708 28228
rect 120496 28158 120502 28222
rect 120566 28158 120708 28222
rect 120496 28086 120708 28158
rect 120496 28022 120638 28086
rect 120702 28022 120708 28086
rect 120496 28016 120708 28022
rect 116960 27956 117036 28016
rect 28288 27820 28364 27880
rect 110296 27820 110372 27880
rect 22168 27814 22380 27820
rect 22168 27750 22310 27814
rect 22374 27750 22380 27814
rect 22168 27608 22380 27750
rect 22576 27814 22788 27820
rect 22576 27750 22718 27814
rect 22782 27750 22788 27814
rect 22576 27608 22788 27750
rect 22984 27814 23196 27820
rect 22984 27750 22990 27814
rect 23054 27750 23196 27814
rect 22984 27678 23196 27750
rect 22984 27614 23126 27678
rect 23190 27614 23196 27678
rect 22984 27608 23196 27614
rect 23392 27814 23604 27820
rect 23392 27750 23398 27814
rect 23462 27750 23604 27814
rect 23392 27678 23604 27750
rect 23392 27614 23534 27678
rect 23598 27614 23604 27678
rect 23392 27608 23604 27614
rect 28288 27678 28636 27820
rect 28288 27614 28294 27678
rect 28358 27614 28636 27678
rect 18360 27548 18436 27608
rect 21896 27548 21972 27608
rect 22304 27548 22380 27608
rect 22712 27548 22788 27608
rect 18088 27542 18436 27548
rect 18088 27478 18094 27542
rect 18158 27478 18436 27542
rect 18088 27472 18436 27478
rect 1224 27406 1980 27412
rect 1224 27342 1230 27406
rect 1294 27342 1980 27406
rect 1224 27336 1980 27342
rect 1768 27288 1980 27336
rect 1768 27232 1798 27288
rect 1854 27232 1980 27288
rect 1768 27200 1980 27232
rect 18088 27270 18300 27472
rect 18088 27206 18094 27270
rect 18158 27206 18300 27270
rect 18088 27200 18300 27206
rect 18496 27276 18708 27548
rect 18904 27542 19116 27548
rect 18904 27478 19046 27542
rect 19110 27478 19116 27542
rect 18904 27276 19116 27478
rect 18496 27270 19116 27276
rect 18496 27206 18502 27270
rect 18566 27206 19116 27270
rect 18496 27200 19116 27206
rect 19312 27406 19524 27412
rect 19312 27342 19318 27406
rect 19382 27342 19454 27406
rect 19518 27342 19524 27406
rect 19312 27270 19524 27342
rect 19312 27206 19318 27270
rect 19382 27206 19524 27270
rect 19312 27200 19524 27206
rect 19720 27406 19932 27412
rect 19720 27342 19726 27406
rect 19790 27342 19932 27406
rect 19720 27270 19932 27342
rect 19720 27206 19862 27270
rect 19926 27206 19932 27270
rect 19720 27200 19932 27206
rect 21760 27200 21972 27548
rect 22168 27270 22380 27548
rect 22168 27206 22310 27270
rect 22374 27206 22380 27270
rect 22168 27200 22380 27206
rect 22576 27200 22788 27548
rect 22984 27406 23196 27412
rect 22984 27342 23126 27406
rect 23190 27342 23196 27406
rect 22984 27200 23196 27342
rect 23392 27406 23604 27412
rect 23392 27342 23534 27406
rect 23598 27342 23604 27406
rect 23392 27200 23604 27342
rect 28288 27406 28636 27614
rect 28288 27342 28430 27406
rect 28494 27342 28636 27406
rect 28288 27336 28636 27342
rect 110160 27406 110508 27820
rect 115192 27814 115404 27820
rect 115192 27750 115334 27814
rect 115398 27750 115404 27814
rect 115192 27678 115404 27750
rect 115192 27614 115334 27678
rect 115398 27614 115404 27678
rect 115192 27608 115404 27614
rect 115600 27814 115812 27820
rect 115600 27750 115742 27814
rect 115806 27750 115812 27814
rect 115600 27678 115812 27750
rect 115600 27614 115742 27678
rect 115806 27614 115812 27678
rect 115600 27608 115812 27614
rect 116008 27814 116220 27820
rect 116008 27750 116014 27814
rect 116078 27750 116220 27814
rect 116008 27608 116220 27750
rect 116416 27608 116628 27820
rect 116824 27608 117036 27956
rect 119544 27956 119620 28016
rect 120496 27956 120572 28016
rect 119544 27880 120572 27956
rect 116008 27548 116084 27608
rect 116416 27548 116492 27608
rect 116824 27548 116900 27608
rect 116008 27412 116220 27548
rect 116416 27412 116628 27548
rect 110160 27342 110166 27406
rect 110230 27342 110508 27406
rect 110160 27336 110508 27342
rect 110432 27276 110508 27336
rect 18632 27140 18708 27200
rect 21896 27140 21972 27200
rect 18632 27134 18980 27140
rect 18632 27070 18910 27134
rect 18974 27070 18980 27134
rect 18632 27064 18980 27070
rect 21760 26998 21972 27140
rect 22984 27140 23060 27200
rect 23392 27140 23468 27200
rect 21760 26934 21902 26998
rect 21966 26934 21972 26998
rect 21760 26928 21972 26934
rect 22168 26998 22380 27004
rect 22168 26934 22310 26998
rect 22374 26934 22380 26998
rect 22168 26868 22380 26934
rect 16864 26792 18164 26868
rect 22168 26792 22516 26868
rect 22576 26792 22788 27004
rect 16864 26732 16940 26792
rect 18088 26732 18164 26792
rect 22304 26732 22380 26792
rect 16592 26726 16940 26732
rect 16592 26662 16598 26726
rect 16662 26662 16940 26726
rect 16592 26656 16940 26662
rect 16592 26384 16804 26656
rect 17000 26460 17212 26732
rect 18088 26726 18300 26732
rect 18088 26662 18094 26726
rect 18158 26662 18300 26726
rect 18088 26520 18300 26662
rect 18496 26726 19116 26732
rect 18496 26662 18910 26726
rect 18974 26662 19116 26726
rect 18496 26656 19116 26662
rect 18496 26520 18708 26656
rect 18904 26520 19116 26656
rect 19312 26726 19524 26732
rect 19312 26662 19318 26726
rect 19382 26662 19524 26726
rect 17000 26454 18572 26460
rect 17000 26390 18502 26454
rect 18566 26390 18572 26454
rect 17000 26384 18572 26390
rect 19312 26454 19524 26662
rect 19312 26390 19454 26454
rect 19518 26390 19524 26454
rect 19312 26384 19524 26390
rect 19720 26726 19932 26732
rect 19720 26662 19862 26726
rect 19926 26662 19932 26726
rect 19720 26454 19932 26662
rect 21760 26726 21972 26732
rect 21760 26662 21902 26726
rect 21966 26662 21972 26726
rect 21760 26590 21972 26662
rect 21760 26526 21766 26590
rect 21830 26526 21972 26590
rect 21760 26520 21972 26526
rect 22168 26520 22380 26732
rect 22440 26732 22516 26792
rect 22712 26732 22788 26792
rect 22440 26656 22788 26732
rect 22576 26590 22788 26656
rect 22576 26526 22718 26590
rect 22782 26526 22788 26590
rect 22576 26520 22788 26526
rect 22984 26792 23196 27140
rect 23392 26792 23604 27140
rect 22984 26732 23060 26792
rect 23528 26732 23604 26792
rect 19720 26390 19726 26454
rect 19790 26390 19932 26454
rect 19720 26384 19932 26390
rect 22984 26384 23196 26732
rect 23392 26384 23604 26732
rect 28288 27134 28636 27276
rect 28288 27070 28430 27134
rect 28494 27070 28566 27134
rect 28630 27070 28636 27134
rect 28288 26862 28636 27070
rect 28288 26798 28566 26862
rect 28630 26798 28636 26862
rect 28288 26726 28636 26798
rect 28288 26662 28294 26726
rect 28358 26662 28636 26726
rect 28288 26656 28636 26662
rect 110160 27134 110508 27276
rect 110160 27070 110166 27134
rect 110230 27070 110302 27134
rect 110366 27070 110508 27134
rect 110160 26862 110508 27070
rect 110160 26798 110302 26862
rect 110366 26798 110508 26862
rect 110160 26726 110508 26798
rect 115192 27406 115404 27412
rect 115192 27342 115334 27406
rect 115398 27342 115404 27406
rect 115192 27200 115404 27342
rect 115600 27406 115812 27412
rect 115600 27342 115742 27406
rect 115806 27342 115812 27406
rect 115600 27200 115812 27342
rect 116008 27336 116628 27412
rect 116008 27200 116220 27336
rect 116416 27270 116628 27336
rect 116416 27206 116558 27270
rect 116622 27206 116628 27270
rect 116416 27200 116628 27206
rect 116824 27200 117036 27548
rect 119136 27472 119892 27548
rect 119990 27542 120300 27548
rect 119952 27478 119958 27542
rect 120022 27478 120300 27542
rect 119990 27472 120300 27478
rect 119136 27412 119212 27472
rect 118864 27406 119212 27412
rect 118864 27342 119006 27406
rect 119070 27342 119212 27406
rect 118864 27336 119212 27342
rect 119272 27406 119484 27412
rect 119272 27342 119414 27406
rect 119478 27342 119484 27406
rect 118864 27200 119076 27336
rect 119272 27270 119484 27342
rect 119272 27206 119278 27270
rect 119342 27206 119484 27270
rect 119272 27200 119484 27206
rect 119680 27276 119892 27472
rect 120088 27276 120300 27472
rect 119680 27270 120300 27276
rect 119680 27206 120094 27270
rect 120158 27206 120300 27270
rect 119680 27200 120300 27206
rect 120496 27542 120708 27548
rect 120496 27478 120638 27542
rect 120702 27478 120708 27542
rect 120496 27270 120708 27478
rect 120496 27206 120502 27270
rect 120566 27206 120708 27270
rect 120496 27200 120708 27206
rect 136816 27288 137028 27412
rect 136816 27232 136944 27288
rect 137000 27276 137028 27288
rect 137000 27270 137572 27276
rect 137000 27232 137502 27270
rect 136816 27206 137502 27232
rect 137566 27206 137572 27270
rect 136816 27200 137572 27206
rect 115192 27140 115268 27200
rect 115600 27140 115676 27200
rect 116824 27140 116900 27200
rect 115192 26792 115404 27140
rect 115328 26732 115404 26792
rect 110160 26662 110302 26726
rect 110366 26662 110508 26726
rect 110160 26656 110508 26662
rect 28288 26454 28636 26460
rect 28288 26390 28294 26454
rect 28358 26390 28636 26454
rect 22984 26324 23060 26384
rect 23392 26324 23468 26384
rect 21760 26318 21972 26324
rect 21760 26254 21766 26318
rect 21830 26254 21972 26318
rect 21760 26182 21972 26254
rect 21760 26118 21902 26182
rect 21966 26118 21972 26182
rect 21760 26112 21972 26118
rect 22168 26052 22380 26324
rect 22576 26318 22788 26324
rect 22576 26254 22718 26318
rect 22782 26254 22788 26318
rect 3128 25976 4156 26052
rect 22168 26046 22516 26052
rect 22168 25982 22446 26046
rect 22510 25982 22516 26046
rect 22168 25976 22516 25982
rect 22576 25976 22788 26254
rect 22984 26182 23196 26324
rect 22984 26118 22990 26182
rect 23054 26118 23196 26182
rect 22984 26112 23196 26118
rect 23392 26182 23604 26324
rect 23392 26118 23398 26182
rect 23462 26118 23604 26182
rect 23392 26112 23604 26118
rect 28288 26112 28636 26390
rect 110160 26454 110508 26460
rect 110160 26390 110302 26454
rect 110366 26390 110508 26454
rect 110160 26318 110508 26390
rect 110160 26254 110438 26318
rect 110502 26254 110508 26318
rect 110160 26112 110508 26254
rect 115192 26384 115404 26732
rect 115600 26792 115812 27140
rect 116008 26868 116220 27004
rect 116416 26998 116628 27004
rect 116416 26934 116558 26998
rect 116622 26934 116628 26998
rect 116008 26792 116356 26868
rect 116416 26792 116628 26934
rect 116824 26998 117036 27140
rect 116824 26934 116830 26998
rect 116894 26934 117036 26998
rect 116824 26928 117036 26934
rect 115600 26732 115676 26792
rect 116008 26732 116084 26792
rect 116280 26732 116356 26792
rect 116552 26732 116628 26792
rect 119136 26792 119756 26868
rect 119136 26732 119212 26792
rect 119680 26732 119756 26792
rect 121448 26792 122068 26868
rect 121448 26732 121524 26792
rect 121992 26732 122068 26792
rect 115600 26384 115812 26732
rect 116008 26590 116220 26732
rect 116280 26656 116628 26732
rect 116008 26526 116014 26590
rect 116078 26526 116220 26590
rect 116008 26520 116220 26526
rect 116416 26520 116628 26656
rect 116824 26726 117036 26732
rect 116824 26662 116830 26726
rect 116894 26662 117036 26726
rect 116824 26590 117036 26662
rect 116824 26526 116830 26590
rect 116894 26526 117036 26590
rect 116824 26520 117036 26526
rect 118864 26656 119212 26732
rect 119272 26726 119484 26732
rect 119272 26662 119278 26726
rect 119342 26662 119484 26726
rect 118864 26384 119076 26656
rect 119272 26454 119484 26662
rect 119680 26726 120300 26732
rect 119680 26662 120094 26726
rect 120158 26662 120300 26726
rect 119680 26656 120300 26662
rect 119680 26590 119892 26656
rect 119680 26526 119822 26590
rect 119886 26526 119892 26590
rect 119680 26520 119892 26526
rect 120088 26596 120300 26656
rect 120496 26726 121524 26732
rect 120496 26662 120502 26726
rect 120566 26662 121524 26726
rect 120496 26656 121524 26662
rect 120088 26520 120436 26596
rect 120496 26520 120708 26656
rect 119272 26390 119414 26454
rect 119478 26390 119484 26454
rect 119272 26384 119484 26390
rect 120360 26460 120436 26520
rect 121584 26460 121796 26732
rect 120360 26384 121796 26460
rect 121992 26384 122204 26732
rect 115192 26324 115268 26384
rect 115736 26324 115812 26384
rect 115192 26182 115404 26324
rect 115192 26118 115198 26182
rect 115262 26118 115404 26182
rect 115192 26112 115404 26118
rect 115600 26182 115812 26324
rect 115600 26118 115606 26182
rect 115670 26118 115812 26182
rect 115600 26112 115812 26118
rect 116008 26318 116628 26324
rect 116008 26254 116014 26318
rect 116078 26254 116628 26318
rect 116008 26248 116628 26254
rect 28288 26052 28364 26112
rect 110432 26052 110508 26112
rect 3128 25916 3340 25976
rect 3944 25916 4156 25976
rect 22576 25916 22652 25976
rect 544 25910 3340 25916
rect 3846 25910 4156 25916
rect 544 25846 550 25910
rect 614 25846 3340 25910
rect 3808 25846 3814 25910
rect 3878 25846 4156 25910
rect 544 25840 3340 25846
rect 3846 25840 4156 25846
rect 21760 25910 21972 25916
rect 21760 25846 21902 25910
rect 21966 25846 21972 25910
rect 21760 25774 21972 25846
rect 21760 25710 21902 25774
rect 21966 25710 21972 25774
rect 21760 25704 21972 25710
rect 22168 25910 22788 25916
rect 22168 25846 22582 25910
rect 22646 25846 22788 25910
rect 22168 25840 22788 25846
rect 22168 25780 22380 25840
rect 22168 25774 22516 25780
rect 22168 25710 22446 25774
rect 22510 25710 22516 25774
rect 22168 25704 22516 25710
rect 22576 25704 22788 25840
rect 22984 25910 23196 25916
rect 22984 25846 22990 25910
rect 23054 25846 23196 25910
rect 22984 25774 23196 25846
rect 22984 25710 23126 25774
rect 23190 25710 23196 25774
rect 22984 25704 23196 25710
rect 23392 25910 23604 25916
rect 23392 25846 23398 25910
rect 23462 25846 23604 25910
rect 23392 25774 23604 25846
rect 28288 25910 28636 26052
rect 28288 25846 28566 25910
rect 28630 25846 28636 25910
rect 28288 25840 28636 25846
rect 110160 26046 110508 26052
rect 110160 25982 110438 26046
rect 110502 25982 110508 26046
rect 110160 25840 110508 25982
rect 116008 25976 116220 26248
rect 116416 25976 116628 26248
rect 116824 26318 117036 26324
rect 116824 26254 116830 26318
rect 116894 26254 117036 26318
rect 116824 26182 117036 26254
rect 116824 26118 116966 26182
rect 117030 26118 117036 26182
rect 116824 26112 117036 26118
rect 116552 25916 116628 25976
rect 115192 25910 115404 25916
rect 115192 25846 115198 25910
rect 115262 25846 115404 25910
rect 28560 25780 28636 25840
rect 110296 25780 110372 25840
rect 23392 25710 23534 25774
rect 23598 25710 23604 25774
rect 23392 25704 23604 25710
rect 1224 25638 1980 25644
rect 1224 25574 1230 25638
rect 1294 25608 1980 25638
rect 1294 25574 1798 25608
rect 1224 25568 1798 25574
rect 1768 25552 1798 25568
rect 1854 25552 1980 25608
rect 1768 25432 1980 25552
rect 21760 25502 21972 25508
rect 21760 25438 21902 25502
rect 21966 25438 21972 25502
rect 21760 25372 21972 25438
rect 19622 25366 21972 25372
rect 2540 25365 2606 25366
rect 2498 25301 2541 25365
rect 2605 25301 2648 25365
rect 19584 25302 19590 25366
rect 19654 25302 21766 25366
rect 21830 25302 21972 25366
rect 2540 25300 2606 25301
rect 19622 25296 21972 25302
rect 22168 25366 22380 25508
rect 22478 25502 22788 25508
rect 22440 25438 22446 25502
rect 22510 25438 22788 25502
rect 22478 25432 22788 25438
rect 22168 25302 22174 25366
rect 22238 25302 22380 25366
rect 22168 25296 22380 25302
rect 22576 25366 22788 25432
rect 22576 25302 22718 25366
rect 22782 25302 22788 25366
rect 22576 25296 22788 25302
rect 22984 25502 23196 25508
rect 22984 25438 23126 25502
rect 23190 25438 23196 25502
rect 22984 25366 23196 25438
rect 22984 25302 22990 25366
rect 23054 25302 23196 25366
rect 22984 25296 23196 25302
rect 23392 25502 23604 25508
rect 23392 25438 23534 25502
rect 23598 25438 23604 25502
rect 23392 25366 23604 25438
rect 23392 25302 23534 25366
rect 23598 25302 23604 25366
rect 23392 25296 23604 25302
rect 28288 25502 28636 25780
rect 28288 25438 28566 25502
rect 28630 25438 28636 25502
rect 28288 25296 28636 25438
rect 110160 25296 110508 25780
rect 115192 25774 115404 25846
rect 115192 25710 115334 25774
rect 115398 25710 115404 25774
rect 115192 25704 115404 25710
rect 115600 25910 115812 25916
rect 115600 25846 115606 25910
rect 115670 25846 115812 25910
rect 115600 25774 115812 25846
rect 115600 25710 115742 25774
rect 115806 25710 115812 25774
rect 115600 25704 115812 25710
rect 116008 25840 116628 25916
rect 116008 25704 116220 25840
rect 116416 25780 116628 25840
rect 116318 25774 116628 25780
rect 116280 25710 116286 25774
rect 116350 25710 116422 25774
rect 116486 25710 116628 25774
rect 116318 25704 116628 25710
rect 116824 25910 117036 25916
rect 116824 25846 116966 25910
rect 117030 25846 117036 25910
rect 116824 25780 117036 25846
rect 116824 25774 119348 25780
rect 116824 25710 116966 25774
rect 117030 25710 119278 25774
rect 119342 25710 119348 25774
rect 116824 25704 119348 25710
rect 136816 25638 137572 25644
rect 136816 25608 137502 25638
rect 136816 25552 136944 25608
rect 137000 25574 137502 25608
rect 137566 25574 137572 25638
rect 137000 25568 137572 25574
rect 137000 25552 137028 25568
rect 115192 25502 115404 25508
rect 115192 25438 115334 25502
rect 115398 25438 115404 25502
rect 115192 25366 115404 25438
rect 115192 25302 115198 25366
rect 115262 25302 115404 25366
rect 115192 25296 115404 25302
rect 115600 25502 115812 25508
rect 115600 25438 115742 25502
rect 115806 25438 115812 25502
rect 115600 25366 115812 25438
rect 115600 25302 115742 25366
rect 115806 25302 115812 25366
rect 115600 25296 115812 25302
rect 116008 25502 116356 25508
rect 116008 25438 116286 25502
rect 116350 25438 116356 25502
rect 116008 25432 116356 25438
rect 116416 25502 116628 25508
rect 116416 25438 116422 25502
rect 116486 25438 116628 25502
rect 116008 25296 116220 25432
rect 116416 25366 116628 25438
rect 116416 25302 116558 25366
rect 116622 25302 116628 25366
rect 116416 25296 116628 25302
rect 116824 25502 117036 25508
rect 116824 25438 116966 25502
rect 117030 25438 117036 25502
rect 116824 25366 117036 25438
rect 136816 25432 137028 25552
rect 116824 25302 116966 25366
rect 117030 25302 117036 25366
rect 116824 25296 117036 25302
rect 28424 25236 28500 25296
rect 110296 25236 110372 25296
rect 18088 24958 18300 25100
rect 18088 24894 18230 24958
rect 18294 24894 18300 24958
rect 18088 24888 18300 24894
rect 18496 25024 19116 25100
rect 18496 24888 18708 25024
rect 18904 24964 19116 25024
rect 19312 25094 19660 25100
rect 19312 25030 19454 25094
rect 19518 25030 19590 25094
rect 19654 25030 19660 25094
rect 19312 25024 19660 25030
rect 19720 25094 19932 25100
rect 19720 25030 19726 25094
rect 19790 25030 19932 25094
rect 18904 24958 19252 24964
rect 18904 24894 18910 24958
rect 18974 24894 19252 24958
rect 18904 24888 19252 24894
rect 19312 24958 19524 25024
rect 19312 24894 19318 24958
rect 19382 24894 19524 24958
rect 19312 24888 19524 24894
rect 19720 24888 19932 25030
rect 21760 25094 21972 25100
rect 21760 25030 21766 25094
rect 21830 25030 21972 25094
rect 21760 24958 21972 25030
rect 21760 24894 21902 24958
rect 21966 24894 21972 24958
rect 21760 24888 21972 24894
rect 22168 25094 22380 25100
rect 22168 25030 22174 25094
rect 22238 25030 22380 25094
rect 22168 24964 22380 25030
rect 22576 25094 22788 25100
rect 22576 25030 22718 25094
rect 22782 25030 22788 25094
rect 22576 24964 22788 25030
rect 22168 24958 22788 24964
rect 22168 24894 22174 24958
rect 22238 24894 22788 24958
rect 22168 24888 22788 24894
rect 22984 25094 23196 25100
rect 22984 25030 22990 25094
rect 23054 25030 23196 25094
rect 22984 24958 23196 25030
rect 22984 24894 23126 24958
rect 23190 24894 23196 24958
rect 22984 24888 23196 24894
rect 23392 25094 23604 25100
rect 23392 25030 23534 25094
rect 23598 25030 23604 25094
rect 23392 24958 23604 25030
rect 28288 25024 28636 25236
rect 110160 25024 110508 25236
rect 115192 25094 115404 25100
rect 115192 25030 115198 25094
rect 115262 25030 115404 25094
rect 28560 24964 28636 25024
rect 110296 24964 110372 25024
rect 23392 24894 23398 24958
rect 23462 24894 23604 24958
rect 23392 24888 23604 24894
rect 19176 24828 19252 24888
rect 19720 24828 19796 24888
rect 19176 24752 19796 24828
rect 22304 24828 22380 24888
rect 22304 24752 22652 24828
rect 28288 24752 28636 24964
rect 110160 24752 110508 24964
rect 115192 24958 115404 25030
rect 115192 24894 115198 24958
rect 115262 24894 115404 24958
rect 115192 24888 115404 24894
rect 115600 25094 115812 25100
rect 115600 25030 115742 25094
rect 115806 25030 115812 25094
rect 115600 24958 115812 25030
rect 115600 24894 115606 24958
rect 115670 24894 115812 24958
rect 115600 24888 115812 24894
rect 116008 24964 116220 25100
rect 116416 25094 116628 25100
rect 116416 25030 116558 25094
rect 116622 25030 116628 25094
rect 116416 24964 116628 25030
rect 116008 24958 116628 24964
rect 116008 24894 116150 24958
rect 116214 24894 116628 24958
rect 116008 24888 116628 24894
rect 116824 25094 117036 25100
rect 116824 25030 116966 25094
rect 117030 25030 117036 25094
rect 116824 24958 117036 25030
rect 116824 24894 116966 24958
rect 117030 24894 117036 24958
rect 116824 24888 117036 24894
rect 118864 24958 119076 25100
rect 118864 24894 119006 24958
rect 119070 24894 119076 24958
rect 118864 24888 119076 24894
rect 119272 25094 119484 25100
rect 119272 25030 119278 25094
rect 119342 25030 119414 25094
rect 119478 25030 119484 25094
rect 119272 24958 119484 25030
rect 119272 24894 119414 24958
rect 119478 24894 119484 24958
rect 119272 24888 119484 24894
rect 119680 25094 120300 25100
rect 119680 25030 119822 25094
rect 119886 25030 120300 25094
rect 119680 25024 120300 25030
rect 119680 24888 119892 25024
rect 120088 24958 120300 25024
rect 120088 24894 120094 24958
rect 120158 24894 120300 24958
rect 120088 24888 120300 24894
rect 120496 24958 120708 25100
rect 120496 24894 120638 24958
rect 120702 24894 120708 24958
rect 120496 24888 120708 24894
rect 22576 24692 22652 24752
rect 28424 24692 28500 24752
rect 110432 24692 110508 24752
rect 3128 24556 3340 24692
rect 3944 24556 4156 24692
rect 2350 24550 4156 24556
rect 2312 24486 2318 24550
rect 2382 24486 4156 24550
rect 2350 24480 4156 24486
rect 21760 24686 21972 24692
rect 21760 24622 21902 24686
rect 21966 24622 21972 24686
rect 21760 24550 21972 24622
rect 21760 24486 21766 24550
rect 21830 24486 21972 24550
rect 21760 24480 21972 24486
rect 22168 24686 22380 24692
rect 22168 24622 22174 24686
rect 22238 24622 22380 24686
rect 22168 24550 22380 24622
rect 22168 24486 22310 24550
rect 22374 24486 22380 24550
rect 22168 24480 22380 24486
rect 22576 24480 22788 24692
rect 22984 24686 23196 24692
rect 22984 24622 23126 24686
rect 23190 24622 23196 24686
rect 22984 24550 23196 24622
rect 22984 24486 23126 24550
rect 23190 24486 23196 24550
rect 22984 24480 23196 24486
rect 23392 24686 23604 24692
rect 23392 24622 23398 24686
rect 23462 24622 23604 24686
rect 23392 24550 23604 24622
rect 23392 24486 23534 24550
rect 23598 24486 23604 24550
rect 23392 24480 23604 24486
rect 28288 24480 28636 24692
rect 110160 24480 110508 24692
rect 115192 24686 115404 24692
rect 115192 24622 115198 24686
rect 115262 24622 115404 24686
rect 115192 24550 115404 24622
rect 115192 24486 115198 24550
rect 115262 24486 115404 24550
rect 115192 24480 115404 24486
rect 115600 24686 115812 24692
rect 115600 24622 115606 24686
rect 115670 24622 115812 24686
rect 115600 24550 115812 24622
rect 115600 24486 115742 24550
rect 115806 24486 115812 24550
rect 115600 24480 115812 24486
rect 116008 24686 116220 24692
rect 116008 24622 116150 24686
rect 116214 24622 116220 24686
rect 116008 24556 116220 24622
rect 116416 24556 116628 24692
rect 116008 24550 116628 24556
rect 116008 24486 116014 24550
rect 116078 24486 116628 24550
rect 116008 24480 116628 24486
rect 116824 24686 117036 24692
rect 116824 24622 116966 24686
rect 117030 24622 117036 24686
rect 116824 24550 117036 24622
rect 116824 24486 116830 24550
rect 116894 24486 117036 24550
rect 116824 24480 117036 24486
rect 28424 24420 28500 24480
rect 110432 24420 110508 24480
rect 18088 24278 18300 24284
rect 18088 24214 18230 24278
rect 18294 24214 18300 24278
rect 18088 24142 18300 24214
rect 18088 24078 18230 24142
rect 18294 24078 18300 24142
rect 18088 24072 18300 24078
rect 18496 24278 19116 24284
rect 18496 24214 18910 24278
rect 18974 24214 19116 24278
rect 18496 24208 19116 24214
rect 18496 24142 18708 24208
rect 18496 24078 18502 24142
rect 18566 24078 18708 24142
rect 18496 24072 18708 24078
rect 18904 24072 19116 24208
rect 19312 24278 19524 24284
rect 19312 24214 19318 24278
rect 19382 24214 19524 24278
rect 19312 24142 19524 24214
rect 19312 24078 19318 24142
rect 19382 24078 19524 24142
rect 19312 24072 19524 24078
rect 19720 24142 19932 24284
rect 19720 24078 19862 24142
rect 19926 24078 19932 24142
rect 19720 24072 19932 24078
rect 21760 24278 21972 24284
rect 21760 24214 21766 24278
rect 21830 24214 21972 24278
rect 21760 24072 21972 24214
rect 22168 24278 22380 24284
rect 22168 24214 22310 24278
rect 22374 24214 22380 24278
rect 22168 24142 22380 24214
rect 22168 24078 22310 24142
rect 22374 24078 22380 24142
rect 22168 24072 22380 24078
rect 22576 24142 22788 24284
rect 22576 24078 22582 24142
rect 22646 24078 22788 24142
rect 22576 24072 22788 24078
rect 22984 24278 23196 24284
rect 22984 24214 23126 24278
rect 23190 24214 23196 24278
rect 22984 24142 23196 24214
rect 22984 24078 22990 24142
rect 23054 24078 23196 24142
rect 22984 24072 23196 24078
rect 23392 24278 23604 24284
rect 23392 24214 23534 24278
rect 23598 24214 23604 24278
rect 23392 24142 23604 24214
rect 23392 24078 23398 24142
rect 23462 24078 23604 24142
rect 23392 24072 23604 24078
rect 28288 24208 28636 24420
rect 110160 24208 110508 24420
rect 119136 24344 119756 24420
rect 119136 24284 119212 24344
rect 119680 24284 119756 24344
rect 115192 24278 115404 24284
rect 115192 24214 115198 24278
rect 115262 24214 115404 24278
rect 28288 24148 28364 24208
rect 110296 24148 110372 24208
rect 21760 24012 21836 24072
rect 1224 24006 2388 24012
rect 1224 23942 1230 24006
rect 1294 23942 2318 24006
rect 2382 23942 2388 24006
rect 1224 23936 2388 23942
rect 1768 23928 1980 23936
rect 1768 23872 1798 23928
rect 1854 23872 1980 23928
rect 1768 23800 1980 23872
rect 21760 23664 21972 24012
rect 28288 24006 28636 24148
rect 28288 23942 28430 24006
rect 28494 23942 28636 24006
rect 28288 23936 28636 23942
rect 110160 24006 110508 24148
rect 115192 24142 115404 24214
rect 115192 24078 115334 24142
rect 115398 24078 115404 24142
rect 115192 24072 115404 24078
rect 115600 24278 115812 24284
rect 115600 24214 115742 24278
rect 115806 24214 115812 24278
rect 115600 24142 115812 24214
rect 115600 24078 115742 24142
rect 115806 24078 115812 24142
rect 115600 24072 115812 24078
rect 116008 24278 116220 24284
rect 116008 24214 116014 24278
rect 116078 24214 116220 24278
rect 116008 24142 116220 24214
rect 116008 24078 116150 24142
rect 116214 24078 116220 24142
rect 116008 24072 116220 24078
rect 116416 24142 116628 24284
rect 116416 24078 116558 24142
rect 116622 24078 116628 24142
rect 116416 24072 116628 24078
rect 116824 24278 117036 24284
rect 116824 24214 116830 24278
rect 116894 24214 117036 24278
rect 116824 24072 117036 24214
rect 118864 24278 119212 24284
rect 118864 24214 119006 24278
rect 119070 24214 119212 24278
rect 118864 24208 119212 24214
rect 119272 24278 119484 24284
rect 119272 24214 119414 24278
rect 119478 24214 119484 24278
rect 118864 24142 119076 24208
rect 118864 24078 119006 24142
rect 119070 24078 119076 24142
rect 118864 24072 119076 24078
rect 119272 24148 119484 24214
rect 119680 24278 120300 24284
rect 119680 24214 120094 24278
rect 120158 24214 120300 24278
rect 119680 24208 120300 24214
rect 119272 24142 119620 24148
rect 119272 24078 119278 24142
rect 119342 24078 119620 24142
rect 119272 24072 119620 24078
rect 119680 24142 119892 24208
rect 119680 24078 119686 24142
rect 119750 24078 119892 24142
rect 119680 24072 119892 24078
rect 120088 24072 120300 24208
rect 120496 24278 120708 24284
rect 120496 24214 120638 24278
rect 120702 24214 120708 24278
rect 120496 24142 120708 24214
rect 120496 24078 120638 24142
rect 120702 24078 120708 24142
rect 120496 24072 120708 24078
rect 110160 23942 110438 24006
rect 110502 23942 110508 24006
rect 110160 23936 110508 23942
rect 28560 23876 28636 23936
rect 110432 23876 110508 23936
rect 116824 24012 116900 24072
rect 119544 24012 119620 24072
rect 22168 23870 22788 23876
rect 22168 23806 22310 23870
rect 22374 23806 22582 23870
rect 22646 23806 22788 23870
rect 22168 23800 22788 23806
rect 22168 23740 22380 23800
rect 22168 23664 22516 23740
rect 22576 23664 22788 23800
rect 22984 23870 23196 23876
rect 22984 23806 22990 23870
rect 23054 23806 23196 23870
rect 22984 23734 23196 23806
rect 22984 23670 22990 23734
rect 23054 23670 23196 23734
rect 22984 23664 23196 23670
rect 23392 23870 23604 23876
rect 23392 23806 23398 23870
rect 23462 23806 23604 23870
rect 23392 23734 23604 23806
rect 23392 23670 23398 23734
rect 23462 23670 23604 23734
rect 23392 23664 23604 23670
rect 28288 23734 28636 23876
rect 28288 23670 28430 23734
rect 28494 23670 28636 23734
rect 21896 23604 21972 23664
rect 22304 23604 22380 23664
rect 18088 23598 18300 23604
rect 18088 23534 18230 23598
rect 18294 23534 18300 23598
rect 3128 23326 3884 23332
rect 3128 23262 3814 23326
rect 3878 23262 3884 23326
rect 3128 23256 3884 23262
rect 3128 23196 3340 23256
rect 3944 23196 4156 23332
rect 18088 23326 18300 23534
rect 18088 23262 18230 23326
rect 18294 23262 18300 23326
rect 18088 23256 18300 23262
rect 18496 23598 18708 23604
rect 18496 23534 18502 23598
rect 18566 23534 18708 23598
rect 18496 23332 18708 23534
rect 18904 23332 19116 23604
rect 18496 23326 19116 23332
rect 18496 23262 18638 23326
rect 18702 23262 19116 23326
rect 18496 23256 19116 23262
rect 19312 23462 19524 23468
rect 19312 23398 19318 23462
rect 19382 23398 19524 23462
rect 19312 23326 19524 23398
rect 19312 23262 19318 23326
rect 19382 23262 19524 23326
rect 19312 23256 19524 23262
rect 19720 23462 19932 23468
rect 19720 23398 19862 23462
rect 19926 23398 19932 23462
rect 19720 23326 19932 23398
rect 19720 23262 19726 23326
rect 19790 23262 19932 23326
rect 19720 23256 19932 23262
rect 21760 23256 21972 23604
rect 22168 23326 22380 23604
rect 22440 23604 22516 23664
rect 22440 23528 22788 23604
rect 22168 23262 22174 23326
rect 22238 23262 22380 23326
rect 22168 23256 22380 23262
rect 22576 23326 22788 23528
rect 22576 23262 22582 23326
rect 22646 23262 22788 23326
rect 22576 23256 22788 23262
rect 22984 23462 23196 23468
rect 22984 23398 22990 23462
rect 23054 23398 23196 23462
rect 22984 23326 23196 23398
rect 22984 23262 23126 23326
rect 23190 23262 23196 23326
rect 22984 23256 23196 23262
rect 23392 23462 23604 23468
rect 23392 23398 23398 23462
rect 23462 23398 23604 23462
rect 23392 23326 23604 23398
rect 28288 23392 28636 23670
rect 110160 23734 110508 23876
rect 110160 23670 110438 23734
rect 110502 23670 110508 23734
rect 110160 23392 110508 23670
rect 115192 23870 115404 23876
rect 115192 23806 115334 23870
rect 115398 23806 115404 23870
rect 115192 23734 115404 23806
rect 115192 23670 115334 23734
rect 115398 23670 115404 23734
rect 115192 23664 115404 23670
rect 115600 23870 115812 23876
rect 115600 23806 115742 23870
rect 115806 23806 115812 23870
rect 115600 23734 115812 23806
rect 115600 23670 115742 23734
rect 115806 23670 115812 23734
rect 115600 23664 115812 23670
rect 116008 23870 116628 23876
rect 116008 23806 116150 23870
rect 116214 23806 116558 23870
rect 116622 23806 116628 23870
rect 116008 23800 116628 23806
rect 116008 23740 116220 23800
rect 116008 23664 116356 23740
rect 116416 23664 116628 23800
rect 116824 23664 117036 24012
rect 119544 24006 120572 24012
rect 119544 23942 120502 24006
rect 120566 23942 120572 24006
rect 119544 23936 120572 23942
rect 136816 24006 137572 24012
rect 136816 23942 137502 24006
rect 137566 23942 137572 24006
rect 136816 23936 137572 23942
rect 136816 23928 137028 23936
rect 136816 23872 136944 23928
rect 137000 23872 137028 23928
rect 136816 23800 137028 23872
rect 116144 23604 116220 23664
rect 115192 23462 115404 23468
rect 115192 23398 115334 23462
rect 115398 23398 115404 23462
rect 28424 23332 28500 23392
rect 110296 23332 110372 23392
rect 23392 23262 23534 23326
rect 23598 23262 23604 23326
rect 23392 23256 23604 23262
rect 19312 23196 19388 23256
rect 3128 23120 4156 23196
rect 18398 23190 19388 23196
rect 18360 23126 18366 23190
rect 18430 23126 19388 23190
rect 18398 23120 19388 23126
rect 21760 23196 21836 23256
rect 21760 23054 21972 23196
rect 28288 23120 28636 23332
rect 110160 23190 110508 23332
rect 115192 23326 115404 23398
rect 115192 23262 115334 23326
rect 115398 23262 115404 23326
rect 115192 23256 115404 23262
rect 115600 23462 115812 23468
rect 115600 23398 115742 23462
rect 115806 23398 115812 23462
rect 115600 23326 115812 23398
rect 115600 23262 115742 23326
rect 115806 23262 115812 23326
rect 115600 23256 115812 23262
rect 116008 23256 116220 23604
rect 116280 23604 116356 23664
rect 116824 23604 116900 23664
rect 116280 23528 116628 23604
rect 116416 23332 116628 23528
rect 116318 23326 116628 23332
rect 116280 23262 116286 23326
rect 116350 23262 116628 23326
rect 116318 23256 116628 23262
rect 116824 23256 117036 23604
rect 119680 23598 119892 23604
rect 119680 23534 119686 23598
rect 119750 23534 119892 23598
rect 119680 23468 119892 23534
rect 120088 23468 120300 23604
rect 118864 23462 119076 23468
rect 118864 23398 119006 23462
rect 119070 23398 119076 23462
rect 118864 23326 119076 23398
rect 118864 23262 119006 23326
rect 119070 23262 119076 23326
rect 118864 23256 119076 23262
rect 119272 23462 119484 23468
rect 119272 23398 119278 23462
rect 119342 23398 119484 23462
rect 119272 23326 119484 23398
rect 119272 23262 119278 23326
rect 119342 23262 119484 23326
rect 119272 23256 119484 23262
rect 119680 23392 120300 23468
rect 119680 23326 119892 23392
rect 119680 23262 119686 23326
rect 119750 23262 119892 23326
rect 119680 23256 119892 23262
rect 120088 23256 120300 23392
rect 120496 23598 120708 23604
rect 120496 23534 120502 23598
rect 120566 23534 120638 23598
rect 120702 23534 120708 23598
rect 120496 23326 120708 23534
rect 120496 23262 120638 23326
rect 120702 23262 120708 23326
rect 120496 23256 120708 23262
rect 110160 23126 110438 23190
rect 110502 23126 110508 23190
rect 110160 23120 110508 23126
rect 116824 23196 116900 23256
rect 28288 23060 28364 23120
rect 110296 23060 110372 23120
rect 21760 22990 21766 23054
rect 21830 22990 21972 23054
rect 21760 22984 21972 22990
rect 22168 23054 22380 23060
rect 22168 22990 22174 23054
rect 22238 22990 22380 23054
rect 16864 22848 18164 22924
rect 16864 22788 16940 22848
rect 18088 22788 18164 22848
rect 19176 22848 19796 22924
rect 22168 22848 22380 22990
rect 22576 23054 22788 23060
rect 22576 22990 22582 23054
rect 22646 22990 22788 23054
rect 22576 22924 22788 22990
rect 22440 22848 22788 22924
rect 22984 23054 23196 23060
rect 22984 22990 23126 23054
rect 23190 22990 23196 23054
rect 22984 22848 23196 22990
rect 19176 22788 19252 22848
rect 19720 22788 19796 22848
rect 22440 22788 22516 22848
rect 23120 22788 23196 22848
rect 16592 22712 16940 22788
rect 16592 22440 16804 22712
rect 17000 22516 17212 22788
rect 18088 22782 18436 22788
rect 18088 22718 18230 22782
rect 18294 22718 18366 22782
rect 18430 22718 18436 22782
rect 18088 22712 18436 22718
rect 18496 22782 19252 22788
rect 18496 22718 18638 22782
rect 18702 22718 19252 22782
rect 18496 22712 19252 22718
rect 19312 22782 19524 22788
rect 19312 22718 19318 22782
rect 19382 22718 19524 22782
rect 18088 22576 18300 22712
rect 18496 22576 18708 22712
rect 18904 22576 19116 22712
rect 18496 22516 18572 22576
rect 19312 22516 19524 22718
rect 17000 22440 18572 22516
rect 18670 22510 19524 22516
rect 18632 22446 18638 22510
rect 18702 22446 19524 22510
rect 18670 22440 19524 22446
rect 19720 22782 19932 22788
rect 19720 22718 19726 22782
rect 19790 22718 19932 22782
rect 19720 22510 19932 22718
rect 21760 22782 21972 22788
rect 21760 22718 21766 22782
rect 21830 22718 21972 22782
rect 21760 22646 21972 22718
rect 21760 22582 21766 22646
rect 21830 22582 21972 22646
rect 21760 22576 21972 22582
rect 22168 22712 22516 22788
rect 22168 22652 22380 22712
rect 22168 22646 22516 22652
rect 22168 22582 22446 22646
rect 22510 22582 22516 22646
rect 22168 22576 22516 22582
rect 22576 22576 22788 22788
rect 19720 22446 19862 22510
rect 19926 22446 19932 22510
rect 19720 22440 19932 22446
rect 22304 22516 22380 22576
rect 22576 22516 22652 22576
rect 22304 22440 22652 22516
rect 22984 22440 23196 22788
rect 23392 23054 23604 23060
rect 23392 22990 23534 23054
rect 23598 22990 23604 23054
rect 23392 22848 23604 22990
rect 23392 22788 23468 22848
rect 23392 22440 23604 22788
rect 28288 22782 28636 23060
rect 28288 22718 28566 22782
rect 28630 22718 28636 22782
rect 28288 22712 28636 22718
rect 110160 22918 110508 23060
rect 110160 22854 110438 22918
rect 110502 22854 110508 22918
rect 110160 22782 110508 22854
rect 110160 22718 110166 22782
rect 110230 22718 110508 22782
rect 110160 22712 110508 22718
rect 115192 23054 115404 23060
rect 115192 22990 115334 23054
rect 115398 22990 115404 23054
rect 115192 22848 115404 22990
rect 115600 23054 115812 23060
rect 115600 22990 115742 23054
rect 115806 22990 115812 23054
rect 115600 22848 115812 22990
rect 116008 23054 116356 23060
rect 116008 22990 116286 23054
rect 116350 22990 116356 23054
rect 116008 22984 116356 22990
rect 116008 22924 116220 22984
rect 116008 22848 116356 22924
rect 116416 22848 116628 23060
rect 116824 23054 117036 23196
rect 116824 22990 116830 23054
rect 116894 22990 117036 23054
rect 116824 22984 117036 22990
rect 115192 22788 115268 22848
rect 115600 22788 115676 22848
rect 116008 22788 116084 22848
rect 116280 22788 116356 22848
rect 116552 22788 116628 22848
rect 121448 22848 122068 22924
rect 121448 22788 121524 22848
rect 121992 22788 122068 22848
rect 23120 22380 23196 22440
rect 23528 22380 23604 22440
rect 1224 22374 1980 22380
rect 1224 22310 1230 22374
rect 1294 22310 1980 22374
rect 1224 22304 1980 22310
rect 1768 22248 1980 22304
rect 1768 22192 1798 22248
rect 1854 22244 1980 22248
rect 21760 22374 21972 22380
rect 21760 22310 21766 22374
rect 21830 22310 21972 22374
rect 1854 22238 3204 22244
rect 1854 22192 3134 22238
rect 1768 22174 3134 22192
rect 3198 22174 3204 22238
rect 1768 22168 3204 22174
rect 21760 22238 21972 22310
rect 21760 22174 21766 22238
rect 21830 22174 21972 22238
rect 21760 22168 21972 22174
rect 22168 22032 22380 22380
rect 22478 22374 22788 22380
rect 22440 22310 22446 22374
rect 22510 22310 22788 22374
rect 22478 22304 22788 22310
rect 22576 22032 22788 22304
rect 22984 22032 23196 22380
rect 23392 22032 23604 22380
rect 28288 22374 28636 22516
rect 28288 22310 28294 22374
rect 28358 22310 28566 22374
rect 28630 22310 28636 22374
rect 28288 22102 28636 22310
rect 28288 22038 28294 22102
rect 28358 22038 28430 22102
rect 28494 22038 28636 22102
rect 22168 21972 22244 22032
rect 22576 21972 22652 22032
rect 22984 21972 23060 22032
rect 23392 21972 23468 22032
rect 21760 21966 21972 21972
rect 21760 21902 21766 21966
rect 21830 21902 21972 21966
rect 3128 21830 3340 21836
rect 3128 21766 3134 21830
rect 3198 21766 3340 21830
rect 3128 21700 3340 21766
rect 3944 21700 4156 21836
rect 21760 21830 21972 21902
rect 21760 21766 21902 21830
rect 21966 21766 21972 21830
rect 21760 21760 21972 21766
rect 22168 21836 22380 21972
rect 22576 21836 22788 21972
rect 22168 21830 22788 21836
rect 22168 21766 22310 21830
rect 22374 21766 22788 21830
rect 22168 21760 22788 21766
rect 22984 21830 23196 21972
rect 22984 21766 23126 21830
rect 23190 21766 23196 21830
rect 22984 21760 23196 21766
rect 23392 21830 23604 21972
rect 28288 21896 28636 22038
rect 110160 22510 110508 22516
rect 110160 22446 110166 22510
rect 110230 22446 110508 22510
rect 110160 21896 110508 22446
rect 115192 22440 115404 22788
rect 115328 22380 115404 22440
rect 28424 21836 28500 21896
rect 110432 21836 110508 21896
rect 23392 21766 23398 21830
rect 23462 21766 23604 21830
rect 23392 21760 23604 21766
rect 28288 21830 28636 21836
rect 28288 21766 28430 21830
rect 28494 21766 28636 21830
rect 3128 21624 4156 21700
rect 21760 21558 21972 21564
rect 21760 21494 21902 21558
rect 21966 21494 21972 21558
rect 21760 21422 21972 21494
rect 21760 21358 21902 21422
rect 21966 21358 21972 21422
rect 21760 21352 21972 21358
rect 22168 21558 22788 21564
rect 22168 21494 22310 21558
rect 22374 21494 22788 21558
rect 22168 21488 22788 21494
rect 22168 21428 22380 21488
rect 22168 21422 22516 21428
rect 22168 21358 22310 21422
rect 22374 21358 22446 21422
rect 22510 21358 22516 21422
rect 22168 21352 22516 21358
rect 22576 21352 22788 21488
rect 22984 21558 23196 21564
rect 22984 21494 23126 21558
rect 23190 21494 23196 21558
rect 22984 21422 23196 21494
rect 22984 21358 22990 21422
rect 23054 21358 23196 21422
rect 22984 21352 23196 21358
rect 23392 21558 23604 21564
rect 23392 21494 23398 21558
rect 23462 21494 23604 21558
rect 23392 21422 23604 21494
rect 23392 21358 23398 21422
rect 23462 21358 23604 21422
rect 23392 21352 23604 21358
rect 28288 21352 28636 21766
rect 28560 21292 28636 21352
rect 18768 21216 19388 21292
rect 18768 21156 18844 21216
rect 19312 21156 19388 21216
rect 18496 21150 18844 21156
rect 18496 21086 18638 21150
rect 18702 21086 18844 21150
rect 18496 21080 18844 21086
rect 18496 20944 18708 21080
rect 18904 21014 19116 21156
rect 18904 20950 18910 21014
rect 18974 20950 19116 21014
rect 18904 20944 19116 20950
rect 19312 21014 19524 21156
rect 19312 20950 19318 21014
rect 19382 20950 19524 21014
rect 19312 20944 19524 20950
rect 19720 21150 19932 21156
rect 19720 21086 19862 21150
rect 19926 21086 19932 21150
rect 19720 21014 19932 21086
rect 19720 20950 19862 21014
rect 19926 20950 19932 21014
rect 19720 20944 19932 20950
rect 21760 21150 21972 21156
rect 21760 21086 21902 21150
rect 21966 21086 21972 21150
rect 21760 21014 21972 21086
rect 21760 20950 21766 21014
rect 21830 20950 21972 21014
rect 21760 20944 21972 20950
rect 22168 21150 22380 21156
rect 22478 21150 22788 21156
rect 22168 21086 22310 21150
rect 22374 21086 22380 21150
rect 22440 21086 22446 21150
rect 22510 21086 22788 21150
rect 22168 20944 22380 21086
rect 22478 21080 22788 21086
rect 22576 21014 22788 21080
rect 22576 20950 22718 21014
rect 22782 20950 22788 21014
rect 22576 20944 22788 20950
rect 22984 21150 23196 21156
rect 22984 21086 22990 21150
rect 23054 21086 23196 21150
rect 22984 21014 23196 21086
rect 22984 20950 22990 21014
rect 23054 20950 23196 21014
rect 22984 20944 23196 20950
rect 23392 21150 23604 21156
rect 23392 21086 23398 21150
rect 23462 21086 23604 21150
rect 23392 21014 23604 21086
rect 28288 21080 28636 21292
rect 110160 21352 110508 21836
rect 115192 22032 115404 22380
rect 115600 22440 115812 22788
rect 116008 22652 116220 22788
rect 116280 22712 116628 22788
rect 116008 22646 116356 22652
rect 116008 22582 116286 22646
rect 116350 22582 116356 22646
rect 116008 22576 116356 22582
rect 116416 22576 116628 22712
rect 116824 22782 117036 22788
rect 116824 22718 116830 22782
rect 116894 22718 117036 22782
rect 116824 22646 117036 22718
rect 116824 22582 116830 22646
rect 116894 22582 117036 22646
rect 116824 22576 117036 22582
rect 118864 22782 119076 22788
rect 118864 22718 119006 22782
rect 119070 22718 119076 22782
rect 116824 22516 116900 22576
rect 115872 22440 116900 22516
rect 118864 22510 119076 22718
rect 118864 22446 119006 22510
rect 119070 22446 119076 22510
rect 118864 22440 119076 22446
rect 119272 22782 119484 22788
rect 119272 22718 119278 22782
rect 119342 22718 119484 22782
rect 119272 22440 119484 22718
rect 119680 22782 120300 22788
rect 119680 22718 119686 22782
rect 119750 22718 120300 22782
rect 119680 22712 120300 22718
rect 119680 22576 119892 22712
rect 120088 22652 120300 22712
rect 120496 22782 121524 22788
rect 120496 22718 120638 22782
rect 120702 22718 121524 22782
rect 120496 22712 121524 22718
rect 120088 22576 120436 22652
rect 120496 22646 120708 22712
rect 120496 22582 120502 22646
rect 120566 22582 120708 22646
rect 120496 22576 120708 22582
rect 120360 22516 120436 22576
rect 121584 22516 121796 22788
rect 120360 22440 121796 22516
rect 121992 22440 122204 22788
rect 115600 22380 115676 22440
rect 115872 22380 115948 22440
rect 115600 22304 115948 22380
rect 115600 22032 115812 22304
rect 116008 22032 116220 22380
rect 116318 22374 116628 22380
rect 116280 22310 116286 22374
rect 116350 22310 116628 22374
rect 116318 22304 116628 22310
rect 116416 22108 116628 22304
rect 116824 22374 117036 22380
rect 116824 22310 116830 22374
rect 116894 22310 117036 22374
rect 116824 22238 117036 22310
rect 116824 22174 116830 22238
rect 116894 22174 117036 22238
rect 116824 22168 117036 22174
rect 136816 22374 137572 22380
rect 136816 22310 137502 22374
rect 137566 22310 137572 22374
rect 136816 22304 137572 22310
rect 136816 22248 137028 22304
rect 136816 22192 136944 22248
rect 137000 22192 137028 22248
rect 136816 22168 137028 22192
rect 115192 21972 115268 22032
rect 115736 21972 115812 22032
rect 116144 21972 116220 22032
rect 116280 22032 116628 22108
rect 116280 21972 116356 22032
rect 115192 21830 115404 21972
rect 115192 21766 115198 21830
rect 115262 21766 115404 21830
rect 115192 21760 115404 21766
rect 115600 21830 115812 21972
rect 115600 21766 115606 21830
rect 115670 21766 115812 21830
rect 115600 21760 115812 21766
rect 116008 21896 116356 21972
rect 116008 21836 116220 21896
rect 116416 21836 116628 21972
rect 116008 21830 116628 21836
rect 116008 21766 116558 21830
rect 116622 21766 116628 21830
rect 116008 21760 116628 21766
rect 116824 21966 117036 21972
rect 116824 21902 116830 21966
rect 116894 21902 117036 21966
rect 116824 21830 117036 21902
rect 116824 21766 116966 21830
rect 117030 21766 117036 21830
rect 116824 21760 117036 21766
rect 115192 21558 115404 21564
rect 115192 21494 115198 21558
rect 115262 21494 115404 21558
rect 115192 21422 115404 21494
rect 115192 21358 115334 21422
rect 115398 21358 115404 21422
rect 115192 21352 115404 21358
rect 115600 21558 115812 21564
rect 115600 21494 115606 21558
rect 115670 21494 115812 21558
rect 115600 21422 115812 21494
rect 115600 21358 115606 21422
rect 115670 21358 115812 21422
rect 115600 21352 115812 21358
rect 116008 21428 116220 21564
rect 116416 21558 116628 21564
rect 116416 21494 116558 21558
rect 116622 21494 116628 21558
rect 116416 21428 116628 21494
rect 116824 21558 117036 21564
rect 116824 21494 116966 21558
rect 117030 21494 117036 21558
rect 116008 21422 116764 21428
rect 116008 21358 116014 21422
rect 116078 21358 116764 21422
rect 116008 21352 116764 21358
rect 116824 21422 117036 21494
rect 116824 21358 116966 21422
rect 117030 21358 117036 21422
rect 116824 21352 117036 21358
rect 110160 21292 110236 21352
rect 116144 21292 116220 21352
rect 116688 21292 116764 21352
rect 110160 21080 110508 21292
rect 116144 21216 116492 21292
rect 116688 21216 118940 21292
rect 116416 21156 116492 21216
rect 118864 21156 118940 21216
rect 119544 21216 120164 21292
rect 119544 21156 119620 21216
rect 120088 21156 120164 21216
rect 115192 21150 115404 21156
rect 115192 21086 115334 21150
rect 115398 21086 115404 21150
rect 28560 21020 28636 21080
rect 110296 21020 110372 21080
rect 23392 20950 23534 21014
rect 23598 20950 23604 21014
rect 23392 20944 23604 20950
rect 28288 20808 28636 21020
rect 28560 20748 28636 20808
rect 21760 20742 21972 20748
rect 21760 20678 21766 20742
rect 21830 20678 21972 20742
rect 1768 20568 1980 20612
rect 1768 20512 1798 20568
rect 1854 20512 1980 20568
rect 21760 20606 21972 20678
rect 21760 20542 21902 20606
rect 21966 20542 21972 20606
rect 21760 20536 21972 20542
rect 22168 20612 22380 20748
rect 22576 20742 22788 20748
rect 22576 20678 22718 20742
rect 22782 20678 22788 20742
rect 22576 20612 22788 20678
rect 22168 20606 22788 20612
rect 22168 20542 22310 20606
rect 22374 20542 22718 20606
rect 22782 20542 22788 20606
rect 22168 20536 22788 20542
rect 22984 20742 23196 20748
rect 22984 20678 22990 20742
rect 23054 20678 23196 20742
rect 22984 20606 23196 20678
rect 22984 20542 22990 20606
rect 23054 20542 23196 20606
rect 22984 20536 23196 20542
rect 23392 20742 23604 20748
rect 23392 20678 23534 20742
rect 23598 20678 23604 20742
rect 23392 20606 23604 20678
rect 23392 20542 23398 20606
rect 23462 20542 23604 20606
rect 23392 20536 23604 20542
rect 28288 20536 28636 20748
rect 110160 20808 110508 21020
rect 115192 21014 115404 21086
rect 115192 20950 115198 21014
rect 115262 20950 115404 21014
rect 115192 20944 115404 20950
rect 115600 21150 115812 21156
rect 115600 21086 115606 21150
rect 115670 21086 115812 21150
rect 115600 21014 115812 21086
rect 115600 20950 115606 21014
rect 115670 20950 115812 21014
rect 115600 20944 115812 20950
rect 116008 21150 116220 21156
rect 116008 21086 116014 21150
rect 116078 21086 116220 21150
rect 116008 21014 116220 21086
rect 116008 20950 116014 21014
rect 116078 20950 116220 21014
rect 116008 20944 116220 20950
rect 116416 20944 116628 21156
rect 116824 21150 117036 21156
rect 116824 21086 116966 21150
rect 117030 21086 117036 21150
rect 116824 21014 117036 21086
rect 116824 20950 116830 21014
rect 116894 20950 117036 21014
rect 116824 20944 117036 20950
rect 118864 21150 119076 21156
rect 118864 21086 119006 21150
rect 119070 21086 119076 21150
rect 118864 21020 119076 21086
rect 119272 21080 119620 21156
rect 118864 21014 119212 21020
rect 118864 20950 118870 21014
rect 118934 20950 119212 21014
rect 118864 20944 119212 20950
rect 119272 21014 119484 21080
rect 119272 20950 119414 21014
rect 119478 20950 119484 21014
rect 119272 20944 119484 20950
rect 119680 21014 119892 21156
rect 119680 20950 119822 21014
rect 119886 20950 119892 21014
rect 119680 20944 119892 20950
rect 120088 21150 120572 21156
rect 120088 21086 120502 21150
rect 120566 21086 120572 21150
rect 120088 21080 120572 21086
rect 120088 20944 120300 21080
rect 119136 20884 119212 20944
rect 119680 20884 119756 20944
rect 119136 20808 119756 20884
rect 110160 20748 110236 20808
rect 110160 20536 110508 20748
rect 115192 20742 115404 20748
rect 115192 20678 115198 20742
rect 115262 20678 115404 20742
rect 115192 20606 115404 20678
rect 115192 20542 115198 20606
rect 115262 20542 115404 20606
rect 115192 20536 115404 20542
rect 115600 20742 115812 20748
rect 115600 20678 115606 20742
rect 115670 20678 115812 20742
rect 115600 20606 115812 20678
rect 115600 20542 115606 20606
rect 115670 20542 115812 20606
rect 115600 20536 115812 20542
rect 116008 20742 116220 20748
rect 116008 20678 116014 20742
rect 116078 20678 116220 20742
rect 116008 20612 116220 20678
rect 116416 20612 116628 20748
rect 116008 20606 116628 20612
rect 116008 20542 116014 20606
rect 116078 20542 116628 20606
rect 116008 20536 116628 20542
rect 116824 20742 117036 20748
rect 116824 20678 116830 20742
rect 116894 20678 117036 20742
rect 116824 20606 117036 20678
rect 116824 20542 116966 20606
rect 117030 20542 117036 20606
rect 116824 20536 117036 20542
rect 136816 20568 137028 20612
rect 1768 20476 1980 20512
rect 28424 20476 28500 20536
rect 110296 20476 110372 20536
rect 136816 20512 136944 20568
rect 137000 20512 137028 20568
rect 136816 20476 137028 20512
rect 1224 20470 1980 20476
rect 1224 20406 1230 20470
rect 1294 20406 1980 20470
rect 1224 20400 1980 20406
rect 3128 20340 3340 20476
rect 3944 20340 4156 20476
rect 18360 20400 18980 20476
rect 18360 20340 18436 20400
rect 18904 20340 18980 20400
rect 19176 20400 19796 20476
rect 19176 20340 19252 20400
rect 19720 20340 19796 20400
rect 544 20334 4156 20340
rect 544 20270 550 20334
rect 614 20270 3950 20334
rect 4014 20270 4156 20334
rect 544 20264 4156 20270
rect 17136 20204 17348 20340
rect 17544 20264 18436 20340
rect 17136 20198 17484 20204
rect 17136 20134 17142 20198
rect 17206 20134 17484 20198
rect 17136 20128 17484 20134
rect 17544 20198 17756 20264
rect 17544 20134 17550 20198
rect 17614 20134 17756 20198
rect 17544 20128 17756 20134
rect 18496 20204 18708 20340
rect 18904 20334 19252 20340
rect 18904 20270 18910 20334
rect 18974 20270 19252 20334
rect 18904 20264 19252 20270
rect 19312 20334 19524 20340
rect 19312 20270 19318 20334
rect 19382 20270 19524 20334
rect 18496 20128 18844 20204
rect 18904 20128 19116 20264
rect 19312 20128 19524 20270
rect 19720 20334 19932 20340
rect 19720 20270 19862 20334
rect 19926 20270 19932 20334
rect 19720 20128 19932 20270
rect 21760 20334 21972 20340
rect 21760 20270 21902 20334
rect 21966 20270 21972 20334
rect 21760 20198 21972 20270
rect 21760 20134 21766 20198
rect 21830 20134 21972 20198
rect 21760 20128 21972 20134
rect 22168 20334 22380 20340
rect 22168 20270 22310 20334
rect 22374 20270 22380 20334
rect 22168 20128 22380 20270
rect 22576 20334 22788 20340
rect 22576 20270 22718 20334
rect 22782 20270 22788 20334
rect 22576 20128 22788 20270
rect 22984 20334 23196 20340
rect 22984 20270 22990 20334
rect 23054 20270 23196 20334
rect 22984 20128 23196 20270
rect 23392 20334 23604 20340
rect 23392 20270 23398 20334
rect 23462 20270 23604 20334
rect 23392 20204 23604 20270
rect 28288 20264 28636 20476
rect 110160 20264 110508 20476
rect 119952 20400 121116 20476
rect 136816 20470 137572 20476
rect 136816 20406 137502 20470
rect 137566 20406 137572 20470
rect 136816 20400 137572 20406
rect 119952 20340 120028 20400
rect 121040 20340 121116 20400
rect 28424 20204 28500 20264
rect 110432 20204 110508 20264
rect 23392 20198 24284 20204
rect 23392 20134 23534 20198
rect 23598 20134 24214 20198
rect 24278 20134 24284 20198
rect 23392 20128 24284 20134
rect 17408 20068 17484 20128
rect 18496 20068 18572 20128
rect 17408 19992 18572 20068
rect 18768 20068 18844 20128
rect 19312 20068 19388 20128
rect 18768 19992 19388 20068
rect 28288 20062 28636 20204
rect 28288 19998 28294 20062
rect 28358 19998 28636 20062
rect 28288 19992 28636 19998
rect 110160 19992 110508 20204
rect 115192 20334 115404 20340
rect 115192 20270 115198 20334
rect 115262 20270 115404 20334
rect 115192 20128 115404 20270
rect 115600 20334 115812 20340
rect 115600 20270 115606 20334
rect 115670 20270 115812 20334
rect 115600 20128 115812 20270
rect 116008 20334 116220 20340
rect 116008 20270 116014 20334
rect 116078 20270 116220 20334
rect 116008 20204 116220 20270
rect 116416 20204 116628 20340
rect 116008 20128 116628 20204
rect 116824 20334 117036 20340
rect 116824 20270 116966 20334
rect 117030 20270 117036 20334
rect 116824 20128 117036 20270
rect 118864 20334 119076 20340
rect 118864 20270 118870 20334
rect 118934 20270 119076 20334
rect 118864 20128 119076 20270
rect 119272 20334 119484 20340
rect 119272 20270 119414 20334
rect 119478 20270 119484 20334
rect 119272 20204 119484 20270
rect 119680 20334 120028 20340
rect 119680 20270 119822 20334
rect 119886 20270 120028 20334
rect 119680 20264 120028 20270
rect 119272 20128 119620 20204
rect 119680 20128 119892 20264
rect 120088 20204 120300 20340
rect 121040 20204 121252 20340
rect 121448 20204 121660 20340
rect 120088 20128 120980 20204
rect 121040 20198 121388 20204
rect 121040 20134 121318 20198
rect 121382 20134 121388 20198
rect 121040 20128 121388 20134
rect 121448 20198 124244 20204
rect 121448 20134 124174 20198
rect 124238 20134 124244 20198
rect 121448 20128 124244 20134
rect 119544 20068 119620 20128
rect 120088 20068 120164 20128
rect 119544 19992 120164 20068
rect 120904 20068 120980 20128
rect 121448 20068 121524 20128
rect 120904 19992 121524 20068
rect 28288 19932 28364 19992
rect 110432 19932 110508 19992
rect 23392 19790 23604 19796
rect 23392 19726 23534 19790
rect 23598 19726 23604 19790
rect 23392 19654 23604 19726
rect 23392 19590 23398 19654
rect 23462 19590 23604 19654
rect 23392 19584 23604 19590
rect 24208 19790 27140 19796
rect 24208 19726 24214 19790
rect 24278 19726 27140 19790
rect 24208 19720 27140 19726
rect 24208 19584 24556 19720
rect 26928 19660 27140 19720
rect 28016 19660 28228 19796
rect 28288 19720 28636 19932
rect 110160 19796 110508 19932
rect 124168 19926 124380 19932
rect 124168 19862 124174 19926
rect 124238 19862 124380 19926
rect 110160 19790 110780 19796
rect 110160 19726 110166 19790
rect 110230 19726 110780 19790
rect 110160 19720 110780 19726
rect 124168 19790 124380 19862
rect 124168 19726 124310 19790
rect 124374 19726 124380 19790
rect 124168 19720 124380 19726
rect 26928 19654 27956 19660
rect 26928 19590 27886 19654
rect 27950 19590 27956 19654
rect 26928 19584 27956 19590
rect 28016 19654 28364 19660
rect 28016 19590 28294 19654
rect 28358 19590 28364 19654
rect 28016 19584 28364 19590
rect 110568 19584 110780 19720
rect 123560 19571 123644 19575
rect 123527 19566 123644 19571
rect 123527 19510 123532 19566
rect 123588 19510 123644 19566
rect 123527 19505 123644 19510
rect 123560 19501 123644 19505
rect 27918 19382 30540 19388
rect 27880 19318 27886 19382
rect 27950 19318 30540 19382
rect 27918 19312 30540 19318
rect 28968 19246 29316 19312
rect 28968 19182 29110 19246
rect 29174 19182 29316 19246
rect 28968 19176 29316 19182
rect 29648 19176 29860 19312
rect 30328 19252 30540 19312
rect 30872 19252 31084 19388
rect 31552 19312 32444 19388
rect 31552 19252 31764 19312
rect 30328 19246 31764 19252
rect 30328 19182 30470 19246
rect 30534 19182 31764 19246
rect 30328 19176 31764 19182
rect 32096 19246 32444 19312
rect 32096 19182 32238 19246
rect 32302 19182 32444 19246
rect 32096 19176 32444 19182
rect 32776 19252 32988 19388
rect 33456 19312 34212 19388
rect 33456 19252 33668 19312
rect 32776 19246 33668 19252
rect 32776 19182 32782 19246
rect 32846 19182 32918 19246
rect 32982 19182 33668 19246
rect 32776 19176 33668 19182
rect 34000 19246 34212 19312
rect 34000 19182 34142 19246
rect 34206 19182 34212 19246
rect 34000 19176 34212 19182
rect 34680 19252 34892 19388
rect 35224 19252 35572 19388
rect 34680 19246 35572 19252
rect 34680 19182 34686 19246
rect 34750 19182 35502 19246
rect 35566 19182 35572 19246
rect 34680 19176 35572 19182
rect 35904 19312 36796 19388
rect 35904 19246 36116 19312
rect 35904 19182 35910 19246
rect 35974 19182 36116 19246
rect 35904 19176 36116 19182
rect 36584 19252 36796 19312
rect 37128 19252 37340 19388
rect 37808 19312 39244 19388
rect 37808 19252 38020 19312
rect 36584 19246 38020 19252
rect 36584 19182 36726 19246
rect 36790 19182 38020 19246
rect 36584 19176 38020 19182
rect 38352 19246 38564 19312
rect 38352 19182 38494 19246
rect 38558 19182 38564 19246
rect 38352 19176 38564 19182
rect 39032 19246 39244 19312
rect 39032 19182 39174 19246
rect 39238 19182 39244 19246
rect 39032 19176 39244 19182
rect 39576 19252 39924 19388
rect 40256 19312 41148 19388
rect 40256 19252 40468 19312
rect 39576 19246 40468 19252
rect 39576 19182 39582 19246
rect 39646 19182 40468 19246
rect 39576 19176 40468 19182
rect 40936 19252 41148 19312
rect 41480 19252 41692 19388
rect 42160 19312 43052 19388
rect 42160 19252 42372 19312
rect 40936 19246 42372 19252
rect 40936 19182 40942 19246
rect 41006 19182 41622 19246
rect 41686 19182 42372 19246
rect 40936 19176 42372 19182
rect 42704 19246 43052 19312
rect 42704 19182 42846 19246
rect 42910 19182 43052 19246
rect 42704 19176 43052 19182
rect 43384 19252 43596 19388
rect 44064 19312 46180 19388
rect 44064 19252 44276 19312
rect 43384 19246 44276 19252
rect 43384 19182 43390 19246
rect 43454 19182 44070 19246
rect 44134 19182 44276 19246
rect 43384 19176 44276 19182
rect 44608 19176 44820 19312
rect 45288 19252 45500 19312
rect 45832 19252 46180 19312
rect 46512 19252 46724 19388
rect 45288 19246 45772 19252
rect 45288 19182 45702 19246
rect 45766 19182 45772 19246
rect 45288 19176 45772 19182
rect 45832 19246 46724 19252
rect 45832 19182 46654 19246
rect 46718 19182 46724 19246
rect 45832 19176 46724 19182
rect 47192 19252 47404 19388
rect 47736 19252 47948 19388
rect 47192 19246 47948 19252
rect 47192 19182 47198 19246
rect 47262 19182 47878 19246
rect 47942 19182 47948 19246
rect 47192 19176 47948 19182
rect 48416 19312 49172 19388
rect 48416 19246 48628 19312
rect 48416 19182 48422 19246
rect 48486 19182 48628 19246
rect 48416 19176 48628 19182
rect 48960 19246 49172 19312
rect 48960 19182 49102 19246
rect 49166 19182 49172 19246
rect 48960 19176 49172 19182
rect 49640 19252 49852 19388
rect 50184 19252 50532 19388
rect 50864 19312 51756 19388
rect 50864 19252 51076 19312
rect 49640 19246 51076 19252
rect 49640 19182 49646 19246
rect 49710 19182 50462 19246
rect 50526 19182 51076 19246
rect 49640 19176 51076 19182
rect 51544 19252 51756 19312
rect 52088 19252 52300 19388
rect 52768 19312 54204 19388
rect 52768 19252 52980 19312
rect 51544 19246 52980 19252
rect 51544 19182 52094 19246
rect 52158 19182 52910 19246
rect 52974 19182 52980 19246
rect 51544 19176 52980 19182
rect 53312 19176 53660 19312
rect 53992 19246 54204 19312
rect 53992 19182 54134 19246
rect 54198 19182 54204 19246
rect 53992 19176 54204 19182
rect 54672 19312 55428 19388
rect 54672 19246 54884 19312
rect 54672 19182 54678 19246
rect 54742 19182 54884 19246
rect 54672 19176 54884 19182
rect 55216 19246 55428 19312
rect 55216 19182 55358 19246
rect 55422 19182 55428 19246
rect 55216 19176 55428 19182
rect 55896 19252 56108 19388
rect 56440 19252 56788 19388
rect 55896 19246 56788 19252
rect 55896 19182 55902 19246
rect 55966 19182 56718 19246
rect 56782 19182 56788 19246
rect 55896 19176 56788 19182
rect 57120 19252 57332 19388
rect 57800 19252 58012 19388
rect 58344 19252 58556 19388
rect 59024 19252 59236 19388
rect 57120 19246 57740 19252
rect 57120 19182 57126 19246
rect 57190 19182 57670 19246
rect 57734 19182 57740 19246
rect 57120 19176 57740 19182
rect 57800 19246 59236 19252
rect 57800 19182 58350 19246
rect 58414 19182 59166 19246
rect 59230 19182 59236 19246
rect 57800 19176 59236 19182
rect 59568 19312 60460 19388
rect 60558 19382 61140 19388
rect 60520 19318 60526 19382
rect 60590 19318 61140 19382
rect 60558 19312 61140 19318
rect 59568 19246 59780 19312
rect 59568 19182 59710 19246
rect 59774 19182 59780 19246
rect 59568 19176 59780 19182
rect 60248 19252 60460 19312
rect 60792 19252 61140 19312
rect 61472 19252 61684 19388
rect 60248 19246 61684 19252
rect 60248 19182 61614 19246
rect 61678 19182 61684 19246
rect 60248 19176 61684 19182
rect 62152 19252 62364 19388
rect 62696 19252 62908 19388
rect 62152 19246 62908 19252
rect 62152 19182 62158 19246
rect 62222 19182 62838 19246
rect 62902 19182 62908 19246
rect 62152 19176 62908 19182
rect 63376 19312 64268 19388
rect 63376 19246 63588 19312
rect 63376 19182 63382 19246
rect 63446 19182 63588 19246
rect 63376 19176 63588 19182
rect 63920 19246 64268 19312
rect 63920 19182 64198 19246
rect 64262 19182 64268 19246
rect 63920 19176 64268 19182
rect 64600 19252 64812 19388
rect 65280 19312 66716 19388
rect 65280 19252 65492 19312
rect 64600 19246 65492 19252
rect 64600 19182 64606 19246
rect 64670 19182 65492 19246
rect 64600 19176 65492 19182
rect 65824 19246 66036 19312
rect 65824 19182 65830 19246
rect 65894 19182 66036 19246
rect 65824 19176 66036 19182
rect 66504 19252 66716 19312
rect 67048 19252 67396 19388
rect 67728 19252 67940 19388
rect 66504 19246 67940 19252
rect 66504 19182 67190 19246
rect 67254 19182 67870 19246
rect 67934 19182 67940 19246
rect 66504 19176 67940 19182
rect 68408 19252 68620 19388
rect 68952 19252 69164 19388
rect 69632 19312 70388 19388
rect 69632 19252 69844 19312
rect 68408 19246 69844 19252
rect 68408 19182 68414 19246
rect 68478 19182 69094 19246
rect 69158 19182 69844 19246
rect 68408 19176 69844 19182
rect 70176 19246 70388 19312
rect 70176 19182 70318 19246
rect 70382 19182 70388 19246
rect 70176 19176 70388 19182
rect 70856 19252 71068 19388
rect 71400 19252 71748 19388
rect 72080 19312 72972 19388
rect 72080 19252 72292 19312
rect 70856 19246 72292 19252
rect 70856 19182 70862 19246
rect 70926 19182 71542 19246
rect 71606 19182 72292 19246
rect 70856 19176 72292 19182
rect 72760 19252 72972 19312
rect 73304 19252 73516 19388
rect 73984 19312 74876 19388
rect 73984 19252 74196 19312
rect 72760 19246 74196 19252
rect 72760 19182 73310 19246
rect 73374 19182 74196 19246
rect 72760 19176 74196 19182
rect 74528 19246 74876 19312
rect 74528 19182 74670 19246
rect 74734 19182 74876 19246
rect 74528 19176 74876 19182
rect 75208 19246 75420 19388
rect 75208 19182 75214 19246
rect 75278 19182 75350 19246
rect 75414 19182 75420 19246
rect 75208 19176 75420 19182
rect 75888 19312 76644 19388
rect 75888 19246 76100 19312
rect 75888 19182 75894 19246
rect 75958 19182 76100 19246
rect 75888 19176 76100 19182
rect 76432 19246 76644 19312
rect 76432 19182 76574 19246
rect 76638 19182 76644 19246
rect 76432 19176 76644 19182
rect 77112 19252 77324 19388
rect 77656 19252 78004 19388
rect 77112 19246 78004 19252
rect 77112 19182 77118 19246
rect 77182 19182 77934 19246
rect 77998 19182 78004 19246
rect 77112 19176 78004 19182
rect 78336 19312 79228 19388
rect 78336 19246 78548 19312
rect 78336 19182 78342 19246
rect 78406 19182 78548 19246
rect 78336 19176 78548 19182
rect 79016 19252 79228 19312
rect 79560 19252 79772 19388
rect 80240 19312 80996 19388
rect 80240 19252 80452 19312
rect 80784 19252 80996 19312
rect 79016 19246 80452 19252
rect 80550 19246 80996 19252
rect 79016 19182 79158 19246
rect 79222 19182 80452 19246
rect 80512 19182 80518 19246
rect 80582 19182 80996 19246
rect 79016 19176 80452 19182
rect 80550 19176 80996 19182
rect 81464 19246 81676 19388
rect 81464 19182 81470 19246
rect 81534 19182 81606 19246
rect 81670 19182 81676 19246
rect 81464 19176 81676 19182
rect 82008 19252 82356 19388
rect 82688 19252 82900 19388
rect 82008 19246 82900 19252
rect 82008 19182 82014 19246
rect 82078 19182 82830 19246
rect 82894 19182 82900 19246
rect 82008 19176 82900 19182
rect 83368 19252 83580 19388
rect 83912 19252 84124 19388
rect 83368 19246 84124 19252
rect 83368 19182 83374 19246
rect 83438 19182 84054 19246
rect 84118 19182 84124 19246
rect 83368 19176 84124 19182
rect 84592 19312 85484 19388
rect 84592 19246 84804 19312
rect 84592 19182 84598 19246
rect 84662 19182 84804 19246
rect 84592 19176 84804 19182
rect 85136 19246 85484 19312
rect 85136 19182 85278 19246
rect 85342 19182 85484 19246
rect 85136 19176 85484 19182
rect 85816 19252 86028 19388
rect 86496 19252 86708 19388
rect 87040 19312 89836 19388
rect 87040 19252 87252 19312
rect 85816 19246 86708 19252
rect 86806 19246 87252 19252
rect 85816 19182 85822 19246
rect 85886 19182 86502 19246
rect 86566 19182 86708 19246
rect 86768 19182 86774 19246
rect 86838 19182 87252 19246
rect 85816 19176 86708 19182
rect 86806 19176 87252 19182
rect 87720 19252 87932 19312
rect 87720 19246 88204 19252
rect 87720 19182 88134 19246
rect 88198 19182 88204 19246
rect 87720 19176 88204 19182
rect 88264 19176 88612 19312
rect 88944 19176 89156 19312
rect 89624 19252 89836 19312
rect 90168 19252 90380 19388
rect 89624 19246 90380 19252
rect 89624 19182 89630 19246
rect 89694 19182 90310 19246
rect 90374 19182 90380 19246
rect 89624 19176 90380 19182
rect 90848 19312 92284 19388
rect 90848 19246 91060 19312
rect 90848 19182 90854 19246
rect 90918 19182 91060 19246
rect 90848 19176 91060 19182
rect 91392 19176 91604 19312
rect 92072 19252 92284 19312
rect 92616 19312 94188 19388
rect 94286 19382 94732 19388
rect 94248 19318 94254 19382
rect 94318 19318 94732 19382
rect 94286 19312 94732 19318
rect 92616 19252 92964 19312
rect 92072 19246 92964 19252
rect 92072 19182 92078 19246
rect 92142 19182 92758 19246
rect 92822 19182 92964 19246
rect 92072 19176 92964 19182
rect 93296 19176 93508 19312
rect 93976 19252 94188 19312
rect 94520 19252 94732 19312
rect 95200 19252 95412 19388
rect 93976 19246 94460 19252
rect 93976 19182 94390 19246
rect 94454 19182 94460 19246
rect 93976 19176 94460 19182
rect 94520 19246 95412 19252
rect 94520 19182 95342 19246
rect 95406 19182 95412 19246
rect 94520 19176 95412 19182
rect 95744 19252 96092 19388
rect 96424 19252 96636 19388
rect 97104 19312 98540 19388
rect 97104 19252 97316 19312
rect 95744 19246 97316 19252
rect 95744 19182 95750 19246
rect 95814 19182 96566 19246
rect 96630 19182 97316 19246
rect 95744 19176 97316 19182
rect 97648 19176 97860 19312
rect 98328 19252 98540 19312
rect 98872 19252 99220 19388
rect 98328 19246 99220 19252
rect 98328 19182 98334 19246
rect 98398 19182 99150 19246
rect 99214 19182 99220 19246
rect 98328 19176 99220 19182
rect 99552 19312 100444 19388
rect 99552 19246 99764 19312
rect 99552 19182 99558 19246
rect 99622 19182 99764 19246
rect 99552 19176 99764 19182
rect 100232 19252 100444 19312
rect 100776 19252 100988 19388
rect 101456 19252 101668 19388
rect 100232 19246 101668 19252
rect 100232 19182 100374 19246
rect 100438 19182 101598 19246
rect 101662 19182 101668 19246
rect 100232 19176 101668 19182
rect 102000 19312 102892 19388
rect 102990 19382 103572 19388
rect 102952 19318 102958 19382
rect 103022 19318 103572 19382
rect 102990 19312 103572 19318
rect 102000 19246 102212 19312
rect 102000 19182 102006 19246
rect 102070 19182 102212 19246
rect 102000 19176 102212 19182
rect 102680 19252 102892 19312
rect 103224 19252 103572 19312
rect 102680 19176 103572 19252
rect 103904 19246 104116 19388
rect 103904 19182 104046 19246
rect 104110 19182 104116 19246
rect 103904 19176 104116 19182
rect 104584 19252 104796 19388
rect 105128 19252 105340 19388
rect 104584 19246 105340 19252
rect 104584 19182 104590 19246
rect 104654 19182 105270 19246
rect 105334 19182 105340 19246
rect 104584 19176 105340 19182
rect 105808 19312 106700 19388
rect 105808 19246 106020 19312
rect 105808 19182 105814 19246
rect 105878 19182 106020 19246
rect 105808 19176 106020 19182
rect 106352 19246 106700 19312
rect 106352 19182 106630 19246
rect 106694 19182 106700 19246
rect 106352 19176 106700 19182
rect 107032 19252 107244 19388
rect 107712 19312 109148 19388
rect 107712 19252 107924 19312
rect 107032 19246 107924 19252
rect 107032 19182 107038 19246
rect 107102 19182 107924 19246
rect 107032 19176 107924 19182
rect 108256 19246 108468 19312
rect 108256 19182 108262 19246
rect 108326 19182 108468 19246
rect 108256 19176 108468 19182
rect 108936 19252 109148 19312
rect 109480 19252 109828 19388
rect 108936 19246 109828 19252
rect 108936 19182 109078 19246
rect 109142 19182 109828 19246
rect 124576 19312 138796 19388
rect 124576 19310 124788 19312
rect 124576 19254 124614 19310
rect 124670 19254 124788 19310
rect 108936 19176 109828 19182
rect 123326 19241 123392 19244
rect 123664 19241 123730 19244
rect 123326 19239 123730 19241
rect 123326 19183 123331 19239
rect 123387 19183 123669 19239
rect 123725 19183 123730 19239
rect 123326 19181 123730 19183
rect 123326 19178 123392 19181
rect 123664 19178 123730 19181
rect 124576 19176 124788 19254
rect 3128 18980 3340 19116
rect 1224 18974 3340 18980
rect 1224 18910 1230 18974
rect 1294 18910 3340 18974
rect 1224 18904 3340 18910
rect 1768 18888 1980 18904
rect 1768 18832 1798 18888
rect 1854 18832 1980 18888
rect 1768 18768 1980 18832
rect 3128 18844 3340 18904
rect 3944 18844 4156 19116
rect 3128 18768 4156 18844
rect 15096 19110 17212 19116
rect 15096 19046 17142 19110
rect 17206 19046 17212 19110
rect 15096 19040 17212 19046
rect 15096 18838 15308 19040
rect 35496 18974 35980 18980
rect 35496 18910 35910 18974
rect 35974 18910 35980 18974
rect 35496 18904 35980 18910
rect 77928 18974 78412 18980
rect 77928 18910 78342 18974
rect 78406 18910 78412 18974
rect 77928 18904 78412 18910
rect 35496 18844 35572 18904
rect 77928 18844 78004 18904
rect 136816 18888 137028 18980
rect 15096 18774 15238 18838
rect 15302 18774 15308 18838
rect 15096 18768 15308 18774
rect 29104 18838 29724 18844
rect 29104 18774 29110 18838
rect 29174 18774 29724 18838
rect 29104 18768 29724 18774
rect 29104 18632 29452 18768
rect 29512 18632 29724 18768
rect 30464 18838 31084 18844
rect 30464 18774 30470 18838
rect 30534 18774 31084 18838
rect 30464 18768 31084 18774
rect 30464 18632 30676 18768
rect 30736 18632 31084 18768
rect 31688 18708 31900 18844
rect 32096 18838 32852 18844
rect 32096 18774 32238 18838
rect 32302 18774 32782 18838
rect 32846 18774 32852 18838
rect 32096 18768 32852 18774
rect 32912 18838 33532 18844
rect 32912 18774 32918 18838
rect 32982 18774 33532 18838
rect 32912 18768 33532 18774
rect 32096 18708 32308 18768
rect 31688 18632 32308 18708
rect 32912 18632 33124 18768
rect 33320 18632 33532 18768
rect 34136 18838 34348 18844
rect 34136 18774 34142 18838
rect 34206 18774 34348 18838
rect 34136 18708 34348 18774
rect 34544 18838 34756 18844
rect 34544 18774 34686 18838
rect 34750 18774 34756 18838
rect 34544 18708 34756 18774
rect 34136 18632 34756 18708
rect 35360 18838 35980 18844
rect 35360 18774 35502 18838
rect 35566 18774 35980 18838
rect 35360 18768 35980 18774
rect 35360 18632 35572 18768
rect 35768 18632 35980 18768
rect 36584 18838 36932 18844
rect 36584 18774 36726 18838
rect 36790 18774 36932 18838
rect 36584 18708 36932 18774
rect 36992 18708 37204 18844
rect 36584 18632 37204 18708
rect 37944 18708 38156 18844
rect 38216 18838 38564 18844
rect 38216 18774 38494 18838
rect 38558 18774 38564 18838
rect 38216 18708 38564 18774
rect 37944 18632 38564 18708
rect 39168 18838 39788 18844
rect 39168 18774 39174 18838
rect 39238 18774 39582 18838
rect 39646 18774 39788 18838
rect 39168 18768 39788 18774
rect 39168 18632 39380 18768
rect 39576 18632 39788 18768
rect 40392 18708 40604 18844
rect 40800 18838 41012 18844
rect 40800 18774 40942 18838
rect 41006 18774 41012 18838
rect 40800 18708 41012 18774
rect 40392 18632 41012 18708
rect 41616 18838 42236 18844
rect 41616 18774 41622 18838
rect 41686 18774 42236 18838
rect 41616 18768 42236 18774
rect 41616 18632 41828 18768
rect 42024 18632 42236 18768
rect 42840 18838 43052 18844
rect 42840 18774 42846 18838
rect 42910 18774 43052 18838
rect 42840 18708 43052 18774
rect 43248 18838 43460 18844
rect 43248 18774 43390 18838
rect 43454 18774 43460 18838
rect 43248 18708 43460 18774
rect 42840 18632 43460 18708
rect 44064 18838 44684 18844
rect 44064 18774 44070 18838
rect 44134 18774 44684 18838
rect 44064 18768 44684 18774
rect 44064 18632 44412 18768
rect 44472 18632 44684 18768
rect 45424 18838 46044 18844
rect 45424 18774 45702 18838
rect 45766 18774 46044 18838
rect 45424 18768 46044 18774
rect 45424 18632 45636 18768
rect 45696 18632 46044 18768
rect 46648 18838 46860 18844
rect 46648 18774 46654 18838
rect 46718 18774 46860 18838
rect 46648 18708 46860 18774
rect 47056 18838 47268 18844
rect 47056 18774 47198 18838
rect 47262 18774 47268 18838
rect 47056 18708 47268 18774
rect 46648 18632 47268 18708
rect 47872 18838 48492 18844
rect 47872 18774 47878 18838
rect 47942 18774 48422 18838
rect 48486 18774 48492 18838
rect 47872 18768 48492 18774
rect 47872 18632 48084 18768
rect 48280 18632 48492 18768
rect 49096 18838 49308 18844
rect 49096 18774 49102 18838
rect 49166 18774 49308 18838
rect 49096 18708 49308 18774
rect 49504 18838 49716 18844
rect 49504 18774 49646 18838
rect 49710 18774 49716 18838
rect 49504 18708 49716 18774
rect 49096 18632 49716 18708
rect 50320 18838 50940 18844
rect 50320 18774 50462 18838
rect 50526 18774 50940 18838
rect 50320 18768 50940 18774
rect 50320 18632 50668 18768
rect 50728 18632 50940 18768
rect 51680 18838 52300 18844
rect 51680 18774 52094 18838
rect 52158 18774 52300 18838
rect 51680 18768 52300 18774
rect 51680 18632 51892 18768
rect 51952 18632 52300 18768
rect 52904 18838 53116 18844
rect 52904 18774 52910 18838
rect 52974 18774 53116 18838
rect 52904 18708 53116 18774
rect 53312 18708 53524 18844
rect 52904 18632 53524 18708
rect 54128 18838 54748 18844
rect 54128 18774 54134 18838
rect 54198 18774 54678 18838
rect 54742 18774 54748 18838
rect 54128 18768 54748 18774
rect 54128 18632 54340 18768
rect 54536 18632 54748 18768
rect 55352 18838 55564 18844
rect 55352 18774 55358 18838
rect 55422 18774 55564 18838
rect 55352 18708 55564 18774
rect 55760 18838 55972 18844
rect 55760 18774 55902 18838
rect 55966 18774 55972 18838
rect 55760 18708 55972 18774
rect 55352 18632 55972 18708
rect 56576 18838 57196 18844
rect 57702 18838 58148 18844
rect 56576 18774 56718 18838
rect 56782 18774 57126 18838
rect 57190 18774 57196 18838
rect 57664 18774 57670 18838
rect 57734 18774 58148 18838
rect 56576 18768 57196 18774
rect 57702 18768 58148 18774
rect 56576 18632 56788 18768
rect 56984 18632 57196 18768
rect 57800 18708 58148 18768
rect 58208 18838 58420 18844
rect 58208 18774 58350 18838
rect 58414 18774 58420 18838
rect 58208 18708 58420 18774
rect 57800 18632 58420 18708
rect 59160 18838 59372 18844
rect 59160 18774 59166 18838
rect 59230 18774 59372 18838
rect 59160 18708 59372 18774
rect 59432 18838 59780 18844
rect 59432 18774 59710 18838
rect 59774 18774 59780 18838
rect 59432 18708 59780 18774
rect 59160 18632 59780 18708
rect 60384 18838 61004 18844
rect 60384 18774 60526 18838
rect 60590 18774 61004 18838
rect 60384 18768 61004 18774
rect 60384 18632 60596 18768
rect 60792 18632 61004 18768
rect 61608 18838 61820 18844
rect 61608 18774 61614 18838
rect 61678 18774 61820 18838
rect 61608 18708 61820 18774
rect 62016 18838 62228 18844
rect 62016 18774 62158 18838
rect 62222 18774 62228 18838
rect 62016 18708 62228 18774
rect 61608 18632 62228 18708
rect 62832 18838 63452 18844
rect 62832 18774 62838 18838
rect 62902 18774 63382 18838
rect 63446 18774 63452 18838
rect 62832 18768 63452 18774
rect 62832 18632 63044 18768
rect 63240 18632 63452 18768
rect 64056 18838 64268 18844
rect 64056 18774 64198 18838
rect 64262 18774 64268 18838
rect 64056 18708 64268 18774
rect 64464 18838 64676 18844
rect 64464 18774 64606 18838
rect 64670 18774 64676 18838
rect 64464 18708 64676 18774
rect 64056 18632 64676 18708
rect 65280 18838 65900 18844
rect 65280 18774 65830 18838
rect 65894 18774 65900 18838
rect 65280 18768 65900 18774
rect 65280 18632 65628 18768
rect 65688 18632 65900 18768
rect 66640 18838 67260 18844
rect 66640 18774 67190 18838
rect 67254 18774 67260 18838
rect 66640 18768 67260 18774
rect 66640 18632 66852 18768
rect 66912 18632 67260 18768
rect 67864 18838 68076 18844
rect 67864 18774 67870 18838
rect 67934 18774 68076 18838
rect 67864 18708 68076 18774
rect 68272 18838 68484 18844
rect 68272 18774 68414 18838
rect 68478 18774 68484 18838
rect 68272 18708 68484 18774
rect 67864 18632 68484 18708
rect 69088 18838 69708 18844
rect 69088 18774 69094 18838
rect 69158 18774 69708 18838
rect 69088 18768 69708 18774
rect 69088 18632 69300 18768
rect 69496 18632 69708 18768
rect 70312 18838 70524 18844
rect 70312 18774 70318 18838
rect 70382 18774 70524 18838
rect 70312 18708 70524 18774
rect 70720 18838 70932 18844
rect 70720 18774 70862 18838
rect 70926 18774 70932 18838
rect 70720 18708 70932 18774
rect 70312 18632 70932 18708
rect 71536 18838 72156 18844
rect 71536 18774 71542 18838
rect 71606 18774 72156 18838
rect 71536 18768 72156 18774
rect 71536 18632 71884 18768
rect 71944 18632 72156 18768
rect 72896 18838 73516 18844
rect 72896 18774 73310 18838
rect 73374 18774 73516 18838
rect 72896 18768 73516 18774
rect 72896 18632 73108 18768
rect 73168 18632 73516 18768
rect 74120 18708 74332 18844
rect 74528 18838 75284 18844
rect 74528 18774 74670 18838
rect 74734 18774 75214 18838
rect 75278 18774 75284 18838
rect 74528 18768 75284 18774
rect 75344 18838 75964 18844
rect 75344 18774 75350 18838
rect 75414 18774 75894 18838
rect 75958 18774 75964 18838
rect 75344 18768 75964 18774
rect 74528 18708 74740 18768
rect 74120 18632 74740 18708
rect 75344 18632 75556 18768
rect 75752 18632 75964 18768
rect 76568 18838 76780 18844
rect 76568 18774 76574 18838
rect 76638 18774 76780 18838
rect 76568 18708 76780 18774
rect 76976 18838 77188 18844
rect 76976 18774 77118 18838
rect 77182 18774 77188 18838
rect 76976 18708 77188 18774
rect 76568 18702 77188 18708
rect 76568 18638 77118 18702
rect 77182 18638 77188 18702
rect 76568 18632 77188 18638
rect 77792 18838 78412 18844
rect 77792 18774 77934 18838
rect 77998 18774 78412 18838
rect 77792 18768 78412 18774
rect 77792 18632 78004 18768
rect 78200 18632 78412 18768
rect 79016 18838 79636 18844
rect 79016 18774 79158 18838
rect 79222 18774 79636 18838
rect 79016 18768 79636 18774
rect 79016 18632 79364 18768
rect 79424 18632 79636 18768
rect 80376 18838 80588 18844
rect 80376 18774 80518 18838
rect 80582 18774 80588 18838
rect 80376 18708 80588 18774
rect 80648 18838 81540 18844
rect 80648 18774 81470 18838
rect 81534 18774 81540 18838
rect 80648 18768 81540 18774
rect 81600 18838 82220 18844
rect 81600 18774 81606 18838
rect 81670 18774 82014 18838
rect 82078 18774 82220 18838
rect 81600 18768 82220 18774
rect 80648 18708 80996 18768
rect 80376 18632 80996 18708
rect 81600 18632 81812 18768
rect 82008 18632 82220 18768
rect 82824 18838 83036 18844
rect 82824 18774 82830 18838
rect 82894 18774 83036 18838
rect 82824 18708 83036 18774
rect 83232 18838 83444 18844
rect 83232 18774 83374 18838
rect 83438 18774 83444 18838
rect 83232 18708 83444 18774
rect 82824 18632 83444 18708
rect 84048 18838 84668 18844
rect 84048 18774 84054 18838
rect 84118 18774 84598 18838
rect 84662 18774 84668 18838
rect 84048 18768 84668 18774
rect 84048 18632 84260 18768
rect 84456 18632 84668 18768
rect 85272 18838 85484 18844
rect 85272 18774 85278 18838
rect 85342 18774 85484 18838
rect 85272 18708 85484 18774
rect 85680 18838 85892 18844
rect 85680 18774 85822 18838
rect 85886 18774 85892 18838
rect 85680 18708 85892 18774
rect 85272 18632 85892 18708
rect 86496 18838 87116 18844
rect 86496 18774 86502 18838
rect 86566 18774 86774 18838
rect 86838 18774 87116 18838
rect 86496 18768 87116 18774
rect 86496 18632 86844 18768
rect 86904 18632 87116 18768
rect 87856 18838 88476 18844
rect 87856 18774 88134 18838
rect 88198 18774 88476 18838
rect 87856 18768 88476 18774
rect 87856 18632 88068 18768
rect 88128 18632 88476 18768
rect 89080 18708 89292 18844
rect 89488 18838 89700 18844
rect 89488 18774 89630 18838
rect 89694 18774 89700 18838
rect 89488 18708 89700 18774
rect 89080 18632 89700 18708
rect 90304 18838 90924 18844
rect 90304 18774 90310 18838
rect 90374 18774 90854 18838
rect 90918 18774 90924 18838
rect 90304 18768 90924 18774
rect 90304 18632 90516 18768
rect 90712 18632 90924 18768
rect 91528 18708 91740 18844
rect 91936 18838 92148 18844
rect 91936 18774 92078 18838
rect 92142 18774 92148 18838
rect 91936 18708 92148 18774
rect 91528 18632 92148 18708
rect 92752 18838 93372 18844
rect 92752 18774 92758 18838
rect 92822 18774 93372 18838
rect 92752 18768 93372 18774
rect 92752 18632 93100 18768
rect 93160 18632 93372 18768
rect 94112 18838 94732 18844
rect 94112 18774 94254 18838
rect 94318 18774 94390 18838
rect 94454 18774 94732 18838
rect 94112 18768 94732 18774
rect 94112 18632 94324 18768
rect 94384 18632 94732 18768
rect 95336 18838 95548 18844
rect 95336 18774 95342 18838
rect 95406 18774 95548 18838
rect 95336 18708 95548 18774
rect 95744 18838 95956 18844
rect 95744 18774 95750 18838
rect 95814 18774 95956 18838
rect 95744 18708 95956 18774
rect 95336 18632 95956 18708
rect 96560 18838 97180 18844
rect 96560 18774 96566 18838
rect 96630 18774 97180 18838
rect 96560 18768 97180 18774
rect 96560 18632 96772 18768
rect 96968 18632 97180 18768
rect 97784 18708 97996 18844
rect 98192 18838 98404 18844
rect 98192 18774 98334 18838
rect 98398 18774 98404 18838
rect 98192 18708 98404 18774
rect 97784 18632 98404 18708
rect 99008 18838 99628 18844
rect 99008 18774 99150 18838
rect 99214 18774 99558 18838
rect 99622 18774 99628 18838
rect 99008 18768 99628 18774
rect 99008 18632 99220 18768
rect 99416 18632 99628 18768
rect 100232 18838 100580 18844
rect 100232 18774 100374 18838
rect 100438 18774 100580 18838
rect 100232 18708 100580 18774
rect 100640 18708 100852 18844
rect 100232 18632 100852 18708
rect 101592 18838 101804 18844
rect 101592 18774 101598 18838
rect 101662 18774 101804 18838
rect 101592 18708 101804 18774
rect 101864 18838 102212 18844
rect 101864 18774 102006 18838
rect 102070 18774 102212 18838
rect 101864 18708 102212 18774
rect 101592 18632 102212 18708
rect 102816 18838 103436 18844
rect 102816 18774 102958 18838
rect 103022 18774 103436 18838
rect 102816 18768 103436 18774
rect 102816 18632 103028 18768
rect 103224 18708 103436 18768
rect 104040 18838 104252 18844
rect 104040 18774 104046 18838
rect 104110 18774 104252 18838
rect 104040 18708 104252 18774
rect 104448 18838 104660 18844
rect 104448 18774 104590 18838
rect 104654 18774 104660 18838
rect 104448 18708 104660 18774
rect 103224 18632 104660 18708
rect 105264 18838 105884 18844
rect 105264 18774 105270 18838
rect 105334 18774 105814 18838
rect 105878 18774 105884 18838
rect 105264 18768 105884 18774
rect 105264 18632 105476 18768
rect 105672 18632 105884 18768
rect 106488 18838 106700 18844
rect 106488 18774 106630 18838
rect 106694 18774 106700 18838
rect 106488 18708 106700 18774
rect 106896 18838 107108 18844
rect 106896 18774 107038 18838
rect 107102 18774 107108 18838
rect 106896 18708 107108 18774
rect 106488 18632 107108 18708
rect 107712 18838 108332 18844
rect 107712 18774 108262 18838
rect 108326 18774 108332 18838
rect 107712 18768 108332 18774
rect 107712 18632 108060 18768
rect 108120 18632 108332 18768
rect 109072 18838 109284 18844
rect 109072 18774 109078 18838
rect 109142 18774 109284 18838
rect 109072 18632 109284 18774
rect 136816 18832 136944 18888
rect 137000 18844 137028 18888
rect 137000 18838 137572 18844
rect 137000 18832 137502 18838
rect 136816 18774 137502 18832
rect 137566 18774 137572 18838
rect 136816 18768 137572 18774
rect 121350 18566 124380 18572
rect 121312 18502 121318 18566
rect 121382 18502 124380 18566
rect 121350 18496 124380 18502
rect 124168 18430 124380 18496
rect 124168 18366 124174 18430
rect 124238 18366 124380 18430
rect 124168 18360 124380 18366
rect 15205 18255 15271 18258
rect 23747 18255 23813 18258
rect 15205 18253 23813 18255
rect 15205 18197 15210 18253
rect 15266 18197 23752 18253
rect 23808 18197 23813 18253
rect 15205 18195 23813 18197
rect 15205 18192 15271 18195
rect 23747 18192 23813 18195
rect 2535 17894 2541 17958
rect 2605 17956 2611 17958
rect 2605 17896 29383 17956
rect 2605 17894 2611 17896
rect 123246 17683 123312 17686
rect 123664 17683 123730 17686
rect 123246 17681 123730 17683
rect 123246 17625 123251 17681
rect 123307 17625 123669 17681
rect 123725 17625 123730 17681
rect 123246 17623 123730 17625
rect 123246 17620 123312 17623
rect 123664 17620 123730 17623
rect 3128 17614 3884 17620
rect 3128 17550 3814 17614
rect 3878 17550 3884 17614
rect 3128 17544 3884 17550
rect 3128 17484 3340 17544
rect 3944 17484 4156 17620
rect 3128 17408 4156 17484
rect 15096 17614 17620 17620
rect 15096 17550 17550 17614
rect 17614 17550 17620 17614
rect 15096 17544 17620 17550
rect 124576 17610 124788 17756
rect 124576 17554 124614 17610
rect 124670 17554 124788 17610
rect 15096 17478 15308 17544
rect 15096 17414 15102 17478
rect 15166 17414 15308 17478
rect 15096 17408 15308 17414
rect 124576 17484 124788 17554
rect 124576 17408 138796 17484
rect 1768 17208 1980 17348
rect 1768 17152 1798 17208
rect 1854 17152 1980 17208
rect 1768 17076 1980 17152
rect 21080 17342 21836 17348
rect 21080 17278 21766 17342
rect 21830 17278 21836 17342
rect 21080 17272 21836 17278
rect 21080 17212 21292 17272
rect 22168 17212 22380 17348
rect 21080 17206 22380 17212
rect 21080 17142 21086 17206
rect 21150 17142 22380 17206
rect 21080 17136 22380 17142
rect 29920 17136 32716 17212
rect 1224 17070 1980 17076
rect 1224 17006 1230 17070
rect 1294 17006 1980 17070
rect 1224 17000 1980 17006
rect 29920 17070 30268 17136
rect 29920 17006 29926 17070
rect 29990 17006 30268 17070
rect 29920 17000 30268 17006
rect 31280 17000 31492 17136
rect 32504 17076 32716 17136
rect 33728 17136 35164 17212
rect 33728 17076 33940 17136
rect 32504 17070 33940 17076
rect 32504 17006 32646 17070
rect 32710 17006 33940 17070
rect 32504 17000 33940 17006
rect 34952 17076 35164 17136
rect 36176 17136 37748 17212
rect 36176 17076 36388 17136
rect 34952 17070 36388 17076
rect 34952 17006 35094 17070
rect 35158 17006 36388 17070
rect 34952 17000 36388 17006
rect 37400 17076 37748 17136
rect 38760 17076 38972 17212
rect 39984 17136 41420 17212
rect 39984 17076 40196 17136
rect 37400 17070 40196 17076
rect 37400 17006 37406 17070
rect 37470 17006 40126 17070
rect 40190 17006 40196 17070
rect 37400 17000 40196 17006
rect 41208 17076 41420 17136
rect 42432 17136 43868 17212
rect 42432 17076 42644 17136
rect 41208 17070 42644 17076
rect 41208 17006 42438 17070
rect 42502 17006 42644 17070
rect 41208 17000 42644 17006
rect 43656 17076 43868 17136
rect 44880 17136 47676 17212
rect 44880 17076 45228 17136
rect 43656 17070 45228 17076
rect 43656 17006 44886 17070
rect 44950 17006 45228 17070
rect 43656 17000 45228 17006
rect 46240 17000 46452 17136
rect 47464 17076 47676 17136
rect 48688 17136 50124 17212
rect 48688 17076 48900 17136
rect 47464 17070 48900 17076
rect 47464 17006 47606 17070
rect 47670 17006 48900 17070
rect 47464 17000 48900 17006
rect 49912 17076 50124 17136
rect 51136 17136 53932 17212
rect 51136 17076 51484 17136
rect 49912 17070 51484 17076
rect 49912 17006 49918 17070
rect 49982 17006 51484 17070
rect 49912 17000 51484 17006
rect 52496 17070 52708 17136
rect 52496 17006 52502 17070
rect 52566 17006 52708 17070
rect 52496 17000 52708 17006
rect 53720 17076 53932 17136
rect 54944 17136 56380 17212
rect 54944 17076 55156 17136
rect 53720 17070 55156 17076
rect 53720 17006 55086 17070
rect 55150 17006 55156 17070
rect 53720 17000 55156 17006
rect 56168 17076 56380 17136
rect 57392 17136 58964 17212
rect 57392 17076 57604 17136
rect 56168 17070 57604 17076
rect 56168 17006 57398 17070
rect 57462 17006 57604 17070
rect 56168 17000 57604 17006
rect 58616 17076 58964 17136
rect 59976 17076 60188 17212
rect 61200 17136 62636 17212
rect 61200 17076 61412 17136
rect 58616 17070 61412 17076
rect 58616 17006 59982 17070
rect 60046 17006 61412 17070
rect 58616 17000 61412 17006
rect 62424 17076 62636 17136
rect 63648 17136 65084 17212
rect 63648 17076 63860 17136
rect 62424 17070 63860 17076
rect 62424 17006 62566 17070
rect 62630 17006 63860 17070
rect 62424 17000 63860 17006
rect 64872 17076 65084 17136
rect 66096 17136 68892 17212
rect 66096 17076 66444 17136
rect 64872 17070 66444 17076
rect 64872 17006 64878 17070
rect 64942 17006 66444 17070
rect 64872 17000 66444 17006
rect 67456 17070 67668 17136
rect 67456 17006 67598 17070
rect 67662 17006 67668 17070
rect 67456 17000 67668 17006
rect 68680 17076 68892 17136
rect 69904 17136 71340 17212
rect 69904 17076 70116 17136
rect 68680 17070 70116 17076
rect 68680 17006 69910 17070
rect 69974 17006 70116 17070
rect 68680 17000 70116 17006
rect 71128 17076 71340 17136
rect 72352 17076 72700 17212
rect 73712 17136 75148 17212
rect 73712 17076 73924 17136
rect 71128 17070 73924 17076
rect 71128 17006 72358 17070
rect 72422 17006 73924 17070
rect 71128 17000 73924 17006
rect 74936 17076 75148 17136
rect 76160 17136 77596 17212
rect 76160 17076 76372 17136
rect 74936 17070 76372 17076
rect 74936 17006 75078 17070
rect 75142 17006 76372 17070
rect 74936 17000 76372 17006
rect 77384 17076 77596 17136
rect 78608 17136 80180 17212
rect 78608 17076 78820 17136
rect 77384 17070 78820 17076
rect 77384 17006 77526 17070
rect 77590 17006 78820 17070
rect 77384 17000 78820 17006
rect 79832 17076 80180 17136
rect 81192 17076 81404 17212
rect 82416 17136 83852 17212
rect 82416 17076 82628 17136
rect 79832 17070 82628 17076
rect 79832 17006 79838 17070
rect 79902 17006 82558 17070
rect 82622 17006 82628 17070
rect 79832 17000 82628 17006
rect 83640 17076 83852 17136
rect 84864 17136 86300 17212
rect 84864 17076 85076 17136
rect 83640 17070 85076 17076
rect 83640 17006 84870 17070
rect 84934 17006 85076 17070
rect 83640 17000 85076 17006
rect 86088 17076 86300 17136
rect 87312 17136 90108 17212
rect 87312 17076 87660 17136
rect 86088 17070 87660 17076
rect 86088 17006 87318 17070
rect 87382 17006 87660 17070
rect 86088 17000 87660 17006
rect 88672 17000 88884 17136
rect 89896 17076 90108 17136
rect 91120 17136 92556 17212
rect 91120 17076 91332 17136
rect 89896 17070 91332 17076
rect 89896 17006 90038 17070
rect 90102 17006 91332 17070
rect 89896 17000 91332 17006
rect 92344 17076 92556 17136
rect 93568 17076 93916 17212
rect 94928 17136 96364 17212
rect 94928 17076 95140 17136
rect 92344 17070 95140 17076
rect 92344 17006 92350 17070
rect 92414 17006 94934 17070
rect 94998 17006 95140 17070
rect 92344 17000 95140 17006
rect 96152 17076 96364 17136
rect 97376 17136 98812 17212
rect 97376 17076 97588 17136
rect 96152 17070 97588 17076
rect 96152 17006 97518 17070
rect 97582 17006 97588 17070
rect 96152 17000 97588 17006
rect 98600 17076 98812 17136
rect 99824 17136 101396 17212
rect 99824 17076 100036 17136
rect 98600 17070 100036 17076
rect 98600 17006 99830 17070
rect 99894 17006 100036 17070
rect 98600 17000 100036 17006
rect 101048 17076 101396 17136
rect 102408 17076 102620 17212
rect 103632 17136 105068 17212
rect 103632 17076 103844 17136
rect 101048 17070 103844 17076
rect 101048 17006 102414 17070
rect 102478 17006 103844 17070
rect 101048 17000 103844 17006
rect 104856 17076 105068 17136
rect 106080 17136 107516 17212
rect 106080 17076 106292 17136
rect 104856 17070 106292 17076
rect 104856 17006 104998 17070
rect 105062 17006 106292 17070
rect 104856 17000 106292 17006
rect 107304 17076 107516 17136
rect 108528 17206 110236 17212
rect 108528 17142 110166 17206
rect 110230 17142 110236 17206
rect 108528 17136 110236 17142
rect 136816 17208 137028 17348
rect 136816 17152 136944 17208
rect 137000 17152 137028 17208
rect 108528 17076 108876 17136
rect 136816 17076 137028 17152
rect 107304 17070 108876 17076
rect 107304 17006 107310 17070
rect 107374 17006 108876 17070
rect 107304 17000 108876 17006
rect 124168 17070 124380 17076
rect 124168 17006 124310 17070
rect 124374 17006 124380 17070
rect 124168 16940 124380 17006
rect 136816 17070 137572 17076
rect 136816 17006 137502 17070
rect 137566 17006 137572 17070
rect 136816 17000 137572 17006
rect 124168 16934 124478 16940
rect 124168 16870 124446 16934
rect 124510 16870 124516 16934
rect 124168 16864 124478 16870
rect 124576 16482 138796 16532
rect 124576 16426 124614 16482
rect 124670 16456 138796 16482
rect 124670 16426 124788 16456
rect 123166 16413 123232 16416
rect 123664 16413 123730 16416
rect 123166 16411 123730 16413
rect 123166 16355 123171 16411
rect 123227 16355 123669 16411
rect 123725 16355 123730 16411
rect 123166 16353 123730 16355
rect 123166 16350 123232 16353
rect 123664 16350 123730 16353
rect 124576 16320 124788 16426
rect 3128 16184 4156 16260
rect 3128 16118 3340 16184
rect 3128 16054 3134 16118
rect 3198 16054 3340 16118
rect 3128 16048 3340 16054
rect 3944 16048 4156 16184
rect 15096 16254 15308 16260
rect 15096 16190 15238 16254
rect 15302 16190 15308 16254
rect 15096 16118 15308 16190
rect 15096 16054 15238 16118
rect 15302 16054 15308 16118
rect 15096 16048 15308 16054
rect 21080 15912 22380 15988
rect 21080 15776 21292 15912
rect 22168 15852 22380 15912
rect 22168 15846 23468 15852
rect 22168 15782 22310 15846
rect 22374 15782 23398 15846
rect 23462 15782 23468 15846
rect 22168 15776 23468 15782
rect 124168 15710 124380 15716
rect 124168 15646 124174 15710
rect 124238 15646 124380 15710
rect 1224 15574 3204 15580
rect 1224 15510 1230 15574
rect 1294 15528 3134 15574
rect 1294 15510 1798 15528
rect 1224 15504 1798 15510
rect 1768 15472 1798 15504
rect 1854 15510 3134 15528
rect 3198 15510 3204 15574
rect 1854 15504 3204 15510
rect 124168 15574 124380 15646
rect 124168 15510 124310 15574
rect 124374 15510 124380 15574
rect 124168 15504 124380 15510
rect 136816 15574 137572 15580
rect 136816 15528 137502 15574
rect 1854 15472 1980 15504
rect 1768 15368 1980 15472
rect 136816 15472 136944 15528
rect 137000 15510 137502 15528
rect 137566 15510 137572 15574
rect 137000 15504 137572 15510
rect 137000 15472 137028 15504
rect 15205 15427 15271 15430
rect 27450 15427 27516 15430
rect 15205 15425 27516 15427
rect 15205 15369 15210 15425
rect 15266 15369 27455 15425
rect 27511 15369 27516 15425
rect 15205 15367 27516 15369
rect 136816 15368 137028 15472
rect 15205 15364 15271 15367
rect 27450 15364 27516 15367
rect 29865 15172 29963 15197
rect 32361 15172 32459 15197
rect 34857 15172 34955 15197
rect 37353 15172 37451 15197
rect 39849 15172 39947 15197
rect 42345 15172 42443 15197
rect 44841 15172 44939 15197
rect 47337 15172 47435 15197
rect 49833 15172 49931 15197
rect 52329 15172 52427 15197
rect 54825 15172 54923 15197
rect 57321 15172 57419 15197
rect 59817 15172 59915 15197
rect 62313 15172 62411 15197
rect 64809 15172 64907 15197
rect 67305 15172 67403 15197
rect 69801 15172 69899 15197
rect 72297 15172 72395 15197
rect 74793 15172 74891 15197
rect 77289 15172 77387 15197
rect 79785 15172 79883 15197
rect 82281 15172 82379 15197
rect 84777 15172 84875 15197
rect 87273 15172 87371 15197
rect 89769 15172 89867 15197
rect 92265 15172 92363 15197
rect 94761 15172 94859 15197
rect 97257 15172 97355 15197
rect 99753 15172 99851 15197
rect 102249 15172 102347 15197
rect 104745 15172 104843 15197
rect 107241 15172 107339 15197
rect 29784 15166 30094 15172
rect 32232 15166 32716 15172
rect 29784 15102 29926 15166
rect 29990 15102 30062 15166
rect 30126 15102 30132 15166
rect 32232 15102 32510 15166
rect 32574 15102 32646 15166
rect 32710 15102 32716 15166
rect 29784 15096 30094 15102
rect 32232 15096 32716 15102
rect 34816 15166 35164 15172
rect 34816 15102 34958 15166
rect 35022 15102 35094 15166
rect 35158 15102 35164 15166
rect 34816 15096 35164 15102
rect 37264 15166 37574 15172
rect 39848 15166 40196 15172
rect 37264 15102 37406 15166
rect 37470 15102 37542 15166
rect 37606 15102 37612 15166
rect 39848 15102 39990 15166
rect 40054 15102 40126 15166
rect 40190 15102 40196 15166
rect 37264 15096 37574 15102
rect 39848 15096 40196 15102
rect 42296 15166 42606 15172
rect 44744 15166 45054 15172
rect 47328 15166 47676 15172
rect 42296 15102 42438 15166
rect 42502 15102 42574 15166
rect 42638 15102 42644 15166
rect 44744 15102 44886 15166
rect 44950 15102 45022 15166
rect 45086 15102 45092 15166
rect 47328 15102 47470 15166
rect 47534 15102 47606 15166
rect 47670 15102 47676 15166
rect 42296 15096 42606 15102
rect 44744 15096 45054 15102
rect 47328 15096 47676 15102
rect 49776 15166 50222 15172
rect 52224 15166 52572 15172
rect 49776 15102 49918 15166
rect 49982 15102 50190 15166
rect 50254 15102 50260 15166
rect 52224 15102 52366 15166
rect 52430 15102 52502 15166
rect 52566 15102 52572 15166
rect 49776 15096 50222 15102
rect 52224 15096 52572 15102
rect 54808 15166 55156 15172
rect 54808 15102 54950 15166
rect 55014 15102 55086 15166
rect 55150 15102 55156 15166
rect 54808 15096 55156 15102
rect 57256 15166 57566 15172
rect 59704 15166 60014 15172
rect 62288 15166 62636 15172
rect 57256 15102 57398 15166
rect 57462 15102 57534 15166
rect 57598 15102 57604 15166
rect 59704 15102 59846 15166
rect 59910 15102 59982 15166
rect 60046 15102 60052 15166
rect 62288 15102 62430 15166
rect 62494 15102 62566 15166
rect 62630 15102 62636 15166
rect 57256 15096 57566 15102
rect 59704 15096 60014 15102
rect 62288 15096 62636 15102
rect 64736 15166 65046 15172
rect 67184 15166 67668 15172
rect 64736 15102 64878 15166
rect 64942 15102 65014 15166
rect 65078 15102 65084 15166
rect 67184 15102 67462 15166
rect 67526 15102 67598 15166
rect 67662 15102 67668 15166
rect 64736 15096 65046 15102
rect 67184 15096 67668 15102
rect 69768 15166 70078 15172
rect 72216 15166 72526 15172
rect 74664 15166 75148 15172
rect 69768 15102 69910 15166
rect 69974 15102 70046 15166
rect 70110 15102 70116 15166
rect 72216 15102 72358 15166
rect 72422 15102 72494 15166
rect 72558 15102 72564 15166
rect 74664 15102 74942 15166
rect 75006 15102 75078 15166
rect 75142 15102 75148 15166
rect 69768 15096 70078 15102
rect 72216 15096 72526 15102
rect 74664 15096 75148 15102
rect 77248 15166 77596 15172
rect 77248 15102 77390 15166
rect 77454 15102 77526 15166
rect 77590 15102 77596 15166
rect 77248 15096 77596 15102
rect 79696 15166 80006 15172
rect 82280 15166 82628 15172
rect 79696 15102 79838 15166
rect 79902 15102 79974 15166
rect 80038 15102 80044 15166
rect 82280 15102 82422 15166
rect 82486 15102 82558 15166
rect 82622 15102 82628 15166
rect 79696 15096 80006 15102
rect 82280 15096 82628 15102
rect 84728 15166 85038 15172
rect 87176 15166 87486 15172
rect 89760 15166 90108 15172
rect 84728 15102 84870 15166
rect 84934 15102 85006 15166
rect 85070 15102 85076 15166
rect 87176 15102 87318 15166
rect 87382 15102 87454 15166
rect 87518 15102 87524 15166
rect 89760 15102 89902 15166
rect 89966 15102 90038 15166
rect 90102 15102 90108 15166
rect 84728 15096 85038 15102
rect 87176 15096 87486 15102
rect 89760 15096 90108 15102
rect 92208 15166 92518 15172
rect 94656 15166 94966 15172
rect 97240 15166 97588 15172
rect 92208 15102 92350 15166
rect 92414 15102 92486 15166
rect 92550 15102 92556 15166
rect 94656 15102 94798 15166
rect 94862 15102 94934 15166
rect 94998 15102 95004 15166
rect 97240 15102 97382 15166
rect 97446 15102 97518 15166
rect 97582 15102 97588 15166
rect 92208 15096 92518 15102
rect 94656 15096 94966 15102
rect 97240 15096 97588 15102
rect 99688 15166 99998 15172
rect 102136 15166 102446 15172
rect 104720 15166 105068 15172
rect 99688 15102 99830 15166
rect 99894 15102 99966 15166
rect 100030 15102 100036 15166
rect 102136 15102 102278 15166
rect 102342 15102 102414 15166
rect 102478 15102 102484 15166
rect 104720 15102 104862 15166
rect 104926 15102 104998 15166
rect 105062 15102 105068 15166
rect 99688 15096 99998 15102
rect 102136 15096 102446 15102
rect 104720 15096 105068 15102
rect 107168 15166 107478 15172
rect 107168 15102 107310 15166
rect 107374 15102 107446 15166
rect 107510 15102 107516 15166
rect 107168 15096 107478 15102
rect 123086 14855 123152 14858
rect 123664 14855 123730 14858
rect 123086 14853 123730 14855
rect 123086 14797 123091 14853
rect 123147 14797 123669 14853
rect 123725 14797 123730 14853
rect 123086 14795 123730 14797
rect 123086 14792 123152 14795
rect 123664 14792 123730 14795
rect 124576 14782 124788 14900
rect 544 14758 3340 14764
rect 544 14694 550 14758
rect 614 14694 3340 14758
rect 544 14688 3340 14694
rect 3128 14628 3340 14688
rect 3944 14628 4156 14764
rect 3128 14552 4156 14628
rect 15096 14758 15308 14764
rect 15096 14694 15102 14758
rect 15166 14694 15308 14758
rect 15096 14622 15308 14694
rect 124576 14726 124614 14782
rect 124670 14764 124788 14782
rect 124670 14726 138796 14764
rect 124576 14688 138796 14726
rect 15096 14558 15102 14622
rect 15166 14558 15308 14622
rect 15096 14552 15308 14558
rect 21080 14622 21292 14628
rect 21080 14558 21086 14622
rect 21150 14558 21292 14622
rect 21080 14356 21292 14558
rect 22168 14356 22380 14628
rect 21080 14350 22380 14356
rect 21080 14286 22174 14350
rect 22238 14286 22380 14350
rect 21080 14280 22380 14286
rect 29648 14350 29996 14492
rect 29648 14286 29926 14350
rect 29990 14286 29996 14350
rect 29648 14280 29996 14286
rect 32232 14356 32444 14492
rect 34680 14356 34892 14492
rect 32232 14350 34892 14356
rect 32232 14286 32374 14350
rect 32438 14286 34822 14350
rect 34886 14286 34892 14350
rect 32232 14280 34892 14286
rect 37264 14416 42372 14492
rect 37264 14350 37476 14416
rect 37264 14286 37406 14350
rect 37470 14286 37476 14350
rect 37264 14280 37476 14286
rect 39712 14350 39924 14416
rect 39712 14286 39854 14350
rect 39918 14286 39924 14350
rect 39712 14280 39924 14286
rect 42160 14350 42372 14416
rect 42160 14286 42166 14350
rect 42230 14286 42372 14350
rect 42160 14280 42372 14286
rect 44744 14350 44956 14492
rect 44744 14286 44886 14350
rect 44950 14286 44956 14350
rect 44744 14280 44956 14286
rect 47192 14350 47404 14492
rect 47192 14286 47198 14350
rect 47262 14286 47404 14350
rect 47192 14280 47404 14286
rect 49640 14350 49852 14492
rect 49640 14286 49782 14350
rect 49846 14286 49852 14350
rect 49640 14280 49852 14286
rect 52224 14350 52436 14492
rect 52224 14286 52230 14350
rect 52294 14286 52436 14350
rect 52224 14280 52436 14286
rect 54672 14350 54884 14492
rect 54672 14286 54814 14350
rect 54878 14286 54884 14350
rect 54672 14280 54884 14286
rect 57120 14416 59916 14492
rect 57120 14350 57468 14416
rect 57120 14286 57398 14350
rect 57462 14286 57468 14350
rect 57120 14280 57468 14286
rect 59704 14350 59916 14416
rect 59704 14286 59846 14350
rect 59910 14286 59916 14350
rect 59704 14280 59916 14286
rect 62152 14356 62364 14492
rect 64600 14356 64948 14492
rect 62152 14350 64948 14356
rect 62152 14286 62294 14350
rect 62358 14286 64878 14350
rect 64942 14286 64948 14350
rect 62152 14280 64948 14286
rect 67184 14350 67396 14492
rect 67184 14286 67190 14350
rect 67254 14286 67396 14350
rect 67184 14280 67396 14286
rect 69632 14350 69844 14492
rect 69632 14286 69638 14350
rect 69702 14286 69844 14350
rect 69632 14280 69844 14286
rect 72080 14350 72428 14492
rect 72080 14286 72086 14350
rect 72150 14286 72222 14350
rect 72286 14286 72428 14350
rect 72080 14280 72428 14286
rect 74664 14356 74876 14492
rect 77112 14486 77324 14492
rect 77112 14422 77118 14486
rect 77182 14422 77324 14486
rect 74664 14350 77052 14356
rect 74664 14286 74806 14350
rect 74870 14286 76982 14350
rect 77046 14286 77052 14350
rect 74664 14280 77052 14286
rect 77112 14350 77324 14422
rect 77112 14286 77254 14350
rect 77318 14286 77324 14350
rect 77112 14280 77324 14286
rect 79696 14350 79908 14492
rect 79696 14286 79838 14350
rect 79902 14286 79908 14350
rect 79696 14280 79908 14286
rect 82144 14350 82356 14492
rect 82144 14286 82286 14350
rect 82350 14286 82356 14350
rect 82144 14280 82356 14286
rect 84592 14350 84804 14492
rect 84592 14286 84598 14350
rect 84662 14286 84804 14350
rect 84592 14280 84804 14286
rect 87176 14356 87388 14492
rect 89624 14356 89836 14492
rect 87176 14350 89836 14356
rect 87176 14286 87318 14350
rect 87382 14286 89630 14350
rect 89694 14286 89836 14350
rect 87176 14280 89836 14286
rect 92072 14350 92284 14492
rect 92072 14286 92214 14350
rect 92278 14286 92284 14350
rect 92072 14280 92284 14286
rect 94656 14350 94868 14492
rect 94656 14286 94662 14350
rect 94726 14286 94868 14350
rect 94656 14280 94868 14286
rect 97104 14350 97316 14492
rect 97104 14286 97246 14350
rect 97310 14286 97316 14350
rect 97104 14280 97316 14286
rect 99552 14350 99900 14492
rect 99552 14286 99694 14350
rect 99758 14286 99900 14350
rect 99552 14280 99900 14286
rect 102136 14350 102348 14492
rect 102136 14286 102278 14350
rect 102342 14286 102348 14350
rect 102136 14280 102348 14286
rect 104584 14356 104796 14492
rect 107032 14356 107380 14492
rect 104584 14350 107380 14356
rect 104584 14286 104726 14350
rect 104790 14286 107310 14350
rect 107374 14286 107380 14350
rect 104584 14280 107380 14286
rect 124168 14350 124516 14356
rect 124168 14286 124446 14350
rect 124510 14286 124516 14350
rect 124168 14280 124516 14286
rect 124168 14078 124380 14280
rect 15205 14013 15271 14016
rect 27698 14013 27764 14016
rect 15205 14011 27764 14013
rect 15205 13955 15210 14011
rect 15266 13955 27703 14011
rect 27759 13955 27764 14011
rect 124168 14014 124174 14078
rect 124238 14014 124380 14078
rect 124168 14008 124380 14014
rect 15205 13953 27764 13955
rect 15205 13950 15271 13953
rect 27698 13950 27764 13953
rect 1224 13942 1980 13948
rect 1224 13878 1230 13942
rect 1294 13878 1980 13942
rect 1224 13872 1980 13878
rect 1768 13848 1980 13872
rect 1768 13792 1798 13848
rect 1854 13812 1980 13848
rect 136816 13942 137572 13948
rect 136816 13878 137502 13942
rect 137566 13878 137572 13942
rect 136816 13872 137572 13878
rect 136816 13848 137028 13872
rect 1854 13806 3204 13812
rect 1854 13792 3134 13806
rect 1768 13742 3134 13792
rect 3198 13742 3204 13806
rect 1768 13736 3204 13742
rect 136816 13792 136944 13848
rect 137000 13792 137028 13848
rect 136816 13736 137028 13792
rect 29784 13670 29996 13676
rect 29784 13606 29926 13670
rect 29990 13606 29996 13670
rect 29784 13600 29996 13606
rect 32232 13670 32444 13676
rect 32232 13606 32374 13670
rect 32438 13606 32444 13670
rect 32232 13600 32444 13606
rect 34680 13670 34892 13676
rect 34680 13606 34686 13670
rect 34750 13606 34822 13670
rect 34886 13606 34892 13670
rect 34680 13600 34892 13606
rect 37264 13670 37476 13676
rect 37264 13606 37406 13670
rect 37470 13606 37476 13670
rect 29795 13534 29996 13600
rect 29795 13487 29926 13534
rect 29920 13470 29926 13487
rect 29990 13470 29996 13534
rect 32291 13534 32444 13600
rect 32291 13487 32374 13534
rect 29920 13464 29996 13470
rect 32368 13470 32374 13487
rect 32438 13470 32444 13534
rect 34787 13487 34885 13600
rect 37264 13534 37476 13606
rect 32368 13464 32444 13470
rect 37264 13470 37270 13534
rect 37334 13470 37476 13534
rect 37264 13464 37476 13470
rect 39712 13670 39924 13676
rect 39712 13606 39854 13670
rect 39918 13606 39924 13670
rect 39712 13534 39924 13606
rect 42160 13670 42508 13676
rect 42160 13606 42166 13670
rect 42230 13606 42508 13670
rect 42160 13600 42508 13606
rect 44744 13670 44956 13676
rect 44744 13606 44886 13670
rect 44950 13606 44956 13670
rect 44744 13600 44956 13606
rect 47192 13670 47404 13676
rect 47192 13606 47198 13670
rect 47262 13606 47404 13670
rect 47192 13600 47404 13606
rect 49640 13670 49988 13676
rect 49640 13606 49646 13670
rect 49710 13606 49782 13670
rect 49846 13606 49988 13670
rect 49640 13600 49988 13606
rect 52224 13670 52436 13676
rect 52224 13606 52230 13670
rect 52294 13606 52436 13670
rect 39712 13470 39718 13534
rect 39782 13470 39924 13534
rect 42275 13534 42508 13600
rect 42275 13487 42438 13534
rect 39712 13464 39924 13470
rect 42432 13470 42438 13487
rect 42502 13470 42508 13534
rect 44771 13534 44956 13600
rect 44771 13487 44886 13534
rect 42432 13464 42508 13470
rect 44880 13470 44886 13487
rect 44950 13470 44956 13534
rect 47267 13534 47404 13600
rect 47267 13487 47334 13534
rect 44880 13464 44956 13470
rect 47328 13470 47334 13487
rect 47398 13470 47404 13534
rect 49763 13487 49861 13600
rect 52224 13534 52436 13606
rect 54672 13670 54884 13676
rect 54672 13606 54814 13670
rect 54878 13606 54884 13670
rect 54672 13600 54884 13606
rect 57120 13670 57468 13676
rect 57120 13606 57398 13670
rect 57462 13606 57468 13670
rect 57120 13600 57468 13606
rect 59704 13670 59916 13676
rect 59704 13606 59846 13670
rect 59910 13606 59916 13670
rect 59704 13600 59916 13606
rect 62152 13670 62364 13676
rect 62152 13606 62294 13670
rect 62358 13606 62364 13670
rect 62152 13600 62364 13606
rect 47328 13464 47404 13470
rect 52224 13470 52230 13534
rect 52294 13470 52436 13534
rect 54755 13534 54884 13600
rect 54755 13487 54814 13534
rect 52224 13464 52436 13470
rect 54808 13470 54814 13487
rect 54878 13470 54884 13534
rect 57251 13534 57468 13600
rect 57251 13487 57398 13534
rect 54808 13464 54884 13470
rect 57392 13470 57398 13487
rect 57462 13470 57468 13534
rect 59747 13534 59916 13600
rect 59747 13487 59846 13534
rect 57392 13464 57468 13470
rect 59840 13470 59846 13487
rect 59910 13470 59916 13534
rect 62243 13534 62364 13600
rect 62243 13487 62294 13534
rect 59840 13464 59916 13470
rect 62288 13470 62294 13487
rect 62358 13470 62364 13534
rect 62288 13464 62364 13470
rect 64736 13670 64948 13676
rect 64736 13606 64878 13670
rect 64942 13606 64948 13670
rect 64736 13534 64948 13606
rect 67184 13670 67396 13676
rect 67184 13606 67190 13670
rect 67254 13606 67396 13670
rect 67184 13600 67396 13606
rect 69632 13670 72156 13676
rect 69632 13606 69638 13670
rect 69702 13606 69774 13670
rect 69838 13606 72086 13670
rect 72150 13606 72156 13670
rect 69632 13600 72156 13606
rect 72216 13670 72428 13676
rect 72216 13606 72222 13670
rect 72286 13606 72428 13670
rect 72216 13600 72428 13606
rect 74664 13670 74876 13676
rect 77014 13670 77324 13676
rect 74664 13606 74806 13670
rect 74870 13606 74876 13670
rect 76976 13606 76982 13670
rect 77046 13606 77118 13670
rect 77182 13606 77254 13670
rect 77318 13606 77324 13670
rect 74664 13600 74876 13606
rect 77014 13600 77324 13606
rect 79696 13670 82356 13676
rect 79696 13606 79838 13670
rect 79902 13606 82286 13670
rect 82350 13606 82356 13670
rect 79696 13600 82356 13606
rect 84592 13670 84940 13676
rect 84592 13606 84598 13670
rect 84662 13606 84940 13670
rect 84592 13600 84940 13606
rect 87176 13670 87388 13676
rect 87176 13606 87318 13670
rect 87382 13606 87388 13670
rect 87176 13600 87388 13606
rect 89624 13670 89836 13676
rect 89624 13606 89630 13670
rect 89694 13606 89836 13670
rect 89624 13600 89836 13606
rect 92072 13670 92420 13676
rect 92072 13606 92214 13670
rect 92278 13606 92420 13670
rect 92072 13600 92420 13606
rect 94656 13670 94868 13676
rect 94656 13606 94662 13670
rect 94726 13606 94868 13670
rect 94656 13600 94868 13606
rect 97104 13670 99900 13676
rect 97104 13606 97246 13670
rect 97310 13606 99694 13670
rect 99758 13606 99900 13670
rect 97104 13600 99900 13606
rect 102136 13670 104796 13676
rect 102136 13606 102278 13670
rect 102342 13606 104726 13670
rect 104790 13606 104796 13670
rect 102136 13600 104796 13606
rect 107168 13670 107380 13676
rect 107168 13606 107310 13670
rect 107374 13606 107380 13670
rect 107168 13600 107380 13606
rect 64736 13470 64742 13534
rect 64806 13470 64948 13534
rect 67235 13534 67396 13600
rect 67235 13487 67326 13534
rect 64736 13464 64948 13470
rect 67320 13470 67326 13487
rect 67390 13470 67396 13534
rect 69731 13487 69829 13600
rect 72227 13534 72428 13600
rect 72227 13487 72358 13534
rect 67320 13464 67396 13470
rect 72352 13470 72358 13487
rect 72422 13470 72428 13534
rect 74723 13534 74876 13600
rect 74723 13487 74806 13534
rect 72352 13464 72428 13470
rect 74800 13470 74806 13487
rect 74870 13470 74876 13534
rect 77219 13487 77317 13600
rect 79715 13534 79908 13600
rect 79715 13487 79838 13534
rect 74800 13464 74876 13470
rect 79832 13470 79838 13487
rect 79902 13470 79908 13534
rect 82211 13534 82356 13600
rect 82211 13487 82286 13534
rect 79832 13464 79908 13470
rect 82280 13470 82286 13487
rect 82350 13470 82356 13534
rect 84707 13534 84940 13600
rect 84707 13487 84870 13534
rect 82280 13464 82356 13470
rect 84864 13470 84870 13487
rect 84934 13470 84940 13534
rect 87203 13534 87388 13600
rect 87203 13487 87318 13534
rect 84864 13464 84940 13470
rect 87312 13470 87318 13487
rect 87382 13470 87388 13534
rect 89699 13534 89836 13600
rect 89699 13487 89766 13534
rect 87312 13464 87388 13470
rect 89760 13470 89766 13487
rect 89830 13470 89836 13534
rect 92195 13534 92420 13600
rect 92195 13487 92350 13534
rect 89760 13464 89836 13470
rect 92344 13470 92350 13487
rect 92414 13470 92420 13534
rect 94691 13534 94868 13600
rect 94691 13487 94798 13534
rect 92344 13464 92420 13470
rect 94792 13470 94798 13487
rect 94862 13470 94868 13534
rect 97187 13534 97316 13600
rect 97187 13487 97246 13534
rect 94792 13464 94868 13470
rect 97240 13470 97246 13487
rect 97310 13470 97316 13534
rect 99683 13534 99900 13600
rect 99683 13487 99830 13534
rect 97240 13464 97316 13470
rect 99824 13470 99830 13487
rect 99894 13470 99900 13534
rect 102179 13534 102348 13600
rect 102179 13487 102278 13534
rect 99824 13464 99900 13470
rect 102272 13470 102278 13487
rect 102342 13470 102348 13534
rect 104675 13534 104796 13600
rect 104675 13487 104726 13534
rect 102272 13464 102348 13470
rect 104720 13470 104726 13487
rect 104790 13470 104796 13534
rect 107171 13534 107380 13600
rect 124576 13654 124788 13676
rect 124576 13598 124614 13654
rect 124670 13598 124788 13654
rect 107171 13487 107310 13534
rect 104720 13464 104796 13470
rect 107304 13470 107310 13487
rect 107374 13470 107380 13534
rect 123006 13585 123072 13588
rect 123664 13585 123730 13588
rect 123006 13583 123730 13585
rect 123006 13527 123011 13583
rect 123067 13527 123669 13583
rect 123725 13527 123730 13583
rect 123006 13525 123730 13527
rect 123006 13522 123072 13525
rect 123664 13522 123730 13525
rect 124576 13540 124788 13598
rect 124576 13534 124924 13540
rect 107304 13464 107380 13470
rect 124576 13470 124854 13534
rect 124918 13470 124924 13534
rect 124576 13464 124924 13470
rect 3128 13398 3340 13404
rect 3128 13334 3134 13398
rect 3198 13334 3340 13398
rect 3128 13268 3340 13334
rect 3944 13268 4156 13404
rect 3128 13192 4156 13268
rect 15096 13398 15308 13404
rect 15096 13334 15238 13398
rect 15302 13334 15308 13398
rect 15096 13262 15308 13334
rect 15096 13198 15238 13262
rect 15302 13198 15308 13262
rect 15096 13192 15308 13198
rect 29512 13261 29724 13404
rect 29920 13263 30132 13268
rect 29512 13205 29562 13261
rect 29618 13205 29724 13261
rect 29512 13132 29724 13205
rect 29795 13262 30132 13263
rect 29795 13198 30062 13262
rect 30126 13198 30132 13262
rect 29795 13192 30132 13198
rect 31960 13261 32172 13404
rect 34408 13328 34756 13404
rect 32368 13263 32580 13268
rect 31960 13205 32058 13261
rect 32114 13205 32172 13261
rect 29795 13165 29996 13192
rect 21080 12996 21292 13132
rect 22168 13126 22380 13132
rect 22168 13062 22310 13126
rect 22374 13062 22380 13126
rect 22168 12996 22380 13062
rect 28968 13126 29724 13132
rect 28968 13062 28974 13126
rect 29038 13062 29724 13126
rect 28968 13056 29724 13062
rect 29920 13132 29996 13165
rect 29920 13126 30094 13132
rect 31960 13126 32172 13205
rect 32291 13262 32580 13263
rect 32291 13198 32510 13262
rect 32574 13198 32580 13262
rect 32291 13192 32580 13198
rect 34408 13261 34631 13328
rect 34408 13205 34554 13261
rect 34610 13205 34631 13261
rect 32291 13165 32444 13192
rect 29920 13062 30062 13126
rect 30126 13062 30132 13126
rect 31960 13062 31966 13126
rect 32030 13062 32172 13126
rect 29920 13056 30094 13062
rect 31960 13056 32172 13062
rect 32368 13132 32444 13165
rect 34408 13184 34631 13205
rect 32368 13126 32542 13132
rect 34408 13126 34620 13184
rect 32368 13062 32510 13126
rect 32574 13062 32580 13126
rect 34408 13062 34414 13126
rect 34478 13062 34620 13126
rect 34787 13132 34885 13263
rect 36992 13261 37204 13404
rect 36992 13205 37050 13261
rect 37106 13205 37204 13261
rect 34787 13126 35028 13132
rect 34787 13094 34822 13126
rect 32368 13056 32542 13062
rect 34408 13056 34620 13062
rect 34816 13062 34822 13094
rect 34886 13062 34958 13126
rect 35022 13062 35028 13126
rect 34816 13056 35028 13062
rect 36992 13126 37204 13205
rect 36992 13062 36998 13126
rect 37062 13062 37204 13126
rect 36992 13056 37204 13062
rect 37264 13262 37612 13268
rect 37264 13198 37542 13262
rect 37606 13198 37612 13262
rect 37264 13192 37612 13198
rect 39440 13261 39652 13404
rect 41888 13328 42236 13404
rect 39440 13205 39546 13261
rect 39602 13205 39652 13261
rect 37264 13126 37476 13192
rect 37264 13062 37406 13126
rect 37470 13062 37476 13126
rect 37264 13056 37476 13062
rect 39440 13126 39652 13205
rect 39440 13062 39446 13126
rect 39510 13062 39652 13126
rect 39440 13056 39652 13062
rect 39712 13262 40060 13268
rect 39712 13198 39990 13262
rect 40054 13198 40060 13262
rect 39712 13192 40060 13198
rect 41888 13261 42119 13328
rect 42432 13263 42644 13268
rect 41888 13205 42042 13261
rect 42098 13205 42119 13261
rect 39712 13126 39924 13192
rect 41888 13184 42119 13205
rect 42275 13262 42644 13263
rect 42275 13198 42574 13262
rect 42638 13198 42644 13262
rect 42275 13192 42644 13198
rect 44472 13261 44684 13404
rect 44880 13263 45092 13268
rect 44472 13205 44538 13261
rect 44594 13205 44684 13261
rect 41888 13132 42100 13184
rect 42275 13165 42508 13192
rect 42432 13132 42508 13165
rect 44472 13132 44684 13205
rect 44771 13262 45092 13263
rect 44771 13198 45022 13262
rect 45086 13198 45092 13262
rect 44771 13192 45092 13198
rect 46920 13261 47132 13404
rect 49504 13398 49988 13404
rect 49504 13334 49918 13398
rect 49982 13334 49988 13398
rect 49504 13328 49988 13334
rect 47328 13263 47540 13268
rect 46920 13205 47034 13261
rect 47090 13205 47132 13261
rect 44771 13165 44956 13192
rect 39712 13062 39854 13126
rect 39918 13062 39924 13126
rect 39712 13056 39924 13062
rect 41752 13126 42100 13132
rect 41752 13062 41758 13126
rect 41822 13062 42100 13126
rect 41752 13056 42100 13062
rect 42296 13126 42508 13132
rect 42296 13062 42302 13126
rect 42366 13062 42508 13126
rect 42296 13056 42508 13062
rect 44200 13126 44684 13132
rect 44200 13062 44206 13126
rect 44270 13062 44684 13126
rect 44200 13056 44684 13062
rect 44880 13132 44956 13165
rect 46920 13132 47132 13205
rect 47267 13262 47540 13263
rect 47267 13198 47470 13262
rect 47534 13198 47540 13262
rect 47267 13192 47540 13198
rect 49504 13261 49607 13328
rect 49504 13205 49530 13261
rect 49586 13205 49607 13261
rect 47267 13165 47404 13192
rect 44880 13126 45054 13132
rect 46512 13126 47132 13132
rect 44880 13062 45022 13126
rect 45086 13062 45092 13126
rect 46512 13062 46518 13126
rect 46582 13062 47132 13126
rect 44880 13056 45054 13062
rect 46512 13056 47132 13062
rect 47328 13132 47404 13165
rect 49504 13184 49607 13205
rect 47328 13126 47502 13132
rect 47328 13062 47470 13126
rect 47534 13062 47540 13126
rect 47328 13056 47502 13062
rect 49504 13056 49580 13184
rect 49763 13132 49861 13263
rect 51952 13261 52164 13404
rect 51952 13205 52026 13261
rect 52082 13205 52164 13261
rect 49763 13126 50260 13132
rect 49763 13094 49782 13126
rect 49776 13062 49782 13094
rect 49846 13062 50190 13126
rect 50254 13062 50260 13126
rect 49776 13056 50260 13062
rect 51952 13126 52164 13205
rect 51952 13062 51958 13126
rect 52022 13062 52164 13126
rect 51952 13056 52164 13062
rect 52224 13262 52436 13268
rect 52224 13198 52366 13262
rect 52430 13198 52436 13262
rect 52224 13126 52436 13198
rect 52224 13062 52366 13126
rect 52430 13062 52436 13126
rect 52224 13056 52436 13062
rect 54400 13261 54612 13404
rect 56984 13328 57196 13404
rect 54808 13263 55020 13268
rect 54400 13205 54522 13261
rect 54578 13205 54612 13261
rect 54400 13126 54612 13205
rect 54755 13262 55020 13263
rect 54755 13198 54950 13262
rect 55014 13198 55020 13262
rect 54755 13192 55020 13198
rect 56984 13261 57095 13328
rect 57392 13263 57604 13268
rect 56984 13205 57018 13261
rect 57074 13205 57095 13261
rect 54755 13165 54884 13192
rect 54400 13062 54542 13126
rect 54606 13062 54612 13126
rect 54400 13056 54612 13062
rect 54808 13132 54884 13165
rect 56984 13184 57095 13205
rect 57251 13262 57604 13263
rect 57251 13198 57534 13262
rect 57598 13198 57604 13262
rect 57251 13192 57604 13198
rect 59432 13261 59644 13404
rect 59840 13263 60052 13268
rect 59432 13205 59514 13261
rect 59570 13205 59644 13261
rect 54808 13126 54982 13132
rect 56984 13126 57060 13184
rect 57251 13165 57468 13192
rect 57392 13132 57468 13165
rect 59432 13132 59644 13205
rect 59747 13262 60052 13263
rect 59747 13198 59982 13262
rect 60046 13198 60052 13262
rect 59747 13192 60052 13198
rect 61880 13261 62092 13404
rect 62288 13263 62500 13268
rect 61880 13205 62010 13261
rect 62066 13205 62092 13261
rect 59747 13165 59916 13192
rect 54808 13062 54950 13126
rect 55014 13062 55020 13126
rect 56984 13062 56990 13126
rect 57054 13062 57060 13126
rect 54808 13056 54982 13062
rect 56984 13056 57060 13062
rect 57256 13126 57468 13132
rect 57256 13062 57262 13126
rect 57326 13062 57468 13126
rect 57256 13056 57468 13062
rect 59296 13126 59644 13132
rect 59296 13062 59302 13126
rect 59366 13062 59644 13126
rect 59296 13056 59644 13062
rect 59840 13132 59916 13165
rect 59840 13126 60014 13132
rect 61880 13126 62092 13205
rect 62243 13262 62500 13263
rect 62243 13198 62430 13262
rect 62494 13198 62500 13262
rect 62243 13192 62500 13198
rect 64464 13261 64676 13404
rect 64464 13205 64506 13261
rect 64562 13205 64676 13261
rect 62243 13165 62364 13192
rect 59840 13062 59982 13126
rect 60046 13062 60052 13126
rect 61880 13062 61886 13126
rect 61950 13062 62092 13126
rect 59840 13056 60014 13062
rect 61880 13056 62092 13062
rect 62288 13132 62364 13165
rect 62288 13126 62462 13132
rect 64464 13126 64676 13205
rect 62288 13062 62430 13126
rect 62494 13062 62500 13126
rect 64464 13062 64470 13126
rect 64534 13062 64676 13126
rect 62288 13056 62462 13062
rect 64464 13056 64676 13062
rect 64736 13262 65084 13268
rect 64736 13198 65014 13262
rect 65078 13198 65084 13262
rect 64736 13192 65084 13198
rect 66912 13261 67124 13404
rect 69360 13328 69708 13404
rect 67320 13263 67532 13268
rect 66912 13205 67002 13261
rect 67058 13205 67124 13261
rect 64736 13126 64948 13192
rect 64736 13062 64878 13126
rect 64942 13062 64948 13126
rect 64736 13056 64948 13062
rect 66912 13126 67124 13205
rect 67235 13262 67532 13263
rect 67235 13198 67462 13262
rect 67526 13198 67532 13262
rect 67235 13192 67532 13198
rect 69360 13261 69575 13328
rect 69360 13205 69498 13261
rect 69554 13205 69575 13261
rect 67235 13165 67396 13192
rect 66912 13062 66918 13126
rect 66982 13062 67124 13126
rect 66912 13056 67124 13062
rect 67320 13132 67396 13165
rect 69360 13184 69575 13205
rect 67320 13126 67494 13132
rect 69360 13126 69572 13184
rect 67320 13062 67462 13126
rect 67526 13062 67532 13126
rect 69360 13062 69502 13126
rect 69566 13062 69572 13126
rect 69731 13132 69829 13263
rect 71944 13261 72156 13404
rect 72352 13263 72564 13268
rect 71944 13205 71994 13261
rect 72050 13205 72156 13261
rect 69731 13126 69942 13132
rect 71944 13126 72156 13205
rect 72227 13262 72564 13263
rect 72227 13198 72494 13262
rect 72558 13198 72564 13262
rect 72227 13192 72564 13198
rect 74392 13261 74604 13404
rect 76840 13328 77188 13404
rect 74800 13263 75012 13268
rect 74392 13205 74490 13261
rect 74546 13205 74604 13261
rect 72227 13165 72428 13192
rect 69731 13094 69910 13126
rect 67320 13056 67494 13062
rect 69360 13056 69572 13062
rect 69768 13062 69910 13094
rect 69974 13062 69980 13126
rect 71944 13062 71950 13126
rect 72014 13062 72156 13126
rect 69768 13056 69942 13062
rect 71944 13056 72156 13062
rect 72352 13132 72428 13165
rect 72352 13126 72526 13132
rect 74392 13126 74604 13205
rect 74723 13262 75012 13263
rect 74723 13198 74942 13262
rect 75006 13198 75012 13262
rect 74723 13192 75012 13198
rect 76840 13261 77063 13328
rect 76840 13205 76986 13261
rect 77042 13205 77063 13261
rect 74723 13165 74876 13192
rect 72352 13062 72494 13126
rect 72558 13062 72564 13126
rect 74392 13062 74398 13126
rect 74462 13062 74604 13126
rect 72352 13056 72526 13062
rect 74392 13056 74604 13062
rect 74800 13132 74876 13165
rect 76840 13184 77063 13205
rect 74800 13126 74974 13132
rect 76840 13126 77052 13184
rect 74800 13062 74942 13126
rect 75006 13062 75012 13126
rect 76840 13062 76846 13126
rect 76910 13062 77052 13126
rect 77219 13132 77317 13263
rect 79424 13261 79636 13404
rect 79832 13263 80044 13268
rect 79424 13205 79482 13261
rect 79538 13205 79636 13261
rect 77219 13126 77460 13132
rect 77219 13094 77254 13126
rect 74800 13056 74974 13062
rect 76840 13056 77052 13062
rect 77248 13062 77254 13094
rect 77318 13062 77390 13126
rect 77454 13062 77460 13126
rect 77248 13056 77460 13062
rect 79424 13126 79636 13205
rect 79715 13262 80044 13263
rect 79715 13198 79974 13262
rect 80038 13198 80044 13262
rect 79715 13192 80044 13198
rect 81872 13261 82084 13404
rect 84320 13328 84668 13404
rect 82280 13263 82492 13268
rect 81872 13205 81978 13261
rect 82034 13205 82084 13261
rect 79715 13165 79908 13192
rect 79424 13062 79430 13126
rect 79494 13062 79636 13126
rect 79424 13056 79636 13062
rect 79832 13132 79908 13165
rect 79832 13126 80006 13132
rect 81872 13126 82084 13205
rect 82211 13262 82492 13263
rect 82211 13198 82422 13262
rect 82486 13198 82492 13262
rect 82211 13192 82492 13198
rect 84320 13261 84551 13328
rect 84864 13263 85076 13268
rect 84320 13205 84474 13261
rect 84530 13205 84551 13261
rect 82211 13165 82356 13192
rect 79832 13062 79974 13126
rect 80038 13062 80044 13126
rect 81872 13062 81878 13126
rect 81942 13062 82084 13126
rect 79832 13056 80006 13062
rect 81872 13056 82084 13062
rect 82280 13132 82356 13165
rect 84320 13184 84551 13205
rect 84707 13262 85076 13263
rect 84707 13198 85006 13262
rect 85070 13198 85076 13262
rect 84707 13192 85076 13198
rect 86904 13261 87116 13404
rect 87312 13263 87524 13268
rect 86904 13205 86970 13261
rect 87026 13205 87116 13261
rect 82280 13126 82454 13132
rect 84320 13126 84532 13184
rect 84707 13165 84940 13192
rect 84864 13132 84940 13165
rect 82280 13062 82422 13126
rect 82486 13062 82492 13126
rect 84320 13062 84326 13126
rect 84390 13062 84532 13126
rect 82280 13056 82454 13062
rect 84320 13056 84532 13062
rect 84728 13126 84940 13132
rect 84728 13062 84734 13126
rect 84798 13062 84940 13126
rect 84728 13056 84940 13062
rect 86904 13126 87116 13205
rect 87203 13262 87524 13263
rect 87203 13198 87454 13262
rect 87518 13198 87524 13262
rect 87203 13192 87524 13198
rect 89352 13261 89564 13404
rect 91936 13328 92148 13404
rect 89760 13263 89972 13268
rect 89352 13205 89466 13261
rect 89522 13205 89564 13261
rect 87203 13165 87388 13192
rect 86904 13062 86910 13126
rect 86974 13062 87116 13126
rect 86904 13056 87116 13062
rect 87312 13132 87388 13165
rect 89352 13132 89564 13205
rect 89699 13262 89972 13263
rect 89699 13198 89902 13262
rect 89966 13198 89972 13262
rect 89699 13192 89972 13198
rect 91936 13261 92039 13328
rect 92344 13263 92556 13268
rect 91936 13205 91962 13261
rect 92018 13205 92039 13261
rect 89699 13165 89836 13192
rect 87312 13126 87486 13132
rect 89080 13126 89564 13132
rect 87312 13062 87454 13126
rect 87518 13062 87524 13126
rect 89080 13062 89086 13126
rect 89150 13062 89564 13126
rect 87312 13056 87486 13062
rect 89080 13056 89564 13062
rect 89760 13132 89836 13165
rect 91936 13184 92039 13205
rect 92195 13262 92556 13263
rect 92195 13198 92486 13262
rect 92550 13198 92556 13262
rect 92195 13192 92556 13198
rect 94384 13261 94596 13404
rect 94792 13263 95004 13268
rect 94384 13205 94458 13261
rect 94514 13205 94596 13261
rect 89760 13126 89934 13132
rect 91936 13126 92012 13184
rect 92195 13165 92420 13192
rect 92344 13132 92420 13165
rect 89760 13062 89902 13126
rect 89966 13062 89972 13126
rect 91936 13062 91942 13126
rect 92006 13062 92012 13126
rect 89760 13056 89934 13062
rect 91936 13056 92012 13062
rect 92208 13126 92420 13132
rect 92208 13062 92214 13126
rect 92278 13062 92420 13126
rect 92208 13056 92420 13062
rect 94384 13126 94596 13205
rect 94691 13262 95004 13263
rect 94691 13198 94934 13262
rect 94998 13198 95004 13262
rect 94691 13192 95004 13198
rect 96832 13261 97044 13404
rect 99416 13328 99628 13404
rect 97240 13263 97452 13268
rect 96832 13205 96954 13261
rect 97010 13205 97044 13261
rect 94691 13165 94868 13192
rect 94384 13062 94390 13126
rect 94454 13062 94596 13126
rect 94384 13056 94596 13062
rect 94792 13132 94868 13165
rect 94792 13126 94966 13132
rect 96832 13126 97044 13205
rect 97187 13262 97452 13263
rect 97187 13198 97382 13262
rect 97446 13198 97452 13262
rect 97187 13192 97452 13198
rect 99416 13261 99527 13328
rect 99824 13263 100036 13268
rect 99416 13205 99450 13261
rect 99506 13205 99527 13261
rect 97187 13165 97316 13192
rect 94792 13062 94934 13126
rect 94998 13062 95004 13126
rect 96832 13062 96838 13126
rect 96902 13062 97044 13126
rect 94792 13056 94966 13062
rect 96832 13056 97044 13062
rect 97240 13132 97316 13165
rect 99416 13184 99527 13205
rect 99683 13262 100036 13263
rect 99683 13198 99966 13262
rect 100030 13198 100036 13262
rect 99683 13192 100036 13198
rect 101864 13261 102076 13404
rect 102272 13263 102484 13268
rect 101864 13205 101946 13261
rect 102002 13205 102076 13261
rect 97240 13126 97414 13132
rect 99416 13126 99492 13184
rect 99683 13165 99900 13192
rect 99824 13132 99900 13165
rect 97240 13062 97382 13126
rect 97446 13062 97452 13126
rect 99416 13062 99422 13126
rect 99486 13062 99492 13126
rect 97240 13056 97414 13062
rect 99416 13056 99492 13062
rect 99688 13126 99900 13132
rect 99688 13062 99694 13126
rect 99758 13062 99900 13126
rect 99688 13056 99900 13062
rect 101864 13126 102076 13205
rect 102179 13262 102484 13263
rect 102179 13198 102414 13262
rect 102478 13198 102484 13262
rect 102179 13192 102484 13198
rect 104312 13261 104524 13404
rect 104720 13263 104932 13268
rect 104312 13205 104442 13261
rect 104498 13205 104524 13261
rect 102179 13165 102348 13192
rect 101864 13062 101870 13126
rect 101934 13062 102076 13126
rect 101864 13056 102076 13062
rect 102272 13132 102348 13165
rect 102272 13126 102446 13132
rect 104312 13126 104524 13205
rect 104675 13262 104932 13263
rect 104675 13198 104862 13262
rect 104926 13198 104932 13262
rect 104675 13192 104932 13198
rect 106896 13261 107108 13404
rect 107304 13263 107516 13268
rect 106896 13205 106938 13261
rect 106994 13205 107108 13261
rect 104675 13165 104796 13192
rect 102272 13062 102414 13126
rect 102478 13062 102484 13126
rect 104312 13062 104318 13126
rect 104382 13062 104524 13126
rect 102272 13056 102446 13062
rect 104312 13056 104524 13062
rect 104720 13132 104796 13165
rect 104720 13126 104894 13132
rect 106896 13126 107108 13205
rect 107171 13262 107516 13263
rect 107171 13198 107446 13262
rect 107510 13198 107516 13262
rect 107171 13192 107516 13198
rect 107171 13165 107380 13192
rect 104720 13062 104862 13126
rect 104926 13062 104932 13126
rect 106896 13062 106902 13126
rect 106966 13062 107108 13126
rect 104720 13056 104894 13062
rect 106896 13056 107108 13062
rect 107304 13132 107380 13165
rect 107304 13126 107478 13132
rect 107304 13062 107446 13126
rect 107510 13062 107516 13126
rect 107304 13056 107478 13062
rect 21080 12920 22380 12996
rect 69768 12996 69844 13056
rect 69768 12990 70116 12996
rect 69768 12926 70046 12990
rect 70110 12926 70116 12990
rect 69768 12920 70116 12926
rect 124168 12854 124380 12860
rect 124168 12790 124310 12854
rect 124374 12790 124380 12854
rect 124168 12718 124380 12790
rect 124168 12654 124310 12718
rect 124374 12654 124380 12718
rect 124168 12648 124380 12654
rect 15205 12599 15271 12602
rect 27574 12599 27640 12602
rect 15205 12597 27640 12599
rect 15205 12541 15210 12597
rect 15266 12541 27579 12597
rect 27635 12541 27640 12597
rect 15205 12539 27640 12541
rect 15205 12536 15271 12539
rect 27574 12536 27640 12539
rect 29648 12582 30132 12588
rect 29648 12518 30062 12582
rect 30126 12518 30132 12582
rect 29648 12512 30132 12518
rect 32096 12582 32580 12588
rect 32096 12518 32510 12582
rect 32574 12518 32580 12582
rect 32096 12512 32580 12518
rect 34544 12582 34892 12588
rect 34544 12518 34822 12582
rect 34886 12518 34892 12582
rect 1768 12180 1980 12316
rect 29648 12310 29860 12512
rect 29648 12246 29790 12310
rect 29854 12246 29860 12310
rect 29648 12240 29860 12246
rect 32096 12310 32308 12512
rect 32096 12246 32238 12310
rect 32302 12246 32308 12310
rect 32096 12240 32308 12246
rect 34544 12310 34892 12518
rect 34544 12246 34822 12310
rect 34886 12246 34892 12310
rect 34544 12240 34892 12246
rect 37128 12582 37476 12588
rect 37128 12518 37406 12582
rect 37470 12518 37476 12582
rect 37128 12512 37476 12518
rect 39576 12582 39924 12588
rect 39576 12518 39854 12582
rect 39918 12518 39924 12582
rect 39576 12512 39924 12518
rect 42160 12582 42372 12588
rect 42160 12518 42302 12582
rect 42366 12518 42372 12582
rect 37128 12316 37340 12512
rect 39576 12316 39788 12512
rect 37128 12310 37476 12316
rect 37128 12246 37406 12310
rect 37470 12246 37476 12310
rect 37128 12240 37476 12246
rect 39576 12310 39924 12316
rect 39576 12246 39854 12310
rect 39918 12246 39924 12310
rect 39576 12240 39924 12246
rect 42160 12310 42372 12518
rect 42160 12246 42166 12310
rect 42230 12246 42372 12310
rect 42160 12240 42372 12246
rect 44608 12582 45092 12588
rect 44608 12518 45022 12582
rect 45086 12518 45092 12582
rect 44608 12512 45092 12518
rect 47056 12582 47540 12588
rect 47056 12518 47470 12582
rect 47534 12518 47540 12582
rect 47056 12512 47540 12518
rect 49640 12582 49852 12588
rect 49640 12518 49782 12582
rect 49846 12518 49852 12582
rect 44608 12310 44820 12512
rect 44608 12246 44614 12310
rect 44678 12246 44820 12310
rect 44608 12240 44820 12246
rect 47056 12310 47268 12512
rect 49640 12316 49852 12518
rect 47056 12246 47198 12310
rect 47262 12246 47268 12310
rect 47056 12240 47268 12246
rect 49504 12310 49852 12316
rect 49504 12246 49510 12310
rect 49574 12246 49852 12310
rect 49504 12240 49852 12246
rect 52088 12582 52436 12588
rect 52088 12518 52366 12582
rect 52430 12518 52436 12582
rect 52088 12512 52436 12518
rect 54536 12582 55020 12588
rect 54536 12518 54950 12582
rect 55014 12518 55020 12582
rect 54536 12512 55020 12518
rect 57120 12582 57332 12588
rect 57120 12518 57262 12582
rect 57326 12518 57332 12582
rect 52088 12316 52300 12512
rect 54536 12316 54748 12512
rect 52088 12310 52436 12316
rect 54438 12310 54748 12316
rect 52088 12246 52366 12310
rect 52430 12246 52436 12310
rect 54400 12246 54406 12310
rect 54470 12246 54748 12310
rect 52088 12240 52436 12246
rect 54438 12240 54748 12246
rect 57120 12316 57332 12518
rect 59568 12582 60052 12588
rect 59568 12518 59982 12582
rect 60046 12518 60052 12582
rect 59568 12512 60052 12518
rect 62016 12582 62500 12588
rect 62016 12518 62430 12582
rect 62494 12518 62500 12582
rect 62016 12512 62500 12518
rect 64600 12582 64948 12588
rect 64600 12518 64878 12582
rect 64942 12518 64948 12582
rect 64600 12512 64948 12518
rect 67048 12582 67532 12588
rect 67048 12518 67462 12582
rect 67526 12518 67532 12582
rect 67048 12512 67532 12518
rect 69496 12582 69980 12588
rect 69496 12518 69910 12582
rect 69974 12518 69980 12582
rect 69496 12512 69980 12518
rect 72080 12582 72564 12588
rect 72080 12518 72494 12582
rect 72558 12518 72564 12582
rect 72080 12512 72564 12518
rect 74528 12582 75012 12588
rect 74528 12518 74942 12582
rect 75006 12518 75012 12582
rect 74528 12512 75012 12518
rect 76976 12582 77324 12588
rect 76976 12518 77254 12582
rect 77318 12518 77324 12582
rect 57120 12310 57604 12316
rect 57120 12246 57534 12310
rect 57598 12246 57604 12310
rect 57120 12240 57604 12246
rect 59568 12310 59780 12512
rect 59568 12246 59574 12310
rect 59638 12246 59780 12310
rect 59568 12240 59780 12246
rect 62016 12316 62228 12512
rect 64600 12316 64812 12512
rect 67048 12316 67260 12512
rect 69496 12316 69844 12512
rect 72080 12316 72292 12512
rect 62016 12310 62500 12316
rect 62016 12246 62430 12310
rect 62494 12246 62500 12310
rect 62016 12240 62500 12246
rect 64600 12310 64948 12316
rect 64600 12246 64878 12310
rect 64942 12246 64948 12310
rect 64600 12240 64948 12246
rect 67048 12310 67532 12316
rect 67048 12246 67462 12310
rect 67526 12246 67532 12310
rect 67048 12240 67532 12246
rect 69496 12310 69980 12316
rect 69496 12246 69910 12310
rect 69974 12246 69980 12310
rect 69496 12240 69980 12246
rect 72080 12310 72564 12316
rect 72080 12246 72494 12310
rect 72558 12246 72564 12310
rect 72080 12240 72564 12246
rect 74528 12310 74740 12512
rect 74528 12246 74670 12310
rect 74734 12246 74740 12310
rect 74528 12240 74740 12246
rect 76976 12310 77324 12518
rect 76976 12246 76982 12310
rect 77046 12246 77324 12310
rect 76976 12240 77324 12246
rect 79560 12582 80044 12588
rect 79560 12518 79974 12582
rect 80038 12518 80044 12582
rect 79560 12512 80044 12518
rect 82008 12582 82492 12588
rect 82008 12518 82422 12582
rect 82486 12518 82492 12582
rect 82008 12512 82492 12518
rect 84592 12582 84804 12588
rect 84592 12518 84734 12582
rect 84798 12518 84804 12582
rect 79560 12316 79772 12512
rect 82008 12316 82220 12512
rect 79560 12310 80044 12316
rect 79560 12246 79974 12310
rect 80038 12246 80044 12310
rect 79560 12240 80044 12246
rect 82008 12310 82492 12316
rect 82008 12246 82422 12310
rect 82486 12246 82492 12310
rect 82008 12240 82492 12246
rect 84592 12310 84804 12518
rect 84592 12246 84734 12310
rect 84798 12246 84804 12310
rect 84592 12240 84804 12246
rect 87040 12582 87524 12588
rect 87040 12518 87454 12582
rect 87518 12518 87524 12582
rect 87040 12512 87524 12518
rect 89488 12582 89972 12588
rect 89488 12518 89902 12582
rect 89966 12518 89972 12582
rect 89488 12512 89972 12518
rect 92072 12582 92284 12588
rect 92072 12518 92214 12582
rect 92278 12518 92284 12582
rect 87040 12310 87252 12512
rect 87040 12246 87046 12310
rect 87110 12246 87252 12310
rect 87040 12240 87252 12246
rect 89488 12310 89700 12512
rect 89488 12246 89630 12310
rect 89694 12246 89700 12310
rect 89488 12240 89700 12246
rect 92072 12316 92284 12518
rect 94520 12582 95004 12588
rect 94520 12518 94934 12582
rect 94998 12518 95004 12582
rect 94520 12512 95004 12518
rect 96968 12582 97452 12588
rect 96968 12518 97382 12582
rect 97446 12518 97452 12582
rect 96968 12512 97452 12518
rect 99552 12582 99764 12588
rect 99552 12518 99694 12582
rect 99758 12518 99764 12582
rect 94520 12316 94732 12512
rect 96968 12316 97180 12512
rect 92072 12310 92556 12316
rect 92072 12246 92486 12310
rect 92550 12246 92556 12310
rect 92072 12240 92556 12246
rect 94520 12310 95004 12316
rect 94520 12246 94934 12310
rect 94998 12246 95004 12310
rect 94520 12240 95004 12246
rect 96968 12310 97452 12316
rect 96968 12246 97382 12310
rect 97446 12246 97452 12310
rect 96968 12240 97452 12246
rect 99552 12310 99764 12518
rect 99552 12246 99694 12310
rect 99758 12246 99764 12310
rect 99552 12240 99764 12246
rect 102000 12582 102484 12588
rect 102000 12518 102414 12582
rect 102478 12518 102484 12582
rect 102000 12512 102484 12518
rect 104448 12582 104932 12588
rect 104448 12518 104862 12582
rect 104926 12518 104932 12582
rect 104448 12512 104932 12518
rect 107032 12582 107516 12588
rect 107032 12518 107446 12582
rect 107510 12518 107516 12582
rect 107032 12512 107516 12518
rect 102000 12310 102212 12512
rect 102000 12246 102006 12310
rect 102070 12246 102212 12310
rect 102000 12240 102212 12246
rect 104448 12310 104660 12512
rect 104448 12246 104454 12310
rect 104518 12246 104660 12310
rect 104448 12240 104660 12246
rect 107032 12316 107244 12512
rect 107032 12310 107516 12316
rect 107032 12246 107446 12310
rect 107510 12246 107516 12310
rect 107032 12240 107516 12246
rect 1224 12174 1980 12180
rect 1224 12110 1230 12174
rect 1294 12168 1980 12174
rect 1294 12112 1798 12168
rect 1854 12112 1980 12168
rect 1294 12110 1980 12112
rect 1224 12104 1980 12110
rect 1768 11968 1980 12104
rect 136816 12168 137028 12316
rect 136816 12112 136944 12168
rect 137000 12112 137028 12168
rect 136816 12044 137028 12112
rect 15096 12038 15308 12044
rect 15096 11974 15102 12038
rect 15166 11974 15308 12038
rect 15096 11766 15308 11974
rect 29648 12038 29996 12044
rect 29648 11974 29926 12038
rect 29990 11974 29996 12038
rect 29648 11968 29996 11974
rect 32096 12038 32444 12044
rect 32096 11974 32374 12038
rect 32438 11974 32444 12038
rect 32096 11968 32444 11974
rect 34544 12038 34892 12044
rect 34544 11974 34686 12038
rect 34750 11974 34892 12038
rect 29648 11902 29860 11968
rect 29648 11838 29654 11902
rect 29718 11838 29860 11902
rect 29648 11832 29860 11838
rect 32096 11902 32308 11968
rect 32096 11838 32102 11902
rect 32166 11838 32308 11902
rect 32096 11832 32308 11838
rect 34544 11902 34892 11974
rect 34544 11838 34686 11902
rect 34750 11838 34892 11902
rect 34544 11832 34892 11838
rect 37128 12038 37340 12044
rect 37128 11974 37270 12038
rect 37334 11974 37340 12038
rect 37128 11902 37340 11974
rect 37128 11838 37270 11902
rect 37334 11838 37340 11902
rect 37128 11832 37340 11838
rect 39576 12038 39788 12044
rect 39576 11974 39718 12038
rect 39782 11974 39788 12038
rect 39576 11902 39788 11974
rect 39576 11838 39718 11902
rect 39782 11838 39788 11902
rect 39576 11832 39788 11838
rect 42024 12038 42508 12044
rect 42024 11974 42438 12038
rect 42502 11974 42508 12038
rect 42024 11968 42508 11974
rect 44608 12038 44956 12044
rect 44608 11974 44886 12038
rect 44950 11974 44956 12038
rect 44608 11968 44956 11974
rect 47056 12038 47404 12044
rect 47056 11974 47334 12038
rect 47398 11974 47404 12038
rect 47056 11968 47404 11974
rect 49504 12038 49852 12044
rect 49504 11974 49646 12038
rect 49710 11974 49852 12038
rect 42024 11908 42372 11968
rect 44608 11908 44820 11968
rect 47056 11908 47268 11968
rect 49504 11908 49852 11974
rect 42024 11902 49852 11908
rect 42024 11838 42302 11902
rect 42366 11838 44750 11902
rect 44814 11838 47062 11902
rect 47126 11838 49782 11902
rect 49846 11838 49852 11902
rect 42024 11832 49852 11838
rect 52088 12038 52300 12044
rect 52088 11974 52230 12038
rect 52294 11974 52300 12038
rect 52088 11902 52300 11974
rect 52088 11838 52230 11902
rect 52294 11838 52300 11902
rect 52088 11832 52300 11838
rect 54536 12038 54884 12044
rect 54536 11974 54814 12038
rect 54878 11974 54884 12038
rect 54536 11968 54884 11974
rect 57120 12038 57468 12044
rect 57120 11974 57398 12038
rect 57462 11974 57468 12038
rect 57120 11968 57468 11974
rect 59568 12038 59916 12044
rect 59568 11974 59846 12038
rect 59910 11974 59916 12038
rect 59568 11968 59916 11974
rect 62016 12038 62364 12044
rect 62016 11974 62294 12038
rect 62358 11974 62364 12038
rect 62016 11968 62364 11974
rect 64600 12038 64812 12044
rect 64600 11974 64742 12038
rect 64806 11974 64812 12038
rect 54536 11908 54748 11968
rect 54536 11902 54884 11908
rect 54536 11838 54814 11902
rect 54878 11838 54884 11902
rect 54536 11832 54884 11838
rect 57120 11902 57332 11968
rect 57120 11838 57262 11902
rect 57326 11838 57332 11902
rect 57120 11832 57332 11838
rect 59568 11908 59780 11968
rect 62016 11908 62228 11968
rect 59568 11902 62228 11908
rect 59568 11838 59710 11902
rect 59774 11838 62158 11902
rect 62222 11838 62228 11902
rect 59568 11832 62228 11838
rect 64600 11908 64812 11974
rect 67048 12038 67396 12044
rect 67048 11974 67326 12038
rect 67390 11974 67396 12038
rect 67048 11968 67396 11974
rect 69496 12038 69844 12044
rect 69496 11974 69774 12038
rect 69838 11974 69844 12038
rect 69496 11968 69844 11974
rect 72080 12038 72428 12044
rect 72080 11974 72358 12038
rect 72422 11974 72428 12038
rect 72080 11968 72428 11974
rect 74528 12038 74876 12044
rect 74528 11974 74806 12038
rect 74870 11974 74876 12038
rect 74528 11968 74876 11974
rect 76976 12038 77324 12044
rect 76976 11974 77118 12038
rect 77182 11974 77324 12038
rect 67048 11908 67260 11968
rect 64600 11902 67260 11908
rect 64600 11838 64742 11902
rect 64806 11838 67190 11902
rect 67254 11838 67260 11902
rect 64600 11832 67260 11838
rect 69496 11908 69708 11968
rect 69496 11902 69844 11908
rect 69496 11838 69774 11902
rect 69838 11838 69844 11902
rect 69496 11832 69844 11838
rect 72080 11902 72292 11968
rect 72080 11838 72222 11902
rect 72286 11838 72292 11902
rect 72080 11832 72292 11838
rect 74528 11902 74740 11968
rect 74528 11838 74534 11902
rect 74598 11838 74740 11902
rect 74528 11832 74740 11838
rect 76976 11902 77324 11974
rect 76976 11838 77254 11902
rect 77318 11838 77324 11902
rect 76976 11832 77324 11838
rect 79560 12038 79908 12044
rect 79560 11974 79838 12038
rect 79902 11974 79908 12038
rect 79560 11968 79908 11974
rect 82008 12038 82356 12044
rect 82008 11974 82286 12038
rect 82350 11974 82356 12038
rect 82008 11968 82356 11974
rect 84456 12038 84940 12044
rect 84456 11974 84870 12038
rect 84934 11974 84940 12038
rect 84456 11968 84940 11974
rect 87040 12038 87388 12044
rect 87040 11974 87318 12038
rect 87382 11974 87388 12038
rect 87040 11968 87388 11974
rect 89488 12038 89836 12044
rect 89488 11974 89766 12038
rect 89830 11974 89836 12038
rect 89488 11968 89836 11974
rect 91936 12038 92420 12044
rect 91936 11974 92350 12038
rect 92414 11974 92420 12038
rect 91936 11968 92420 11974
rect 94520 12038 94868 12044
rect 94520 11974 94798 12038
rect 94862 11974 94868 12038
rect 94520 11968 94868 11974
rect 96968 12038 97316 12044
rect 96968 11974 97246 12038
rect 97310 11974 97316 12038
rect 96968 11968 97316 11974
rect 99552 12038 99900 12044
rect 99552 11974 99830 12038
rect 99894 11974 99900 12038
rect 99552 11968 99900 11974
rect 102000 12038 102348 12044
rect 102000 11974 102278 12038
rect 102342 11974 102348 12038
rect 102000 11968 102348 11974
rect 104448 12038 104796 12044
rect 104448 11974 104726 12038
rect 104790 11974 104796 12038
rect 104448 11968 104796 11974
rect 107032 12038 107380 12044
rect 107032 11974 107310 12038
rect 107374 11974 107380 12038
rect 107032 11968 107380 11974
rect 122926 12027 122992 12030
rect 123664 12027 123730 12030
rect 122926 12025 123730 12027
rect 122926 11969 122931 12025
rect 122987 11969 123669 12025
rect 123725 11969 123730 12025
rect 79560 11902 79772 11968
rect 79560 11838 79702 11902
rect 79766 11838 79772 11902
rect 79560 11832 79772 11838
rect 82008 11908 82220 11968
rect 84456 11908 84804 11968
rect 87040 11908 87252 11968
rect 82008 11902 87252 11908
rect 82008 11838 82150 11902
rect 82214 11838 84598 11902
rect 84662 11838 87182 11902
rect 87246 11838 87252 11902
rect 82008 11832 87252 11838
rect 89488 11908 89700 11968
rect 91936 11908 92284 11968
rect 89488 11902 92284 11908
rect 89488 11838 89494 11902
rect 89558 11838 92214 11902
rect 92278 11838 92284 11902
rect 89488 11832 92284 11838
rect 94520 11902 94732 11968
rect 94520 11838 94662 11902
rect 94726 11838 94732 11902
rect 94520 11832 94732 11838
rect 96968 11902 97180 11968
rect 96968 11838 97110 11902
rect 97174 11838 97180 11902
rect 96968 11832 97180 11838
rect 99552 11902 99764 11968
rect 99552 11838 99558 11902
rect 99622 11838 99764 11902
rect 99552 11832 99764 11838
rect 102000 11902 102212 11968
rect 102000 11838 102142 11902
rect 102206 11838 102212 11902
rect 102000 11832 102212 11838
rect 104448 11902 104660 11968
rect 104448 11838 104590 11902
rect 104654 11838 104660 11902
rect 104448 11832 104660 11838
rect 107032 11902 107244 11968
rect 122926 11967 123730 11969
rect 122926 11964 122992 11967
rect 123664 11964 123730 11967
rect 124576 11954 124788 12044
rect 136816 12038 137572 12044
rect 136816 11974 137502 12038
rect 137566 11974 137572 12038
rect 136816 11968 137572 11974
rect 124576 11908 124614 11954
rect 107032 11838 107174 11902
rect 107238 11838 107244 11902
rect 107032 11832 107244 11838
rect 124440 11902 124614 11908
rect 124440 11838 124446 11902
rect 124510 11898 124614 11902
rect 124670 11898 124788 11954
rect 124510 11838 124788 11898
rect 124440 11832 124788 11838
rect 15096 11702 15102 11766
rect 15166 11702 15308 11766
rect 15096 11696 15308 11702
rect 21080 11636 21292 11772
rect 22168 11766 22380 11772
rect 22168 11702 22174 11766
rect 22238 11702 22380 11766
rect 22168 11636 22380 11702
rect 21080 11560 22380 11636
rect 29784 11766 29996 11772
rect 29784 11702 29790 11766
rect 29854 11702 29996 11766
rect 29784 11560 29996 11702
rect 32232 11766 32444 11772
rect 32232 11702 32238 11766
rect 32302 11702 32444 11766
rect 32232 11560 32444 11702
rect 34680 11766 34892 11772
rect 34680 11702 34822 11766
rect 34886 11702 34892 11766
rect 34680 11560 34892 11702
rect 29784 11500 29860 11560
rect 32232 11500 32308 11560
rect 34816 11500 34892 11560
rect 37264 11766 37476 11772
rect 37264 11702 37406 11766
rect 37470 11702 37476 11766
rect 37264 11560 37476 11702
rect 39712 11766 39924 11772
rect 39712 11702 39854 11766
rect 39918 11702 39924 11766
rect 39712 11560 39924 11702
rect 42160 11766 42372 11772
rect 44646 11766 44956 11772
rect 42160 11702 42166 11766
rect 42230 11702 42372 11766
rect 44608 11702 44614 11766
rect 44678 11702 44956 11766
rect 42160 11560 42372 11702
rect 44646 11696 44956 11702
rect 44744 11560 44956 11696
rect 47192 11766 47404 11772
rect 49542 11766 49988 11772
rect 47192 11702 47198 11766
rect 47262 11702 47404 11766
rect 49504 11702 49510 11766
rect 49574 11702 49988 11766
rect 47192 11560 47404 11702
rect 49542 11696 49988 11702
rect 49640 11560 49988 11696
rect 52224 11766 52436 11772
rect 52224 11702 52366 11766
rect 52430 11702 52436 11766
rect 52224 11560 52436 11702
rect 54672 11560 54884 11772
rect 57120 11766 57566 11772
rect 59606 11766 59916 11772
rect 57120 11702 57534 11766
rect 57598 11702 57604 11766
rect 59568 11702 59574 11766
rect 59638 11702 59916 11766
rect 57120 11696 57566 11702
rect 59606 11696 59916 11702
rect 57120 11560 57468 11696
rect 59704 11560 59916 11696
rect 62152 11766 62462 11772
rect 64600 11766 64948 11772
rect 62152 11702 62430 11766
rect 62494 11702 62500 11766
rect 64600 11702 64878 11766
rect 64942 11702 64948 11766
rect 62152 11696 62462 11702
rect 62152 11560 62364 11696
rect 64600 11560 64948 11702
rect 67184 11766 67494 11772
rect 69632 11766 69942 11772
rect 72216 11766 72526 11772
rect 74664 11766 74876 11772
rect 77014 11766 77324 11772
rect 67184 11702 67462 11766
rect 67526 11702 67532 11766
rect 69632 11702 69910 11766
rect 69974 11702 69980 11766
rect 72216 11702 72494 11766
rect 72558 11702 72564 11766
rect 74664 11702 74670 11766
rect 74734 11702 74876 11766
rect 76976 11702 76982 11766
rect 77046 11702 77324 11766
rect 67184 11696 67494 11702
rect 69632 11696 69942 11702
rect 72216 11696 72526 11702
rect 67184 11560 67396 11696
rect 69632 11560 69844 11696
rect 72216 11560 72428 11696
rect 74664 11560 74876 11702
rect 77014 11696 77324 11702
rect 77112 11560 77324 11696
rect 79696 11766 80006 11772
rect 82144 11766 82454 11772
rect 84592 11766 84804 11772
rect 87078 11766 87388 11772
rect 79696 11702 79974 11766
rect 80038 11702 80044 11766
rect 82144 11702 82422 11766
rect 82486 11702 82492 11766
rect 84592 11702 84734 11766
rect 84798 11702 84804 11766
rect 87040 11702 87046 11766
rect 87110 11702 87388 11766
rect 79696 11696 80006 11702
rect 82144 11696 82454 11702
rect 79696 11560 79908 11696
rect 82144 11560 82356 11696
rect 84592 11560 84804 11702
rect 87078 11696 87388 11702
rect 37264 11500 37340 11560
rect 39712 11500 39788 11560
rect 42160 11500 42236 11560
rect 44744 11500 44820 11560
rect 47192 11500 47268 11560
rect 29648 11364 29860 11500
rect 29278 11358 29860 11364
rect 29240 11294 29246 11358
rect 29310 11294 29860 11358
rect 29278 11288 29860 11294
rect 32096 11288 32308 11500
rect 34544 11288 34892 11500
rect 37128 11288 37340 11500
rect 39576 11288 39788 11500
rect 42024 11288 42372 11500
rect 44608 11288 44820 11500
rect 47056 11288 47268 11500
rect 49640 11500 49716 11560
rect 52224 11500 52300 11560
rect 54672 11500 54748 11560
rect 57256 11500 57332 11560
rect 59704 11500 59780 11560
rect 62152 11500 62228 11560
rect 49640 11288 49852 11500
rect 52088 11288 52300 11500
rect 54400 11494 54748 11500
rect 54400 11430 54406 11494
rect 54470 11430 54748 11494
rect 54400 11424 54748 11430
rect 54536 11288 54748 11424
rect 57120 11288 57332 11500
rect 59568 11288 59780 11500
rect 62016 11288 62228 11500
rect 64600 11500 64676 11560
rect 67184 11500 67260 11560
rect 69632 11500 69708 11560
rect 72216 11500 72292 11560
rect 74664 11500 74740 11560
rect 77112 11500 77188 11560
rect 79696 11500 79772 11560
rect 82144 11500 82220 11560
rect 84728 11500 84804 11560
rect 87176 11560 87388 11696
rect 89624 11766 89836 11772
rect 89624 11702 89630 11766
rect 89694 11702 89836 11766
rect 89624 11560 89836 11702
rect 92072 11766 92518 11772
rect 94656 11766 94966 11772
rect 97104 11766 97414 11772
rect 99552 11766 99900 11772
rect 102038 11766 102348 11772
rect 104486 11766 104796 11772
rect 92072 11702 92486 11766
rect 92550 11702 92556 11766
rect 94656 11702 94934 11766
rect 94998 11702 95004 11766
rect 97104 11702 97382 11766
rect 97446 11702 97452 11766
rect 99552 11702 99694 11766
rect 99758 11702 99900 11766
rect 102000 11702 102006 11766
rect 102070 11702 102348 11766
rect 104448 11702 104454 11766
rect 104518 11702 104796 11766
rect 92072 11696 92518 11702
rect 94656 11696 94966 11702
rect 97104 11696 97414 11702
rect 92072 11560 92420 11696
rect 94656 11560 94868 11696
rect 97104 11560 97316 11696
rect 99552 11560 99900 11702
rect 102038 11696 102348 11702
rect 104486 11696 104796 11702
rect 102136 11560 102348 11696
rect 104584 11560 104796 11696
rect 107032 11766 107478 11772
rect 107032 11702 107446 11766
rect 107510 11702 107516 11766
rect 107032 11696 107478 11702
rect 107032 11560 107380 11696
rect 87176 11500 87252 11560
rect 89624 11500 89700 11560
rect 64600 11288 64812 11500
rect 67048 11288 67260 11500
rect 69496 11288 69844 11500
rect 72080 11288 72292 11500
rect 74528 11288 74740 11500
rect 76976 11288 77324 11500
rect 79560 11288 79772 11500
rect 82008 11288 82220 11500
rect 84456 11288 84804 11500
rect 87040 11288 87252 11500
rect 89488 11288 89700 11500
rect 92072 11500 92148 11560
rect 94656 11500 94732 11560
rect 97104 11500 97180 11560
rect 99688 11500 99764 11560
rect 102136 11500 102212 11560
rect 104584 11500 104660 11560
rect 92072 11288 92284 11500
rect 94520 11288 94732 11500
rect 96968 11288 97180 11500
rect 99552 11288 99764 11500
rect 102000 11288 102212 11500
rect 104448 11288 104660 11500
rect 107032 11500 107108 11560
rect 107032 11364 107244 11500
rect 124168 11494 124380 11500
rect 124168 11430 124174 11494
rect 124238 11430 124380 11494
rect 107032 11358 109420 11364
rect 107032 11294 109350 11358
rect 109414 11294 109420 11358
rect 107032 11288 109420 11294
rect 124168 11358 124380 11430
rect 124168 11294 124174 11358
rect 124238 11294 124380 11358
rect 124168 11288 124380 11294
rect 29550 11086 32308 11092
rect 29512 11022 29518 11086
rect 29582 11022 29654 11086
rect 29718 11022 32102 11086
rect 32166 11022 32308 11086
rect 29550 11016 32308 11022
rect 34680 11086 37340 11092
rect 34680 11022 34686 11086
rect 34750 11022 37270 11086
rect 37334 11022 37340 11086
rect 34680 11016 37340 11022
rect 39576 11086 39788 11092
rect 39576 11022 39718 11086
rect 39782 11022 39788 11086
rect 39576 11016 39788 11022
rect 42160 11086 42372 11092
rect 42160 11022 42302 11086
rect 42366 11022 42372 11086
rect 42160 11016 42372 11022
rect 44608 11086 44820 11092
rect 44608 11022 44750 11086
rect 44814 11022 44820 11086
rect 44608 11016 44820 11022
rect 47056 11086 47268 11092
rect 47056 11022 47062 11086
rect 47126 11022 47268 11086
rect 47056 11016 47268 11022
rect 49640 11086 57332 11092
rect 49640 11022 49782 11086
rect 49846 11022 52230 11086
rect 52294 11022 54814 11086
rect 54878 11022 57262 11086
rect 57326 11022 57332 11086
rect 49640 11016 57332 11022
rect 59568 11086 59780 11092
rect 59568 11022 59710 11086
rect 59774 11022 59780 11086
rect 59568 11016 59780 11022
rect 62016 11086 62364 11092
rect 62016 11022 62158 11086
rect 62222 11022 62364 11086
rect 62016 11016 62364 11022
rect 64600 11086 64812 11092
rect 64600 11022 64742 11086
rect 64806 11022 64812 11086
rect 64600 11016 64812 11022
rect 67048 11086 69844 11092
rect 67048 11022 67190 11086
rect 67254 11022 69774 11086
rect 69838 11022 69844 11086
rect 67048 11016 69844 11022
rect 72080 11086 74740 11092
rect 72080 11022 72222 11086
rect 72286 11022 74534 11086
rect 74598 11022 74740 11086
rect 72080 11016 74740 11022
rect 77112 11086 79772 11092
rect 77112 11022 77254 11086
rect 77318 11022 79702 11086
rect 79766 11022 79772 11086
rect 77112 11016 79772 11022
rect 82008 11086 82220 11092
rect 82008 11022 82150 11086
rect 82214 11022 82220 11086
rect 82008 11016 82220 11022
rect 84592 11086 84804 11092
rect 84592 11022 84598 11086
rect 84662 11022 84804 11086
rect 84592 11016 84804 11022
rect 87040 11086 87252 11092
rect 87040 11022 87182 11086
rect 87246 11022 87252 11086
rect 87040 11016 87252 11022
rect 89488 11086 89700 11092
rect 89488 11022 89494 11086
rect 89558 11022 89700 11086
rect 89488 11016 89700 11022
rect 92072 11086 97316 11092
rect 92072 11022 92214 11086
rect 92278 11022 94662 11086
rect 94726 11022 97110 11086
rect 97174 11022 97316 11086
rect 92072 11016 97316 11022
rect 99552 11086 102212 11092
rect 99552 11022 99558 11086
rect 99622 11022 102142 11086
rect 102206 11022 102212 11086
rect 99552 11016 102212 11022
rect 104448 11086 104796 11092
rect 104448 11022 104590 11086
rect 104654 11022 104796 11086
rect 104448 11016 104796 11022
rect 107032 11086 109284 11092
rect 107032 11022 107174 11086
rect 107238 11022 109214 11086
rect 109278 11022 109284 11086
rect 107032 11016 109284 11022
rect 29690 10985 29788 11016
rect 32186 10985 32284 11016
rect 34682 10985 34780 11016
rect 37178 10985 37276 11016
rect 39674 10985 39772 11016
rect 42170 10985 42268 11016
rect 44666 10985 44764 11016
rect 47162 10985 47260 11016
rect 49658 10985 49756 11016
rect 52154 10985 52252 11016
rect 54650 10985 54748 11016
rect 57146 10985 57244 11016
rect 59642 10985 59740 11016
rect 62138 10985 62236 11016
rect 64634 10985 64732 11016
rect 67130 10985 67228 11016
rect 69626 10985 69724 11016
rect 72122 10985 72220 11016
rect 74618 10985 74716 11016
rect 77114 10985 77212 11016
rect 79610 10985 79708 11016
rect 82106 10985 82204 11016
rect 84602 10985 84700 11016
rect 87098 10985 87196 11016
rect 89594 10985 89692 11016
rect 92090 10985 92188 11016
rect 94586 10985 94684 11016
rect 97082 10985 97180 11016
rect 99578 10985 99676 11016
rect 102074 10985 102172 11016
rect 104570 10985 104668 11016
rect 107066 10985 107164 11016
rect 124576 10826 124788 10956
rect 124576 10814 124614 10826
rect 122846 10757 122912 10760
rect 123664 10757 123730 10760
rect 122846 10755 123730 10757
rect 122846 10699 122851 10755
rect 122907 10699 123669 10755
rect 123725 10699 123730 10755
rect 124576 10750 124582 10814
rect 124670 10770 124788 10826
rect 124646 10750 124788 10770
rect 124576 10744 124788 10750
rect 122846 10697 123730 10699
rect 122846 10694 122912 10697
rect 123664 10694 123730 10697
rect 28016 10678 29588 10684
rect 28016 10614 29518 10678
rect 29582 10614 29588 10678
rect 28016 10608 29588 10614
rect 109208 10678 109420 10684
rect 109208 10614 109214 10678
rect 109278 10614 109420 10678
rect 1768 10488 1980 10548
rect 1768 10432 1798 10488
rect 1854 10432 1980 10488
rect 1768 10412 1980 10432
rect 2448 10412 2796 10548
rect 1224 10406 1980 10412
rect 1224 10342 1230 10406
rect 1294 10342 1980 10406
rect 1224 10336 1980 10342
rect 2040 10336 2796 10412
rect 15096 10542 15308 10548
rect 15096 10478 15238 10542
rect 15302 10478 15308 10542
rect 15096 10406 15308 10478
rect 28016 10472 28228 10608
rect 109208 10472 109420 10614
rect 136816 10542 137572 10548
rect 136816 10488 137502 10542
rect 15096 10342 15238 10406
rect 15302 10342 15308 10406
rect 15096 10336 15308 10342
rect 136816 10432 136944 10488
rect 137000 10478 137502 10488
rect 137566 10478 137572 10542
rect 137000 10472 137572 10478
rect 137000 10432 137028 10472
rect 136816 10336 137028 10432
rect 2040 10276 2116 10336
rect 544 10270 2116 10276
rect 544 10206 550 10270
rect 614 10206 2116 10270
rect 544 10200 2116 10206
rect 2720 9912 2932 10004
rect 2720 9868 2758 9912
rect 0 9856 2758 9868
rect 2814 9856 2932 9912
rect 0 9792 2932 9856
rect 124168 9998 124380 10004
rect 124168 9934 124310 9998
rect 124374 9934 124380 9998
rect 124168 9792 124380 9934
rect 28016 9590 29316 9596
rect 28016 9526 29246 9590
rect 29310 9526 29316 9590
rect 28016 9520 29316 9526
rect 109208 9590 109420 9596
rect 109208 9526 109350 9590
rect 109414 9526 109420 9590
rect 28016 9384 28228 9520
rect 109208 9384 109420 9526
rect 122766 9199 122832 9202
rect 123664 9199 123730 9202
rect 122766 9197 123730 9199
rect 2448 8976 2796 9188
rect 15096 9182 15308 9188
rect 15096 9118 15102 9182
rect 15166 9118 15308 9182
rect 122766 9141 122771 9197
rect 122827 9141 123669 9197
rect 123725 9141 123730 9197
rect 122766 9139 123730 9141
rect 122766 9136 122832 9139
rect 123664 9136 123730 9139
rect 15096 9052 15308 9118
rect 124576 9126 124788 9188
rect 124576 9070 124614 9126
rect 124670 9070 124788 9126
rect 15096 9046 16940 9052
rect 15096 8982 16870 9046
rect 16934 8982 16940 9046
rect 15096 8976 16940 8982
rect 124576 9046 124788 9070
rect 124576 8982 124718 9046
rect 124782 8982 124788 9046
rect 124576 8976 124788 8982
rect 2448 8916 2524 8976
rect 1224 8910 2524 8916
rect 1224 8846 1230 8910
rect 1294 8846 2524 8910
rect 1224 8840 2524 8846
rect 1768 8808 1980 8840
rect 1768 8752 1798 8808
rect 1854 8752 1980 8808
rect 1768 8704 1980 8752
rect 136816 8808 137028 8916
rect 136816 8752 136944 8808
rect 137000 8780 137028 8808
rect 137000 8774 137572 8780
rect 137000 8752 137502 8774
rect 136816 8710 137502 8752
rect 137566 8710 137572 8774
rect 136816 8704 137572 8710
rect 124168 8638 124380 8644
rect 124168 8574 124174 8638
rect 124238 8574 124380 8638
rect 124168 8432 124380 8574
rect 0 8317 6060 8372
rect 0 8296 5979 8317
rect 5848 8261 5979 8296
rect 6035 8261 6060 8317
rect 2720 8212 2932 8236
rect 2720 8156 2758 8212
rect 2814 8156 2932 8212
rect 5848 8160 6060 8261
rect 2720 8100 2932 8156
rect 0 8024 2932 8100
rect 544 7686 2796 7692
rect 544 7622 550 7686
rect 614 7622 2796 7686
rect 544 7616 2796 7622
rect 2448 7480 2796 7616
rect 15096 7686 15308 7692
rect 15096 7622 15238 7686
rect 15302 7622 15308 7686
rect 15096 7480 15308 7622
rect 1768 7128 1980 7284
rect 1768 7072 1798 7128
rect 1854 7072 1980 7128
rect 1768 7012 1980 7072
rect 1224 7006 1980 7012
rect 1224 6942 1230 7006
rect 1294 6942 1980 7006
rect 1224 6936 1980 6942
rect 136816 7148 137028 7284
rect 136816 7142 137572 7148
rect 136816 7128 137502 7142
rect 136816 7072 136944 7128
rect 137000 7078 137502 7128
rect 137566 7078 137572 7142
rect 137000 7072 137572 7078
rect 136816 6936 137028 7072
rect 1224 5510 1980 5516
rect 1224 5446 1230 5510
rect 1294 5448 1980 5510
rect 1294 5446 1798 5448
rect 1224 5440 1798 5446
rect 1768 5392 1798 5440
rect 1854 5392 1980 5448
rect 1768 5304 1980 5392
rect 136816 5510 137572 5516
rect 136816 5448 137502 5510
rect 136816 5392 136944 5448
rect 137000 5446 137502 5448
rect 137566 5446 137572 5510
rect 137000 5440 137572 5446
rect 137000 5392 137028 5440
rect 136816 5304 137028 5392
rect 1224 3878 1980 3884
rect 1224 3814 1230 3878
rect 1294 3814 1980 3878
rect 1224 3808 1980 3814
rect 1768 3768 1980 3808
rect 1768 3712 1798 3768
rect 1854 3712 1980 3768
rect 1768 3672 1980 3712
rect 16864 3878 18300 3884
rect 16864 3814 16870 3878
rect 16934 3814 18300 3878
rect 16864 3808 18300 3814
rect 16864 3672 17076 3808
rect 18088 3748 18300 3808
rect 19176 3748 19388 3884
rect 20400 3808 21836 3884
rect 20400 3748 20612 3808
rect 18088 3672 20612 3748
rect 21488 3748 21836 3808
rect 22712 3748 22924 3884
rect 23936 3808 26460 3884
rect 23936 3748 24148 3808
rect 21488 3672 24148 3748
rect 25024 3672 25236 3808
rect 26248 3748 26460 3808
rect 27336 3748 27684 3884
rect 28560 3808 29996 3884
rect 28560 3748 28772 3808
rect 26248 3672 28772 3748
rect 29784 3748 29996 3808
rect 30872 3748 31084 3884
rect 32096 3808 34620 3884
rect 32096 3748 32308 3808
rect 29784 3672 32308 3748
rect 33184 3672 33396 3808
rect 34408 3748 34620 3808
rect 35496 3808 38156 3884
rect 35496 3748 35844 3808
rect 34408 3672 35844 3748
rect 36720 3742 36932 3808
rect 36720 3678 36726 3742
rect 36790 3678 36932 3742
rect 36720 3672 36932 3678
rect 37944 3748 38156 3808
rect 39032 3748 39244 3884
rect 40256 3808 41692 3884
rect 40256 3748 40468 3808
rect 37944 3672 40468 3748
rect 41344 3748 41692 3808
rect 42568 3748 42780 3884
rect 43792 3808 46316 3884
rect 43792 3748 44004 3808
rect 41344 3672 44004 3748
rect 44880 3672 45092 3808
rect 46104 3748 46316 3808
rect 47192 3748 47540 3884
rect 48416 3808 49852 3884
rect 48416 3748 48628 3808
rect 46104 3672 48628 3748
rect 49640 3748 49852 3808
rect 50728 3748 50940 3884
rect 51952 3808 54476 3884
rect 51952 3748 52164 3808
rect 49640 3672 52164 3748
rect 53040 3672 53252 3808
rect 54264 3748 54476 3808
rect 55352 3748 55700 3884
rect 56576 3808 58012 3884
rect 56576 3748 56788 3808
rect 54264 3672 56788 3748
rect 57800 3748 58012 3808
rect 58888 3748 59100 3884
rect 60112 3748 60324 3884
rect 57800 3672 60324 3748
rect 136816 3878 137572 3884
rect 136816 3814 137502 3878
rect 137566 3814 137572 3878
rect 136816 3808 137572 3814
rect 136816 3768 137028 3808
rect 136816 3712 136944 3768
rect 137000 3712 137028 3768
rect 136816 3672 137028 3712
rect 16456 2988 16668 3068
rect 16456 2932 16548 2988
rect 16604 2932 16668 2988
rect 16456 2926 16668 2932
rect 16456 2862 16598 2926
rect 16662 2862 16668 2926
rect 16456 2856 16668 2862
rect 17680 2988 17892 3068
rect 17680 2932 17716 2988
rect 17772 2932 17892 2988
rect 17680 2926 17892 2932
rect 17680 2862 17686 2926
rect 17750 2862 17892 2926
rect 17680 2856 17892 2862
rect 18768 2988 18980 3068
rect 20128 3009 20204 3068
rect 21216 3009 21428 3068
rect 22440 3009 22516 3068
rect 18768 2932 18884 2988
rect 18940 2932 18980 2988
rect 20031 2988 20204 3009
rect 20031 2932 20052 2988
rect 20108 2932 20204 2988
rect 21199 2988 21428 3009
rect 21199 2932 21220 2988
rect 21276 2932 21428 2988
rect 22367 2988 22516 3009
rect 22367 2932 22388 2988
rect 22444 2932 22516 2988
rect 18768 2926 18980 2932
rect 18768 2862 18774 2926
rect 18838 2862 18980 2926
rect 18768 2856 18980 2862
rect 19992 2926 20204 2932
rect 19992 2862 20134 2926
rect 20198 2862 20204 2926
rect 19992 2856 20204 2862
rect 21080 2926 21428 2932
rect 21080 2862 21086 2926
rect 21150 2862 21428 2926
rect 21080 2856 21428 2862
rect 22304 2926 22516 2932
rect 22304 2862 22310 2926
rect 22374 2862 22516 2926
rect 22304 2856 22516 2862
rect 23528 2988 23740 3068
rect 24752 3009 24828 3068
rect 23528 2932 23556 2988
rect 23612 2932 23740 2988
rect 24703 2988 24828 3009
rect 24703 2932 24724 2988
rect 24780 2932 24828 2988
rect 23528 2926 23740 2932
rect 23528 2862 23670 2926
rect 23734 2862 23740 2926
rect 23528 2856 23740 2862
rect 24616 2926 24828 2932
rect 24616 2862 24758 2926
rect 24822 2862 24828 2926
rect 24616 2856 24828 2862
rect 25840 2988 26052 3068
rect 27064 3009 27140 3068
rect 28288 3009 28364 3068
rect 29376 3009 29588 3068
rect 30600 3009 30676 3068
rect 25840 2932 25892 2988
rect 25948 2932 26052 2988
rect 27039 2988 27140 3009
rect 27039 2932 27060 2988
rect 27116 2932 27140 2988
rect 28207 2988 28364 3009
rect 28207 2932 28228 2988
rect 28284 2932 28364 2988
rect 29375 2988 29588 3009
rect 29375 2932 29396 2988
rect 29452 2932 29588 2988
rect 30543 2988 30676 3009
rect 30543 2932 30564 2988
rect 30620 2932 30676 2988
rect 25840 2926 26052 2932
rect 25840 2862 25982 2926
rect 26046 2862 26052 2926
rect 25840 2856 26052 2862
rect 26928 2926 27140 2932
rect 26928 2862 27070 2926
rect 27134 2862 27140 2926
rect 26928 2856 27140 2862
rect 28152 2926 28364 2932
rect 28152 2862 28158 2926
rect 28222 2862 28364 2926
rect 28152 2856 28364 2862
rect 29240 2926 29588 2932
rect 29240 2862 29246 2926
rect 29310 2862 29588 2926
rect 29240 2856 29588 2862
rect 30464 2926 30676 2932
rect 30464 2862 30606 2926
rect 30670 2862 30676 2926
rect 30464 2856 30676 2862
rect 31688 2988 31900 3068
rect 32912 3009 32988 3068
rect 34136 3009 34212 3068
rect 35224 3009 35436 3068
rect 36448 3009 36524 3068
rect 31688 2932 31732 2988
rect 31788 2932 31900 2988
rect 32879 2988 32988 3009
rect 32879 2932 32900 2988
rect 32956 2932 32988 2988
rect 34047 2988 34212 3009
rect 34047 2932 34068 2988
rect 34124 2932 34212 2988
rect 35215 2988 35436 3009
rect 35215 2932 35236 2988
rect 35292 2932 35436 2988
rect 36383 2988 36524 3009
rect 36383 2932 36404 2988
rect 36460 2932 36524 2988
rect 31688 2926 31900 2932
rect 31688 2862 31830 2926
rect 31894 2862 31900 2926
rect 31688 2856 31900 2862
rect 32776 2926 32988 2932
rect 32776 2862 32918 2926
rect 32982 2862 32988 2926
rect 32776 2856 32988 2862
rect 34000 2926 34212 2932
rect 34000 2862 34006 2926
rect 34070 2862 34212 2926
rect 34000 2856 34212 2862
rect 35088 2926 35436 2932
rect 35088 2862 35094 2926
rect 35158 2862 35436 2926
rect 35088 2856 35436 2862
rect 36312 2926 36524 2932
rect 36312 2862 36454 2926
rect 36518 2862 36524 2926
rect 36312 2856 36524 2862
rect 37536 2988 37748 3068
rect 38760 3009 38836 3068
rect 39984 3009 40060 3068
rect 41072 3009 41284 3068
rect 42296 3009 42372 3068
rect 37536 2932 37572 2988
rect 37628 2932 37748 2988
rect 38719 2988 38836 3009
rect 38719 2932 38740 2988
rect 38796 2932 38836 2988
rect 39887 2988 40060 3009
rect 39887 2932 39908 2988
rect 39964 2932 40060 2988
rect 41055 2988 41284 3009
rect 41055 2932 41076 2988
rect 41132 2932 41284 2988
rect 42223 2988 42372 3009
rect 42223 2932 42244 2988
rect 42300 2932 42372 2988
rect 37536 2926 37748 2932
rect 37536 2862 37542 2926
rect 37606 2862 37748 2926
rect 37536 2856 37748 2862
rect 38624 2926 38836 2932
rect 38624 2862 38630 2926
rect 38694 2862 38836 2926
rect 38624 2856 38836 2862
rect 39848 2926 40060 2932
rect 39848 2862 39990 2926
rect 40054 2862 40060 2926
rect 39848 2856 40060 2862
rect 40936 2926 41284 2932
rect 40936 2862 41214 2926
rect 41278 2862 41284 2926
rect 40936 2856 41284 2862
rect 42160 2926 42372 2932
rect 42160 2862 42302 2926
rect 42366 2862 42372 2926
rect 42160 2856 42372 2862
rect 43384 2988 43596 3068
rect 44608 3009 44684 3068
rect 43384 2932 43412 2988
rect 43468 2932 43596 2988
rect 44559 2988 44684 3009
rect 44559 2932 44580 2988
rect 44636 2932 44684 2988
rect 43384 2926 43596 2932
rect 43384 2862 43390 2926
rect 43454 2862 43596 2926
rect 43384 2856 43596 2862
rect 44472 2926 44684 2932
rect 44472 2862 44478 2926
rect 44542 2862 44684 2926
rect 44472 2856 44684 2862
rect 45696 2988 45908 3068
rect 46920 3009 46996 3068
rect 48144 3009 48220 3068
rect 49232 3009 49444 3068
rect 50456 3009 50532 3068
rect 45696 2932 45748 2988
rect 45804 2932 45908 2988
rect 46895 2988 46996 3009
rect 46895 2932 46916 2988
rect 46972 2932 46996 2988
rect 48063 2988 48220 3009
rect 48063 2932 48084 2988
rect 48140 2932 48220 2988
rect 49231 2988 49444 3009
rect 49231 2932 49252 2988
rect 49308 2932 49444 2988
rect 50399 2988 50532 3009
rect 50399 2932 50420 2988
rect 50476 2932 50532 2988
rect 45696 2926 45908 2932
rect 45696 2862 45838 2926
rect 45902 2862 45908 2926
rect 45696 2856 45908 2862
rect 46784 2926 46996 2932
rect 46784 2862 46926 2926
rect 46990 2862 46996 2926
rect 46784 2856 46996 2862
rect 48008 2926 48220 2932
rect 48008 2862 48150 2926
rect 48214 2862 48220 2926
rect 48008 2856 48220 2862
rect 49096 2926 49444 2932
rect 49096 2862 49238 2926
rect 49302 2862 49444 2926
rect 49096 2856 49444 2862
rect 50320 2926 50532 2932
rect 50320 2862 50326 2926
rect 50390 2862 50532 2926
rect 50320 2856 50532 2862
rect 51544 2988 51756 3068
rect 52768 3009 52844 3068
rect 53992 3009 54068 3068
rect 55080 3009 55292 3068
rect 56304 3009 56380 3068
rect 51544 2932 51588 2988
rect 51644 2932 51756 2988
rect 52735 2988 52844 3009
rect 52735 2932 52756 2988
rect 52812 2932 52844 2988
rect 53903 2988 54068 3009
rect 53903 2932 53924 2988
rect 53980 2932 54068 2988
rect 55071 2988 55292 3009
rect 55071 2932 55092 2988
rect 55148 2932 55292 2988
rect 56239 2988 56380 3009
rect 56239 2932 56260 2988
rect 56316 2932 56380 2988
rect 51544 2926 51756 2932
rect 51544 2862 51686 2926
rect 51750 2862 51756 2926
rect 51544 2856 51756 2862
rect 52632 2926 52844 2932
rect 52632 2862 52774 2926
rect 52838 2862 52844 2926
rect 52632 2856 52844 2862
rect 53856 2926 54068 2932
rect 53856 2862 53862 2926
rect 53926 2862 54068 2926
rect 53856 2856 54068 2862
rect 54944 2926 55292 2932
rect 54944 2862 54950 2926
rect 55014 2862 55292 2926
rect 54944 2856 55292 2862
rect 56168 2926 56380 2932
rect 56168 2862 56310 2926
rect 56374 2862 56380 2926
rect 56168 2856 56380 2862
rect 57392 2988 57604 3068
rect 58616 3009 58692 3068
rect 59840 3009 59916 3068
rect 57392 2932 57428 2988
rect 57484 2932 57604 2988
rect 58575 2988 58692 3009
rect 58575 2932 58596 2988
rect 58652 2932 58692 2988
rect 59743 2988 59916 3009
rect 59743 2932 59764 2988
rect 59820 2932 59916 2988
rect 57392 2926 57604 2932
rect 57392 2862 57534 2926
rect 57598 2862 57604 2926
rect 57392 2856 57604 2862
rect 58480 2926 58692 2932
rect 58480 2862 58622 2926
rect 58686 2862 58692 2926
rect 58480 2856 58692 2862
rect 59704 2926 59916 2932
rect 59704 2862 59710 2926
rect 59774 2862 59916 2926
rect 59704 2856 59916 2862
rect 15289 2734 15355 2737
rect 15289 2732 17574 2734
rect 15289 2676 15294 2732
rect 15350 2676 17574 2732
rect 15289 2674 17574 2676
rect 15289 2671 15355 2674
rect 16864 2448 18300 2524
rect 16864 2312 17076 2448
rect 18088 2388 18300 2448
rect 19176 2388 19388 2524
rect 20400 2448 22924 2524
rect 20400 2388 20612 2448
rect 18088 2382 20612 2388
rect 18088 2318 19318 2382
rect 19382 2318 20612 2382
rect 18088 2312 20612 2318
rect 21488 2312 21836 2448
rect 22712 2388 22924 2448
rect 23936 2448 26460 2524
rect 23936 2388 24148 2448
rect 22712 2312 24148 2388
rect 25024 2312 25236 2448
rect 26248 2388 26460 2448
rect 27336 2388 27684 2524
rect 28560 2448 29996 2524
rect 28560 2388 28772 2448
rect 26248 2312 28772 2388
rect 29784 2388 29996 2448
rect 30872 2388 31084 2524
rect 32096 2448 34620 2524
rect 32096 2388 32308 2448
rect 29784 2312 32308 2388
rect 33184 2312 33396 2448
rect 34408 2388 34620 2448
rect 35496 2388 35844 2524
rect 36720 2448 38156 2524
rect 36720 2388 36932 2448
rect 34408 2312 36932 2388
rect 37944 2388 38156 2448
rect 39032 2388 39244 2524
rect 40256 2448 42780 2524
rect 40256 2388 40468 2448
rect 37944 2312 40468 2388
rect 41344 2312 41692 2448
rect 42568 2388 42780 2448
rect 43792 2448 46316 2524
rect 43792 2388 44004 2448
rect 42568 2312 44004 2388
rect 44880 2312 45092 2448
rect 46104 2388 46316 2448
rect 47192 2388 47540 2524
rect 48416 2448 49852 2524
rect 48416 2388 48628 2448
rect 46104 2312 48628 2388
rect 49640 2388 49852 2448
rect 50728 2388 50940 2524
rect 51952 2448 54476 2524
rect 51952 2388 52164 2448
rect 49640 2312 52164 2388
rect 53040 2312 53252 2448
rect 54264 2388 54476 2448
rect 55352 2448 58012 2524
rect 55352 2388 55700 2448
rect 54264 2312 55700 2388
rect 56576 2312 56788 2448
rect 57800 2388 58012 2448
rect 58888 2388 59100 2524
rect 60112 2388 60324 2524
rect 57800 2312 60324 2388
rect 1768 2088 1980 2116
rect 1768 2032 1798 2088
rect 1854 2032 1980 2088
rect 1768 1980 1980 2032
rect 136816 2088 137028 2116
rect 136816 2032 136944 2088
rect 137000 2032 137028 2088
rect 1768 1904 2116 1980
rect 2040 1844 2116 1904
rect 136816 1904 137028 2032
rect 136816 1844 136892 1904
rect 2040 1752 2252 1844
rect 2040 1702 2134 1752
rect 2040 1638 2046 1702
rect 2110 1696 2134 1702
rect 2190 1696 2252 1752
rect 2110 1638 2252 1696
rect 2040 1632 2252 1638
rect 3672 1752 4020 1844
rect 3672 1638 3814 1752
rect 3870 1702 4020 1752
rect 3878 1638 4020 1702
rect 3672 1632 4020 1638
rect 5440 1752 5652 1844
rect 5440 1702 5494 1752
rect 5440 1638 5446 1702
rect 5550 1696 5652 1752
rect 5510 1638 5652 1696
rect 5440 1632 5652 1638
rect 7072 1752 7284 1844
rect 7072 1696 7174 1752
rect 7230 1702 7284 1752
rect 7072 1638 7214 1696
rect 7278 1638 7284 1702
rect 7072 1632 7284 1638
rect 8704 1752 9052 1844
rect 8704 1702 8854 1752
rect 8704 1638 8710 1702
rect 8774 1696 8854 1702
rect 8910 1696 9052 1752
rect 8774 1638 9052 1696
rect 8704 1632 9052 1638
rect 10472 1752 10684 1844
rect 10472 1702 10534 1752
rect 10472 1638 10478 1702
rect 10590 1696 10684 1752
rect 10542 1638 10684 1696
rect 10472 1632 10684 1638
rect 12104 1752 12316 1844
rect 12104 1702 12214 1752
rect 12104 1638 12110 1702
rect 12174 1696 12214 1702
rect 12270 1696 12316 1752
rect 12174 1638 12316 1696
rect 12104 1632 12316 1638
rect 13872 1752 14084 1844
rect 13872 1702 13894 1752
rect 13872 1638 13878 1702
rect 13950 1696 14084 1752
rect 13942 1638 14084 1696
rect 13872 1632 14084 1638
rect 15504 1752 15716 1844
rect 15504 1696 15574 1752
rect 15630 1702 15716 1752
rect 15630 1696 15646 1702
rect 15504 1638 15646 1696
rect 15710 1638 15716 1702
rect 15504 1632 15716 1638
rect 17136 1752 17348 1844
rect 17136 1702 17254 1752
rect 17136 1638 17142 1702
rect 17206 1696 17254 1702
rect 17310 1696 17348 1752
rect 17206 1638 17348 1696
rect 17136 1632 17348 1638
rect 18904 1752 19116 1844
rect 18904 1696 18934 1752
rect 18990 1702 19116 1752
rect 18990 1696 19046 1702
rect 18904 1638 19046 1696
rect 19110 1638 19116 1702
rect 18904 1632 19116 1638
rect 20536 1752 20748 1844
rect 20536 1702 20614 1752
rect 20536 1638 20542 1702
rect 20606 1696 20614 1702
rect 20670 1696 20748 1752
rect 20606 1638 20748 1696
rect 20536 1632 20748 1638
rect 22168 1752 22380 1844
rect 22168 1702 22294 1752
rect 22168 1638 22174 1702
rect 22238 1696 22294 1702
rect 22350 1696 22380 1752
rect 22238 1638 22380 1696
rect 22168 1632 22380 1638
rect 23936 1752 24148 1844
rect 23936 1702 23974 1752
rect 23936 1638 23942 1702
rect 24030 1696 24148 1752
rect 24006 1638 24148 1696
rect 23936 1632 24148 1638
rect 25568 1752 25780 1844
rect 25568 1696 25654 1752
rect 25710 1702 25780 1752
rect 25568 1638 25710 1696
rect 25774 1638 25780 1702
rect 25568 1632 25780 1638
rect 27200 1752 27412 1844
rect 27200 1702 27334 1752
rect 27200 1638 27206 1702
rect 27270 1696 27334 1702
rect 27390 1696 27412 1752
rect 28968 1752 29180 1844
rect 28968 1708 29014 1752
rect 27270 1638 27412 1696
rect 27200 1632 27412 1638
rect 28832 1702 29014 1708
rect 28832 1638 28838 1702
rect 28902 1696 29014 1702
rect 29070 1696 29180 1752
rect 30600 1752 30812 1844
rect 30600 1708 30694 1752
rect 28902 1638 29180 1696
rect 28832 1632 29180 1638
rect 30464 1702 30694 1708
rect 30464 1638 30470 1702
rect 30534 1696 30694 1702
rect 30750 1696 30812 1752
rect 30534 1638 30812 1696
rect 30464 1632 30812 1638
rect 32232 1752 32580 1844
rect 32232 1702 32374 1752
rect 32232 1638 32238 1702
rect 32302 1696 32374 1702
rect 32430 1696 32580 1752
rect 32302 1638 32580 1696
rect 32232 1632 32580 1638
rect 34000 1752 34212 1844
rect 34000 1696 34054 1752
rect 34110 1708 34212 1752
rect 35632 1752 35844 1844
rect 36758 1838 37612 1844
rect 36720 1774 36726 1838
rect 36790 1774 37612 1838
rect 36758 1768 37612 1774
rect 34110 1702 34348 1708
rect 34110 1696 34278 1702
rect 34000 1638 34278 1696
rect 34342 1638 34348 1702
rect 34000 1632 34348 1638
rect 35632 1702 35734 1752
rect 35632 1638 35638 1702
rect 35702 1696 35734 1702
rect 35790 1696 35844 1752
rect 35702 1638 35844 1696
rect 35632 1632 35844 1638
rect 37264 1752 37612 1768
rect 37264 1702 37414 1752
rect 37264 1638 37270 1702
rect 37334 1696 37414 1702
rect 37470 1696 37612 1752
rect 37334 1638 37612 1696
rect 37264 1632 37612 1638
rect 39032 1752 39244 1844
rect 39032 1702 39094 1752
rect 39032 1638 39038 1702
rect 39150 1696 39244 1752
rect 39102 1638 39244 1696
rect 39032 1632 39244 1638
rect 40664 1752 40876 1844
rect 40664 1702 40774 1752
rect 40664 1638 40670 1702
rect 40734 1696 40774 1702
rect 40830 1696 40876 1752
rect 40734 1638 40876 1696
rect 40664 1632 40876 1638
rect 42432 1752 42644 1844
rect 42432 1702 42454 1752
rect 42432 1638 42438 1702
rect 42510 1696 42644 1752
rect 42502 1638 42644 1696
rect 42432 1632 42644 1638
rect 44064 1752 44276 1844
rect 44064 1702 44134 1752
rect 44064 1638 44070 1702
rect 44190 1696 44276 1752
rect 44134 1638 44276 1696
rect 44064 1632 44276 1638
rect 45696 1752 45908 1844
rect 45696 1702 45814 1752
rect 45696 1638 45702 1702
rect 45766 1696 45814 1702
rect 45870 1696 45908 1752
rect 45766 1638 45908 1696
rect 45696 1632 45908 1638
rect 47464 1752 47676 1844
rect 47464 1702 47494 1752
rect 47464 1638 47470 1702
rect 47550 1696 47676 1752
rect 49096 1752 49308 1844
rect 49096 1708 49174 1752
rect 47534 1638 47676 1696
rect 47464 1632 47676 1638
rect 48960 1702 49174 1708
rect 48960 1638 48966 1702
rect 49030 1696 49174 1702
rect 49230 1696 49308 1752
rect 49030 1638 49308 1696
rect 48960 1632 49308 1638
rect 50728 1752 50940 1844
rect 50728 1702 50854 1752
rect 50728 1638 50734 1702
rect 50798 1696 50854 1702
rect 50910 1696 50940 1752
rect 50798 1638 50940 1696
rect 50728 1632 50940 1638
rect 52496 1752 52708 1844
rect 52496 1702 52534 1752
rect 52496 1638 52502 1702
rect 52590 1696 52708 1752
rect 52566 1638 52708 1696
rect 52496 1632 52708 1638
rect 54128 1752 54340 1844
rect 54128 1702 54214 1752
rect 54128 1638 54134 1702
rect 54198 1696 54214 1702
rect 54270 1696 54340 1752
rect 54198 1638 54340 1696
rect 54128 1632 54340 1638
rect 55760 1752 55972 1844
rect 55760 1696 55894 1752
rect 55950 1702 55972 1752
rect 57528 1752 57740 1844
rect 57528 1708 57574 1752
rect 55760 1638 55902 1696
rect 55966 1638 55972 1702
rect 55760 1632 55972 1638
rect 57392 1702 57574 1708
rect 57392 1638 57398 1702
rect 57462 1696 57574 1702
rect 57630 1696 57740 1752
rect 57462 1638 57740 1696
rect 57392 1632 57740 1638
rect 59160 1752 59372 1844
rect 59160 1702 59254 1752
rect 59160 1638 59166 1702
rect 59230 1696 59254 1702
rect 59310 1696 59372 1752
rect 59230 1638 59372 1696
rect 59160 1632 59372 1638
rect 60792 1752 61140 1844
rect 60792 1638 60934 1752
rect 60990 1702 61140 1752
rect 60998 1638 61140 1702
rect 60792 1632 61140 1638
rect 62560 1752 62772 1844
rect 62560 1696 62614 1752
rect 62670 1702 62772 1752
rect 62670 1696 62702 1702
rect 62560 1638 62702 1696
rect 62766 1638 62772 1702
rect 62560 1632 62772 1638
rect 64192 1752 64404 1844
rect 64192 1702 64294 1752
rect 64192 1638 64198 1702
rect 64262 1696 64294 1702
rect 64350 1696 64404 1752
rect 64262 1638 64404 1696
rect 64192 1632 64404 1638
rect 65824 1752 66172 1844
rect 65824 1702 65974 1752
rect 65824 1638 65830 1702
rect 65894 1696 65974 1702
rect 66030 1696 66172 1752
rect 65894 1638 66172 1696
rect 65824 1632 66172 1638
rect 67592 1752 67804 1844
rect 67592 1702 67654 1752
rect 67592 1638 67598 1702
rect 67710 1696 67804 1752
rect 67662 1638 67804 1696
rect 67592 1632 67804 1638
rect 69224 1752 69436 1844
rect 69224 1702 69334 1752
rect 69224 1638 69230 1702
rect 69294 1696 69334 1702
rect 69390 1696 69436 1752
rect 69294 1638 69436 1696
rect 69224 1632 69436 1638
rect 70992 1752 71204 1844
rect 70992 1696 71014 1752
rect 71070 1702 71204 1752
rect 71070 1696 71134 1702
rect 70992 1638 71134 1696
rect 71198 1638 71204 1702
rect 70992 1632 71204 1638
rect 72624 1752 72836 1844
rect 72624 1702 72694 1752
rect 72624 1638 72630 1702
rect 72750 1696 72836 1752
rect 72694 1638 72836 1696
rect 72624 1632 72836 1638
rect 74256 1752 74468 1844
rect 74256 1702 74374 1752
rect 74256 1638 74262 1702
rect 74326 1696 74374 1702
rect 74430 1696 74468 1752
rect 74326 1638 74468 1696
rect 74256 1632 74468 1638
rect 76024 1752 76236 1844
rect 76024 1702 76054 1752
rect 76024 1638 76030 1702
rect 76110 1696 76236 1752
rect 76094 1638 76236 1696
rect 76024 1632 76236 1638
rect 77656 1752 77868 1844
rect 77656 1702 77734 1752
rect 77656 1638 77662 1702
rect 77726 1696 77734 1702
rect 77790 1696 77868 1752
rect 77726 1638 77868 1696
rect 77656 1632 77868 1638
rect 79288 1752 79500 1844
rect 79288 1702 79414 1752
rect 79288 1638 79294 1702
rect 79358 1696 79414 1702
rect 79470 1696 79500 1752
rect 79358 1638 79500 1696
rect 79288 1632 79500 1638
rect 81056 1752 81268 1844
rect 81056 1696 81094 1752
rect 81150 1702 81268 1752
rect 81150 1696 81198 1702
rect 81056 1638 81198 1696
rect 81262 1638 81268 1702
rect 81056 1632 81268 1638
rect 82688 1752 82900 1844
rect 82688 1702 82774 1752
rect 82688 1638 82694 1702
rect 82758 1696 82774 1702
rect 82830 1696 82900 1752
rect 82758 1638 82900 1696
rect 82688 1632 82900 1638
rect 84320 1752 84532 1844
rect 84320 1696 84454 1752
rect 84510 1708 84532 1752
rect 86088 1752 86300 1844
rect 84510 1702 84668 1708
rect 84510 1696 84598 1702
rect 84320 1638 84598 1696
rect 84662 1638 84668 1702
rect 84320 1632 84668 1638
rect 86088 1702 86134 1752
rect 86088 1638 86094 1702
rect 86190 1696 86300 1752
rect 86158 1638 86300 1696
rect 86088 1632 86300 1638
rect 87720 1752 87932 1844
rect 87720 1702 87814 1752
rect 87720 1638 87726 1702
rect 87790 1696 87814 1702
rect 87870 1696 87932 1752
rect 87790 1638 87932 1696
rect 87720 1632 87932 1638
rect 89352 1752 89700 1844
rect 89352 1702 89494 1752
rect 89352 1638 89358 1702
rect 89422 1696 89494 1702
rect 89550 1696 89700 1752
rect 89422 1638 89700 1696
rect 89352 1632 89700 1638
rect 91120 1752 91332 1844
rect 91120 1702 91174 1752
rect 91120 1638 91126 1702
rect 91230 1696 91332 1752
rect 91190 1638 91332 1696
rect 91120 1632 91332 1638
rect 92752 1752 92964 1844
rect 92752 1696 92854 1752
rect 92910 1702 92964 1752
rect 92752 1638 92894 1696
rect 92958 1638 92964 1702
rect 92752 1632 92964 1638
rect 94384 1752 94732 1844
rect 94384 1696 94534 1752
rect 94590 1702 94732 1752
rect 94590 1696 94662 1702
rect 94384 1638 94662 1696
rect 94726 1638 94732 1702
rect 94384 1632 94732 1638
rect 96152 1752 96364 1844
rect 96152 1702 96214 1752
rect 96152 1638 96158 1702
rect 96270 1696 96364 1752
rect 96222 1638 96364 1696
rect 96152 1632 96364 1638
rect 97784 1752 97996 1844
rect 97784 1696 97894 1752
rect 97950 1702 97996 1752
rect 97784 1638 97926 1696
rect 97990 1638 97996 1702
rect 97784 1632 97996 1638
rect 99552 1752 99764 1844
rect 99552 1696 99574 1752
rect 99630 1702 99764 1752
rect 99630 1696 99694 1702
rect 99552 1638 99694 1696
rect 99758 1638 99764 1702
rect 99552 1632 99764 1638
rect 101184 1752 101396 1844
rect 101184 1702 101254 1752
rect 101184 1638 101190 1702
rect 101310 1696 101396 1752
rect 101254 1638 101396 1696
rect 101184 1632 101396 1638
rect 102816 1752 103028 1844
rect 102816 1696 102934 1752
rect 102990 1702 103028 1752
rect 102816 1638 102958 1696
rect 103022 1638 103028 1702
rect 102816 1632 103028 1638
rect 104584 1752 104796 1844
rect 104584 1702 104614 1752
rect 104584 1638 104590 1702
rect 104670 1696 104796 1752
rect 104654 1638 104796 1696
rect 104584 1632 104796 1638
rect 106216 1752 106428 1844
rect 106216 1702 106294 1752
rect 106216 1638 106222 1702
rect 106286 1696 106294 1702
rect 106350 1696 106428 1752
rect 106286 1638 106428 1696
rect 106216 1632 106428 1638
rect 107848 1752 108060 1844
rect 107848 1702 107974 1752
rect 107848 1638 107854 1702
rect 107918 1696 107974 1702
rect 108030 1696 108060 1752
rect 107918 1638 108060 1696
rect 107848 1632 108060 1638
rect 109616 1752 109828 1844
rect 109616 1702 109654 1752
rect 109616 1638 109622 1702
rect 109710 1696 109828 1752
rect 109686 1638 109828 1696
rect 109616 1632 109828 1638
rect 111248 1752 111460 1844
rect 111248 1696 111334 1752
rect 111390 1702 111460 1752
rect 111248 1638 111390 1696
rect 111454 1638 111460 1702
rect 111248 1632 111460 1638
rect 112880 1752 113092 1844
rect 112880 1702 113014 1752
rect 112880 1638 112886 1702
rect 112950 1696 113014 1702
rect 113070 1696 113092 1752
rect 112950 1638 113092 1696
rect 112880 1632 113092 1638
rect 114648 1752 114860 1844
rect 114648 1702 114694 1752
rect 114648 1638 114654 1702
rect 114750 1696 114860 1752
rect 114718 1638 114860 1696
rect 114648 1632 114860 1638
rect 116280 1752 116492 1844
rect 116280 1702 116374 1752
rect 116280 1638 116286 1702
rect 116350 1696 116374 1702
rect 116430 1696 116492 1752
rect 116350 1638 116492 1696
rect 116280 1632 116492 1638
rect 117912 1752 118260 1844
rect 117912 1638 118054 1752
rect 118110 1702 118260 1752
rect 118118 1638 118260 1702
rect 117912 1632 118260 1638
rect 119680 1752 119892 1844
rect 119680 1702 119734 1752
rect 119680 1638 119686 1702
rect 119790 1696 119892 1752
rect 119750 1638 119892 1696
rect 119680 1632 119892 1638
rect 121312 1752 121524 1844
rect 121312 1696 121414 1752
rect 121470 1702 121524 1752
rect 121312 1638 121454 1696
rect 121518 1638 121524 1702
rect 121312 1632 121524 1638
rect 122944 1752 123292 1844
rect 122944 1702 123094 1752
rect 122944 1638 122950 1702
rect 123014 1696 123094 1702
rect 123150 1696 123292 1752
rect 123014 1638 123292 1696
rect 122944 1632 123292 1638
rect 124712 1752 124924 1844
rect 124712 1696 124774 1752
rect 124830 1708 124924 1752
rect 126344 1752 126556 1844
rect 124830 1702 125196 1708
rect 124830 1696 125126 1702
rect 124712 1638 125126 1696
rect 125190 1638 125196 1702
rect 124712 1632 125196 1638
rect 126344 1702 126454 1752
rect 126344 1638 126350 1702
rect 126414 1696 126454 1702
rect 126510 1696 126556 1752
rect 126414 1638 126556 1696
rect 126344 1632 126556 1638
rect 128112 1752 128324 1844
rect 128112 1702 128134 1752
rect 128112 1638 128118 1702
rect 128190 1696 128324 1752
rect 128182 1638 128324 1696
rect 128112 1632 128324 1638
rect 129744 1752 129956 1844
rect 129744 1696 129814 1752
rect 129870 1702 129956 1752
rect 129870 1696 129886 1702
rect 129744 1638 129886 1696
rect 129950 1638 129956 1702
rect 129744 1632 129956 1638
rect 131376 1752 131588 1844
rect 131376 1702 131494 1752
rect 131376 1638 131382 1702
rect 131446 1696 131494 1702
rect 131550 1696 131588 1752
rect 131446 1638 131588 1696
rect 131376 1632 131588 1638
rect 133144 1752 133356 1844
rect 133144 1702 133174 1752
rect 133144 1638 133150 1702
rect 133230 1696 133356 1752
rect 133214 1638 133356 1696
rect 133144 1632 133356 1638
rect 134776 1752 134988 1844
rect 134776 1702 134854 1752
rect 134776 1638 134782 1702
rect 134846 1696 134854 1702
rect 134910 1696 134988 1752
rect 134846 1638 134988 1696
rect 134776 1632 134988 1638
rect 136408 1768 136892 1844
rect 136408 1752 136620 1768
rect 136408 1696 136534 1752
rect 136590 1702 136620 1752
rect 136408 1638 136550 1696
rect 136614 1638 136620 1702
rect 136408 1632 136620 1638
rect 952 1294 137844 1300
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 2046 1294
rect 2110 1230 3814 1294
rect 3878 1230 5446 1294
rect 5510 1230 7214 1294
rect 7278 1230 8710 1294
rect 8774 1230 10478 1294
rect 10542 1230 12110 1294
rect 12174 1230 13878 1294
rect 13942 1230 15646 1294
rect 15710 1230 17142 1294
rect 17206 1230 19046 1294
rect 19110 1230 20542 1294
rect 20606 1230 22174 1294
rect 22238 1230 23942 1294
rect 24006 1230 25710 1294
rect 25774 1230 27206 1294
rect 27270 1230 28838 1294
rect 28902 1230 30470 1294
rect 30534 1230 32238 1294
rect 32302 1230 34278 1294
rect 34342 1230 35638 1294
rect 35702 1230 37270 1294
rect 37334 1230 39038 1294
rect 39102 1230 40670 1294
rect 40734 1230 42438 1294
rect 42502 1230 44070 1294
rect 44134 1230 45702 1294
rect 45766 1230 47470 1294
rect 47534 1230 48966 1294
rect 49030 1230 50734 1294
rect 50798 1230 52502 1294
rect 52566 1230 54134 1294
rect 54198 1230 55902 1294
rect 55966 1230 57398 1294
rect 57462 1230 59166 1294
rect 59230 1230 60934 1294
rect 60998 1230 62702 1294
rect 62766 1230 64198 1294
rect 64262 1230 65830 1294
rect 65894 1230 67598 1294
rect 67662 1230 69230 1294
rect 69294 1230 71134 1294
rect 71198 1230 72630 1294
rect 72694 1230 74262 1294
rect 74326 1230 76030 1294
rect 76094 1230 77662 1294
rect 77726 1230 79294 1294
rect 79358 1230 81198 1294
rect 81262 1230 82694 1294
rect 82758 1230 84598 1294
rect 84662 1230 86094 1294
rect 86158 1230 87726 1294
rect 87790 1230 89358 1294
rect 89422 1230 91126 1294
rect 91190 1230 92894 1294
rect 92958 1230 94662 1294
rect 94726 1230 96158 1294
rect 96222 1230 97926 1294
rect 97990 1230 99694 1294
rect 99758 1230 101190 1294
rect 101254 1230 102958 1294
rect 103022 1230 104590 1294
rect 104654 1230 106222 1294
rect 106286 1230 107854 1294
rect 107918 1230 109622 1294
rect 109686 1230 111390 1294
rect 111454 1230 112886 1294
rect 112950 1230 114654 1294
rect 114718 1230 116286 1294
rect 116350 1230 118054 1294
rect 118118 1230 119686 1294
rect 119750 1230 121454 1294
rect 121518 1230 122950 1294
rect 123014 1230 125126 1294
rect 125190 1230 126350 1294
rect 126414 1230 128118 1294
rect 128182 1230 129886 1294
rect 129950 1230 131382 1294
rect 131446 1230 133150 1294
rect 133214 1230 134782 1294
rect 134846 1230 136550 1294
rect 136614 1230 137502 1294
rect 137566 1230 137638 1294
rect 137702 1230 137774 1294
rect 137838 1230 137844 1294
rect 952 1158 137844 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 137502 1158
rect 137566 1094 137638 1158
rect 137702 1094 137774 1158
rect 137838 1094 137844 1158
rect 952 1022 137844 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 137502 1022
rect 137566 958 137638 1022
rect 137702 958 137774 1022
rect 137838 958 137844 1022
rect 952 952 137844 958
rect 272 614 138524 620
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 19318 614
rect 19382 550 138182 614
rect 138246 550 138318 614
rect 138382 550 138454 614
rect 138518 550 138524 614
rect 272 478 138524 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 138182 478
rect 138246 414 138318 478
rect 138382 414 138454 478
rect 138518 414 138524 478
rect 272 342 138524 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 138182 342
rect 138246 278 138318 342
rect 138382 278 138454 342
rect 138518 278 138524 342
rect 272 272 138524 278
<< via3 >>
rect 278 133422 342 133486
rect 414 133422 478 133486
rect 550 133422 614 133486
rect 138182 133422 138246 133486
rect 138318 133422 138382 133486
rect 138454 133422 138518 133486
rect 278 133286 342 133350
rect 414 133286 478 133350
rect 550 133286 614 133350
rect 138182 133286 138246 133350
rect 138318 133286 138382 133350
rect 138454 133286 138518 133350
rect 278 133150 342 133214
rect 414 133150 478 133214
rect 550 133150 614 133214
rect 120638 133150 120702 133214
rect 123630 133150 123694 133214
rect 138182 133150 138246 133214
rect 138318 133150 138382 133214
rect 138454 133150 138518 133214
rect 958 132742 1022 132806
rect 1094 132742 1158 132806
rect 1230 132742 1294 132806
rect 137502 132742 137566 132806
rect 137638 132742 137702 132806
rect 137774 132742 137838 132806
rect 958 132606 1022 132670
rect 1094 132606 1158 132670
rect 1230 132606 1294 132670
rect 137502 132606 137566 132670
rect 137638 132606 137702 132670
rect 137774 132606 137838 132670
rect 958 132470 1022 132534
rect 1094 132470 1158 132534
rect 1230 132470 1294 132534
rect 2182 132470 2246 132534
rect 3678 132470 3742 132534
rect 5446 132470 5510 132534
rect 7214 132470 7278 132534
rect 8982 132470 9046 132534
rect 10478 132470 10542 132534
rect 12110 132470 12174 132534
rect 13878 132470 13942 132534
rect 15646 132470 15710 132534
rect 17142 132470 17206 132534
rect 18910 132470 18974 132534
rect 20678 132470 20742 132534
rect 22174 132470 22238 132534
rect 23942 132470 24006 132534
rect 25710 132470 25774 132534
rect 27206 132470 27270 132534
rect 28974 132470 29038 132534
rect 30742 132470 30806 132534
rect 32238 132470 32302 132534
rect 34142 132470 34206 132534
rect 35638 132470 35702 132534
rect 37406 132470 37470 132534
rect 39174 132470 39238 132534
rect 40670 132470 40734 132534
rect 42438 132470 42502 132534
rect 44206 132470 44270 132534
rect 45702 132470 45766 132534
rect 47470 132470 47534 132534
rect 49102 132470 49166 132534
rect 50734 132470 50798 132534
rect 52638 132470 52702 132534
rect 54134 132470 54198 132534
rect 55902 132470 55966 132534
rect 57670 132470 57734 132534
rect 59166 132470 59230 132534
rect 61070 132470 61134 132534
rect 62702 132470 62766 132534
rect 64198 132470 64262 132534
rect 66102 132470 66166 132534
rect 67734 132470 67798 132534
rect 69230 132470 69294 132534
rect 71134 132470 71198 132534
rect 72630 132470 72694 132534
rect 74262 132470 74326 132534
rect 76166 132470 76230 132534
rect 77662 132470 77726 132534
rect 79294 132470 79358 132534
rect 81198 132470 81262 132534
rect 82694 132470 82758 132534
rect 84326 132470 84390 132534
rect 86094 132470 86158 132534
rect 87726 132470 87790 132534
rect 89766 132470 89830 132534
rect 91126 132470 91190 132534
rect 92894 132470 92958 132534
rect 94662 132470 94726 132534
rect 96158 132470 96222 132534
rect 97926 132470 97990 132534
rect 99694 132470 99758 132534
rect 101190 132470 101254 132534
rect 102958 132470 103022 132534
rect 104726 132470 104790 132534
rect 106222 132470 106286 132534
rect 107854 132470 107918 132534
rect 109622 132470 109686 132534
rect 111390 132470 111454 132534
rect 112886 132470 112950 132534
rect 114654 132470 114718 132534
rect 116422 132470 116486 132534
rect 117918 132470 117982 132534
rect 119686 132470 119750 132534
rect 121454 132470 121518 132534
rect 123086 132470 123150 132534
rect 124718 132470 124782 132534
rect 126350 132470 126414 132534
rect 128118 132470 128182 132534
rect 129886 132470 129950 132534
rect 131382 132470 131446 132534
rect 133150 132470 133214 132534
rect 134918 132470 134982 132534
rect 136414 132470 136478 132534
rect 137502 132470 137566 132534
rect 137638 132470 137702 132534
rect 137774 132470 137838 132534
rect 2182 132062 2246 132126
rect 2046 131926 2110 131990
rect 3678 132062 3742 132126
rect 5446 132062 5510 132126
rect 7214 132062 7278 132126
rect 8982 132062 9046 132126
rect 10478 132062 10542 132126
rect 12110 132062 12174 132126
rect 13878 132062 13942 132126
rect 15646 132062 15710 132126
rect 17142 132062 17206 132126
rect 18910 132062 18974 132126
rect 20678 132062 20742 132126
rect 22174 132062 22238 132126
rect 23942 132062 24006 132126
rect 25710 132062 25774 132126
rect 27206 132062 27270 132126
rect 28974 132062 29038 132126
rect 30742 132062 30806 132126
rect 32238 132062 32302 132126
rect 34142 132062 34206 132126
rect 35638 132062 35702 132126
rect 37406 132062 37470 132126
rect 39174 132062 39238 132126
rect 40670 132062 40734 132126
rect 42438 132062 42502 132126
rect 44206 132062 44270 132126
rect 45702 132062 45766 132126
rect 47470 132062 47534 132126
rect 49102 132062 49166 132126
rect 50734 132062 50798 132126
rect 52638 132062 52702 132126
rect 54134 132062 54198 132126
rect 55902 132062 55966 132126
rect 57670 132062 57734 132126
rect 59166 132062 59230 132126
rect 61070 132062 61134 132126
rect 62702 132062 62766 132126
rect 64198 132062 64262 132126
rect 66102 132062 66166 132126
rect 67734 132062 67798 132126
rect 69230 132062 69294 132126
rect 71134 132062 71198 132126
rect 72630 132062 72694 132126
rect 74262 132062 74326 132126
rect 76166 132062 76230 132126
rect 77662 132062 77726 132126
rect 79294 132062 79358 132126
rect 81198 132062 81262 132126
rect 82694 132062 82758 132126
rect 84326 132062 84390 132126
rect 86094 132062 86158 132126
rect 87726 132062 87790 132126
rect 89766 132062 89830 132126
rect 91126 132062 91190 132126
rect 92894 132062 92958 132126
rect 94662 132062 94726 132126
rect 96158 132062 96222 132126
rect 97926 132062 97990 132126
rect 99694 132062 99758 132126
rect 101190 132062 101254 132126
rect 102958 132062 103022 132126
rect 104726 132062 104790 132126
rect 106222 132062 106286 132126
rect 107854 132062 107918 132126
rect 109622 132062 109686 132126
rect 111390 132062 111454 132126
rect 112886 132062 112950 132126
rect 114654 132062 114718 132126
rect 116422 132062 116486 132126
rect 117918 132062 117982 132126
rect 119686 132062 119750 132126
rect 119686 131926 119750 131990
rect 121454 132062 121518 132126
rect 123086 132062 123150 132126
rect 124718 132062 124782 132126
rect 126350 132062 126414 132126
rect 128118 132062 128182 132126
rect 129886 132062 129950 132126
rect 131382 132062 131446 132126
rect 133150 132062 133214 132126
rect 134918 132062 134982 132126
rect 136414 132062 136478 132126
rect 136822 131926 136886 131990
rect 2046 131518 2110 131582
rect 136822 131518 136886 131582
rect 120638 131382 120702 131446
rect 119550 131246 119614 131310
rect 119958 130838 120022 130902
rect 121182 130838 121246 130902
rect 123630 130430 123694 130494
rect 123766 130294 123830 130358
rect 138182 130430 138246 130494
rect 119686 130022 119750 130086
rect 119414 129886 119478 129950
rect 123630 129886 123694 129950
rect 1230 129750 1294 129814
rect 132742 129750 132806 129814
rect 137502 129750 137566 129814
rect 119550 129206 119614 129270
rect 117510 129070 117574 129134
rect 123630 128934 123694 128998
rect 123630 128798 123694 128862
rect 136822 128798 136886 128862
rect 1230 128118 1294 128182
rect 136822 128118 136886 128182
rect 137502 128118 137566 128182
rect 119414 127846 119478 127910
rect 29654 127574 29718 127638
rect 29926 127438 29990 127502
rect 31966 127574 32030 127638
rect 34550 127607 34614 127638
rect 34550 127574 34554 127607
rect 34554 127574 34610 127607
rect 34610 127574 34614 127607
rect 32510 127438 32574 127502
rect 36998 127607 37062 127638
rect 36998 127574 37050 127607
rect 37050 127574 37062 127607
rect 34958 127438 35022 127502
rect 37270 127438 37334 127502
rect 39582 127607 39646 127638
rect 39582 127574 39602 127607
rect 39602 127574 39646 127607
rect 42030 127607 42094 127638
rect 42030 127574 42042 127607
rect 42042 127574 42094 127607
rect 39990 127438 40054 127502
rect 42438 127438 42502 127502
rect 44614 127574 44678 127638
rect 44886 127438 44950 127502
rect 47062 127607 47126 127638
rect 47062 127574 47090 127607
rect 47090 127574 47126 127607
rect 47334 127438 47398 127502
rect 49510 127607 49574 127638
rect 49510 127574 49530 127607
rect 49530 127574 49574 127607
rect 49918 127438 49982 127502
rect 51958 127574 52022 127638
rect 52366 127438 52430 127502
rect 54406 127574 54470 127638
rect 56990 127607 57054 127638
rect 56990 127574 57018 127607
rect 57018 127574 57054 127607
rect 54950 127438 55014 127502
rect 57398 127438 57462 127502
rect 59574 127574 59638 127638
rect 59846 127438 59910 127502
rect 62022 127607 62086 127638
rect 62022 127574 62066 127607
rect 62066 127574 62086 127607
rect 64606 127574 64670 127638
rect 62430 127438 62494 127502
rect 64742 127438 64806 127502
rect 67054 127607 67118 127638
rect 67054 127574 67058 127607
rect 67058 127574 67118 127607
rect 67326 127438 67390 127502
rect 69366 127574 69430 127638
rect 69774 127438 69838 127502
rect 72086 127574 72150 127638
rect 72358 127438 72422 127502
rect 74398 127574 74462 127638
rect 76982 127607 77046 127638
rect 76982 127574 76986 127607
rect 76986 127574 77042 127607
rect 77042 127574 77046 127607
rect 74942 127438 75006 127502
rect 79430 127607 79494 127638
rect 79430 127574 79482 127607
rect 79482 127574 79494 127607
rect 77390 127438 77454 127502
rect 79838 127438 79902 127502
rect 82014 127607 82078 127638
rect 82014 127574 82034 127607
rect 82034 127574 82078 127607
rect 84462 127607 84526 127638
rect 84462 127574 84474 127607
rect 84474 127574 84526 127607
rect 82422 127438 82486 127502
rect 84870 127438 84934 127502
rect 87046 127574 87110 127638
rect 87318 127438 87382 127502
rect 89494 127607 89558 127638
rect 89494 127574 89522 127607
rect 89522 127574 89558 127607
rect 89766 127438 89830 127502
rect 91942 127607 92006 127638
rect 91942 127574 91962 127607
rect 91962 127574 92006 127607
rect 92350 127438 92414 127502
rect 94390 127574 94454 127638
rect 94798 127438 94862 127502
rect 96838 127574 96902 127638
rect 99422 127607 99486 127638
rect 99422 127574 99450 127607
rect 99450 127574 99486 127607
rect 117374 127710 117438 127774
rect 97382 127438 97446 127502
rect 99830 127438 99894 127502
rect 102006 127574 102070 127638
rect 102278 127438 102342 127502
rect 104454 127607 104518 127638
rect 104454 127574 104498 127607
rect 104498 127574 104518 127607
rect 107038 127574 107102 127638
rect 104862 127438 104926 127502
rect 107310 127438 107374 127502
rect 123766 127574 123830 127638
rect 123902 127438 123966 127502
rect 29790 127166 29854 127230
rect 32102 127166 32166 127230
rect 32374 127166 32438 127230
rect 34822 127166 34886 127230
rect 37134 127166 37198 127230
rect 37406 127166 37470 127230
rect 39854 127166 39918 127230
rect 42166 127166 42230 127230
rect 44886 127166 44950 127230
rect 47198 127166 47262 127230
rect 49510 127166 49574 127230
rect 49782 127166 49846 127230
rect 52230 127166 52294 127230
rect 54814 127166 54878 127230
rect 56990 127166 57054 127230
rect 57262 127166 57326 127230
rect 59574 127166 59638 127230
rect 59846 127166 59910 127230
rect 62294 127166 62358 127230
rect 64878 127166 64942 127230
rect 67054 127166 67118 127230
rect 67190 127166 67254 127230
rect 69638 127166 69702 127230
rect 72222 127166 72286 127230
rect 74534 127166 74598 127230
rect 74806 127166 74870 127230
rect 77254 127166 77318 127230
rect 79566 127166 79630 127230
rect 79838 127166 79902 127230
rect 82014 127166 82078 127230
rect 82286 127166 82350 127230
rect 84462 127166 84526 127230
rect 84598 127166 84662 127230
rect 87318 127166 87382 127230
rect 89630 127166 89694 127230
rect 92214 127166 92278 127230
rect 94662 127166 94726 127230
rect 97246 127166 97310 127230
rect 99422 127166 99486 127230
rect 99694 127166 99758 127230
rect 102278 127166 102342 127230
rect 104726 127166 104790 127230
rect 107174 127166 107238 127230
rect 1230 126350 1294 126414
rect 29790 126486 29854 126550
rect 32102 126486 32166 126550
rect 32374 126486 32438 126550
rect 34822 126486 34886 126550
rect 37134 126486 37198 126550
rect 37406 126486 37470 126550
rect 39854 126486 39918 126550
rect 42166 126486 42230 126550
rect 44886 126486 44950 126550
rect 47198 126486 47262 126550
rect 49510 126486 49574 126550
rect 49782 126486 49846 126550
rect 52230 126486 52294 126550
rect 54814 126486 54878 126550
rect 56990 126486 57054 126550
rect 57262 126486 57326 126550
rect 59574 126486 59638 126550
rect 59846 126486 59910 126550
rect 62294 126486 62358 126550
rect 64878 126486 64942 126550
rect 67054 126486 67118 126550
rect 67190 126486 67254 126550
rect 69638 126486 69702 126550
rect 72222 126486 72286 126550
rect 74534 126486 74598 126550
rect 74806 126486 74870 126550
rect 77254 126486 77318 126550
rect 79566 126486 79630 126550
rect 79838 126486 79902 126550
rect 82014 126486 82078 126550
rect 82286 126486 82350 126550
rect 84462 126486 84526 126550
rect 84598 126486 84662 126550
rect 87318 126486 87382 126550
rect 89630 126486 89694 126550
rect 87862 126350 87926 126414
rect 92214 126486 92278 126550
rect 94662 126486 94726 126550
rect 97246 126486 97310 126550
rect 99422 126486 99486 126550
rect 99694 126486 99758 126550
rect 102278 126486 102342 126550
rect 104726 126486 104790 126550
rect 107174 126486 107238 126550
rect 137502 126486 137566 126550
rect 117510 126350 117574 126414
rect 117238 126214 117302 126278
rect 123630 126214 123694 126278
rect 123766 126078 123830 126142
rect 29926 125670 29990 125734
rect 30062 125670 30126 125734
rect 32510 125670 32574 125734
rect 32646 125670 32710 125734
rect 34958 125670 35022 125734
rect 35094 125670 35158 125734
rect 37270 125670 37334 125734
rect 37406 125670 37470 125734
rect 39990 125670 40054 125734
rect 40126 125670 40190 125734
rect 42438 125670 42502 125734
rect 42574 125670 42638 125734
rect 44750 125670 44814 125734
rect 44886 125670 44950 125734
rect 47334 125670 47398 125734
rect 47470 125670 47534 125734
rect 49918 125670 49982 125734
rect 50054 125670 50118 125734
rect 52366 125670 52430 125734
rect 52502 125670 52566 125734
rect 54950 125670 55014 125734
rect 55086 125670 55150 125734
rect 57398 125670 57462 125734
rect 57534 125670 57598 125734
rect 59710 125670 59774 125734
rect 59982 125670 60046 125734
rect 62430 125670 62494 125734
rect 62566 125670 62630 125734
rect 64742 125670 64806 125734
rect 64878 125670 64942 125734
rect 67326 125670 67390 125734
rect 67462 125670 67526 125734
rect 69774 125670 69838 125734
rect 69910 125670 69974 125734
rect 72358 125670 72422 125734
rect 72494 125670 72558 125734
rect 74942 125670 75006 125734
rect 75078 125670 75142 125734
rect 77390 125670 77454 125734
rect 77526 125670 77590 125734
rect 79702 125670 79766 125734
rect 79838 125670 79902 125734
rect 82422 125670 82486 125734
rect 82558 125670 82622 125734
rect 84870 125670 84934 125734
rect 85006 125670 85070 125734
rect 87182 125670 87246 125734
rect 87318 125670 87382 125734
rect 89766 125670 89830 125734
rect 89902 125670 89966 125734
rect 92350 125670 92414 125734
rect 92486 125670 92550 125734
rect 94798 125670 94862 125734
rect 94934 125670 94998 125734
rect 97382 125670 97446 125734
rect 97518 125670 97582 125734
rect 99830 125670 99894 125734
rect 99966 125670 100030 125734
rect 102142 125670 102206 125734
rect 102414 125670 102478 125734
rect 104862 125670 104926 125734
rect 104998 125670 105062 125734
rect 107310 125670 107374 125734
rect 107446 125670 107510 125734
rect 117374 124990 117438 125054
rect 116286 124854 116350 124918
rect 1230 124582 1294 124646
rect 123902 124718 123966 124782
rect 123630 124582 123694 124646
rect 137502 124718 137566 124782
rect 30062 123766 30126 123830
rect 32646 123766 32710 123830
rect 35094 123766 35158 123830
rect 29926 123494 29990 123558
rect 37406 123766 37470 123830
rect 40126 123766 40190 123830
rect 42574 123766 42638 123830
rect 44886 123766 44950 123830
rect 47470 123766 47534 123830
rect 50054 123766 50118 123830
rect 52502 123766 52566 123830
rect 55086 123766 55150 123830
rect 57534 123766 57598 123830
rect 59982 123766 60046 123830
rect 62566 123766 62630 123830
rect 64878 123766 64942 123830
rect 67462 123766 67526 123830
rect 69910 123766 69974 123830
rect 72494 123766 72558 123830
rect 75078 123766 75142 123830
rect 77526 123766 77590 123830
rect 79838 123766 79902 123830
rect 82558 123766 82622 123830
rect 85006 123766 85070 123830
rect 87318 123766 87382 123830
rect 89902 123766 89966 123830
rect 92486 123766 92550 123830
rect 94934 123766 94998 123830
rect 97518 123766 97582 123830
rect 99966 123766 100030 123830
rect 102414 123766 102478 123830
rect 104998 123766 105062 123830
rect 107446 123766 107510 123830
rect 117374 123630 117438 123694
rect 110166 123494 110230 123558
rect 117374 123358 117438 123422
rect 123766 123358 123830 123422
rect 138182 123358 138246 123422
rect 134646 123222 134710 123286
rect 1230 123086 1294 123150
rect 137502 122950 137566 123014
rect 136193 122854 136257 122918
rect 29654 121998 29718 122062
rect 30334 121998 30398 122062
rect 30470 121998 30534 122062
rect 31694 121998 31758 122062
rect 32782 121998 32846 122062
rect 33462 121998 33526 122062
rect 34142 121998 34206 122062
rect 34686 121998 34750 122062
rect 35366 121998 35430 122062
rect 35910 121998 35974 122062
rect 37134 121998 37198 122062
rect 38494 121998 38558 122062
rect 39174 121998 39238 122062
rect 39582 121998 39646 122062
rect 40398 121998 40462 122062
rect 40942 121998 41006 122062
rect 42166 121998 42230 122062
rect 42846 121998 42910 122062
rect 43390 121998 43454 122062
rect 43934 121998 43998 122062
rect 44070 121998 44134 122062
rect 44614 121998 44678 122062
rect 45702 121998 45766 122062
rect 46654 121998 46718 122062
rect 47878 121998 47942 122062
rect 48422 121998 48486 122062
rect 49102 121998 49166 122062
rect 49238 121998 49302 122062
rect 50326 121998 50390 122062
rect 50870 121998 50934 122062
rect 52230 121998 52294 122062
rect 52910 121998 52974 122062
rect 53318 121998 53382 122062
rect 54134 121998 54198 122062
rect 54678 121998 54742 122062
rect 55358 121998 55422 122062
rect 56718 121998 56782 122062
rect 57126 121998 57190 122062
rect 58078 121998 58142 122062
rect 59166 121998 59230 122062
rect 60934 121998 60998 122062
rect 61614 121998 61678 122062
rect 62158 121998 62222 122062
rect 62838 121998 62902 122062
rect 63382 121998 63446 122062
rect 64062 121998 64126 122062
rect 64606 121998 64670 122062
rect 65694 121998 65758 122062
rect 67190 121998 67254 122062
rect 67870 121998 67934 122062
rect 68414 121998 68478 122062
rect 69094 121998 69158 122062
rect 69638 121998 69702 122062
rect 70318 121998 70382 122062
rect 70862 121998 70926 122062
rect 72086 121998 72150 122062
rect 72766 121998 72830 122062
rect 72902 121998 72966 122062
rect 73310 121998 73374 122062
rect 74126 121998 74190 122062
rect 75214 121998 75278 122062
rect 75350 121998 75414 122062
rect 75894 121998 75958 122062
rect 76574 121998 76638 122062
rect 77118 121998 77182 122062
rect 77798 121998 77862 122062
rect 78342 121998 78406 122062
rect 79566 121998 79630 122062
rect 80518 121998 80582 122062
rect 81470 121998 81534 122062
rect 81606 121998 81670 122062
rect 82830 121998 82894 122062
rect 83374 121998 83438 122062
rect 84054 121998 84118 122062
rect 84598 121998 84662 122062
rect 85414 121998 85478 122062
rect 85822 121998 85886 122062
rect 86502 121998 86566 122062
rect 87046 121998 87110 122062
rect 87862 122134 87926 122198
rect 88406 121998 88470 122062
rect 89086 121998 89150 122062
rect 89222 121998 89286 122062
rect 90310 121998 90374 122062
rect 90854 121998 90918 122062
rect 91534 121998 91598 122062
rect 92758 121998 92822 122062
rect 93302 121998 93366 122062
rect 94254 121998 94318 122062
rect 95478 121998 95542 122062
rect 97110 121998 97174 122062
rect 97790 121998 97854 122062
rect 98334 121998 98398 122062
rect 99014 121998 99078 122062
rect 99558 121998 99622 122062
rect 100782 121998 100846 122062
rect 101598 121998 101662 122062
rect 102006 121998 102070 122062
rect 103366 121998 103430 122062
rect 103910 121998 103974 122062
rect 104046 121998 104110 122062
rect 104590 121998 104654 122062
rect 105814 121998 105878 122062
rect 107038 121998 107102 122062
rect 108126 121998 108190 122062
rect 109486 121998 109550 122062
rect 123630 121862 123694 121926
rect 136822 121726 136886 121790
rect 29654 121590 29718 121654
rect 1230 121454 1294 121518
rect 30334 121590 30398 121654
rect 30470 121590 30534 121654
rect 31694 121590 31758 121654
rect 32782 121590 32846 121654
rect 33462 121590 33526 121654
rect 34142 121590 34206 121654
rect 34686 121590 34750 121654
rect 35366 121590 35430 121654
rect 35910 121590 35974 121654
rect 37134 121590 37198 121654
rect 38494 121590 38558 121654
rect 39174 121590 39238 121654
rect 39582 121590 39646 121654
rect 40398 121590 40462 121654
rect 40942 121590 41006 121654
rect 42166 121590 42230 121654
rect 42846 121590 42910 121654
rect 43390 121590 43454 121654
rect 43934 121590 43998 121654
rect 44070 121590 44134 121654
rect 44614 121590 44678 121654
rect 45702 121590 45766 121654
rect 46654 121590 46718 121654
rect 47878 121590 47942 121654
rect 48422 121590 48486 121654
rect 49102 121590 49166 121654
rect 49238 121590 49302 121654
rect 50326 121590 50390 121654
rect 50870 121590 50934 121654
rect 52230 121590 52294 121654
rect 52910 121590 52974 121654
rect 53318 121590 53382 121654
rect 54134 121590 54198 121654
rect 54678 121590 54742 121654
rect 55358 121590 55422 121654
rect 56718 121590 56782 121654
rect 57126 121590 57190 121654
rect 58078 121590 58142 121654
rect 59166 121590 59230 121654
rect 60934 121590 60998 121654
rect 61614 121590 61678 121654
rect 62158 121590 62222 121654
rect 62838 121590 62902 121654
rect 63382 121590 63446 121654
rect 64062 121590 64126 121654
rect 64606 121590 64670 121654
rect 65694 121590 65758 121654
rect 67190 121590 67254 121654
rect 67870 121590 67934 121654
rect 68414 121590 68478 121654
rect 69094 121590 69158 121654
rect 69638 121590 69702 121654
rect 70318 121590 70382 121654
rect 70862 121590 70926 121654
rect 72086 121590 72150 121654
rect 72766 121590 72830 121654
rect 72902 121590 72966 121654
rect 73310 121590 73374 121654
rect 74126 121590 74190 121654
rect 75214 121590 75278 121654
rect 75350 121590 75414 121654
rect 75894 121590 75958 121654
rect 76574 121590 76638 121654
rect 77118 121590 77182 121654
rect 77798 121590 77862 121654
rect 78342 121590 78406 121654
rect 79566 121590 79630 121654
rect 80518 121454 80582 121518
rect 81470 121590 81534 121654
rect 81606 121590 81670 121654
rect 82830 121590 82894 121654
rect 83374 121590 83438 121654
rect 84054 121590 84118 121654
rect 84598 121590 84662 121654
rect 85414 121590 85478 121654
rect 85822 121590 85886 121654
rect 86502 121590 86566 121654
rect 87046 121590 87110 121654
rect 88406 121590 88470 121654
rect 89086 121590 89150 121654
rect 89222 121590 89286 121654
rect 90310 121590 90374 121654
rect 90854 121590 90918 121654
rect 91534 121590 91598 121654
rect 92758 121590 92822 121654
rect 93302 121590 93366 121654
rect 94254 121590 94318 121654
rect 95478 121454 95542 121518
rect 97110 121590 97174 121654
rect 97790 121590 97854 121654
rect 98334 121590 98398 121654
rect 99014 121590 99078 121654
rect 99558 121590 99622 121654
rect 100782 121590 100846 121654
rect 101598 121590 101662 121654
rect 102006 121590 102070 121654
rect 103366 121590 103430 121654
rect 103910 121590 103974 121654
rect 104046 121590 104110 121654
rect 104590 121590 104654 121654
rect 105814 121590 105878 121654
rect 107038 121590 107102 121654
rect 108126 121590 108190 121654
rect 109486 121590 109550 121654
rect 111662 121454 111726 121518
rect 136822 121454 136886 121518
rect 137502 121454 137566 121518
rect 111662 121182 111726 121246
rect 29926 121046 29990 121110
rect 110166 121046 110230 121110
rect 116286 121182 116350 121246
rect 115334 121046 115398 121110
rect 21766 120502 21830 120566
rect 22310 120502 22374 120566
rect 22582 120502 22646 120566
rect 22990 120502 23054 120566
rect 115334 120638 115398 120702
rect 23398 120502 23462 120566
rect 115198 120502 115262 120566
rect 115742 120502 115806 120566
rect 116014 120502 116078 120566
rect 117374 120638 117438 120702
rect 116966 120502 117030 120566
rect 134646 120502 134710 120566
rect 134646 120366 134710 120430
rect 21766 120230 21830 120294
rect 21766 120094 21830 120158
rect 22310 120230 22374 120294
rect 22582 120230 22646 120294
rect 22582 120094 22646 120158
rect 22990 120230 23054 120294
rect 23126 120094 23190 120158
rect 23398 120230 23462 120294
rect 23534 120094 23598 120158
rect 115198 120230 115262 120294
rect 115334 120094 115398 120158
rect 115742 120230 115806 120294
rect 115742 120094 115806 120158
rect 116014 120230 116078 120294
rect 116966 120230 117030 120294
rect 116830 120094 116894 120158
rect 21766 119822 21830 119886
rect 1230 119686 1294 119750
rect 21902 119686 21966 119750
rect 22582 119822 22646 119886
rect 23126 119822 23190 119886
rect 22990 119686 23054 119750
rect 23534 119822 23598 119886
rect 23398 119686 23462 119750
rect 21902 119414 21966 119478
rect 21766 119278 21830 119342
rect 22310 119278 22374 119342
rect 22446 119278 22510 119342
rect 22990 119414 23054 119478
rect 23126 119278 23190 119342
rect 23398 119414 23462 119478
rect 23398 119278 23462 119342
rect 115334 119822 115398 119886
rect 115198 119686 115262 119750
rect 115742 119822 115806 119886
rect 115606 119686 115670 119750
rect 116558 119686 116622 119750
rect 116830 119822 116894 119886
rect 116966 119686 117030 119750
rect 137502 119686 137566 119750
rect 136822 119550 136886 119614
rect 115198 119414 115262 119478
rect 115334 119278 115398 119342
rect 115606 119414 115670 119478
rect 115742 119278 115806 119342
rect 116558 119414 116622 119478
rect 116014 119278 116078 119342
rect 116286 119278 116350 119342
rect 116966 119414 117030 119478
rect 116966 119278 117030 119342
rect 21766 119006 21830 119070
rect 22310 119006 22374 119070
rect 22446 119006 22510 119070
rect 22582 118870 22646 118934
rect 23126 119006 23190 119070
rect 22990 118870 23054 118934
rect 23398 119006 23462 119070
rect 23398 118870 23462 118934
rect 136822 119142 136886 119206
rect 115334 119006 115398 119070
rect 28566 118734 28630 118798
rect 115198 118870 115262 118934
rect 115742 119006 115806 119070
rect 115606 118870 115670 118934
rect 116014 119006 116078 119070
rect 116286 119006 116350 119070
rect 116286 118870 116350 118934
rect 116966 119006 117030 119070
rect 110302 118734 110366 118798
rect 22582 118598 22646 118662
rect 22990 118598 23054 118662
rect 22990 118462 23054 118526
rect 23398 118598 23462 118662
rect 23398 118462 23462 118526
rect 28430 118462 28494 118526
rect 28566 118462 28630 118526
rect 1230 118054 1294 118118
rect 22174 118054 22238 118118
rect 22990 118190 23054 118254
rect 23398 118190 23462 118254
rect 110302 118462 110366 118526
rect 115198 118598 115262 118662
rect 115198 118462 115262 118526
rect 115606 118598 115670 118662
rect 115606 118462 115670 118526
rect 116286 118598 116350 118662
rect 110302 118190 110366 118254
rect 115198 118190 115262 118254
rect 21766 117782 21830 117846
rect 22174 117782 22238 117846
rect 21766 117510 21830 117574
rect 21902 117374 21966 117438
rect 22446 117374 22510 117438
rect 21902 117102 21966 117166
rect 21766 116966 21830 117030
rect 22446 117102 22510 117166
rect 22990 116966 23054 117030
rect 28430 118054 28494 118118
rect 28430 117918 28494 117982
rect 28430 117646 28494 117710
rect 28566 117510 28630 117574
rect 115606 118190 115670 118254
rect 116286 118054 116350 118118
rect 137502 118054 137566 118118
rect 110302 117918 110366 117982
rect 110438 117918 110502 117982
rect 110438 117646 110502 117710
rect 110166 117510 110230 117574
rect 116286 117782 116350 117846
rect 116830 117782 116894 117846
rect 134646 117646 134710 117710
rect 23534 116966 23598 117030
rect 28430 117102 28494 117166
rect 28566 117102 28630 117166
rect 110166 117238 110230 117302
rect 116558 117374 116622 117438
rect 116830 117510 116894 117574
rect 116966 117374 117030 117438
rect 115334 116966 115398 117030
rect 115742 116966 115806 117030
rect 28430 116830 28494 116894
rect 21766 116694 21830 116758
rect 21902 116558 21966 116622
rect 22990 116694 23054 116758
rect 23126 116558 23190 116622
rect 23534 116694 23598 116758
rect 28566 116694 28630 116758
rect 116558 117102 116622 117166
rect 116966 117102 117030 117166
rect 116830 116966 116894 117030
rect 23398 116558 23462 116622
rect 1230 116286 1294 116350
rect 21902 116286 21966 116350
rect 21902 116150 21966 116214
rect 22446 116150 22510 116214
rect 23126 116286 23190 116350
rect 22990 116150 23054 116214
rect 23398 116286 23462 116350
rect 23398 116150 23462 116214
rect 28566 116286 28630 116350
rect 115334 116694 115398 116758
rect 115198 116558 115262 116622
rect 115742 116694 115806 116758
rect 115742 116558 115806 116622
rect 116558 116558 116622 116622
rect 116830 116694 116894 116758
rect 116966 116558 117030 116622
rect 115198 116286 115262 116350
rect 115198 116150 115262 116214
rect 115742 116286 115806 116350
rect 115742 116150 115806 116214
rect 116558 116286 116622 116350
rect 116014 116150 116078 116214
rect 116286 116150 116350 116214
rect 116966 116286 117030 116350
rect 116966 116150 117030 116214
rect 137502 116150 137566 116214
rect 21902 115878 21966 115942
rect 21766 115742 21830 115806
rect 22446 115878 22510 115942
rect 22174 115742 22238 115806
rect 22582 115742 22646 115806
rect 22990 115878 23054 115942
rect 23126 115742 23190 115806
rect 23398 115878 23462 115942
rect 23534 115742 23598 115806
rect 115198 115878 115262 115942
rect 115334 115742 115398 115806
rect 115742 115878 115806 115942
rect 115742 115742 115806 115806
rect 116014 115878 116078 115942
rect 116286 115878 116350 115942
rect 116966 115878 117030 115942
rect 116830 115742 116894 115806
rect 21766 115470 21830 115534
rect 21902 115334 21966 115398
rect 22174 115470 22238 115534
rect 22582 115470 22646 115534
rect 22718 115334 22782 115398
rect 23126 115470 23190 115534
rect 23126 115334 23190 115398
rect 23534 115470 23598 115534
rect 23398 115334 23462 115398
rect 115334 115470 115398 115534
rect 115334 115334 115398 115398
rect 115742 115470 115806 115534
rect 115606 115334 115670 115398
rect 116558 115334 116622 115398
rect 116830 115470 116894 115534
rect 116966 115334 117030 115398
rect 21902 115062 21966 115126
rect 22718 115062 22782 115126
rect 23126 115062 23190 115126
rect 23126 114926 23190 114990
rect 23398 115062 23462 115126
rect 23534 114926 23598 114990
rect 1230 114654 1294 114718
rect 115334 115062 115398 115126
rect 115334 114926 115398 114990
rect 115606 115062 115670 115126
rect 115742 114926 115806 114990
rect 116558 115062 116622 115126
rect 116150 114926 116214 114990
rect 116966 115062 117030 115126
rect 110302 114790 110366 114854
rect 23126 114654 23190 114718
rect 22990 114518 23054 114582
rect 23534 114654 23598 114718
rect 23398 114518 23462 114582
rect 22446 114110 22510 114174
rect 22990 114246 23054 114310
rect 23126 114110 23190 114174
rect 23398 114246 23462 114310
rect 110302 114518 110366 114582
rect 115334 114654 115398 114718
rect 115198 114518 115262 114582
rect 115742 114654 115806 114718
rect 115742 114518 115806 114582
rect 116150 114654 116214 114718
rect 115198 114246 115262 114310
rect 23398 114110 23462 114174
rect 28566 113974 28630 114038
rect 115198 114110 115262 114174
rect 115742 114246 115806 114310
rect 115606 114110 115670 114174
rect 116422 114110 116486 114174
rect 138182 114790 138246 114854
rect 135326 114654 135390 114718
rect 137502 114518 137566 114582
rect 21766 113838 21830 113902
rect 22446 113838 22510 113902
rect 23126 113838 23190 113902
rect 23398 113838 23462 113902
rect 21766 113566 21830 113630
rect 21902 113430 21966 113494
rect 22174 113430 22238 113494
rect 22446 113430 22510 113494
rect 28294 113702 28358 113766
rect 28566 113702 28630 113766
rect 115198 113838 115262 113902
rect 115606 113838 115670 113902
rect 110438 113566 110502 113630
rect 21902 113158 21966 113222
rect 1230 113022 1294 113086
rect 21902 113022 21966 113086
rect 22174 113158 22238 113222
rect 22446 113158 22510 113222
rect 22990 113022 23054 113086
rect 23398 113022 23462 113086
rect 28294 113294 28358 113358
rect 28294 113158 28358 113222
rect 110438 113294 110502 113358
rect 116422 113838 116486 113902
rect 116830 113838 116894 113902
rect 116830 113566 116894 113630
rect 116830 113430 116894 113494
rect 136822 113294 136886 113358
rect 115198 113022 115262 113086
rect 115606 113022 115670 113086
rect 28294 112886 28358 112950
rect 21902 112750 21966 112814
rect 21766 112614 21830 112678
rect 22174 112614 22238 112678
rect 22990 112750 23054 112814
rect 23126 112614 23190 112678
rect 23398 112750 23462 112814
rect 23534 112614 23598 112678
rect 21766 112342 21830 112406
rect 21902 112206 21966 112270
rect 22174 112342 22238 112406
rect 22310 112206 22374 112270
rect 23126 112342 23190 112406
rect 23126 112206 23190 112270
rect 23534 112342 23598 112406
rect 23398 112206 23462 112270
rect 28430 112342 28494 112406
rect 115198 112750 115262 112814
rect 115198 112614 115262 112678
rect 115606 112750 115670 112814
rect 115742 112614 115806 112678
rect 116150 112614 116214 112678
rect 116830 113158 116894 113222
rect 116966 113022 117030 113086
rect 136822 113022 136886 113086
rect 137502 112886 137566 112950
rect 116966 112750 117030 112814
rect 116830 112614 116894 112678
rect 136193 112679 136257 112683
rect 136193 112623 136197 112679
rect 136197 112623 136253 112679
rect 136253 112623 136257 112679
rect 136193 112619 136257 112623
rect 110302 112342 110366 112406
rect 115198 112342 115262 112406
rect 115198 112206 115262 112270
rect 115742 112342 115806 112406
rect 115742 112206 115806 112270
rect 116150 112342 116214 112406
rect 116014 112206 116078 112270
rect 116422 112206 116486 112270
rect 116830 112342 116894 112406
rect 116830 112206 116894 112270
rect 28430 112070 28494 112134
rect 21902 111934 21966 111998
rect 21902 111798 21966 111862
rect 22310 111934 22374 111998
rect 22174 111798 22238 111862
rect 22718 111798 22782 111862
rect 23126 111934 23190 111998
rect 22990 111798 23054 111862
rect 23398 111934 23462 111998
rect 110302 112070 110366 112134
rect 135326 112070 135390 112134
rect 23398 111798 23462 111862
rect 115198 111934 115262 111998
rect 115334 111798 115398 111862
rect 115742 111934 115806 111998
rect 115606 111798 115670 111862
rect 116014 111934 116078 111998
rect 116422 111934 116486 111998
rect 116014 111798 116078 111862
rect 116830 111934 116894 111998
rect 116966 111798 117030 111862
rect 21902 111526 21966 111590
rect 21766 111390 21830 111454
rect 22174 111526 22238 111590
rect 22718 111526 22782 111590
rect 22582 111390 22646 111454
rect 22990 111526 23054 111590
rect 23126 111390 23190 111454
rect 23398 111526 23462 111590
rect 23534 111390 23598 111454
rect 115334 111526 115398 111590
rect 115334 111390 115398 111454
rect 115606 111526 115670 111590
rect 115742 111390 115806 111454
rect 116014 111526 116078 111590
rect 116422 111390 116486 111454
rect 116966 111526 117030 111590
rect 116830 111390 116894 111454
rect 1230 111254 1294 111318
rect 21766 111118 21830 111182
rect 22582 111118 22646 111182
rect 22310 110982 22374 111046
rect 22446 110982 22510 111046
rect 23126 111118 23190 111182
rect 23126 110982 23190 111046
rect 23534 111118 23598 111182
rect 23398 110982 23462 111046
rect 137502 111254 137566 111318
rect 28294 110846 28358 110910
rect 115334 111118 115398 111182
rect 115198 110982 115262 111046
rect 115742 111118 115806 111182
rect 115606 110982 115670 111046
rect 116422 111118 116486 111182
rect 116558 110982 116622 111046
rect 116830 111118 116894 111182
rect 22310 110710 22374 110774
rect 22446 110710 22510 110774
rect 23126 110710 23190 110774
rect 23126 110574 23190 110638
rect 23398 110710 23462 110774
rect 23398 110574 23462 110638
rect 28294 110574 28358 110638
rect 115198 110710 115262 110774
rect 115198 110574 115262 110638
rect 115606 110710 115670 110774
rect 115742 110574 115806 110638
rect 116558 110710 116622 110774
rect 22446 110166 22510 110230
rect 23126 110302 23190 110366
rect 22990 110166 23054 110230
rect 23398 110302 23462 110366
rect 23534 110166 23598 110230
rect 115198 110302 115262 110366
rect 28566 110030 28630 110094
rect 115198 110166 115262 110230
rect 115742 110302 115806 110366
rect 115742 110166 115806 110230
rect 116014 110166 116078 110230
rect 110166 110030 110230 110094
rect 21902 109894 21966 109958
rect 22446 109894 22510 109958
rect 22310 109758 22374 109822
rect 22990 109894 23054 109958
rect 23534 109894 23598 109958
rect 28566 109758 28630 109822
rect 1230 109622 1294 109686
rect 21902 109622 21966 109686
rect 21766 109486 21830 109550
rect 22446 109622 22510 109686
rect 22446 109486 22510 109550
rect 28294 109622 28358 109686
rect 110166 109758 110230 109822
rect 110166 109622 110230 109686
rect 110302 109622 110366 109686
rect 115198 109894 115262 109958
rect 115742 109894 115806 109958
rect 116014 109894 116078 109958
rect 116966 109894 117030 109958
rect 21766 109214 21830 109278
rect 21902 109078 21966 109142
rect 22446 109214 22510 109278
rect 21902 108806 21966 108870
rect 21902 108670 21966 108734
rect 22310 108670 22374 108734
rect 23126 108670 23190 108734
rect 28294 109350 28358 109414
rect 28294 109214 28358 109278
rect 28294 108942 28358 109006
rect 28430 108806 28494 108870
rect 110166 109350 110230 109414
rect 110302 109214 110366 109278
rect 110438 109214 110502 109278
rect 110438 108942 110502 109006
rect 23398 108670 23462 108734
rect 21902 108398 21966 108462
rect 21766 108262 21830 108326
rect 22310 108398 22374 108462
rect 22174 108262 22238 108326
rect 23126 108398 23190 108462
rect 22990 108262 23054 108326
rect 23398 108398 23462 108462
rect 23534 108262 23598 108326
rect 28430 108398 28494 108462
rect 28566 108398 28630 108462
rect 115198 108670 115262 108734
rect 116150 109486 116214 109550
rect 116286 109486 116350 109550
rect 116966 109622 117030 109686
rect 116966 109486 117030 109550
rect 137502 109622 137566 109686
rect 116150 109214 116214 109278
rect 116286 109214 116350 109278
rect 116966 109214 117030 109278
rect 116966 109078 117030 109142
rect 115606 108670 115670 108734
rect 116014 108670 116078 108734
rect 116966 108806 117030 108870
rect 116966 108670 117030 108734
rect 115198 108398 115262 108462
rect 115334 108262 115398 108326
rect 115606 108398 115670 108462
rect 115742 108262 115806 108326
rect 116014 108398 116078 108462
rect 116286 108262 116350 108326
rect 116966 108398 117030 108462
rect 116830 108262 116894 108326
rect 28566 108126 28630 108190
rect 1230 107990 1294 108054
rect 21766 107990 21830 108054
rect 21902 107854 21966 107918
rect 22174 107990 22238 108054
rect 22310 107854 22374 107918
rect 22582 107854 22646 107918
rect 22990 107990 23054 108054
rect 23126 107854 23190 107918
rect 23534 107990 23598 108054
rect 23398 107854 23462 107918
rect 21902 107582 21966 107646
rect 21902 107446 21966 107510
rect 22310 107582 22374 107646
rect 22582 107582 22646 107646
rect 22446 107446 22510 107510
rect 22582 107446 22646 107510
rect 23126 107582 23190 107646
rect 22990 107446 23054 107510
rect 23398 107582 23462 107646
rect 23534 107446 23598 107510
rect 115334 107990 115398 108054
rect 115198 107854 115262 107918
rect 115742 107990 115806 108054
rect 115606 107854 115670 107918
rect 116286 107990 116350 108054
rect 116150 107854 116214 107918
rect 116422 107854 116486 107918
rect 116830 107990 116894 108054
rect 116966 107854 117030 107918
rect 137502 107990 137566 108054
rect 115198 107582 115262 107646
rect 115198 107446 115262 107510
rect 115606 107582 115670 107646
rect 115606 107446 115670 107510
rect 116150 107582 116214 107646
rect 116014 107446 116078 107510
rect 116422 107582 116486 107646
rect 116966 107582 117030 107646
rect 116966 107446 117030 107510
rect 21902 107174 21966 107238
rect 22446 107174 22510 107238
rect 22582 107174 22646 107238
rect 22174 107038 22238 107102
rect 22582 107038 22646 107102
rect 22990 107174 23054 107238
rect 23126 107038 23190 107102
rect 23534 107174 23598 107238
rect 23534 107038 23598 107102
rect 115198 107174 115262 107238
rect 115198 107038 115262 107102
rect 115606 107174 115670 107238
rect 115742 107038 115806 107102
rect 116014 107174 116078 107238
rect 116014 107038 116078 107102
rect 116966 107174 117030 107238
rect 21902 106630 21966 106694
rect 22174 106766 22238 106830
rect 22582 106766 22646 106830
rect 22718 106630 22782 106694
rect 23126 106766 23190 106830
rect 23126 106630 23190 106694
rect 23534 106766 23598 106830
rect 23398 106630 23462 106694
rect 115198 106766 115262 106830
rect 115198 106630 115262 106694
rect 115742 106766 115806 106830
rect 115606 106630 115670 106694
rect 116014 106766 116078 106830
rect 116558 106630 116622 106694
rect 116966 106630 117030 106694
rect 21902 106358 21966 106422
rect 22718 106358 22782 106422
rect 22446 106222 22510 106286
rect 23126 106358 23190 106422
rect 23126 106222 23190 106286
rect 23398 106358 23462 106422
rect 23534 106222 23598 106286
rect 1230 106086 1294 106150
rect 115198 106358 115262 106422
rect 115334 106222 115398 106286
rect 115606 106358 115670 106422
rect 115742 106222 115806 106286
rect 116558 106358 116622 106422
rect 116966 106358 117030 106422
rect 110302 106086 110366 106150
rect 137502 106222 137566 106286
rect 21766 105950 21830 106014
rect 22446 105950 22510 106014
rect 23126 105950 23190 106014
rect 22990 105814 23054 105878
rect 23534 105950 23598 106014
rect 23534 105814 23598 105878
rect 21766 105678 21830 105742
rect 22310 105406 22374 105470
rect 22446 105406 22510 105470
rect 22990 105542 23054 105606
rect 23534 105542 23598 105606
rect 110302 105814 110366 105878
rect 115334 105950 115398 106014
rect 115334 105814 115398 105878
rect 115742 105950 115806 106014
rect 115742 105814 115806 105878
rect 116830 105950 116894 106014
rect 21902 105134 21966 105198
rect 22310 105134 22374 105198
rect 22446 105134 22510 105198
rect 21902 104862 21966 104926
rect 21902 104726 21966 104790
rect 22582 104726 22646 104790
rect 22990 104726 23054 104790
rect 28294 104998 28358 105062
rect 28566 104862 28630 104926
rect 115334 105542 115398 105606
rect 115742 105542 115806 105606
rect 116422 105406 116486 105470
rect 116830 105678 116894 105742
rect 23534 104726 23598 104790
rect 28294 104726 28358 104790
rect 1230 104590 1294 104654
rect 21902 104454 21966 104518
rect 21902 104318 21966 104382
rect 22582 104454 22646 104518
rect 22990 104454 23054 104518
rect 22990 104318 23054 104382
rect 23534 104454 23598 104518
rect 23398 104318 23462 104382
rect 28430 104454 28494 104518
rect 28566 104454 28630 104518
rect 115198 104726 115262 104790
rect 115606 104726 115670 104790
rect 116422 105134 116486 105198
rect 116966 105134 117030 105198
rect 116014 104726 116078 104790
rect 116966 104862 117030 104926
rect 116966 104726 117030 104790
rect 115198 104454 115262 104518
rect 115198 104318 115262 104382
rect 115606 104454 115670 104518
rect 115606 104318 115670 104382
rect 116014 104454 116078 104518
rect 116150 104318 116214 104382
rect 116966 104454 117030 104518
rect 137502 104454 137566 104518
rect 116966 104318 117030 104382
rect 28430 104182 28494 104246
rect 21902 104046 21966 104110
rect 21766 103910 21830 103974
rect 22174 103910 22238 103974
rect 22990 104046 23054 104110
rect 23126 103910 23190 103974
rect 23398 104046 23462 104110
rect 115198 104046 115262 104110
rect 23534 103910 23598 103974
rect 115334 103910 115398 103974
rect 115606 104046 115670 104110
rect 115742 103910 115806 103974
rect 116150 104046 116214 104110
rect 116014 103910 116078 103974
rect 116966 104046 117030 104110
rect 116830 103910 116894 103974
rect 21766 103638 21830 103702
rect 21766 103502 21830 103566
rect 22174 103638 22238 103702
rect 22310 103502 22374 103566
rect 23126 103638 23190 103702
rect 23126 103502 23190 103566
rect 23534 103638 23598 103702
rect 23398 103502 23462 103566
rect 115334 103638 115398 103702
rect 115334 103502 115398 103566
rect 115742 103638 115806 103702
rect 115742 103502 115806 103566
rect 116014 103638 116078 103702
rect 116286 103502 116350 103566
rect 116830 103638 116894 103702
rect 116830 103502 116894 103566
rect 21766 103230 21830 103294
rect 21902 103094 21966 103158
rect 22310 103230 22374 103294
rect 22174 103094 22238 103158
rect 22446 103094 22510 103158
rect 23126 103230 23190 103294
rect 22990 103094 23054 103158
rect 23398 103230 23462 103294
rect 115334 103230 115398 103294
rect 23398 103094 23462 103158
rect 115334 103094 115398 103158
rect 115742 103230 115806 103294
rect 115742 103094 115806 103158
rect 116286 103230 116350 103294
rect 116830 103230 116894 103294
rect 116966 103094 117030 103158
rect 1230 102686 1294 102750
rect 21902 102822 21966 102886
rect 21766 102686 21830 102750
rect 22174 102822 22238 102886
rect 22446 102822 22510 102886
rect 22582 102686 22646 102750
rect 22990 102822 23054 102886
rect 23126 102686 23190 102750
rect 23398 102822 23462 102886
rect 23534 102686 23598 102750
rect 115334 102822 115398 102886
rect 115198 102686 115262 102750
rect 115742 102822 115806 102886
rect 115742 102686 115806 102750
rect 116150 102686 116214 102750
rect 116422 102686 116486 102750
rect 116966 102822 117030 102886
rect 116830 102686 116894 102750
rect 137502 102822 137566 102886
rect 21766 102414 21830 102478
rect 22310 102278 22374 102342
rect 22582 102414 22646 102478
rect 22718 102278 22782 102342
rect 23126 102414 23190 102478
rect 22990 102278 23054 102342
rect 23534 102414 23598 102478
rect 23398 102278 23462 102342
rect 115198 102414 115262 102478
rect 115198 102278 115262 102342
rect 115742 102414 115806 102478
rect 115606 102278 115670 102342
rect 116150 102414 116214 102478
rect 116422 102414 116486 102478
rect 116558 102278 116622 102342
rect 116830 102414 116894 102478
rect 21766 102006 21830 102070
rect 22310 102006 22374 102070
rect 22446 102006 22510 102070
rect 22718 102006 22782 102070
rect 22990 102006 23054 102070
rect 23126 101870 23190 101934
rect 23398 102006 23462 102070
rect 23534 101870 23598 101934
rect 21766 101734 21830 101798
rect 22446 101734 22510 101798
rect 22718 101462 22782 101526
rect 23126 101598 23190 101662
rect 23534 101598 23598 101662
rect 1230 101190 1294 101254
rect 21902 101190 21966 101254
rect 22718 101190 22782 101254
rect 21902 100918 21966 100982
rect 21766 100782 21830 100846
rect 22446 100782 22510 100846
rect 28294 101598 28358 101662
rect 115198 102006 115262 102070
rect 115198 101870 115262 101934
rect 115606 102006 115670 102070
rect 115606 101870 115670 101934
rect 116558 102006 116622 102070
rect 116966 102006 117030 102070
rect 28294 101326 28358 101390
rect 28566 101326 28630 101390
rect 28566 101054 28630 101118
rect 28294 100918 28358 100982
rect 115198 101598 115262 101662
rect 115606 101598 115670 101662
rect 116286 101462 116350 101526
rect 116966 101734 117030 101798
rect 110166 101326 110230 101390
rect 110166 101054 110230 101118
rect 110302 100918 110366 100982
rect 116286 101190 116350 101254
rect 116966 101190 117030 101254
rect 137502 101190 137566 101254
rect 21766 100510 21830 100574
rect 21766 100374 21830 100438
rect 22446 100510 22510 100574
rect 22990 100374 23054 100438
rect 23398 100374 23462 100438
rect 28294 100646 28358 100710
rect 28430 100374 28494 100438
rect 110302 100646 110366 100710
rect 110302 100510 110366 100574
rect 115334 100374 115398 100438
rect 116150 100782 116214 100846
rect 116422 100782 116486 100846
rect 116966 100918 117030 100982
rect 116966 100782 117030 100846
rect 115742 100374 115806 100438
rect 116150 100510 116214 100574
rect 21766 100102 21830 100166
rect 21902 99966 21966 100030
rect 22174 99966 22238 100030
rect 22990 100102 23054 100166
rect 22990 99966 23054 100030
rect 23398 100102 23462 100166
rect 110302 100238 110366 100302
rect 116422 100510 116486 100574
rect 116966 100510 117030 100574
rect 116966 100374 117030 100438
rect 23398 99966 23462 100030
rect 28430 99966 28494 100030
rect 115334 100102 115398 100166
rect 115198 99966 115262 100030
rect 115742 100102 115806 100166
rect 115606 99966 115670 100030
rect 116014 99966 116078 100030
rect 116966 100102 117030 100166
rect 116830 99966 116894 100030
rect 21902 99694 21966 99758
rect 1230 99558 1294 99622
rect 21766 99558 21830 99622
rect 22174 99694 22238 99758
rect 22174 99558 22238 99622
rect 22446 99558 22510 99622
rect 22990 99694 23054 99758
rect 22990 99558 23054 99622
rect 23398 99694 23462 99758
rect 23534 99558 23598 99622
rect 28566 99694 28630 99758
rect 115198 99694 115262 99758
rect 115198 99558 115262 99622
rect 115606 99694 115670 99758
rect 115742 99558 115806 99622
rect 116014 99694 116078 99758
rect 116286 99558 116350 99622
rect 116422 99558 116486 99622
rect 116830 99694 116894 99758
rect 116830 99558 116894 99622
rect 137502 99558 137566 99622
rect 28566 99422 28630 99486
rect 21766 99286 21830 99350
rect 21902 99150 21966 99214
rect 22174 99286 22238 99350
rect 22446 99286 22510 99350
rect 22582 99150 22646 99214
rect 22990 99286 23054 99350
rect 22990 99150 23054 99214
rect 23534 99286 23598 99350
rect 23398 99150 23462 99214
rect 115198 99286 115262 99350
rect 115198 99150 115262 99214
rect 115742 99286 115806 99350
rect 115606 99150 115670 99214
rect 116286 99286 116350 99350
rect 116422 99286 116486 99350
rect 116150 99150 116214 99214
rect 116558 99150 116622 99214
rect 116830 99286 116894 99350
rect 116966 99150 117030 99214
rect 21902 98878 21966 98942
rect 21902 98742 21966 98806
rect 22582 98878 22646 98942
rect 22174 98742 22238 98806
rect 22990 98878 23054 98942
rect 23126 98742 23190 98806
rect 23398 98878 23462 98942
rect 23398 98742 23462 98806
rect 115198 98878 115262 98942
rect 115198 98742 115262 98806
rect 115606 98878 115670 98942
rect 115606 98742 115670 98806
rect 116150 98878 116214 98942
rect 116558 98878 116622 98942
rect 116014 98742 116078 98806
rect 116966 98878 117030 98942
rect 116966 98742 117030 98806
rect 21902 98470 21966 98534
rect 22174 98470 22238 98534
rect 22174 98334 22238 98398
rect 22582 98334 22646 98398
rect 23126 98470 23190 98534
rect 22990 98334 23054 98398
rect 23398 98470 23462 98534
rect 23534 98334 23598 98398
rect 115198 98470 115262 98534
rect 115334 98334 115398 98398
rect 115606 98470 115670 98534
rect 115742 98334 115806 98398
rect 116014 98470 116078 98534
rect 116014 98334 116078 98398
rect 116422 98334 116486 98398
rect 116966 98470 117030 98534
rect 1230 97790 1294 97854
rect 22174 98062 22238 98126
rect 22582 98062 22646 98126
rect 22990 98062 23054 98126
rect 23126 97926 23190 97990
rect 23534 98062 23598 98126
rect 23398 97926 23462 97990
rect 28294 97926 28358 97990
rect 22582 97518 22646 97582
rect 23126 97654 23190 97718
rect 23126 97518 23190 97582
rect 23398 97654 23462 97718
rect 23398 97518 23462 97582
rect 115334 98062 115398 98126
rect 115198 97926 115262 97990
rect 115742 98062 115806 98126
rect 115606 97926 115670 97990
rect 116014 98062 116078 98126
rect 116422 98062 116486 98126
rect 115198 97654 115262 97718
rect 28294 97518 28358 97582
rect 115334 97518 115398 97582
rect 115606 97654 115670 97718
rect 115742 97518 115806 97582
rect 116286 97518 116350 97582
rect 137502 97790 137566 97854
rect 110166 97382 110230 97446
rect 21766 97246 21830 97310
rect 22582 97246 22646 97310
rect 23126 97246 23190 97310
rect 23398 97246 23462 97310
rect 21766 96974 21830 97038
rect 21902 96838 21966 96902
rect 22718 96838 22782 96902
rect 21902 96566 21966 96630
rect 21766 96430 21830 96494
rect 22718 96566 22782 96630
rect 22990 96430 23054 96494
rect 28430 96974 28494 97038
rect 110166 97110 110230 97174
rect 115334 97246 115398 97310
rect 115742 97246 115806 97310
rect 110302 96974 110366 97038
rect 28430 96702 28494 96766
rect 23534 96430 23598 96494
rect 110302 96702 110366 96766
rect 116286 97246 116350 97310
rect 116830 97246 116894 97310
rect 116558 96838 116622 96902
rect 116830 96974 116894 97038
rect 116966 96838 117030 96902
rect 115334 96430 115398 96494
rect 115742 96430 115806 96494
rect 116558 96566 116622 96630
rect 116286 96430 116350 96494
rect 116966 96566 117030 96630
rect 116966 96430 117030 96494
rect 1230 96158 1294 96222
rect 21766 96158 21830 96222
rect 21902 96022 21966 96086
rect 22174 96022 22238 96086
rect 22718 96022 22782 96086
rect 22990 96158 23054 96222
rect 22990 96022 23054 96086
rect 23534 96158 23598 96222
rect 23398 96022 23462 96086
rect 21902 95750 21966 95814
rect 21902 95614 21966 95678
rect 22174 95750 22238 95814
rect 22718 95750 22782 95814
rect 22990 95750 23054 95814
rect 22990 95614 23054 95678
rect 23398 95750 23462 95814
rect 23398 95614 23462 95678
rect 28430 95750 28494 95814
rect 115334 96158 115398 96222
rect 115334 96022 115398 96086
rect 115742 96158 115806 96222
rect 115742 96022 115806 96086
rect 116286 96158 116350 96222
rect 116558 96022 116622 96086
rect 116966 96158 117030 96222
rect 116966 96022 117030 96086
rect 137502 96022 137566 96086
rect 110166 95750 110230 95814
rect 115334 95750 115398 95814
rect 115198 95614 115262 95678
rect 115742 95750 115806 95814
rect 115606 95614 115670 95678
rect 116558 95750 116622 95814
rect 116150 95614 116214 95678
rect 116966 95750 117030 95814
rect 116966 95614 117030 95678
rect 28430 95478 28494 95542
rect 21902 95342 21966 95406
rect 21766 95206 21830 95270
rect 22174 95206 22238 95270
rect 22582 95206 22646 95270
rect 22990 95342 23054 95406
rect 23126 95206 23190 95270
rect 23398 95342 23462 95406
rect 23534 95206 23598 95270
rect 110166 95478 110230 95542
rect 115198 95342 115262 95406
rect 115334 95206 115398 95270
rect 115606 95342 115670 95406
rect 115742 95206 115806 95270
rect 116150 95342 116214 95406
rect 116014 95206 116078 95270
rect 116422 95206 116486 95270
rect 116966 95342 117030 95406
rect 116830 95206 116894 95270
rect 21766 94934 21830 94998
rect 21902 94798 21966 94862
rect 22174 94934 22238 94998
rect 22310 94798 22374 94862
rect 22582 94934 22646 94998
rect 23126 94934 23190 94998
rect 23126 94798 23190 94862
rect 23534 94934 23598 94998
rect 23534 94798 23598 94862
rect 115334 94934 115398 94998
rect 115198 94798 115262 94862
rect 115742 94934 115806 94998
rect 115606 94798 115670 94862
rect 116014 94934 116078 94998
rect 116422 94934 116486 94998
rect 116830 94934 116894 94998
rect 116830 94798 116894 94862
rect 1230 94526 1294 94590
rect 21902 94526 21966 94590
rect 22310 94526 22374 94590
rect 22582 94390 22646 94454
rect 23126 94526 23190 94590
rect 23126 94390 23190 94454
rect 23534 94526 23598 94590
rect 115198 94526 115262 94590
rect 23398 94390 23462 94454
rect 115334 94390 115398 94454
rect 115606 94526 115670 94590
rect 115606 94390 115670 94454
rect 116014 94390 116078 94454
rect 116286 94390 116350 94454
rect 116830 94526 116894 94590
rect 137502 94390 137566 94454
rect 110166 94254 110230 94318
rect 22582 94118 22646 94182
rect 23126 94118 23190 94182
rect 23126 93982 23190 94046
rect 23398 94118 23462 94182
rect 23534 93982 23598 94046
rect 22446 93574 22510 93638
rect 23126 93710 23190 93774
rect 22990 93574 23054 93638
rect 23534 93710 23598 93774
rect 23398 93574 23462 93638
rect 110166 93982 110230 94046
rect 115334 94118 115398 94182
rect 115334 93982 115398 94046
rect 115606 94118 115670 94182
rect 115742 93982 115806 94046
rect 116014 94118 116078 94182
rect 116286 94118 116350 94182
rect 28566 93438 28630 93502
rect 115334 93710 115398 93774
rect 115198 93574 115262 93638
rect 115742 93710 115806 93774
rect 115606 93574 115670 93638
rect 116422 93574 116486 93638
rect 21902 93302 21966 93366
rect 22446 93302 22510 93366
rect 22990 93302 23054 93366
rect 23398 93302 23462 93366
rect 21902 93030 21966 93094
rect 1230 92894 1294 92958
rect 21766 92894 21830 92958
rect 22582 92894 22646 92958
rect 28566 93166 28630 93230
rect 28294 93030 28358 93094
rect 110302 93030 110366 93094
rect 115198 93302 115262 93366
rect 115606 93302 115670 93366
rect 116422 93302 116486 93366
rect 116830 93302 116894 93366
rect 21766 92622 21830 92686
rect 21902 92486 21966 92550
rect 22582 92622 22646 92686
rect 21902 92214 21966 92278
rect 21766 92078 21830 92142
rect 22446 92078 22510 92142
rect 23126 92078 23190 92142
rect 28294 92758 28358 92822
rect 28566 92622 28630 92686
rect 28430 92350 28494 92414
rect 28566 92350 28630 92414
rect 23534 92078 23598 92142
rect 28430 92078 28494 92142
rect 21766 91806 21830 91870
rect 21766 91670 21830 91734
rect 22446 91806 22510 91870
rect 22310 91670 22374 91734
rect 22718 91670 22782 91734
rect 23126 91806 23190 91870
rect 22990 91670 23054 91734
rect 23534 91806 23598 91870
rect 23534 91670 23598 91734
rect 110302 92758 110366 92822
rect 116422 92894 116486 92958
rect 116830 93030 116894 93094
rect 116830 92894 116894 92958
rect 137502 92894 137566 92958
rect 110302 92622 110366 92686
rect 110302 92350 110366 92414
rect 116422 92622 116486 92686
rect 116830 92622 116894 92686
rect 116966 92486 117030 92550
rect 115334 92078 115398 92142
rect 115606 92078 115670 92142
rect 116286 92078 116350 92142
rect 116966 92214 117030 92278
rect 116966 92078 117030 92142
rect 110438 91806 110502 91870
rect 115334 91806 115398 91870
rect 115334 91670 115398 91734
rect 115606 91806 115670 91870
rect 115606 91670 115670 91734
rect 116286 91806 116350 91870
rect 116150 91670 116214 91734
rect 116966 91806 117030 91870
rect 116966 91670 117030 91734
rect 21766 91398 21830 91462
rect 21902 91262 21966 91326
rect 22310 91398 22374 91462
rect 22718 91398 22782 91462
rect 22174 91262 22238 91326
rect 22718 91262 22782 91326
rect 22990 91398 23054 91462
rect 22990 91262 23054 91326
rect 23534 91398 23598 91462
rect 23398 91262 23462 91326
rect 110438 91534 110502 91598
rect 1230 91126 1294 91190
rect 115334 91398 115398 91462
rect 115198 91262 115262 91326
rect 115606 91398 115670 91462
rect 115606 91262 115670 91326
rect 116150 91398 116214 91462
rect 116150 91262 116214 91326
rect 116966 91398 117030 91462
rect 116966 91262 117030 91326
rect 137502 91126 137566 91190
rect 21902 90990 21966 91054
rect 21766 90854 21830 90918
rect 22174 90990 22238 91054
rect 22174 90854 22238 90918
rect 22718 90990 22782 91054
rect 22582 90854 22646 90918
rect 22990 90990 23054 91054
rect 22990 90854 23054 90918
rect 23398 90990 23462 91054
rect 23534 90854 23598 90918
rect 115198 90990 115262 91054
rect 115334 90854 115398 90918
rect 115606 90990 115670 91054
rect 115742 90854 115806 90918
rect 116150 90990 116214 91054
rect 116422 90854 116486 90918
rect 116966 90990 117030 91054
rect 116830 90854 116894 90918
rect 21766 90582 21830 90646
rect 22174 90582 22238 90646
rect 22582 90582 22646 90646
rect 22446 90446 22510 90510
rect 22990 90582 23054 90646
rect 23126 90446 23190 90510
rect 23534 90582 23598 90646
rect 115334 90582 115398 90646
rect 23534 90446 23598 90510
rect 115334 90446 115398 90510
rect 115742 90582 115806 90646
rect 115742 90446 115806 90510
rect 116422 90582 116486 90646
rect 116150 90446 116214 90510
rect 116286 90446 116350 90510
rect 116830 90582 116894 90646
rect 21766 90038 21830 90102
rect 22446 90174 22510 90238
rect 22174 90038 22238 90102
rect 23126 90174 23190 90238
rect 22990 90038 23054 90102
rect 23534 90174 23598 90238
rect 23534 90038 23598 90102
rect 115334 90174 115398 90238
rect 115198 90038 115262 90102
rect 115742 90174 115806 90238
rect 115742 90038 115806 90102
rect 116150 90174 116214 90238
rect 116286 90174 116350 90238
rect 116014 90038 116078 90102
rect 116286 90038 116350 90102
rect 116830 90038 116894 90102
rect 21766 89766 21830 89830
rect 22174 89766 22238 89830
rect 22582 89630 22646 89694
rect 22990 89766 23054 89830
rect 22990 89630 23054 89694
rect 23534 89766 23598 89830
rect 23534 89630 23598 89694
rect 1230 89494 1294 89558
rect 28294 89494 28358 89558
rect 115198 89766 115262 89830
rect 115198 89630 115262 89694
rect 115742 89766 115806 89830
rect 115742 89630 115806 89694
rect 116014 89766 116078 89830
rect 116286 89766 116350 89830
rect 116830 89766 116894 89830
rect 21766 89358 21830 89422
rect 22582 89358 22646 89422
rect 22446 89222 22510 89286
rect 22990 89358 23054 89422
rect 23534 89358 23598 89422
rect 28294 89222 28358 89286
rect 115198 89358 115262 89422
rect 115742 89358 115806 89422
rect 116966 89358 117030 89422
rect 137502 89494 137566 89558
rect 21766 89086 21830 89150
rect 21902 88950 21966 89014
rect 22174 88950 22238 89014
rect 22446 88950 22510 89014
rect 110166 88950 110230 89014
rect 21902 88678 21966 88742
rect 21766 88542 21830 88606
rect 22174 88542 22238 88606
rect 21766 88270 21830 88334
rect 21902 88134 21966 88198
rect 22718 88134 22782 88198
rect 23126 88134 23190 88198
rect 116558 88950 116622 89014
rect 116966 89086 117030 89150
rect 116830 88950 116894 89014
rect 110166 88678 110230 88742
rect 110302 88678 110366 88742
rect 110302 88406 110366 88470
rect 110438 88406 110502 88470
rect 116830 88678 116894 88742
rect 116558 88542 116622 88606
rect 116830 88542 116894 88606
rect 116286 88406 116350 88470
rect 23398 88134 23462 88198
rect 21902 87862 21966 87926
rect 21766 87726 21830 87790
rect 22718 87862 22782 87926
rect 23126 87862 23190 87926
rect 23126 87726 23190 87790
rect 23398 87862 23462 87926
rect 23534 87726 23598 87790
rect 28294 87862 28358 87926
rect 110438 88134 110502 88198
rect 115198 88134 115262 88198
rect 115606 88134 115670 88198
rect 116286 88134 116350 88198
rect 116558 88134 116622 88198
rect 116830 88270 116894 88334
rect 116966 88134 117030 88198
rect 115198 87862 115262 87926
rect 115334 87726 115398 87790
rect 115606 87862 115670 87926
rect 115742 87726 115806 87790
rect 116558 87862 116622 87926
rect 116150 87726 116214 87790
rect 116286 87726 116350 87790
rect 116422 87726 116486 87790
rect 116966 87862 117030 87926
rect 116966 87726 117030 87790
rect 1230 87590 1294 87654
rect 137502 87726 137566 87790
rect 28294 87590 28358 87654
rect 21766 87454 21830 87518
rect 21766 87318 21830 87382
rect 22174 87318 22238 87382
rect 22582 87318 22646 87382
rect 23126 87454 23190 87518
rect 22990 87318 23054 87382
rect 23534 87454 23598 87518
rect 23534 87318 23598 87382
rect 115334 87454 115398 87518
rect 115198 87318 115262 87382
rect 115742 87454 115806 87518
rect 115742 87318 115806 87382
rect 116150 87454 116214 87518
rect 116286 87454 116350 87518
rect 116422 87454 116486 87518
rect 116014 87318 116078 87382
rect 116286 87318 116350 87382
rect 116966 87454 117030 87518
rect 116966 87318 117030 87382
rect 21766 87046 21830 87110
rect 21902 86910 21966 86974
rect 22174 87046 22238 87110
rect 22582 87046 22646 87110
rect 22990 87046 23054 87110
rect 23126 86910 23190 86974
rect 23534 87046 23598 87110
rect 23398 86910 23462 86974
rect 115198 87046 115262 87110
rect 115198 86910 115262 86974
rect 115742 87046 115806 87110
rect 115606 86910 115670 86974
rect 116014 87046 116078 87110
rect 116286 87046 116350 87110
rect 116150 86910 116214 86974
rect 116966 87046 117030 87110
rect 116966 86910 117030 86974
rect 21902 86638 21966 86702
rect 21766 86502 21830 86566
rect 22446 86502 22510 86566
rect 23126 86638 23190 86702
rect 22990 86502 23054 86566
rect 23398 86638 23462 86702
rect 23534 86502 23598 86566
rect 115198 86638 115262 86702
rect 115334 86502 115398 86566
rect 115606 86638 115670 86702
rect 115742 86502 115806 86566
rect 116150 86638 116214 86702
rect 116014 86502 116078 86566
rect 116422 86502 116486 86566
rect 116966 86638 117030 86702
rect 116830 86502 116894 86566
rect 21766 86230 21830 86294
rect 1230 86094 1294 86158
rect 21766 86094 21830 86158
rect 22446 86230 22510 86294
rect 22310 86094 22374 86158
rect 22990 86230 23054 86294
rect 22990 86094 23054 86158
rect 23534 86230 23598 86294
rect 23534 86094 23598 86158
rect 21766 85822 21830 85886
rect 22310 85822 22374 85886
rect 22446 85686 22510 85750
rect 22718 85686 22782 85750
rect 22990 85822 23054 85886
rect 22990 85686 23054 85750
rect 23534 85822 23598 85886
rect 115334 86230 115398 86294
rect 115334 86094 115398 86158
rect 115742 86230 115806 86294
rect 115606 86094 115670 86158
rect 116014 86230 116078 86294
rect 116422 86230 116486 86294
rect 116830 86230 116894 86294
rect 116830 86094 116894 86158
rect 137502 85958 137566 86022
rect 23534 85686 23598 85750
rect 115334 85822 115398 85886
rect 115334 85686 115398 85750
rect 115606 85822 115670 85886
rect 115606 85686 115670 85750
rect 116014 85686 116078 85750
rect 116830 85822 116894 85886
rect 110166 85550 110230 85614
rect 21766 85414 21830 85478
rect 22446 85414 22510 85478
rect 22718 85414 22782 85478
rect 22990 85414 23054 85478
rect 22990 85278 23054 85342
rect 23534 85414 23598 85478
rect 23534 85278 23598 85342
rect 21766 85142 21830 85206
rect 22718 84870 22782 84934
rect 22990 85006 23054 85070
rect 23534 85006 23598 85070
rect 110166 85278 110230 85342
rect 115334 85414 115398 85478
rect 115334 85278 115398 85342
rect 115606 85414 115670 85478
rect 115742 85278 115806 85342
rect 116014 85414 116078 85478
rect 116966 85414 117030 85478
rect 21902 84598 21966 84662
rect 22718 84598 22782 84662
rect 1230 84326 1294 84390
rect 28566 84734 28630 84798
rect 28566 84462 28630 84526
rect 21902 84326 21966 84390
rect 21766 84190 21830 84254
rect 22582 84190 22646 84254
rect 28430 84326 28494 84390
rect 110166 84326 110230 84390
rect 115334 85006 115398 85070
rect 115742 85006 115806 85070
rect 116558 84870 116622 84934
rect 116966 85142 117030 85206
rect 116558 84598 116622 84662
rect 116966 84598 117030 84662
rect 137502 84462 137566 84526
rect 21766 83918 21830 83982
rect 21902 83782 21966 83846
rect 22582 83918 22646 83982
rect 23126 83782 23190 83846
rect 23398 83782 23462 83846
rect 28430 84054 28494 84118
rect 28430 83918 28494 83982
rect 110166 84054 110230 84118
rect 116966 84326 117030 84390
rect 116830 84190 116894 84254
rect 115198 83782 115262 83846
rect 115606 83782 115670 83846
rect 28430 83646 28494 83710
rect 21902 83510 21966 83574
rect 21766 83374 21830 83438
rect 22310 83374 22374 83438
rect 23126 83510 23190 83574
rect 22990 83374 23054 83438
rect 23398 83510 23462 83574
rect 116830 83918 116894 83982
rect 116966 83782 117030 83846
rect 115198 83510 115262 83574
rect 23398 83374 23462 83438
rect 115198 83374 115262 83438
rect 115606 83510 115670 83574
rect 115742 83374 115806 83438
rect 116014 83374 116078 83438
rect 116422 83374 116486 83438
rect 116966 83510 117030 83574
rect 116966 83374 117030 83438
rect 21766 83102 21830 83166
rect 21766 82966 21830 83030
rect 22310 83102 22374 83166
rect 22174 82966 22238 83030
rect 22582 82966 22646 83030
rect 22990 83102 23054 83166
rect 22990 82966 23054 83030
rect 23398 83102 23462 83166
rect 23398 82966 23462 83030
rect 115198 83102 115262 83166
rect 115198 82966 115262 83030
rect 115742 83102 115806 83166
rect 115742 82966 115806 83030
rect 116014 83102 116078 83166
rect 116014 82966 116078 83030
rect 116422 83102 116486 83166
rect 116966 83102 117030 83166
rect 116830 82966 116894 83030
rect 1230 82694 1294 82758
rect 21766 82694 21830 82758
rect 21902 82558 21966 82622
rect 22174 82694 22238 82758
rect 22582 82694 22646 82758
rect 22446 82558 22510 82622
rect 22990 82694 23054 82758
rect 23126 82558 23190 82622
rect 23398 82694 23462 82758
rect 115198 82694 115262 82758
rect 23398 82558 23462 82622
rect 115198 82558 115262 82622
rect 115742 82694 115806 82758
rect 115606 82558 115670 82622
rect 116014 82694 116078 82758
rect 116014 82558 116078 82622
rect 116830 82694 116894 82758
rect 116966 82558 117030 82622
rect 137502 82694 137566 82758
rect 21902 82286 21966 82350
rect 21766 82150 21830 82214
rect 22446 82286 22510 82350
rect 22582 82150 22646 82214
rect 23126 82286 23190 82350
rect 23126 82150 23190 82214
rect 23398 82286 23462 82350
rect 23534 82150 23598 82214
rect 21766 81878 21830 81942
rect 22310 81742 22374 81806
rect 22582 81878 22646 81942
rect 22582 81742 22646 81806
rect 23126 81878 23190 81942
rect 23126 81742 23190 81806
rect 23534 81878 23598 81942
rect 115198 82286 115262 82350
rect 115334 82150 115398 82214
rect 115606 82286 115670 82350
rect 115742 82150 115806 82214
rect 116014 82286 116078 82350
rect 116014 82150 116078 82214
rect 116422 82150 116486 82214
rect 116966 82286 117030 82350
rect 116830 82150 116894 82214
rect 115334 81878 115398 81942
rect 23534 81742 23598 81806
rect 115198 81742 115262 81806
rect 115742 81878 115806 81942
rect 115606 81742 115670 81806
rect 116014 81878 116078 81942
rect 116422 81878 116486 81942
rect 116286 81742 116350 81806
rect 116830 81878 116894 81942
rect 22310 81470 22374 81534
rect 22582 81470 22646 81534
rect 23126 81470 23190 81534
rect 22990 81334 23054 81398
rect 23534 81470 23598 81534
rect 23534 81334 23598 81398
rect 1230 81062 1294 81126
rect 22174 80926 22238 80990
rect 22990 81062 23054 81126
rect 23534 81062 23598 81126
rect 28294 81062 28358 81126
rect 115198 81470 115262 81534
rect 115198 81334 115262 81398
rect 115606 81470 115670 81534
rect 115606 81334 115670 81398
rect 116286 81470 116350 81534
rect 21902 80654 21966 80718
rect 22174 80654 22238 80718
rect 22446 80518 22510 80582
rect 21902 80382 21966 80446
rect 21902 80246 21966 80310
rect 22446 80246 22510 80310
rect 22718 80246 22782 80310
rect 28294 80790 28358 80854
rect 28566 80790 28630 80854
rect 28566 80518 28630 80582
rect 28294 80382 28358 80446
rect 115198 81062 115262 81126
rect 115606 81062 115670 81126
rect 116150 80926 116214 80990
rect 137502 81062 137566 81126
rect 110438 80382 110502 80446
rect 116150 80654 116214 80718
rect 116830 80654 116894 80718
rect 21902 79974 21966 80038
rect 21766 79838 21830 79902
rect 22718 79974 22782 80038
rect 21766 79566 21830 79630
rect 1230 79430 1294 79494
rect 21902 79430 21966 79494
rect 22990 79838 23054 79902
rect 23534 79838 23598 79902
rect 28294 80110 28358 80174
rect 110438 80110 110502 80174
rect 116014 80246 116078 80310
rect 116286 80246 116350 80310
rect 116830 80382 116894 80446
rect 116830 80246 116894 80310
rect 110166 79974 110230 80038
rect 115334 79838 115398 79902
rect 115742 79838 115806 79902
rect 116014 79974 116078 80038
rect 116286 79974 116350 80038
rect 22718 79430 22782 79494
rect 22990 79566 23054 79630
rect 23126 79430 23190 79494
rect 23534 79566 23598 79630
rect 110166 79702 110230 79766
rect 116830 79974 116894 80038
rect 116830 79838 116894 79902
rect 116286 79702 116350 79766
rect 115334 79566 115398 79630
rect 23398 79430 23462 79494
rect 21902 79158 21966 79222
rect 21766 79022 21830 79086
rect 22718 79158 22782 79222
rect 23126 79158 23190 79222
rect 23126 79022 23190 79086
rect 23398 79158 23462 79222
rect 23398 79022 23462 79086
rect 28294 79158 28358 79222
rect 115198 79430 115262 79494
rect 115742 79566 115806 79630
rect 115606 79430 115670 79494
rect 116286 79430 116350 79494
rect 116558 79430 116622 79494
rect 116830 79566 116894 79630
rect 116966 79430 117030 79494
rect 137502 79430 137566 79494
rect 115198 79158 115262 79222
rect 115198 79022 115262 79086
rect 115606 79158 115670 79222
rect 115742 79022 115806 79086
rect 116558 79158 116622 79222
rect 116014 79022 116078 79086
rect 116966 79158 117030 79222
rect 116966 79022 117030 79086
rect 28294 78886 28358 78950
rect 21766 78750 21830 78814
rect 21902 78614 21966 78678
rect 22310 78614 22374 78678
rect 22582 78614 22646 78678
rect 23126 78750 23190 78814
rect 22990 78614 23054 78678
rect 23398 78750 23462 78814
rect 115198 78750 115262 78814
rect 23398 78614 23462 78678
rect 115334 78614 115398 78678
rect 115742 78750 115806 78814
rect 115742 78614 115806 78678
rect 116014 78750 116078 78814
rect 116014 78614 116078 78678
rect 116966 78750 117030 78814
rect 116966 78614 117030 78678
rect 21902 78342 21966 78406
rect 21902 78206 21966 78270
rect 22310 78342 22374 78406
rect 22582 78342 22646 78406
rect 22310 78206 22374 78270
rect 22990 78342 23054 78406
rect 22990 78206 23054 78270
rect 23398 78342 23462 78406
rect 23398 78206 23462 78270
rect 115334 78342 115398 78406
rect 115334 78206 115398 78270
rect 115742 78342 115806 78406
rect 115606 78206 115670 78270
rect 116014 78342 116078 78406
rect 116014 78206 116078 78270
rect 116966 78342 117030 78406
rect 116966 78206 117030 78270
rect 21902 77934 21966 77998
rect 22310 77934 22374 77998
rect 22446 77798 22510 77862
rect 22990 77934 23054 77998
rect 23126 77798 23190 77862
rect 23398 77934 23462 77998
rect 23534 77798 23598 77862
rect 115334 77934 115398 77998
rect 1230 77662 1294 77726
rect 28294 77662 28358 77726
rect 115334 77798 115398 77862
rect 115606 77934 115670 77998
rect 115742 77798 115806 77862
rect 116014 77934 116078 77998
rect 116286 77798 116350 77862
rect 116966 77934 117030 77998
rect 110438 77662 110502 77726
rect 22446 77526 22510 77590
rect 23126 77526 23190 77590
rect 22990 77390 23054 77454
rect 23534 77526 23598 77590
rect 23398 77390 23462 77454
rect 28294 77390 28358 77454
rect 22582 76982 22646 77046
rect 22990 77118 23054 77182
rect 22990 76982 23054 77046
rect 23398 77118 23462 77182
rect 110438 77390 110502 77454
rect 115334 77526 115398 77590
rect 115334 77390 115398 77454
rect 115742 77526 115806 77590
rect 115606 77390 115670 77454
rect 116286 77526 116350 77590
rect 137502 77526 137566 77590
rect 115334 77118 115398 77182
rect 23534 76982 23598 77046
rect 115334 76982 115398 77046
rect 115606 77118 115670 77182
rect 115742 76982 115806 77046
rect 116014 76982 116078 77046
rect 110438 76846 110502 76910
rect 21766 76710 21830 76774
rect 22582 76710 22646 76774
rect 22990 76710 23054 76774
rect 23534 76710 23598 76774
rect 21766 76438 21830 76502
rect 21902 76302 21966 76366
rect 22582 76302 22646 76366
rect 28294 76438 28358 76502
rect 110438 76574 110502 76638
rect 115334 76710 115398 76774
rect 110302 76438 110366 76502
rect 28294 76166 28358 76230
rect 1230 75894 1294 75958
rect 21902 76030 21966 76094
rect 21766 75894 21830 75958
rect 22582 76030 22646 76094
rect 21766 75622 21830 75686
rect 21766 75486 21830 75550
rect 22446 75486 22510 75550
rect 22990 75486 23054 75550
rect 28566 76030 28630 76094
rect 28566 75758 28630 75822
rect 110302 76166 110366 76230
rect 115742 76710 115806 76774
rect 116014 76710 116078 76774
rect 116150 76302 116214 76366
rect 116830 76710 116894 76774
rect 116558 76302 116622 76366
rect 116830 76438 116894 76502
rect 116966 76302 117030 76366
rect 116150 76030 116214 76094
rect 116558 76030 116622 76094
rect 116966 76030 117030 76094
rect 116830 75894 116894 75958
rect 137502 75894 137566 75958
rect 23534 75486 23598 75550
rect 21766 75214 21830 75278
rect 21902 75078 21966 75142
rect 22446 75214 22510 75278
rect 22718 75078 22782 75142
rect 22990 75214 23054 75278
rect 23126 75078 23190 75142
rect 23534 75214 23598 75278
rect 23398 75078 23462 75142
rect 28430 75214 28494 75278
rect 115334 75486 115398 75550
rect 115742 75486 115806 75550
rect 116150 75486 116214 75550
rect 116422 75486 116486 75550
rect 116830 75622 116894 75686
rect 116830 75486 116894 75550
rect 115334 75214 115398 75278
rect 115198 75078 115262 75142
rect 115742 75214 115806 75278
rect 115606 75078 115670 75142
rect 116150 75214 116214 75278
rect 116422 75214 116486 75278
rect 116558 75078 116622 75142
rect 116830 75214 116894 75278
rect 116966 75078 117030 75142
rect 28430 74942 28494 75006
rect 21902 74806 21966 74870
rect 21766 74670 21830 74734
rect 22718 74806 22782 74870
rect 22174 74670 22238 74734
rect 22446 74670 22510 74734
rect 23126 74806 23190 74870
rect 23126 74670 23190 74734
rect 23398 74806 23462 74870
rect 23398 74670 23462 74734
rect 115198 74806 115262 74870
rect 115198 74670 115262 74734
rect 115606 74806 115670 74870
rect 115606 74670 115670 74734
rect 116558 74806 116622 74870
rect 116014 74670 116078 74734
rect 116966 74806 117030 74870
rect 116966 74670 117030 74734
rect 21766 74398 21830 74462
rect 21766 74262 21830 74326
rect 22174 74398 22238 74462
rect 22446 74398 22510 74462
rect 22582 74262 22646 74326
rect 23126 74398 23190 74462
rect 22990 74262 23054 74326
rect 23398 74398 23462 74462
rect 23398 74262 23462 74326
rect 115198 74398 115262 74462
rect 115198 74262 115262 74326
rect 115606 74398 115670 74462
rect 115606 74262 115670 74326
rect 116014 74398 116078 74462
rect 116014 74262 116078 74326
rect 116966 74398 117030 74462
rect 116966 74262 117030 74326
rect 137502 74262 137566 74326
rect 1230 74126 1294 74190
rect 21766 73990 21830 74054
rect 22582 73990 22646 74054
rect 22718 73854 22782 73918
rect 22990 73990 23054 74054
rect 22990 73854 23054 73918
rect 23398 73990 23462 74054
rect 23398 73854 23462 73918
rect 115198 73990 115262 74054
rect 115198 73854 115262 73918
rect 115606 73990 115670 74054
rect 115606 73854 115670 73918
rect 116014 73990 116078 74054
rect 116150 73854 116214 73918
rect 116966 73990 117030 74054
rect 21902 73446 21966 73510
rect 22718 73582 22782 73646
rect 22174 73446 22238 73510
rect 22990 73582 23054 73646
rect 22990 73446 23054 73510
rect 23398 73582 23462 73646
rect 23534 73446 23598 73510
rect 115198 73582 115262 73646
rect 115334 73446 115398 73510
rect 115606 73582 115670 73646
rect 115742 73446 115806 73510
rect 116150 73582 116214 73646
rect 116014 73446 116078 73510
rect 116830 73446 116894 73510
rect 21902 73174 21966 73238
rect 22174 73174 22238 73238
rect 22446 73038 22510 73102
rect 22990 73174 23054 73238
rect 22990 73038 23054 73102
rect 23534 73174 23598 73238
rect 23398 73038 23462 73102
rect 28430 72902 28494 72966
rect 21902 72766 21966 72830
rect 22446 72766 22510 72830
rect 1230 72630 1294 72694
rect 21902 72494 21966 72558
rect 21766 72358 21830 72422
rect 22174 72358 22238 72422
rect 22582 72358 22646 72422
rect 22990 72766 23054 72830
rect 23398 72766 23462 72830
rect 28430 72630 28494 72694
rect 28430 72494 28494 72558
rect 115334 73174 115398 73238
rect 115334 73038 115398 73102
rect 115742 73174 115806 73238
rect 115742 73038 115806 73102
rect 116014 73174 116078 73238
rect 116014 73038 116078 73102
rect 116422 73038 116486 73102
rect 116830 73174 116894 73238
rect 110438 72494 110502 72558
rect 115334 72766 115398 72830
rect 115742 72766 115806 72830
rect 116014 72766 116078 72830
rect 116422 72766 116486 72830
rect 116966 72766 117030 72830
rect 137502 72630 137566 72694
rect 21766 72086 21830 72150
rect 21902 71950 21966 72014
rect 22174 72086 22238 72150
rect 22582 72086 22646 72150
rect 21902 71678 21966 71742
rect 21902 71542 21966 71606
rect 22446 71542 22510 71606
rect 22718 71542 22782 71606
rect 22990 71542 23054 71606
rect 28430 72222 28494 72286
rect 28294 72086 28358 72150
rect 28294 71814 28358 71878
rect 23534 71542 23598 71606
rect 21902 71270 21966 71334
rect 21766 71134 21830 71198
rect 22446 71270 22510 71334
rect 22718 71270 22782 71334
rect 22174 71134 22238 71198
rect 22582 71134 22646 71198
rect 22990 71270 23054 71334
rect 22990 71134 23054 71198
rect 23534 71270 23598 71334
rect 23534 71134 23598 71198
rect 110438 72222 110502 72286
rect 116014 72358 116078 72422
rect 116966 72494 117030 72558
rect 116830 72358 116894 72422
rect 116014 72086 116078 72150
rect 116830 72086 116894 72150
rect 116830 71950 116894 72014
rect 115198 71542 115262 71606
rect 115742 71542 115806 71606
rect 116014 71542 116078 71606
rect 116286 71542 116350 71606
rect 116830 71678 116894 71742
rect 116830 71542 116894 71606
rect 115198 71270 115262 71334
rect 115334 71134 115398 71198
rect 115742 71270 115806 71334
rect 115742 71134 115806 71198
rect 116014 71270 116078 71334
rect 116286 71270 116350 71334
rect 116286 71134 116350 71198
rect 116830 71270 116894 71334
rect 116830 71134 116894 71198
rect 1230 70998 1294 71062
rect 21766 70862 21830 70926
rect 21902 70726 21966 70790
rect 22174 70862 22238 70926
rect 22582 70862 22646 70926
rect 22718 70726 22782 70790
rect 22990 70862 23054 70926
rect 23126 70726 23190 70790
rect 23534 70862 23598 70926
rect 137502 70998 137566 71062
rect 23398 70726 23462 70790
rect 21902 70454 21966 70518
rect 21902 70318 21966 70382
rect 22718 70454 22782 70518
rect 22446 70318 22510 70382
rect 23126 70454 23190 70518
rect 23126 70318 23190 70382
rect 23398 70454 23462 70518
rect 23534 70318 23598 70382
rect 24214 70318 24278 70382
rect 115334 70862 115398 70926
rect 115198 70726 115262 70790
rect 115742 70862 115806 70926
rect 115606 70726 115670 70790
rect 116286 70862 116350 70926
rect 116558 70726 116622 70790
rect 116830 70862 116894 70926
rect 116966 70726 117030 70790
rect 113294 70318 113358 70382
rect 115198 70454 115262 70518
rect 115198 70318 115262 70382
rect 115606 70454 115670 70518
rect 115742 70318 115806 70382
rect 116558 70454 116622 70518
rect 116150 70318 116214 70382
rect 116966 70454 117030 70518
rect 116966 70318 117030 70382
rect 21902 70046 21966 70110
rect 22446 70046 22510 70110
rect 22174 69910 22238 69974
rect 22582 69910 22646 69974
rect 23126 70046 23190 70110
rect 23534 70046 23598 70110
rect 24214 70046 24278 70110
rect 115198 70046 115262 70110
rect 115742 70046 115806 70110
rect 22990 69910 23054 69974
rect 23398 69910 23462 69974
rect 115198 69910 115262 69974
rect 115606 69910 115670 69974
rect 116150 70046 116214 70110
rect 116014 69910 116078 69974
rect 116558 69910 116622 69974
rect 116966 70046 117030 70110
rect 21902 69502 21966 69566
rect 22174 69638 22238 69702
rect 22582 69638 22646 69702
rect 22446 69502 22510 69566
rect 22990 69638 23054 69702
rect 22990 69502 23054 69566
rect 23398 69638 23462 69702
rect 23398 69502 23462 69566
rect 113294 69638 113358 69702
rect 115198 69638 115262 69702
rect 115198 69502 115262 69566
rect 115606 69638 115670 69702
rect 115606 69502 115670 69566
rect 116014 69638 116078 69702
rect 116150 69502 116214 69566
rect 116558 69638 116622 69702
rect 116830 69502 116894 69566
rect 1230 69230 1294 69294
rect 21902 69230 21966 69294
rect 22446 69230 22510 69294
rect 22582 69094 22646 69158
rect 22990 69230 23054 69294
rect 23126 69094 23190 69158
rect 23398 69230 23462 69294
rect 23534 69094 23598 69158
rect 115198 69230 115262 69294
rect 28294 68958 28358 69022
rect 115334 69094 115398 69158
rect 115606 69230 115670 69294
rect 115742 69094 115806 69158
rect 116150 69230 116214 69294
rect 116286 69094 116350 69158
rect 116830 69230 116894 69294
rect 137502 69230 137566 69294
rect 110438 68958 110502 69022
rect 21902 68822 21966 68886
rect 22582 68822 22646 68886
rect 23126 68822 23190 68886
rect 23126 68686 23190 68750
rect 23534 68822 23598 68886
rect 23398 68686 23462 68750
rect 28294 68686 28358 68750
rect 28430 68686 28494 68750
rect 21902 68550 21966 68614
rect 22174 68278 22238 68342
rect 22582 68278 22646 68342
rect 23126 68414 23190 68478
rect 21766 68006 21830 68070
rect 22174 68006 22238 68070
rect 22582 68006 22646 68070
rect 23398 68414 23462 68478
rect 110438 68686 110502 68750
rect 115334 68822 115398 68886
rect 115334 68686 115398 68750
rect 115742 68822 115806 68886
rect 115742 68686 115806 68750
rect 116286 68822 116350 68886
rect 116966 68822 117030 68886
rect 28430 68278 28494 68342
rect 21766 67734 21830 67798
rect 1230 67598 1294 67662
rect 21766 67598 21830 67662
rect 22582 67598 22646 67662
rect 110438 68142 110502 68206
rect 110438 67870 110502 67934
rect 115334 68414 115398 68478
rect 115742 68414 115806 68478
rect 116014 68278 116078 68342
rect 116966 68550 117030 68614
rect 116014 68006 116078 68070
rect 116830 68006 116894 68070
rect 116558 67598 116622 67662
rect 116830 67734 116894 67798
rect 116830 67598 116894 67662
rect 137502 67462 137566 67526
rect 21766 67326 21830 67390
rect 21902 67190 21966 67254
rect 22582 67326 22646 67390
rect 22990 67190 23054 67254
rect 23534 67190 23598 67254
rect 110302 67326 110366 67390
rect 115198 67190 115262 67254
rect 115606 67190 115670 67254
rect 116558 67326 116622 67390
rect 21902 66918 21966 66982
rect 21766 66782 21830 66846
rect 22582 66782 22646 66846
rect 22990 66918 23054 66982
rect 22990 66782 23054 66846
rect 23534 66918 23598 66982
rect 110302 67054 110366 67118
rect 116830 67326 116894 67390
rect 116966 67190 117030 67254
rect 23534 66782 23598 66846
rect 115198 66918 115262 66982
rect 115334 66782 115398 66846
rect 115606 66918 115670 66982
rect 115742 66782 115806 66846
rect 116286 66782 116350 66846
rect 116966 66918 117030 66982
rect 116830 66782 116894 66846
rect 21766 66510 21830 66574
rect 21902 66374 21966 66438
rect 22582 66510 22646 66574
rect 22446 66374 22510 66438
rect 22990 66510 23054 66574
rect 23126 66374 23190 66438
rect 23534 66510 23598 66574
rect 23398 66374 23462 66438
rect 115334 66510 115398 66574
rect 115198 66374 115262 66438
rect 115742 66510 115806 66574
rect 115606 66374 115670 66438
rect 116286 66510 116350 66574
rect 116558 66374 116622 66438
rect 116830 66510 116894 66574
rect 116966 66374 117030 66438
rect 21902 66102 21966 66166
rect 21766 65966 21830 66030
rect 22446 66102 22510 66166
rect 22310 65966 22374 66030
rect 23126 66102 23190 66166
rect 23126 65966 23190 66030
rect 23398 66102 23462 66166
rect 115198 66102 115262 66166
rect 23534 65966 23598 66030
rect 1230 65830 1294 65894
rect 115198 65966 115262 66030
rect 115606 66102 115670 66166
rect 115606 65966 115670 66030
rect 116558 66102 116622 66166
rect 116150 65966 116214 66030
rect 116422 65966 116486 66030
rect 116966 66102 117030 66166
rect 116830 65966 116894 66030
rect 137502 65966 137566 66030
rect 21766 65694 21830 65758
rect 21902 65558 21966 65622
rect 22310 65694 22374 65758
rect 22582 65558 22646 65622
rect 23126 65694 23190 65758
rect 22990 65558 23054 65622
rect 23534 65694 23598 65758
rect 23534 65558 23598 65622
rect 115198 65694 115262 65758
rect 115198 65558 115262 65622
rect 115606 65694 115670 65758
rect 115606 65558 115670 65622
rect 116150 65694 116214 65758
rect 116014 65558 116078 65622
rect 116422 65694 116486 65758
rect 116830 65694 116894 65758
rect 116830 65558 116894 65622
rect 21902 65286 21966 65350
rect 22582 65286 22646 65350
rect 22310 65150 22374 65214
rect 22446 65150 22510 65214
rect 22990 65286 23054 65350
rect 23126 65150 23190 65214
rect 23534 65286 23598 65350
rect 115198 65286 115262 65350
rect 23398 65150 23462 65214
rect 115198 65150 115262 65214
rect 115606 65286 115670 65350
rect 115606 65150 115670 65214
rect 116014 65286 116078 65350
rect 116150 65150 116214 65214
rect 116830 65286 116894 65350
rect 22310 64878 22374 64942
rect 22446 64878 22510 64942
rect 23126 64878 23190 64942
rect 22990 64742 23054 64806
rect 23398 64878 23462 64942
rect 23534 64742 23598 64806
rect 1230 64334 1294 64398
rect 22174 64334 22238 64398
rect 22582 64334 22646 64398
rect 22990 64470 23054 64534
rect 23534 64470 23598 64534
rect 115198 64878 115262 64942
rect 115334 64742 115398 64806
rect 115606 64878 115670 64942
rect 115742 64742 115806 64806
rect 116150 64878 116214 64942
rect 21902 64062 21966 64126
rect 22174 64062 22238 64126
rect 22582 64062 22646 64126
rect 21902 63790 21966 63854
rect 21766 63654 21830 63718
rect 22310 63654 22374 63718
rect 28566 63790 28630 63854
rect 115334 64470 115398 64534
rect 115742 64470 115806 64534
rect 116014 64334 116078 64398
rect 116558 64334 116622 64398
rect 110166 64198 110230 64262
rect 110166 63926 110230 63990
rect 110438 63790 110502 63854
rect 116014 64062 116078 64126
rect 116558 64062 116622 64126
rect 116830 64062 116894 64126
rect 137502 64198 137566 64262
rect 21766 63382 21830 63446
rect 21902 63246 21966 63310
rect 22310 63382 22374 63446
rect 23126 63246 23190 63310
rect 23398 63246 23462 63310
rect 28566 63518 28630 63582
rect 28294 63382 28358 63446
rect 110438 63518 110502 63582
rect 116286 63654 116350 63718
rect 116830 63790 116894 63854
rect 116830 63654 116894 63718
rect 115198 63246 115262 63310
rect 115606 63246 115670 63310
rect 116286 63382 116350 63446
rect 116830 63382 116894 63446
rect 116966 63246 117030 63310
rect 28294 63110 28358 63174
rect 21902 62974 21966 63038
rect 21766 62838 21830 62902
rect 23126 62974 23190 63038
rect 22582 62838 22646 62902
rect 22990 62838 23054 62902
rect 23398 62974 23462 63038
rect 115198 62974 115262 63038
rect 23398 62838 23462 62902
rect 1230 62566 1294 62630
rect 21766 62566 21830 62630
rect 21766 62430 21830 62494
rect 22174 62430 22238 62494
rect 22582 62566 22646 62630
rect 22990 62566 23054 62630
rect 22990 62430 23054 62494
rect 23398 62566 23462 62630
rect 23534 62430 23598 62494
rect 115198 62838 115262 62902
rect 115606 62974 115670 63038
rect 115606 62838 115670 62902
rect 116150 62838 116214 62902
rect 116286 62838 116350 62902
rect 116966 62974 117030 63038
rect 116966 62838 117030 62902
rect 110166 62566 110230 62630
rect 115198 62566 115262 62630
rect 115334 62430 115398 62494
rect 115606 62566 115670 62630
rect 115742 62430 115806 62494
rect 116150 62566 116214 62630
rect 116286 62566 116350 62630
rect 116422 62430 116486 62494
rect 116966 62566 117030 62630
rect 116830 62430 116894 62494
rect 137502 62566 137566 62630
rect 21766 62158 21830 62222
rect 21902 62022 21966 62086
rect 22174 62158 22238 62222
rect 22446 62022 22510 62086
rect 22990 62158 23054 62222
rect 22990 62022 23054 62086
rect 23534 62158 23598 62222
rect 110166 62294 110230 62358
rect 23398 62022 23462 62086
rect 21902 61750 21966 61814
rect 21902 61614 21966 61678
rect 22446 61750 22510 61814
rect 22310 61614 22374 61678
rect 22446 61614 22510 61678
rect 22990 61750 23054 61814
rect 22990 61614 23054 61678
rect 23398 61750 23462 61814
rect 23534 61614 23598 61678
rect 115334 62158 115398 62222
rect 115198 62022 115262 62086
rect 115742 62158 115806 62222
rect 115606 62022 115670 62086
rect 116422 62158 116486 62222
rect 116558 62022 116622 62086
rect 116830 62158 116894 62222
rect 116966 62022 117030 62086
rect 115198 61750 115262 61814
rect 115334 61614 115398 61678
rect 115606 61750 115670 61814
rect 115742 61614 115806 61678
rect 116558 61750 116622 61814
rect 116150 61614 116214 61678
rect 116966 61750 117030 61814
rect 116830 61614 116894 61678
rect 21902 61342 21966 61406
rect 22310 61342 22374 61406
rect 22446 61342 22510 61406
rect 22718 61206 22782 61270
rect 22990 61342 23054 61406
rect 22990 61206 23054 61270
rect 23534 61342 23598 61406
rect 23534 61206 23598 61270
rect 1230 60934 1294 60998
rect 115334 61342 115398 61406
rect 115198 61206 115262 61270
rect 115742 61342 115806 61406
rect 115742 61206 115806 61270
rect 116150 61342 116214 61406
rect 116014 61206 116078 61270
rect 116558 61206 116622 61270
rect 116830 61342 116894 61406
rect 110438 61070 110502 61134
rect 22446 60934 22510 60998
rect 22718 60934 22782 60998
rect 22990 60934 23054 60998
rect 23126 60798 23190 60862
rect 23534 60934 23598 60998
rect 23398 60798 23462 60862
rect 22446 60662 22510 60726
rect 22174 60390 22238 60454
rect 23126 60526 23190 60590
rect 23126 60390 23190 60454
rect 23398 60526 23462 60590
rect 23534 60390 23598 60454
rect 110438 60798 110502 60862
rect 115198 60934 115262 60998
rect 115198 60798 115262 60862
rect 115742 60934 115806 60998
rect 115606 60798 115670 60862
rect 116014 60934 116078 60998
rect 116558 60934 116622 60998
rect 137502 60934 137566 60998
rect 115198 60526 115262 60590
rect 28566 60254 28630 60318
rect 115334 60390 115398 60454
rect 115606 60526 115670 60590
rect 115742 60390 115806 60454
rect 116014 60390 116078 60454
rect 116422 60390 116486 60454
rect 21902 60118 21966 60182
rect 22174 60118 22238 60182
rect 23126 60118 23190 60182
rect 23534 60118 23598 60182
rect 21902 59846 21966 59910
rect 21902 59710 21966 59774
rect 22310 59710 22374 59774
rect 28294 59982 28358 60046
rect 28566 59982 28630 60046
rect 115334 60118 115398 60182
rect 115742 60118 115806 60182
rect 110166 59846 110230 59910
rect 28294 59574 28358 59638
rect 21902 59438 21966 59502
rect 21766 59302 21830 59366
rect 22310 59438 22374 59502
rect 1230 59166 1294 59230
rect 22990 59302 23054 59366
rect 23534 59302 23598 59366
rect 110166 59574 110230 59638
rect 110438 59438 110502 59502
rect 116014 60118 116078 60182
rect 116422 60118 116486 60182
rect 116830 60118 116894 60182
rect 116558 59710 116622 59774
rect 116830 59846 116894 59910
rect 116966 59710 117030 59774
rect 115334 59302 115398 59366
rect 115742 59302 115806 59366
rect 21766 59030 21830 59094
rect 21902 58894 21966 58958
rect 22310 58894 22374 58958
rect 22990 59030 23054 59094
rect 22990 58894 23054 58958
rect 23534 59030 23598 59094
rect 23398 58894 23462 58958
rect 110438 59166 110502 59230
rect 115334 59030 115398 59094
rect 21902 58622 21966 58686
rect 21902 58486 21966 58550
rect 22310 58622 22374 58686
rect 22174 58486 22238 58550
rect 22718 58486 22782 58550
rect 22990 58622 23054 58686
rect 22990 58486 23054 58550
rect 23398 58622 23462 58686
rect 23398 58486 23462 58550
rect 28566 58622 28630 58686
rect 115198 58894 115262 58958
rect 115742 59030 115806 59094
rect 115742 58894 115806 58958
rect 116150 58894 116214 58958
rect 116558 59438 116622 59502
rect 116966 59438 117030 59502
rect 116830 59302 116894 59366
rect 116558 58894 116622 58958
rect 116830 59030 116894 59094
rect 137502 59030 137566 59094
rect 116830 58894 116894 58958
rect 110438 58622 110502 58686
rect 115198 58622 115262 58686
rect 115198 58486 115262 58550
rect 115742 58622 115806 58686
rect 115742 58486 115806 58550
rect 116150 58622 116214 58686
rect 116558 58622 116622 58686
rect 116014 58486 116078 58550
rect 116830 58622 116894 58686
rect 116830 58486 116894 58550
rect 28566 58350 28630 58414
rect 21902 58214 21966 58278
rect 21766 58078 21830 58142
rect 22174 58214 22238 58278
rect 22718 58214 22782 58278
rect 22446 58078 22510 58142
rect 22990 58214 23054 58278
rect 22990 58078 23054 58142
rect 23398 58214 23462 58278
rect 23534 58078 23598 58142
rect 110438 58350 110502 58414
rect 115198 58214 115262 58278
rect 115198 58078 115262 58142
rect 115742 58214 115806 58278
rect 115742 58078 115806 58142
rect 116014 58214 116078 58278
rect 116830 58214 116894 58278
rect 116830 58078 116894 58142
rect 21766 57806 21830 57870
rect 21902 57670 21966 57734
rect 22446 57806 22510 57870
rect 22718 57670 22782 57734
rect 22990 57806 23054 57870
rect 23126 57670 23190 57734
rect 23534 57806 23598 57870
rect 23398 57670 23462 57734
rect 115198 57806 115262 57870
rect 115198 57670 115262 57734
rect 115742 57806 115806 57870
rect 115606 57670 115670 57734
rect 116558 57670 116622 57734
rect 116830 57806 116894 57870
rect 116966 57670 117030 57734
rect 1230 57398 1294 57462
rect 21902 57398 21966 57462
rect 22718 57398 22782 57462
rect 23126 57398 23190 57462
rect 23126 57262 23190 57326
rect 23398 57398 23462 57462
rect 115198 57398 115262 57462
rect 23534 57262 23598 57326
rect 115334 57262 115398 57326
rect 115606 57398 115670 57462
rect 115742 57262 115806 57326
rect 116558 57398 116622 57462
rect 116150 57262 116214 57326
rect 116286 57262 116350 57326
rect 116966 57398 117030 57462
rect 137502 57398 137566 57462
rect 22446 56854 22510 56918
rect 23126 56990 23190 57054
rect 22990 56854 23054 56918
rect 23534 56990 23598 57054
rect 23534 56854 23598 56918
rect 115334 56990 115398 57054
rect 115198 56854 115262 56918
rect 115742 56990 115806 57054
rect 115606 56854 115670 56918
rect 116150 56990 116214 57054
rect 116286 56990 116350 57054
rect 22446 56582 22510 56646
rect 22446 56446 22510 56510
rect 22718 56446 22782 56510
rect 22990 56582 23054 56646
rect 22990 56446 23054 56510
rect 23534 56582 23598 56646
rect 23398 56446 23462 56510
rect 115198 56582 115262 56646
rect 115198 56446 115262 56510
rect 115606 56582 115670 56646
rect 115606 56446 115670 56510
rect 116558 56446 116622 56510
rect 110438 56310 110502 56374
rect 21902 56174 21966 56238
rect 22446 56174 22510 56238
rect 22718 56174 22782 56238
rect 22990 56174 23054 56238
rect 23398 56174 23462 56238
rect 1230 55766 1294 55830
rect 21902 55902 21966 55966
rect 21766 55766 21830 55830
rect 22582 55766 22646 55830
rect 28566 55902 28630 55966
rect 110438 56038 110502 56102
rect 115198 56174 115262 56238
rect 115606 56174 115670 56238
rect 110438 55902 110502 55966
rect 21766 55494 21830 55558
rect 21902 55358 21966 55422
rect 22582 55494 22646 55558
rect 21902 55086 21966 55150
rect 21766 54950 21830 55014
rect 22174 54950 22238 55014
rect 22990 54950 23054 55014
rect 28566 55630 28630 55694
rect 28566 55494 28630 55558
rect 28566 55222 28630 55286
rect 110438 55630 110502 55694
rect 110438 55494 110502 55558
rect 110438 55222 110502 55286
rect 23534 54950 23598 55014
rect 21766 54678 21830 54742
rect 21902 54542 21966 54606
rect 22174 54678 22238 54742
rect 22310 54542 22374 54606
rect 22446 54542 22510 54606
rect 22990 54678 23054 54742
rect 22990 54542 23054 54606
rect 23534 54678 23598 54742
rect 23534 54542 23598 54606
rect 28294 54678 28358 54742
rect 116558 56174 116622 56238
rect 116966 56174 117030 56238
rect 116558 55766 116622 55830
rect 116966 55902 117030 55966
rect 116966 55766 117030 55830
rect 137502 55766 137566 55830
rect 116558 55494 116622 55558
rect 116966 55494 117030 55558
rect 116966 55358 117030 55422
rect 115198 54950 115262 55014
rect 115742 54950 115806 55014
rect 116286 54950 116350 55014
rect 116966 55086 117030 55150
rect 116830 54950 116894 55014
rect 115198 54678 115262 54742
rect 115334 54542 115398 54606
rect 115742 54678 115806 54742
rect 115742 54542 115806 54606
rect 116286 54678 116350 54742
rect 116150 54542 116214 54606
rect 116286 54542 116350 54606
rect 116830 54678 116894 54742
rect 116830 54542 116894 54606
rect 28294 54406 28358 54470
rect 21902 54270 21966 54334
rect 1230 54134 1294 54198
rect 21902 54134 21966 54198
rect 22310 54270 22374 54334
rect 22446 54270 22510 54334
rect 22174 54134 22238 54198
rect 22990 54270 23054 54334
rect 22990 54134 23054 54198
rect 23534 54270 23598 54334
rect 115334 54270 115398 54334
rect 23398 54134 23462 54198
rect 115334 54134 115398 54198
rect 115742 54270 115806 54334
rect 115606 54134 115670 54198
rect 116150 54270 116214 54334
rect 116286 54270 116350 54334
rect 116014 54134 116078 54198
rect 116422 54134 116486 54198
rect 116830 54270 116894 54334
rect 116830 54134 116894 54198
rect 137502 54134 137566 54198
rect 21902 53862 21966 53926
rect 21766 53726 21830 53790
rect 22174 53862 22238 53926
rect 22174 53726 22238 53790
rect 22582 53726 22646 53790
rect 22990 53862 23054 53926
rect 23126 53726 23190 53790
rect 23398 53862 23462 53926
rect 23534 53726 23598 53790
rect 115334 53862 115398 53926
rect 115334 53726 115398 53790
rect 115606 53862 115670 53926
rect 115742 53726 115806 53790
rect 116014 53862 116078 53926
rect 116422 53862 116486 53926
rect 116286 53726 116350 53790
rect 116830 53862 116894 53926
rect 116830 53726 116894 53790
rect 21766 53454 21830 53518
rect 22174 53454 22238 53518
rect 22582 53454 22646 53518
rect 22718 53318 22782 53382
rect 23126 53454 23190 53518
rect 22990 53318 23054 53382
rect 23534 53454 23598 53518
rect 23398 53318 23462 53382
rect 21766 52910 21830 52974
rect 22718 53046 22782 53110
rect 22446 52910 22510 52974
rect 22990 53046 23054 53110
rect 23126 52910 23190 52974
rect 23398 53046 23462 53110
rect 23534 52910 23598 52974
rect 115334 53454 115398 53518
rect 115198 53318 115262 53382
rect 115742 53454 115806 53518
rect 115606 53318 115670 53382
rect 116286 53454 116350 53518
rect 116558 53318 116622 53382
rect 116830 53454 116894 53518
rect 115198 53046 115262 53110
rect 115334 52910 115398 52974
rect 115606 53046 115670 53110
rect 115742 52910 115806 52974
rect 116558 53046 116622 53110
rect 116150 52910 116214 52974
rect 116286 52910 116350 52974
rect 116422 52910 116486 52974
rect 116830 52910 116894 52974
rect 21766 52638 21830 52702
rect 1230 52502 1294 52566
rect 22446 52638 22510 52702
rect 22174 52502 22238 52566
rect 22718 52502 22782 52566
rect 23126 52638 23190 52702
rect 22990 52502 23054 52566
rect 23534 52638 23598 52702
rect 23398 52502 23462 52566
rect 115334 52638 115398 52702
rect 115334 52502 115398 52566
rect 115742 52638 115806 52702
rect 115742 52502 115806 52566
rect 116150 52638 116214 52702
rect 116286 52638 116350 52702
rect 116422 52638 116486 52702
rect 116014 52502 116078 52566
rect 116286 52502 116350 52566
rect 116830 52638 116894 52702
rect 137502 52502 137566 52566
rect 110438 52366 110502 52430
rect 21902 52230 21966 52294
rect 22174 52230 22238 52294
rect 22718 52230 22782 52294
rect 22990 52230 23054 52294
rect 22990 52094 23054 52158
rect 23398 52230 23462 52294
rect 23398 52094 23462 52158
rect 21902 51958 21966 52022
rect 22174 51686 22238 51750
rect 22990 51822 23054 51886
rect 23398 51822 23462 51886
rect 21766 51414 21830 51478
rect 22174 51414 22238 51478
rect 28430 51822 28494 51886
rect 110438 52094 110502 52158
rect 115334 52230 115398 52294
rect 115198 52094 115262 52158
rect 115742 52230 115806 52294
rect 115606 52094 115670 52158
rect 116014 52230 116078 52294
rect 116286 52230 116350 52294
rect 116966 52230 117030 52294
rect 115198 51822 115262 51886
rect 28430 51550 28494 51614
rect 28566 51550 28630 51614
rect 28566 51278 28630 51342
rect 21766 51142 21830 51206
rect 21902 51006 21966 51070
rect 22310 51006 22374 51070
rect 22446 51006 22510 51070
rect 22990 51006 23054 51070
rect 23398 51006 23462 51070
rect 1230 50870 1294 50934
rect 21902 50734 21966 50798
rect 21766 50598 21830 50662
rect 22310 50734 22374 50798
rect 22446 50734 22510 50798
rect 22174 50598 22238 50662
rect 22582 50598 22646 50662
rect 22990 50734 23054 50798
rect 22990 50598 23054 50662
rect 23398 50734 23462 50798
rect 23534 50598 23598 50662
rect 115606 51822 115670 51886
rect 116014 51686 116078 51750
rect 116422 51686 116486 51750
rect 116966 51958 117030 52022
rect 115198 51006 115262 51070
rect 116014 51414 116078 51478
rect 116422 51414 116486 51478
rect 115606 51006 115670 51070
rect 116830 51414 116894 51478
rect 116558 51006 116622 51070
rect 116830 51142 116894 51206
rect 116830 51006 116894 51070
rect 137502 50870 137566 50934
rect 110438 50734 110502 50798
rect 115198 50734 115262 50798
rect 115334 50598 115398 50662
rect 115606 50734 115670 50798
rect 115742 50598 115806 50662
rect 116014 50598 116078 50662
rect 116558 50734 116622 50798
rect 116422 50598 116486 50662
rect 116830 50734 116894 50798
rect 116830 50598 116894 50662
rect 21766 50326 21830 50390
rect 21902 50190 21966 50254
rect 22174 50326 22238 50390
rect 22582 50326 22646 50390
rect 22446 50190 22510 50254
rect 22990 50326 23054 50390
rect 23126 50190 23190 50254
rect 23534 50326 23598 50390
rect 23534 50190 23598 50254
rect 110438 50462 110502 50526
rect 115334 50326 115398 50390
rect 115334 50190 115398 50254
rect 115742 50326 115806 50390
rect 115606 50190 115670 50254
rect 116014 50326 116078 50390
rect 116422 50326 116486 50390
rect 116150 50190 116214 50254
rect 116286 50190 116350 50254
rect 116830 50326 116894 50390
rect 116966 50190 117030 50254
rect 21902 49918 21966 49982
rect 21902 49782 21966 49846
rect 22446 49918 22510 49982
rect 22174 49782 22238 49846
rect 22582 49782 22646 49846
rect 23126 49918 23190 49982
rect 22990 49782 23054 49846
rect 23534 49918 23598 49982
rect 23534 49782 23598 49846
rect 115334 49918 115398 49982
rect 115334 49782 115398 49846
rect 115606 49918 115670 49982
rect 115742 49782 115806 49846
rect 116150 49918 116214 49982
rect 116286 49918 116350 49982
rect 116014 49782 116078 49846
rect 116966 49918 117030 49982
rect 116966 49782 117030 49846
rect 21902 49510 21966 49574
rect 21766 49374 21830 49438
rect 22174 49510 22238 49574
rect 22582 49510 22646 49574
rect 22582 49374 22646 49438
rect 22990 49510 23054 49574
rect 22990 49374 23054 49438
rect 23534 49510 23598 49574
rect 23534 49374 23598 49438
rect 115334 49510 115398 49574
rect 115334 49374 115398 49438
rect 115742 49510 115806 49574
rect 115742 49374 115806 49438
rect 116014 49510 116078 49574
rect 116422 49374 116486 49438
rect 116966 49510 117030 49574
rect 116830 49374 116894 49438
rect 1230 49102 1294 49166
rect 21766 49102 21830 49166
rect 21902 48966 21966 49030
rect 22582 49102 22646 49166
rect 22718 48966 22782 49030
rect 22990 49102 23054 49166
rect 23126 48966 23190 49030
rect 23534 49102 23598 49166
rect 23398 48966 23462 49030
rect 115334 49102 115398 49166
rect 115198 48966 115262 49030
rect 115742 49102 115806 49166
rect 115606 48966 115670 49030
rect 116422 49102 116486 49166
rect 116558 48966 116622 49030
rect 116830 49102 116894 49166
rect 116966 48966 117030 49030
rect 137502 48966 137566 49030
rect 21902 48694 21966 48758
rect 22718 48694 22782 48758
rect 22310 48558 22374 48622
rect 23126 48694 23190 48758
rect 23126 48558 23190 48622
rect 23398 48694 23462 48758
rect 23398 48558 23462 48622
rect 115198 48694 115262 48758
rect 115334 48558 115398 48622
rect 115606 48694 115670 48758
rect 115742 48558 115806 48622
rect 116558 48694 116622 48758
rect 116150 48558 116214 48622
rect 116286 48558 116350 48622
rect 116966 48694 117030 48758
rect 21766 48286 21830 48350
rect 22310 48286 22374 48350
rect 21766 48014 21830 48078
rect 23126 48286 23190 48350
rect 22990 48150 23054 48214
rect 23398 48286 23462 48350
rect 23398 48150 23462 48214
rect 22718 47742 22782 47806
rect 22990 47878 23054 47942
rect 23398 47878 23462 47942
rect 115334 48286 115398 48350
rect 115198 48150 115262 48214
rect 115742 48286 115806 48350
rect 115742 48150 115806 48214
rect 116150 48286 116214 48350
rect 116286 48286 116350 48350
rect 116830 48286 116894 48350
rect 116150 48150 116214 48214
rect 115198 47878 115262 47942
rect 21766 47470 21830 47534
rect 1230 47334 1294 47398
rect 22718 47470 22782 47534
rect 21766 47198 21830 47262
rect 21766 47062 21830 47126
rect 22446 47062 22510 47126
rect 28294 47198 28358 47262
rect 110166 47606 110230 47670
rect 110166 47334 110230 47398
rect 115742 47878 115806 47942
rect 116286 48014 116350 48078
rect 116558 47742 116622 47806
rect 116830 48014 116894 48078
rect 110302 47198 110366 47262
rect 21766 46790 21830 46854
rect 21902 46654 21966 46718
rect 22446 46790 22510 46854
rect 22990 46654 23054 46718
rect 23398 46654 23462 46718
rect 28294 46926 28358 46990
rect 110302 46926 110366 46990
rect 110438 46790 110502 46854
rect 116558 47470 116622 47534
rect 116966 47470 117030 47534
rect 137502 47470 137566 47534
rect 116150 47062 116214 47126
rect 116286 47062 116350 47126
rect 116966 47198 117030 47262
rect 116830 47062 116894 47126
rect 115198 46654 115262 46718
rect 115606 46654 115670 46718
rect 116150 46790 116214 46854
rect 116286 46790 116350 46854
rect 21902 46382 21966 46446
rect 21766 46246 21830 46310
rect 22174 46246 22238 46310
rect 22990 46382 23054 46446
rect 23126 46246 23190 46310
rect 23398 46382 23462 46446
rect 28294 46382 28358 46446
rect 110438 46518 110502 46582
rect 116830 46790 116894 46854
rect 116830 46654 116894 46718
rect 115198 46382 115262 46446
rect 23534 46246 23598 46310
rect 115334 46246 115398 46310
rect 115606 46382 115670 46446
rect 115742 46246 115806 46310
rect 116014 46246 116078 46310
rect 116830 46382 116894 46446
rect 116830 46246 116894 46310
rect 21766 45974 21830 46038
rect 21902 45838 21966 45902
rect 22174 45974 22238 46038
rect 22310 45838 22374 45902
rect 23126 45974 23190 46038
rect 23126 45838 23190 45902
rect 23534 45974 23598 46038
rect 23398 45838 23462 45902
rect 28294 45974 28358 46038
rect 115334 45974 115398 46038
rect 115198 45838 115262 45902
rect 115742 45974 115806 46038
rect 115606 45838 115670 45902
rect 116014 45974 116078 46038
rect 116422 45838 116486 45902
rect 116830 45974 116894 46038
rect 116966 45838 117030 45902
rect 1230 45566 1294 45630
rect 21902 45566 21966 45630
rect 21902 45430 21966 45494
rect 22310 45566 22374 45630
rect 22582 45430 22646 45494
rect 23126 45566 23190 45630
rect 22990 45430 23054 45494
rect 23398 45566 23462 45630
rect 115198 45566 115262 45630
rect 23398 45430 23462 45494
rect 115334 45430 115398 45494
rect 115606 45566 115670 45630
rect 115742 45430 115806 45494
rect 116422 45566 116486 45630
rect 116150 45430 116214 45494
rect 116286 45430 116350 45494
rect 116966 45566 117030 45630
rect 137502 45566 137566 45630
rect 116966 45430 117030 45494
rect 21902 45158 21966 45222
rect 21766 45022 21830 45086
rect 22174 45022 22238 45086
rect 22582 45158 22646 45222
rect 22582 45022 22646 45086
rect 22990 45158 23054 45222
rect 22990 45022 23054 45086
rect 23398 45158 23462 45222
rect 23534 45022 23598 45086
rect 115334 45158 115398 45222
rect 115334 45022 115398 45086
rect 115742 45158 115806 45222
rect 115742 45022 115806 45086
rect 116150 45158 116214 45222
rect 116286 45158 116350 45222
rect 116422 45022 116486 45086
rect 116966 45158 117030 45222
rect 116830 45022 116894 45086
rect 21766 44750 21830 44814
rect 22174 44750 22238 44814
rect 22310 44614 22374 44678
rect 22582 44750 22646 44814
rect 22718 44614 22782 44678
rect 22990 44750 23054 44814
rect 23126 44614 23190 44678
rect 23534 44750 23598 44814
rect 23398 44614 23462 44678
rect 22310 44342 22374 44406
rect 22718 44342 22782 44406
rect 23126 44342 23190 44406
rect 22990 44206 23054 44270
rect 23398 44342 23462 44406
rect 23398 44206 23462 44270
rect 1230 44070 1294 44134
rect 22174 43798 22238 43862
rect 22582 43798 22646 43862
rect 22990 43934 23054 43998
rect 22990 43798 23054 43862
rect 23398 43934 23462 43998
rect 23398 43798 23462 43862
rect 115334 44750 115398 44814
rect 115198 44614 115262 44678
rect 115742 44750 115806 44814
rect 115606 44614 115670 44678
rect 116422 44750 116486 44814
rect 116558 44614 116622 44678
rect 116830 44750 116894 44814
rect 110166 44478 110230 44542
rect 110166 44206 110230 44270
rect 115198 44342 115262 44406
rect 115198 44206 115262 44270
rect 115606 44342 115670 44406
rect 115606 44206 115670 44270
rect 116286 44342 116350 44406
rect 116558 44342 116622 44406
rect 115198 43934 115262 43998
rect 115198 43798 115262 43862
rect 115606 43934 115670 43998
rect 115606 43798 115670 43862
rect 116286 44070 116350 44134
rect 116014 43798 116078 43862
rect 116558 43798 116622 43862
rect 137502 44070 137566 44134
rect 110438 43662 110502 43726
rect 21902 43526 21966 43590
rect 22174 43526 22238 43590
rect 22446 43526 22510 43590
rect 22582 43526 22646 43590
rect 21902 43254 21966 43318
rect 21766 43118 21830 43182
rect 22582 43254 22646 43318
rect 22446 43118 22510 43182
rect 22990 43526 23054 43590
rect 23398 43526 23462 43590
rect 28294 43254 28358 43318
rect 110438 43390 110502 43454
rect 110166 43254 110230 43318
rect 115198 43526 115262 43590
rect 115606 43526 115670 43590
rect 116014 43526 116078 43590
rect 116558 43526 116622 43590
rect 116966 43526 117030 43590
rect 21766 42846 21830 42910
rect 21766 42710 21830 42774
rect 22446 42846 22510 42910
rect 23126 42710 23190 42774
rect 23398 42710 23462 42774
rect 28294 42982 28358 43046
rect 28294 42846 28358 42910
rect 110166 42982 110230 43046
rect 116966 43254 117030 43318
rect 116966 43118 117030 43182
rect 115334 42710 115398 42774
rect 115606 42710 115670 42774
rect 28294 42574 28358 42638
rect 1230 42438 1294 42502
rect 21766 42438 21830 42502
rect 21902 42302 21966 42366
rect 23126 42438 23190 42502
rect 23126 42302 23190 42366
rect 23398 42438 23462 42502
rect 116966 42846 117030 42910
rect 116966 42710 117030 42774
rect 115334 42438 115398 42502
rect 23398 42302 23462 42366
rect 21902 42030 21966 42094
rect 21766 41894 21830 41958
rect 22174 41894 22238 41958
rect 22446 41894 22510 41958
rect 23126 42030 23190 42094
rect 23126 41894 23190 41958
rect 23398 42030 23462 42094
rect 23534 41894 23598 41958
rect 115198 42302 115262 42366
rect 115606 42438 115670 42502
rect 115606 42302 115670 42366
rect 116150 42302 116214 42366
rect 116966 42438 117030 42502
rect 116966 42302 117030 42366
rect 137502 42438 137566 42502
rect 110438 42030 110502 42094
rect 115198 42030 115262 42094
rect 115334 41894 115398 41958
rect 115606 42030 115670 42094
rect 115742 41894 115806 41958
rect 116150 42030 116214 42094
rect 116014 41894 116078 41958
rect 116422 41894 116486 41958
rect 116966 42030 117030 42094
rect 116830 41894 116894 41958
rect 21766 41622 21830 41686
rect 21766 41486 21830 41550
rect 22174 41622 22238 41686
rect 22446 41622 22510 41686
rect 23126 41622 23190 41686
rect 23126 41486 23190 41550
rect 23534 41622 23598 41686
rect 23398 41486 23462 41550
rect 110438 41758 110502 41822
rect 115334 41622 115398 41686
rect 115198 41486 115262 41550
rect 115742 41622 115806 41686
rect 115606 41486 115670 41550
rect 116014 41622 116078 41686
rect 116422 41622 116486 41686
rect 116014 41486 116078 41550
rect 116286 41486 116350 41550
rect 116558 41486 116622 41550
rect 116830 41622 116894 41686
rect 116966 41486 117030 41550
rect 21766 41214 21830 41278
rect 21766 41078 21830 41142
rect 22174 41078 22238 41142
rect 22718 41078 22782 41142
rect 23126 41214 23190 41278
rect 22990 41078 23054 41142
rect 23398 41214 23462 41278
rect 23534 41078 23598 41142
rect 115198 41214 115262 41278
rect 115198 41078 115262 41142
rect 115606 41214 115670 41278
rect 115742 41078 115806 41142
rect 116014 41214 116078 41278
rect 116286 41214 116350 41278
rect 116558 41214 116622 41278
rect 116014 41078 116078 41142
rect 116966 41214 117030 41278
rect 116966 41078 117030 41142
rect 21766 40806 21830 40870
rect 1230 40670 1294 40734
rect 22174 40806 22238 40870
rect 22718 40806 22782 40870
rect 22582 40670 22646 40734
rect 22990 40806 23054 40870
rect 23126 40670 23190 40734
rect 23534 40806 23598 40870
rect 23534 40670 23598 40734
rect 14694 40534 14758 40598
rect 22582 40398 22646 40462
rect 23126 40398 23190 40462
rect 22990 40262 23054 40326
rect 23534 40398 23598 40462
rect 23398 40262 23462 40326
rect 22582 39854 22646 39918
rect 22990 39990 23054 40054
rect 23126 39854 23190 39918
rect 23398 39990 23462 40054
rect 115198 40806 115262 40870
rect 115198 40670 115262 40734
rect 115742 40806 115806 40870
rect 115742 40670 115806 40734
rect 116014 40806 116078 40870
rect 116014 40670 116078 40734
rect 116966 40806 117030 40870
rect 137502 40670 137566 40734
rect 110166 40534 110230 40598
rect 110166 40262 110230 40326
rect 115198 40398 115262 40462
rect 115198 40262 115262 40326
rect 115742 40398 115806 40462
rect 115606 40262 115670 40326
rect 116014 40398 116078 40462
rect 115198 39990 115262 40054
rect 23534 39854 23598 39918
rect 28430 39718 28494 39782
rect 115198 39854 115262 39918
rect 115606 39990 115670 40054
rect 115606 39854 115670 39918
rect 116422 39854 116486 39918
rect 21766 39582 21830 39646
rect 22582 39582 22646 39646
rect 23126 39582 23190 39646
rect 23534 39582 23598 39646
rect 14558 39174 14622 39238
rect 21766 39310 21830 39374
rect 21902 39174 21966 39238
rect 22310 39174 22374 39238
rect 22446 39174 22510 39238
rect 1230 39038 1294 39102
rect 28430 39446 28494 39510
rect 28294 39310 28358 39374
rect 115198 39582 115262 39646
rect 115606 39582 115670 39646
rect 116422 39582 116486 39646
rect 116830 39582 116894 39646
rect 110438 39310 110502 39374
rect 28294 39038 28358 39102
rect 21902 38902 21966 38966
rect 21902 38766 21966 38830
rect 22310 38902 22374 38966
rect 22446 38902 22510 38966
rect 21902 38494 21966 38558
rect 21902 38358 21966 38422
rect 22174 38358 22238 38422
rect 22718 38358 22782 38422
rect 22990 38358 23054 38422
rect 28294 38902 28358 38966
rect 28294 38630 28358 38694
rect 110438 39038 110502 39102
rect 110166 38630 110230 38694
rect 116558 39174 116622 39238
rect 116830 39310 116894 39374
rect 116966 39174 117030 39238
rect 23398 38358 23462 38422
rect 21902 38086 21966 38150
rect 21902 37950 21966 38014
rect 22174 38086 22238 38150
rect 22718 38086 22782 38150
rect 22990 38086 23054 38150
rect 22990 37950 23054 38014
rect 23398 38086 23462 38150
rect 23398 37950 23462 38014
rect 110166 38358 110230 38422
rect 115334 38358 115398 38422
rect 115742 38358 115806 38422
rect 116558 38902 116622 38966
rect 116966 38902 117030 38966
rect 137502 38902 137566 38966
rect 116966 38766 117030 38830
rect 116014 38358 116078 38422
rect 116966 38494 117030 38558
rect 116830 38358 116894 38422
rect 115334 38086 115398 38150
rect 115198 37950 115262 38014
rect 115742 38086 115806 38150
rect 115606 37950 115670 38014
rect 116014 38086 116078 38150
rect 116014 37950 116078 38014
rect 116830 38086 116894 38150
rect 116966 37950 117030 38014
rect 14694 37814 14758 37878
rect 14830 37678 14894 37742
rect 21902 37678 21966 37742
rect 21766 37542 21830 37606
rect 22174 37542 22238 37606
rect 22446 37542 22510 37606
rect 22990 37678 23054 37742
rect 23126 37542 23190 37606
rect 23398 37678 23462 37742
rect 115198 37678 115262 37742
rect 23534 37542 23598 37606
rect 1230 37406 1294 37470
rect 115334 37542 115398 37606
rect 115606 37678 115670 37742
rect 115742 37542 115806 37606
rect 116014 37678 116078 37742
rect 116150 37542 116214 37606
rect 116286 37542 116350 37606
rect 116966 37678 117030 37742
rect 116830 37542 116894 37606
rect 21766 37270 21830 37334
rect 21902 37134 21966 37198
rect 22174 37270 22238 37334
rect 22446 37270 22510 37334
rect 23126 37270 23190 37334
rect 22990 37134 23054 37198
rect 23534 37270 23598 37334
rect 23398 37134 23462 37198
rect 115334 37270 115398 37334
rect 115334 37134 115398 37198
rect 115742 37270 115806 37334
rect 115606 37134 115670 37198
rect 116150 37270 116214 37334
rect 116286 37270 116350 37334
rect 116150 37134 116214 37198
rect 116286 37134 116350 37198
rect 116558 37134 116622 37198
rect 116830 37270 116894 37334
rect 137502 37270 137566 37334
rect 116830 37134 116894 37198
rect 21902 36862 21966 36926
rect 22174 36726 22238 36790
rect 22718 36726 22782 36790
rect 22990 36862 23054 36926
rect 22990 36726 23054 36790
rect 23398 36862 23462 36926
rect 23398 36726 23462 36790
rect 14558 36454 14622 36518
rect 14694 36318 14758 36382
rect 115334 36862 115398 36926
rect 115198 36726 115262 36790
rect 115606 36862 115670 36926
rect 115606 36726 115670 36790
rect 116150 36862 116214 36926
rect 116286 36862 116350 36926
rect 116558 36862 116622 36926
rect 116014 36726 116078 36790
rect 116286 36726 116350 36790
rect 116830 36862 116894 36926
rect 21902 36318 21966 36382
rect 22174 36454 22238 36518
rect 22174 36318 22238 36382
rect 22718 36454 22782 36518
rect 22582 36318 22646 36382
rect 22990 36454 23054 36518
rect 22990 36318 23054 36382
rect 23398 36454 23462 36518
rect 23534 36318 23598 36382
rect 115198 36454 115262 36518
rect 115334 36318 115398 36382
rect 115606 36454 115670 36518
rect 115742 36318 115806 36382
rect 116014 36454 116078 36518
rect 116286 36454 116350 36518
rect 116286 36318 116350 36382
rect 116966 36318 117030 36382
rect 21902 36046 21966 36110
rect 22174 36046 22238 36110
rect 22582 36046 22646 36110
rect 22718 35910 22782 35974
rect 22990 36046 23054 36110
rect 23126 35910 23190 35974
rect 23534 36046 23598 36110
rect 115334 36046 115398 36110
rect 23398 35910 23462 35974
rect 1230 35774 1294 35838
rect 28566 35774 28630 35838
rect 21902 35638 21966 35702
rect 22718 35638 22782 35702
rect 23126 35638 23190 35702
rect 21902 35366 21966 35430
rect 21766 35230 21830 35294
rect 22582 35230 22646 35294
rect 14830 35094 14894 35158
rect 14558 34822 14622 34886
rect 21766 34958 21830 35022
rect 21902 34822 21966 34886
rect 22582 34822 22646 34886
rect 21902 34550 21966 34614
rect 21902 34414 21966 34478
rect 22446 34414 22510 34478
rect 23126 34414 23190 34478
rect 23398 35638 23462 35702
rect 28566 35502 28630 35566
rect 115334 35910 115398 35974
rect 115742 36046 115806 36110
rect 115606 35910 115670 35974
rect 116286 36046 116350 36110
rect 116558 35910 116622 35974
rect 116966 36046 117030 36110
rect 110302 35774 110366 35838
rect 110302 35502 110366 35566
rect 115334 35638 115398 35702
rect 23398 34414 23462 34478
rect 115606 35638 115670 35702
rect 116286 35638 116350 35702
rect 116558 35638 116622 35702
rect 116966 35638 117030 35702
rect 137502 35638 137566 35702
rect 116286 35366 116350 35430
rect 116558 35230 116622 35294
rect 116966 35366 117030 35430
rect 116830 35230 116894 35294
rect 110438 34958 110502 35022
rect 110166 34686 110230 34750
rect 110438 34686 110502 34750
rect 21902 34142 21966 34206
rect 1230 34006 1294 34070
rect 21766 34006 21830 34070
rect 22446 34142 22510 34206
rect 22174 34006 22238 34070
rect 22718 34006 22782 34070
rect 23126 34142 23190 34206
rect 22990 34006 23054 34070
rect 23398 34142 23462 34206
rect 23534 34006 23598 34070
rect 28294 34142 28358 34206
rect 110166 34414 110230 34478
rect 115334 34414 115398 34478
rect 116830 34958 116894 35022
rect 116558 34822 116622 34886
rect 116966 34822 117030 34886
rect 115606 34414 115670 34478
rect 116014 34414 116078 34478
rect 116966 34550 117030 34614
rect 116966 34414 117030 34478
rect 115334 34142 115398 34206
rect 115334 34006 115398 34070
rect 115606 34142 115670 34206
rect 115606 34006 115670 34070
rect 116014 34142 116078 34206
rect 116286 34006 116350 34070
rect 116558 34006 116622 34070
rect 116966 34142 117030 34206
rect 116830 34006 116894 34070
rect 28294 33870 28358 33934
rect 21766 33734 21830 33798
rect 14694 33598 14758 33662
rect 21902 33598 21966 33662
rect 22174 33734 22238 33798
rect 22718 33734 22782 33798
rect 22990 33734 23054 33798
rect 23126 33598 23190 33662
rect 23534 33734 23598 33798
rect 23398 33598 23462 33662
rect 14694 33462 14758 33526
rect 137502 34006 137566 34070
rect 115334 33734 115398 33798
rect 115198 33598 115262 33662
rect 115606 33734 115670 33798
rect 115606 33598 115670 33662
rect 116286 33734 116350 33798
rect 116558 33734 116622 33798
rect 116150 33598 116214 33662
rect 116830 33734 116894 33798
rect 116966 33598 117030 33662
rect 21902 33326 21966 33390
rect 21766 33190 21830 33254
rect 22174 33190 22238 33254
rect 22582 33190 22646 33254
rect 23126 33326 23190 33390
rect 22990 33190 23054 33254
rect 23398 33326 23462 33390
rect 23534 33190 23598 33254
rect 115198 33326 115262 33390
rect 115334 33190 115398 33254
rect 115606 33326 115670 33390
rect 115742 33190 115806 33254
rect 116150 33326 116214 33390
rect 116150 33190 116214 33254
rect 116422 33190 116486 33254
rect 116966 33326 117030 33390
rect 116830 33190 116894 33254
rect 21766 32918 21830 32982
rect 21902 32782 21966 32846
rect 22174 32918 22238 32982
rect 22582 32918 22646 32982
rect 22310 32782 22374 32846
rect 22446 32782 22510 32846
rect 22990 32918 23054 32982
rect 22990 32782 23054 32846
rect 23534 32918 23598 32982
rect 23534 32782 23598 32846
rect 115334 32918 115398 32982
rect 115334 32782 115398 32846
rect 115742 32918 115806 32982
rect 115606 32782 115670 32846
rect 116150 32918 116214 32982
rect 116422 32918 116486 32982
rect 116014 32782 116078 32846
rect 116286 32782 116350 32846
rect 116830 32918 116894 32982
rect 116830 32782 116894 32846
rect 21902 32510 21966 32574
rect 1230 32374 1294 32438
rect 21902 32374 21966 32438
rect 22310 32510 22374 32574
rect 22446 32510 22510 32574
rect 22990 32510 23054 32574
rect 22990 32374 23054 32438
rect 23534 32510 23598 32574
rect 23398 32374 23462 32438
rect 115334 32510 115398 32574
rect 115198 32374 115262 32438
rect 115606 32510 115670 32574
rect 115606 32374 115670 32438
rect 116014 32510 116078 32574
rect 116286 32510 116350 32574
rect 116014 32374 116078 32438
rect 116286 32374 116350 32438
rect 116830 32510 116894 32574
rect 116966 32374 117030 32438
rect 137502 32374 137566 32438
rect 14558 32238 14622 32302
rect 14558 32102 14622 32166
rect 21902 32102 21966 32166
rect 22582 31966 22646 32030
rect 22990 32102 23054 32166
rect 23126 31966 23190 32030
rect 23398 32102 23462 32166
rect 115198 32102 115262 32166
rect 23534 31966 23598 32030
rect 115334 31966 115398 32030
rect 115606 32102 115670 32166
rect 115742 31966 115806 32030
rect 116014 32102 116078 32166
rect 116286 32102 116350 32166
rect 116966 32102 117030 32166
rect 110166 31830 110230 31894
rect 21766 31694 21830 31758
rect 22582 31694 22646 31758
rect 23126 31694 23190 31758
rect 22990 31558 23054 31622
rect 23534 31694 23598 31758
rect 23398 31558 23462 31622
rect 21766 31422 21830 31486
rect 22582 31150 22646 31214
rect 22990 31286 23054 31350
rect 21766 30878 21830 30942
rect 14694 30742 14758 30806
rect 22582 30878 22646 30942
rect 23398 31286 23462 31350
rect 110166 31558 110230 31622
rect 115334 31694 115398 31758
rect 115198 31558 115262 31622
rect 115742 31694 115806 31758
rect 115606 31558 115670 31622
rect 116150 31694 116214 31758
rect 116286 31694 116350 31758
rect 116422 31694 116486 31758
rect 116830 31694 116894 31758
rect 116422 31422 116486 31486
rect 115198 31286 115262 31350
rect 1230 30606 1294 30670
rect 18502 30606 18566 30670
rect 21766 30606 21830 30670
rect 21902 30470 21966 30534
rect 22446 30470 22510 30534
rect 22718 30470 22782 30534
rect 21902 30198 21966 30262
rect 21766 30062 21830 30126
rect 22446 30198 22510 30262
rect 22718 30198 22782 30262
rect 23126 30062 23190 30126
rect 28294 31014 28358 31078
rect 28294 30742 28358 30806
rect 28294 30606 28358 30670
rect 110438 30606 110502 30670
rect 115606 31286 115670 31350
rect 116014 31150 116078 31214
rect 116830 31422 116894 31486
rect 28294 30334 28358 30398
rect 23398 30062 23462 30126
rect 28294 30198 28358 30262
rect 110438 30334 110502 30398
rect 110166 30198 110230 30262
rect 116014 30878 116078 30942
rect 116830 30878 116894 30942
rect 116286 30470 116350 30534
rect 116830 30606 116894 30670
rect 116966 30470 117030 30534
rect 137502 30470 137566 30534
rect 115334 30062 115398 30126
rect 115742 30062 115806 30126
rect 28294 29926 28358 29990
rect 21766 29790 21830 29854
rect 21766 29654 21830 29718
rect 22582 29654 22646 29718
rect 23126 29790 23190 29854
rect 22990 29654 23054 29718
rect 23398 29790 23462 29854
rect 110166 29926 110230 29990
rect 116286 30198 116350 30262
rect 116966 30198 117030 30262
rect 116966 30062 117030 30126
rect 115334 29790 115398 29854
rect 23398 29654 23462 29718
rect 115198 29654 115262 29718
rect 115742 29790 115806 29854
rect 115606 29654 115670 29718
rect 116014 29654 116078 29718
rect 116966 29790 117030 29854
rect 116966 29654 117030 29718
rect 14558 29382 14622 29446
rect 21766 29382 21830 29446
rect 16598 29246 16662 29310
rect 21902 29246 21966 29310
rect 22582 29382 22646 29446
rect 22718 29246 22782 29310
rect 22990 29382 23054 29446
rect 22990 29246 23054 29310
rect 23398 29382 23462 29446
rect 23398 29246 23462 29310
rect 115198 29382 115262 29446
rect 115198 29246 115262 29310
rect 115606 29382 115670 29446
rect 115606 29246 115670 29310
rect 116014 29382 116078 29446
rect 116150 29246 116214 29310
rect 116966 29382 117030 29446
rect 116966 29246 117030 29310
rect 1230 28838 1294 28902
rect 18094 28838 18158 28902
rect 18502 28974 18566 29038
rect 18910 28838 18974 28902
rect 19454 28838 19518 28902
rect 21902 28974 21966 29038
rect 21766 28838 21830 28902
rect 22718 28974 22782 29038
rect 22174 28838 22238 28902
rect 22446 28838 22510 28902
rect 22990 28974 23054 29038
rect 22990 28838 23054 28902
rect 23398 28974 23462 29038
rect 115198 28974 115262 29038
rect 23534 28838 23598 28902
rect 115334 28838 115398 28902
rect 115606 28974 115670 29038
rect 115742 28838 115806 28902
rect 116150 28974 116214 29038
rect 116014 28838 116078 28902
rect 116966 28974 117030 29038
rect 116830 28838 116894 28902
rect 119006 28838 119070 28902
rect 119278 28838 119342 28902
rect 119958 28838 120022 28902
rect 120502 28838 120566 28902
rect 137502 28974 137566 29038
rect 21766 28566 21830 28630
rect 21766 28430 21830 28494
rect 22174 28566 22238 28630
rect 22446 28566 22510 28630
rect 22990 28566 23054 28630
rect 22990 28430 23054 28494
rect 23534 28566 23598 28630
rect 23398 28430 23462 28494
rect 115334 28566 115398 28630
rect 115334 28430 115398 28494
rect 115742 28566 115806 28630
rect 115742 28430 115806 28494
rect 116014 28566 116078 28630
rect 116830 28566 116894 28630
rect 116966 28430 117030 28494
rect 18094 28158 18158 28222
rect 18094 28022 18158 28086
rect 18910 28158 18974 28222
rect 19454 28158 19518 28222
rect 19046 28022 19110 28086
rect 19454 28022 19518 28086
rect 19726 28022 19790 28086
rect 21766 28158 21830 28222
rect 22310 28022 22374 28086
rect 22718 28022 22782 28086
rect 22990 28158 23054 28222
rect 22990 28022 23054 28086
rect 23398 28158 23462 28222
rect 23398 28022 23462 28086
rect 19318 27614 19382 27678
rect 28294 27886 28358 27950
rect 115334 28158 115398 28222
rect 115334 28022 115398 28086
rect 115742 28158 115806 28222
rect 115742 28022 115806 28086
rect 116014 28022 116078 28086
rect 116966 28158 117030 28222
rect 119006 28158 119070 28222
rect 119006 28022 119070 28086
rect 119278 28158 119342 28222
rect 119958 28158 120022 28222
rect 119414 28022 119478 28086
rect 119958 28022 120022 28086
rect 120502 28158 120566 28222
rect 120638 28022 120702 28086
rect 22310 27750 22374 27814
rect 22718 27750 22782 27814
rect 22990 27750 23054 27814
rect 23126 27614 23190 27678
rect 23398 27750 23462 27814
rect 23534 27614 23598 27678
rect 28294 27614 28358 27678
rect 18094 27478 18158 27542
rect 1230 27342 1294 27406
rect 18094 27206 18158 27270
rect 19046 27478 19110 27542
rect 18502 27206 18566 27270
rect 19318 27342 19382 27406
rect 19454 27342 19518 27406
rect 19318 27206 19382 27270
rect 19726 27342 19790 27406
rect 19862 27206 19926 27270
rect 22310 27206 22374 27270
rect 23126 27342 23190 27406
rect 23534 27342 23598 27406
rect 28430 27342 28494 27406
rect 115334 27750 115398 27814
rect 115334 27614 115398 27678
rect 115742 27750 115806 27814
rect 115742 27614 115806 27678
rect 116014 27750 116078 27814
rect 110166 27342 110230 27406
rect 18910 27070 18974 27134
rect 21902 26934 21966 26998
rect 22310 26934 22374 26998
rect 16598 26662 16662 26726
rect 18094 26662 18158 26726
rect 18910 26662 18974 26726
rect 19318 26662 19382 26726
rect 18502 26390 18566 26454
rect 19454 26390 19518 26454
rect 19862 26662 19926 26726
rect 21902 26662 21966 26726
rect 21766 26526 21830 26590
rect 22718 26526 22782 26590
rect 19726 26390 19790 26454
rect 28430 27070 28494 27134
rect 28566 27070 28630 27134
rect 28566 26798 28630 26862
rect 28294 26662 28358 26726
rect 110166 27070 110230 27134
rect 110302 27070 110366 27134
rect 110302 26798 110366 26862
rect 115334 27342 115398 27406
rect 115742 27342 115806 27406
rect 116558 27206 116622 27270
rect 119958 27478 120022 27542
rect 119006 27342 119070 27406
rect 119414 27342 119478 27406
rect 119278 27206 119342 27270
rect 120094 27206 120158 27270
rect 120638 27478 120702 27542
rect 120502 27206 120566 27270
rect 137502 27206 137566 27270
rect 110302 26662 110366 26726
rect 28294 26390 28358 26454
rect 21766 26254 21830 26318
rect 21902 26118 21966 26182
rect 22718 26254 22782 26318
rect 22446 25982 22510 26046
rect 22990 26118 23054 26182
rect 23398 26118 23462 26182
rect 110302 26390 110366 26454
rect 110438 26254 110502 26318
rect 116558 26934 116622 26998
rect 116830 26934 116894 26998
rect 116014 26526 116078 26590
rect 116830 26662 116894 26726
rect 116830 26526 116894 26590
rect 119278 26662 119342 26726
rect 120094 26662 120158 26726
rect 119822 26526 119886 26590
rect 120502 26662 120566 26726
rect 119414 26390 119478 26454
rect 115198 26118 115262 26182
rect 115606 26118 115670 26182
rect 116014 26254 116078 26318
rect 550 25846 614 25910
rect 3814 25846 3878 25910
rect 21902 25846 21966 25910
rect 21902 25710 21966 25774
rect 22582 25846 22646 25910
rect 22446 25710 22510 25774
rect 22990 25846 23054 25910
rect 23126 25710 23190 25774
rect 23398 25846 23462 25910
rect 28566 25846 28630 25910
rect 110438 25982 110502 26046
rect 116830 26254 116894 26318
rect 116966 26118 117030 26182
rect 115198 25846 115262 25910
rect 23534 25710 23598 25774
rect 1230 25574 1294 25638
rect 21902 25438 21966 25502
rect 2541 25361 2605 25365
rect 2541 25305 2545 25361
rect 2545 25305 2601 25361
rect 2601 25305 2605 25361
rect 2541 25301 2605 25305
rect 19590 25302 19654 25366
rect 21766 25302 21830 25366
rect 22446 25438 22510 25502
rect 22174 25302 22238 25366
rect 22718 25302 22782 25366
rect 23126 25438 23190 25502
rect 22990 25302 23054 25366
rect 23534 25438 23598 25502
rect 23534 25302 23598 25366
rect 28566 25438 28630 25502
rect 115334 25710 115398 25774
rect 115606 25846 115670 25910
rect 115742 25710 115806 25774
rect 116286 25710 116350 25774
rect 116422 25710 116486 25774
rect 116966 25846 117030 25910
rect 116966 25710 117030 25774
rect 119278 25710 119342 25774
rect 137502 25574 137566 25638
rect 115334 25438 115398 25502
rect 115198 25302 115262 25366
rect 115742 25438 115806 25502
rect 115742 25302 115806 25366
rect 116286 25438 116350 25502
rect 116422 25438 116486 25502
rect 116558 25302 116622 25366
rect 116966 25438 117030 25502
rect 116966 25302 117030 25366
rect 18230 24894 18294 24958
rect 19454 25030 19518 25094
rect 19590 25030 19654 25094
rect 19726 25030 19790 25094
rect 18910 24894 18974 24958
rect 19318 24894 19382 24958
rect 21766 25030 21830 25094
rect 21902 24894 21966 24958
rect 22174 25030 22238 25094
rect 22718 25030 22782 25094
rect 22174 24894 22238 24958
rect 22990 25030 23054 25094
rect 23126 24894 23190 24958
rect 23534 25030 23598 25094
rect 115198 25030 115262 25094
rect 23398 24894 23462 24958
rect 115198 24894 115262 24958
rect 115742 25030 115806 25094
rect 115606 24894 115670 24958
rect 116558 25030 116622 25094
rect 116150 24894 116214 24958
rect 116966 25030 117030 25094
rect 116966 24894 117030 24958
rect 119006 24894 119070 24958
rect 119278 25030 119342 25094
rect 119414 25030 119478 25094
rect 119414 24894 119478 24958
rect 119822 25030 119886 25094
rect 120094 24894 120158 24958
rect 120638 24894 120702 24958
rect 2318 24486 2382 24550
rect 21902 24622 21966 24686
rect 21766 24486 21830 24550
rect 22174 24622 22238 24686
rect 22310 24486 22374 24550
rect 23126 24622 23190 24686
rect 23126 24486 23190 24550
rect 23398 24622 23462 24686
rect 23534 24486 23598 24550
rect 115198 24622 115262 24686
rect 115198 24486 115262 24550
rect 115606 24622 115670 24686
rect 115742 24486 115806 24550
rect 116150 24622 116214 24686
rect 116014 24486 116078 24550
rect 116966 24622 117030 24686
rect 116830 24486 116894 24550
rect 18230 24214 18294 24278
rect 18230 24078 18294 24142
rect 18910 24214 18974 24278
rect 18502 24078 18566 24142
rect 19318 24214 19382 24278
rect 19318 24078 19382 24142
rect 19862 24078 19926 24142
rect 21766 24214 21830 24278
rect 22310 24214 22374 24278
rect 22310 24078 22374 24142
rect 22582 24078 22646 24142
rect 23126 24214 23190 24278
rect 22990 24078 23054 24142
rect 23534 24214 23598 24278
rect 23398 24078 23462 24142
rect 115198 24214 115262 24278
rect 1230 23942 1294 24006
rect 2318 23942 2382 24006
rect 28430 23942 28494 24006
rect 115334 24078 115398 24142
rect 115742 24214 115806 24278
rect 115742 24078 115806 24142
rect 116014 24214 116078 24278
rect 116150 24078 116214 24142
rect 116558 24078 116622 24142
rect 116830 24214 116894 24278
rect 119006 24214 119070 24278
rect 119414 24214 119478 24278
rect 119006 24078 119070 24142
rect 120094 24214 120158 24278
rect 119278 24078 119342 24142
rect 119686 24078 119750 24142
rect 120638 24214 120702 24278
rect 120638 24078 120702 24142
rect 110438 23942 110502 24006
rect 22310 23806 22374 23870
rect 22582 23806 22646 23870
rect 22990 23806 23054 23870
rect 22990 23670 23054 23734
rect 23398 23806 23462 23870
rect 23398 23670 23462 23734
rect 28430 23670 28494 23734
rect 18230 23534 18294 23598
rect 3814 23262 3878 23326
rect 18230 23262 18294 23326
rect 18502 23534 18566 23598
rect 18638 23262 18702 23326
rect 19318 23398 19382 23462
rect 19318 23262 19382 23326
rect 19862 23398 19926 23462
rect 19726 23262 19790 23326
rect 22174 23262 22238 23326
rect 22582 23262 22646 23326
rect 22990 23398 23054 23462
rect 23126 23262 23190 23326
rect 23398 23398 23462 23462
rect 110438 23670 110502 23734
rect 115334 23806 115398 23870
rect 115334 23670 115398 23734
rect 115742 23806 115806 23870
rect 115742 23670 115806 23734
rect 116150 23806 116214 23870
rect 116558 23806 116622 23870
rect 120502 23942 120566 24006
rect 137502 23942 137566 24006
rect 115334 23398 115398 23462
rect 23534 23262 23598 23326
rect 18366 23126 18430 23190
rect 115334 23262 115398 23326
rect 115742 23398 115806 23462
rect 115742 23262 115806 23326
rect 116286 23262 116350 23326
rect 119686 23534 119750 23598
rect 119006 23398 119070 23462
rect 119006 23262 119070 23326
rect 119278 23398 119342 23462
rect 119278 23262 119342 23326
rect 119686 23262 119750 23326
rect 120502 23534 120566 23598
rect 120638 23534 120702 23598
rect 120638 23262 120702 23326
rect 110438 23126 110502 23190
rect 21766 22990 21830 23054
rect 22174 22990 22238 23054
rect 22582 22990 22646 23054
rect 23126 22990 23190 23054
rect 18230 22718 18294 22782
rect 18366 22718 18430 22782
rect 18638 22718 18702 22782
rect 19318 22718 19382 22782
rect 18638 22446 18702 22510
rect 19726 22718 19790 22782
rect 21766 22718 21830 22782
rect 21766 22582 21830 22646
rect 22446 22582 22510 22646
rect 19862 22446 19926 22510
rect 23534 22990 23598 23054
rect 28566 22718 28630 22782
rect 110438 22854 110502 22918
rect 110166 22718 110230 22782
rect 115334 22990 115398 23054
rect 115742 22990 115806 23054
rect 116286 22990 116350 23054
rect 116830 22990 116894 23054
rect 1230 22310 1294 22374
rect 21766 22310 21830 22374
rect 3134 22174 3198 22238
rect 21766 22174 21830 22238
rect 22446 22310 22510 22374
rect 28294 22310 28358 22374
rect 28566 22310 28630 22374
rect 28294 22038 28358 22102
rect 28430 22038 28494 22102
rect 21766 21902 21830 21966
rect 3134 21766 3198 21830
rect 21902 21766 21966 21830
rect 22310 21766 22374 21830
rect 23126 21766 23190 21830
rect 110166 22446 110230 22510
rect 23398 21766 23462 21830
rect 28430 21766 28494 21830
rect 21902 21494 21966 21558
rect 21902 21358 21966 21422
rect 22310 21494 22374 21558
rect 22310 21358 22374 21422
rect 22446 21358 22510 21422
rect 23126 21494 23190 21558
rect 22990 21358 23054 21422
rect 23398 21494 23462 21558
rect 23398 21358 23462 21422
rect 18638 21086 18702 21150
rect 18910 20950 18974 21014
rect 19318 20950 19382 21014
rect 19862 21086 19926 21150
rect 19862 20950 19926 21014
rect 21902 21086 21966 21150
rect 21766 20950 21830 21014
rect 22310 21086 22374 21150
rect 22446 21086 22510 21150
rect 22718 20950 22782 21014
rect 22990 21086 23054 21150
rect 22990 20950 23054 21014
rect 23398 21086 23462 21150
rect 116286 22582 116350 22646
rect 116830 22718 116894 22782
rect 116830 22582 116894 22646
rect 119006 22718 119070 22782
rect 119006 22446 119070 22510
rect 119278 22718 119342 22782
rect 119686 22718 119750 22782
rect 120638 22718 120702 22782
rect 120502 22582 120566 22646
rect 116286 22310 116350 22374
rect 116830 22310 116894 22374
rect 116830 22174 116894 22238
rect 137502 22310 137566 22374
rect 115198 21766 115262 21830
rect 115606 21766 115670 21830
rect 116558 21766 116622 21830
rect 116830 21902 116894 21966
rect 116966 21766 117030 21830
rect 115198 21494 115262 21558
rect 115334 21358 115398 21422
rect 115606 21494 115670 21558
rect 115606 21358 115670 21422
rect 116558 21494 116622 21558
rect 116966 21494 117030 21558
rect 116014 21358 116078 21422
rect 116966 21358 117030 21422
rect 115334 21086 115398 21150
rect 23534 20950 23598 21014
rect 21766 20678 21830 20742
rect 21902 20542 21966 20606
rect 22718 20678 22782 20742
rect 22310 20542 22374 20606
rect 22718 20542 22782 20606
rect 22990 20678 23054 20742
rect 22990 20542 23054 20606
rect 23534 20678 23598 20742
rect 23398 20542 23462 20606
rect 115198 20950 115262 21014
rect 115606 21086 115670 21150
rect 115606 20950 115670 21014
rect 116014 21086 116078 21150
rect 116014 20950 116078 21014
rect 116966 21086 117030 21150
rect 116830 20950 116894 21014
rect 119006 21086 119070 21150
rect 118870 20950 118934 21014
rect 119414 20950 119478 21014
rect 119822 20950 119886 21014
rect 120502 21086 120566 21150
rect 115198 20678 115262 20742
rect 115198 20542 115262 20606
rect 115606 20678 115670 20742
rect 115606 20542 115670 20606
rect 116014 20678 116078 20742
rect 116014 20542 116078 20606
rect 116830 20678 116894 20742
rect 116966 20542 117030 20606
rect 1230 20406 1294 20470
rect 550 20270 614 20334
rect 3950 20270 4014 20334
rect 17142 20134 17206 20198
rect 17550 20134 17614 20198
rect 18910 20270 18974 20334
rect 19318 20270 19382 20334
rect 19862 20270 19926 20334
rect 21902 20270 21966 20334
rect 21766 20134 21830 20198
rect 22310 20270 22374 20334
rect 22718 20270 22782 20334
rect 22990 20270 23054 20334
rect 23398 20270 23462 20334
rect 137502 20406 137566 20470
rect 23534 20134 23598 20198
rect 24214 20134 24278 20198
rect 28294 19998 28358 20062
rect 115198 20270 115262 20334
rect 115606 20270 115670 20334
rect 116014 20270 116078 20334
rect 116966 20270 117030 20334
rect 118870 20270 118934 20334
rect 119414 20270 119478 20334
rect 119822 20270 119886 20334
rect 121318 20134 121382 20198
rect 124174 20134 124238 20198
rect 23534 19726 23598 19790
rect 23398 19590 23462 19654
rect 24214 19726 24278 19790
rect 124174 19862 124238 19926
rect 110166 19726 110230 19790
rect 124310 19726 124374 19790
rect 27886 19590 27950 19654
rect 28294 19590 28358 19654
rect 27886 19318 27950 19382
rect 29110 19182 29174 19246
rect 30470 19182 30534 19246
rect 32238 19182 32302 19246
rect 32782 19182 32846 19246
rect 32918 19182 32982 19246
rect 34142 19182 34206 19246
rect 34686 19182 34750 19246
rect 35502 19182 35566 19246
rect 35910 19182 35974 19246
rect 36726 19182 36790 19246
rect 38494 19182 38558 19246
rect 39174 19182 39238 19246
rect 39582 19182 39646 19246
rect 40942 19182 41006 19246
rect 41622 19182 41686 19246
rect 42846 19182 42910 19246
rect 43390 19182 43454 19246
rect 44070 19182 44134 19246
rect 45702 19182 45766 19246
rect 46654 19182 46718 19246
rect 47198 19182 47262 19246
rect 47878 19182 47942 19246
rect 48422 19182 48486 19246
rect 49102 19182 49166 19246
rect 49646 19182 49710 19246
rect 50462 19182 50526 19246
rect 52094 19182 52158 19246
rect 52910 19182 52974 19246
rect 54134 19182 54198 19246
rect 54678 19182 54742 19246
rect 55358 19182 55422 19246
rect 55902 19182 55966 19246
rect 56718 19182 56782 19246
rect 57126 19182 57190 19246
rect 57670 19182 57734 19246
rect 58350 19182 58414 19246
rect 59166 19182 59230 19246
rect 60526 19318 60590 19382
rect 59710 19182 59774 19246
rect 61614 19182 61678 19246
rect 62158 19182 62222 19246
rect 62838 19182 62902 19246
rect 63382 19182 63446 19246
rect 64198 19182 64262 19246
rect 64606 19182 64670 19246
rect 65830 19182 65894 19246
rect 67190 19182 67254 19246
rect 67870 19182 67934 19246
rect 68414 19182 68478 19246
rect 69094 19182 69158 19246
rect 70318 19182 70382 19246
rect 70862 19182 70926 19246
rect 71542 19182 71606 19246
rect 73310 19182 73374 19246
rect 74670 19182 74734 19246
rect 75214 19182 75278 19246
rect 75350 19182 75414 19246
rect 75894 19182 75958 19246
rect 76574 19182 76638 19246
rect 77118 19182 77182 19246
rect 77934 19182 77998 19246
rect 78342 19182 78406 19246
rect 79158 19182 79222 19246
rect 80518 19182 80582 19246
rect 81470 19182 81534 19246
rect 81606 19182 81670 19246
rect 82014 19182 82078 19246
rect 82830 19182 82894 19246
rect 83374 19182 83438 19246
rect 84054 19182 84118 19246
rect 84598 19182 84662 19246
rect 85278 19182 85342 19246
rect 85822 19182 85886 19246
rect 86502 19182 86566 19246
rect 86774 19182 86838 19246
rect 88134 19182 88198 19246
rect 89630 19182 89694 19246
rect 90310 19182 90374 19246
rect 90854 19182 90918 19246
rect 94254 19318 94318 19382
rect 92078 19182 92142 19246
rect 92758 19182 92822 19246
rect 94390 19182 94454 19246
rect 95342 19182 95406 19246
rect 95750 19182 95814 19246
rect 96566 19182 96630 19246
rect 98334 19182 98398 19246
rect 99150 19182 99214 19246
rect 99558 19182 99622 19246
rect 100374 19182 100438 19246
rect 101598 19182 101662 19246
rect 102958 19318 103022 19382
rect 102006 19182 102070 19246
rect 104046 19182 104110 19246
rect 104590 19182 104654 19246
rect 105270 19182 105334 19246
rect 105814 19182 105878 19246
rect 106630 19182 106694 19246
rect 107038 19182 107102 19246
rect 108262 19182 108326 19246
rect 109078 19182 109142 19246
rect 1230 18910 1294 18974
rect 17142 19046 17206 19110
rect 35910 18910 35974 18974
rect 78342 18910 78406 18974
rect 15238 18774 15302 18838
rect 29110 18774 29174 18838
rect 30470 18774 30534 18838
rect 32238 18774 32302 18838
rect 32782 18774 32846 18838
rect 32918 18774 32982 18838
rect 34142 18774 34206 18838
rect 34686 18774 34750 18838
rect 35502 18774 35566 18838
rect 36726 18774 36790 18838
rect 38494 18774 38558 18838
rect 39174 18774 39238 18838
rect 39582 18774 39646 18838
rect 40942 18774 41006 18838
rect 41622 18774 41686 18838
rect 42846 18774 42910 18838
rect 43390 18774 43454 18838
rect 44070 18774 44134 18838
rect 45702 18774 45766 18838
rect 46654 18774 46718 18838
rect 47198 18774 47262 18838
rect 47878 18774 47942 18838
rect 48422 18774 48486 18838
rect 49102 18774 49166 18838
rect 49646 18774 49710 18838
rect 50462 18774 50526 18838
rect 52094 18774 52158 18838
rect 52910 18774 52974 18838
rect 54134 18774 54198 18838
rect 54678 18774 54742 18838
rect 55358 18774 55422 18838
rect 55902 18774 55966 18838
rect 56718 18774 56782 18838
rect 57126 18774 57190 18838
rect 57670 18774 57734 18838
rect 58350 18774 58414 18838
rect 59166 18774 59230 18838
rect 59710 18774 59774 18838
rect 60526 18774 60590 18838
rect 61614 18774 61678 18838
rect 62158 18774 62222 18838
rect 62838 18774 62902 18838
rect 63382 18774 63446 18838
rect 64198 18774 64262 18838
rect 64606 18774 64670 18838
rect 65830 18774 65894 18838
rect 67190 18774 67254 18838
rect 67870 18774 67934 18838
rect 68414 18774 68478 18838
rect 69094 18774 69158 18838
rect 70318 18774 70382 18838
rect 70862 18774 70926 18838
rect 71542 18774 71606 18838
rect 73310 18774 73374 18838
rect 74670 18774 74734 18838
rect 75214 18774 75278 18838
rect 75350 18774 75414 18838
rect 75894 18774 75958 18838
rect 76574 18774 76638 18838
rect 77118 18774 77182 18838
rect 77118 18638 77182 18702
rect 77934 18774 77998 18838
rect 79158 18774 79222 18838
rect 80518 18774 80582 18838
rect 81470 18774 81534 18838
rect 81606 18774 81670 18838
rect 82014 18774 82078 18838
rect 82830 18774 82894 18838
rect 83374 18774 83438 18838
rect 84054 18774 84118 18838
rect 84598 18774 84662 18838
rect 85278 18774 85342 18838
rect 85822 18774 85886 18838
rect 86502 18774 86566 18838
rect 86774 18774 86838 18838
rect 88134 18774 88198 18838
rect 89630 18774 89694 18838
rect 90310 18774 90374 18838
rect 90854 18774 90918 18838
rect 92078 18774 92142 18838
rect 92758 18774 92822 18838
rect 94254 18774 94318 18838
rect 94390 18774 94454 18838
rect 95342 18774 95406 18838
rect 95750 18774 95814 18838
rect 96566 18774 96630 18838
rect 98334 18774 98398 18838
rect 99150 18774 99214 18838
rect 99558 18774 99622 18838
rect 100374 18774 100438 18838
rect 101598 18774 101662 18838
rect 102006 18774 102070 18838
rect 102958 18774 103022 18838
rect 104046 18774 104110 18838
rect 104590 18774 104654 18838
rect 105270 18774 105334 18838
rect 105814 18774 105878 18838
rect 106630 18774 106694 18838
rect 107038 18774 107102 18838
rect 108262 18774 108326 18838
rect 109078 18774 109142 18838
rect 137502 18774 137566 18838
rect 121318 18502 121382 18566
rect 124174 18366 124238 18430
rect 2541 17894 2605 17958
rect 3814 17550 3878 17614
rect 17550 17550 17614 17614
rect 15102 17414 15166 17478
rect 21766 17278 21830 17342
rect 21086 17142 21150 17206
rect 1230 17006 1294 17070
rect 29926 17006 29990 17070
rect 32646 17006 32710 17070
rect 35094 17006 35158 17070
rect 37406 17006 37470 17070
rect 40126 17006 40190 17070
rect 42438 17006 42502 17070
rect 44886 17006 44950 17070
rect 47606 17006 47670 17070
rect 49918 17006 49982 17070
rect 52502 17006 52566 17070
rect 55086 17006 55150 17070
rect 57398 17006 57462 17070
rect 59982 17006 60046 17070
rect 62566 17006 62630 17070
rect 64878 17006 64942 17070
rect 67598 17006 67662 17070
rect 69910 17006 69974 17070
rect 72358 17006 72422 17070
rect 75078 17006 75142 17070
rect 77526 17006 77590 17070
rect 79838 17006 79902 17070
rect 82558 17006 82622 17070
rect 84870 17006 84934 17070
rect 87318 17006 87382 17070
rect 90038 17006 90102 17070
rect 92350 17006 92414 17070
rect 94934 17006 94998 17070
rect 97518 17006 97582 17070
rect 99830 17006 99894 17070
rect 102414 17006 102478 17070
rect 104998 17006 105062 17070
rect 110166 17142 110230 17206
rect 107310 17006 107374 17070
rect 124310 17006 124374 17070
rect 137502 17006 137566 17070
rect 124446 16870 124510 16934
rect 3134 16054 3198 16118
rect 15238 16190 15302 16254
rect 15238 16054 15302 16118
rect 22310 15782 22374 15846
rect 23398 15782 23462 15846
rect 124174 15646 124238 15710
rect 1230 15510 1294 15574
rect 3134 15510 3198 15574
rect 124310 15510 124374 15574
rect 137502 15510 137566 15574
rect 29926 15102 29990 15166
rect 30062 15102 30126 15166
rect 32510 15102 32574 15166
rect 32646 15102 32710 15166
rect 34958 15102 35022 15166
rect 35094 15102 35158 15166
rect 37406 15102 37470 15166
rect 37542 15102 37606 15166
rect 39990 15102 40054 15166
rect 40126 15102 40190 15166
rect 42438 15102 42502 15166
rect 42574 15102 42638 15166
rect 44886 15102 44950 15166
rect 45022 15102 45086 15166
rect 47470 15102 47534 15166
rect 47606 15102 47670 15166
rect 49918 15102 49982 15166
rect 50190 15102 50254 15166
rect 52366 15102 52430 15166
rect 52502 15102 52566 15166
rect 54950 15102 55014 15166
rect 55086 15102 55150 15166
rect 57398 15102 57462 15166
rect 57534 15102 57598 15166
rect 59846 15102 59910 15166
rect 59982 15102 60046 15166
rect 62430 15102 62494 15166
rect 62566 15102 62630 15166
rect 64878 15102 64942 15166
rect 65014 15102 65078 15166
rect 67462 15102 67526 15166
rect 67598 15102 67662 15166
rect 69910 15102 69974 15166
rect 70046 15102 70110 15166
rect 72358 15102 72422 15166
rect 72494 15102 72558 15166
rect 74942 15102 75006 15166
rect 75078 15102 75142 15166
rect 77390 15102 77454 15166
rect 77526 15102 77590 15166
rect 79838 15102 79902 15166
rect 79974 15102 80038 15166
rect 82422 15102 82486 15166
rect 82558 15102 82622 15166
rect 84870 15102 84934 15166
rect 85006 15102 85070 15166
rect 87318 15102 87382 15166
rect 87454 15102 87518 15166
rect 89902 15102 89966 15166
rect 90038 15102 90102 15166
rect 92350 15102 92414 15166
rect 92486 15102 92550 15166
rect 94798 15102 94862 15166
rect 94934 15102 94998 15166
rect 97382 15102 97446 15166
rect 97518 15102 97582 15166
rect 99830 15102 99894 15166
rect 99966 15102 100030 15166
rect 102278 15102 102342 15166
rect 102414 15102 102478 15166
rect 104862 15102 104926 15166
rect 104998 15102 105062 15166
rect 107310 15102 107374 15166
rect 107446 15102 107510 15166
rect 550 14694 614 14758
rect 15102 14694 15166 14758
rect 15102 14558 15166 14622
rect 21086 14558 21150 14622
rect 22174 14286 22238 14350
rect 29926 14286 29990 14350
rect 32374 14286 32438 14350
rect 34822 14286 34886 14350
rect 37406 14286 37470 14350
rect 39854 14286 39918 14350
rect 42166 14286 42230 14350
rect 44886 14286 44950 14350
rect 47198 14286 47262 14350
rect 49782 14286 49846 14350
rect 52230 14286 52294 14350
rect 54814 14286 54878 14350
rect 57398 14286 57462 14350
rect 59846 14286 59910 14350
rect 62294 14286 62358 14350
rect 64878 14286 64942 14350
rect 67190 14286 67254 14350
rect 69638 14286 69702 14350
rect 72086 14286 72150 14350
rect 72222 14286 72286 14350
rect 77118 14422 77182 14486
rect 74806 14286 74870 14350
rect 76982 14286 77046 14350
rect 77254 14286 77318 14350
rect 79838 14286 79902 14350
rect 82286 14286 82350 14350
rect 84598 14286 84662 14350
rect 87318 14286 87382 14350
rect 89630 14286 89694 14350
rect 92214 14286 92278 14350
rect 94662 14286 94726 14350
rect 97246 14286 97310 14350
rect 99694 14286 99758 14350
rect 102278 14286 102342 14350
rect 104726 14286 104790 14350
rect 107310 14286 107374 14350
rect 124446 14286 124510 14350
rect 124174 14014 124238 14078
rect 1230 13878 1294 13942
rect 137502 13878 137566 13942
rect 3134 13742 3198 13806
rect 29926 13606 29990 13670
rect 32374 13606 32438 13670
rect 34686 13606 34750 13670
rect 34822 13606 34886 13670
rect 37406 13606 37470 13670
rect 29926 13470 29990 13534
rect 32374 13470 32438 13534
rect 37270 13470 37334 13534
rect 39854 13606 39918 13670
rect 42166 13606 42230 13670
rect 44886 13606 44950 13670
rect 47198 13606 47262 13670
rect 49646 13606 49710 13670
rect 49782 13606 49846 13670
rect 52230 13606 52294 13670
rect 39718 13470 39782 13534
rect 42438 13470 42502 13534
rect 44886 13470 44950 13534
rect 47334 13470 47398 13534
rect 54814 13606 54878 13670
rect 57398 13606 57462 13670
rect 59846 13606 59910 13670
rect 62294 13606 62358 13670
rect 52230 13470 52294 13534
rect 54814 13470 54878 13534
rect 57398 13470 57462 13534
rect 59846 13470 59910 13534
rect 62294 13470 62358 13534
rect 64878 13606 64942 13670
rect 67190 13606 67254 13670
rect 69638 13606 69702 13670
rect 69774 13606 69838 13670
rect 72086 13606 72150 13670
rect 72222 13606 72286 13670
rect 74806 13606 74870 13670
rect 76982 13606 77046 13670
rect 77118 13606 77182 13670
rect 77254 13606 77318 13670
rect 79838 13606 79902 13670
rect 82286 13606 82350 13670
rect 84598 13606 84662 13670
rect 87318 13606 87382 13670
rect 89630 13606 89694 13670
rect 92214 13606 92278 13670
rect 94662 13606 94726 13670
rect 97246 13606 97310 13670
rect 99694 13606 99758 13670
rect 102278 13606 102342 13670
rect 104726 13606 104790 13670
rect 107310 13606 107374 13670
rect 64742 13470 64806 13534
rect 67326 13470 67390 13534
rect 72358 13470 72422 13534
rect 74806 13470 74870 13534
rect 79838 13470 79902 13534
rect 82286 13470 82350 13534
rect 84870 13470 84934 13534
rect 87318 13470 87382 13534
rect 89766 13470 89830 13534
rect 92350 13470 92414 13534
rect 94798 13470 94862 13534
rect 97246 13470 97310 13534
rect 99830 13470 99894 13534
rect 102278 13470 102342 13534
rect 104726 13470 104790 13534
rect 107310 13470 107374 13534
rect 124854 13470 124918 13534
rect 3134 13334 3198 13398
rect 15238 13334 15302 13398
rect 15238 13198 15302 13262
rect 30062 13198 30126 13262
rect 22310 13062 22374 13126
rect 28974 13062 29038 13126
rect 32510 13198 32574 13262
rect 30062 13062 30126 13126
rect 31966 13062 32030 13126
rect 32510 13062 32574 13126
rect 34414 13062 34478 13126
rect 34822 13062 34886 13126
rect 34958 13062 35022 13126
rect 36998 13062 37062 13126
rect 37542 13198 37606 13262
rect 37406 13062 37470 13126
rect 39446 13062 39510 13126
rect 39990 13198 40054 13262
rect 42574 13198 42638 13262
rect 45022 13198 45086 13262
rect 49918 13334 49982 13398
rect 39854 13062 39918 13126
rect 41758 13062 41822 13126
rect 42302 13062 42366 13126
rect 44206 13062 44270 13126
rect 47470 13198 47534 13262
rect 45022 13062 45086 13126
rect 46518 13062 46582 13126
rect 47470 13062 47534 13126
rect 49782 13062 49846 13126
rect 50190 13062 50254 13126
rect 51958 13062 52022 13126
rect 52366 13198 52430 13262
rect 52366 13062 52430 13126
rect 54950 13198 55014 13262
rect 54542 13062 54606 13126
rect 57534 13198 57598 13262
rect 59982 13198 60046 13262
rect 54950 13062 55014 13126
rect 56990 13062 57054 13126
rect 57262 13062 57326 13126
rect 59302 13062 59366 13126
rect 62430 13198 62494 13262
rect 59982 13062 60046 13126
rect 61886 13062 61950 13126
rect 62430 13062 62494 13126
rect 64470 13062 64534 13126
rect 65014 13198 65078 13262
rect 64878 13062 64942 13126
rect 67462 13198 67526 13262
rect 66918 13062 66982 13126
rect 67462 13062 67526 13126
rect 69502 13062 69566 13126
rect 72494 13198 72558 13262
rect 69910 13062 69974 13126
rect 71950 13062 72014 13126
rect 74942 13198 75006 13262
rect 72494 13062 72558 13126
rect 74398 13062 74462 13126
rect 74942 13062 75006 13126
rect 76846 13062 76910 13126
rect 77254 13062 77318 13126
rect 77390 13062 77454 13126
rect 79974 13198 80038 13262
rect 79430 13062 79494 13126
rect 82422 13198 82486 13262
rect 79974 13062 80038 13126
rect 81878 13062 81942 13126
rect 85006 13198 85070 13262
rect 82422 13062 82486 13126
rect 84326 13062 84390 13126
rect 84734 13062 84798 13126
rect 87454 13198 87518 13262
rect 86910 13062 86974 13126
rect 89902 13198 89966 13262
rect 87454 13062 87518 13126
rect 89086 13062 89150 13126
rect 92486 13198 92550 13262
rect 89902 13062 89966 13126
rect 91942 13062 92006 13126
rect 92214 13062 92278 13126
rect 94934 13198 94998 13262
rect 94390 13062 94454 13126
rect 97382 13198 97446 13262
rect 94934 13062 94998 13126
rect 96838 13062 96902 13126
rect 99966 13198 100030 13262
rect 97382 13062 97446 13126
rect 99422 13062 99486 13126
rect 99694 13062 99758 13126
rect 102414 13198 102478 13262
rect 101870 13062 101934 13126
rect 104862 13198 104926 13262
rect 102414 13062 102478 13126
rect 104318 13062 104382 13126
rect 107446 13198 107510 13262
rect 104862 13062 104926 13126
rect 106902 13062 106966 13126
rect 107446 13062 107510 13126
rect 70046 12926 70110 12990
rect 124310 12790 124374 12854
rect 124310 12654 124374 12718
rect 30062 12518 30126 12582
rect 32510 12518 32574 12582
rect 34822 12518 34886 12582
rect 29790 12246 29854 12310
rect 32238 12246 32302 12310
rect 34822 12246 34886 12310
rect 37406 12518 37470 12582
rect 39854 12518 39918 12582
rect 42302 12518 42366 12582
rect 37406 12246 37470 12310
rect 39854 12246 39918 12310
rect 42166 12246 42230 12310
rect 45022 12518 45086 12582
rect 47470 12518 47534 12582
rect 49782 12518 49846 12582
rect 44614 12246 44678 12310
rect 47198 12246 47262 12310
rect 49510 12246 49574 12310
rect 52366 12518 52430 12582
rect 54950 12518 55014 12582
rect 57262 12518 57326 12582
rect 52366 12246 52430 12310
rect 54406 12246 54470 12310
rect 59982 12518 60046 12582
rect 62430 12518 62494 12582
rect 64878 12518 64942 12582
rect 67462 12518 67526 12582
rect 69910 12518 69974 12582
rect 72494 12518 72558 12582
rect 74942 12518 75006 12582
rect 77254 12518 77318 12582
rect 57534 12246 57598 12310
rect 59574 12246 59638 12310
rect 62430 12246 62494 12310
rect 64878 12246 64942 12310
rect 67462 12246 67526 12310
rect 69910 12246 69974 12310
rect 72494 12246 72558 12310
rect 74670 12246 74734 12310
rect 76982 12246 77046 12310
rect 79974 12518 80038 12582
rect 82422 12518 82486 12582
rect 84734 12518 84798 12582
rect 79974 12246 80038 12310
rect 82422 12246 82486 12310
rect 84734 12246 84798 12310
rect 87454 12518 87518 12582
rect 89902 12518 89966 12582
rect 92214 12518 92278 12582
rect 87046 12246 87110 12310
rect 89630 12246 89694 12310
rect 94934 12518 94998 12582
rect 97382 12518 97446 12582
rect 99694 12518 99758 12582
rect 92486 12246 92550 12310
rect 94934 12246 94998 12310
rect 97382 12246 97446 12310
rect 99694 12246 99758 12310
rect 102414 12518 102478 12582
rect 104862 12518 104926 12582
rect 107446 12518 107510 12582
rect 102006 12246 102070 12310
rect 104454 12246 104518 12310
rect 107446 12246 107510 12310
rect 1230 12110 1294 12174
rect 15102 11974 15166 12038
rect 29926 11974 29990 12038
rect 32374 11974 32438 12038
rect 34686 11974 34750 12038
rect 29654 11838 29718 11902
rect 32102 11838 32166 11902
rect 34686 11838 34750 11902
rect 37270 11974 37334 12038
rect 37270 11838 37334 11902
rect 39718 11974 39782 12038
rect 39718 11838 39782 11902
rect 42438 11974 42502 12038
rect 44886 11974 44950 12038
rect 47334 11974 47398 12038
rect 49646 11974 49710 12038
rect 42302 11838 42366 11902
rect 44750 11838 44814 11902
rect 47062 11838 47126 11902
rect 49782 11838 49846 11902
rect 52230 11974 52294 12038
rect 52230 11838 52294 11902
rect 54814 11974 54878 12038
rect 57398 11974 57462 12038
rect 59846 11974 59910 12038
rect 62294 11974 62358 12038
rect 64742 11974 64806 12038
rect 54814 11838 54878 11902
rect 57262 11838 57326 11902
rect 59710 11838 59774 11902
rect 62158 11838 62222 11902
rect 67326 11974 67390 12038
rect 69774 11974 69838 12038
rect 72358 11974 72422 12038
rect 74806 11974 74870 12038
rect 77118 11974 77182 12038
rect 64742 11838 64806 11902
rect 67190 11838 67254 11902
rect 69774 11838 69838 11902
rect 72222 11838 72286 11902
rect 74534 11838 74598 11902
rect 77254 11838 77318 11902
rect 79838 11974 79902 12038
rect 82286 11974 82350 12038
rect 84870 11974 84934 12038
rect 87318 11974 87382 12038
rect 89766 11974 89830 12038
rect 92350 11974 92414 12038
rect 94798 11974 94862 12038
rect 97246 11974 97310 12038
rect 99830 11974 99894 12038
rect 102278 11974 102342 12038
rect 104726 11974 104790 12038
rect 107310 11974 107374 12038
rect 79702 11838 79766 11902
rect 82150 11838 82214 11902
rect 84598 11838 84662 11902
rect 87182 11838 87246 11902
rect 89494 11838 89558 11902
rect 92214 11838 92278 11902
rect 94662 11838 94726 11902
rect 97110 11838 97174 11902
rect 99558 11838 99622 11902
rect 102142 11838 102206 11902
rect 104590 11838 104654 11902
rect 137502 11974 137566 12038
rect 107174 11838 107238 11902
rect 124446 11838 124510 11902
rect 15102 11702 15166 11766
rect 22174 11702 22238 11766
rect 29790 11702 29854 11766
rect 32238 11702 32302 11766
rect 34822 11702 34886 11766
rect 37406 11702 37470 11766
rect 39854 11702 39918 11766
rect 42166 11702 42230 11766
rect 44614 11702 44678 11766
rect 47198 11702 47262 11766
rect 49510 11702 49574 11766
rect 52366 11702 52430 11766
rect 57534 11702 57598 11766
rect 59574 11702 59638 11766
rect 62430 11702 62494 11766
rect 64878 11702 64942 11766
rect 67462 11702 67526 11766
rect 69910 11702 69974 11766
rect 72494 11702 72558 11766
rect 74670 11702 74734 11766
rect 76982 11702 77046 11766
rect 79974 11702 80038 11766
rect 82422 11702 82486 11766
rect 84734 11702 84798 11766
rect 87046 11702 87110 11766
rect 29246 11294 29310 11358
rect 54406 11430 54470 11494
rect 89630 11702 89694 11766
rect 92486 11702 92550 11766
rect 94934 11702 94998 11766
rect 97382 11702 97446 11766
rect 99694 11702 99758 11766
rect 102006 11702 102070 11766
rect 104454 11702 104518 11766
rect 107446 11702 107510 11766
rect 124174 11430 124238 11494
rect 109350 11294 109414 11358
rect 124174 11294 124238 11358
rect 29518 11022 29582 11086
rect 29654 11022 29718 11086
rect 32102 11022 32166 11086
rect 34686 11022 34750 11086
rect 37270 11022 37334 11086
rect 39718 11022 39782 11086
rect 42302 11022 42366 11086
rect 44750 11022 44814 11086
rect 47062 11022 47126 11086
rect 49782 11022 49846 11086
rect 52230 11022 52294 11086
rect 54814 11022 54878 11086
rect 57262 11022 57326 11086
rect 59710 11022 59774 11086
rect 62158 11022 62222 11086
rect 64742 11022 64806 11086
rect 67190 11022 67254 11086
rect 69774 11022 69838 11086
rect 72222 11022 72286 11086
rect 74534 11022 74598 11086
rect 77254 11022 77318 11086
rect 79702 11022 79766 11086
rect 82150 11022 82214 11086
rect 84598 11022 84662 11086
rect 87182 11022 87246 11086
rect 89494 11022 89558 11086
rect 92214 11022 92278 11086
rect 94662 11022 94726 11086
rect 97110 11022 97174 11086
rect 99558 11022 99622 11086
rect 102142 11022 102206 11086
rect 104590 11022 104654 11086
rect 107174 11022 107238 11086
rect 109214 11022 109278 11086
rect 124582 10770 124614 10814
rect 124614 10770 124646 10814
rect 124582 10750 124646 10770
rect 29518 10614 29582 10678
rect 109214 10614 109278 10678
rect 1230 10342 1294 10406
rect 15238 10478 15302 10542
rect 15238 10342 15302 10406
rect 137502 10478 137566 10542
rect 550 10206 614 10270
rect 124310 9934 124374 9998
rect 29246 9526 29310 9590
rect 109350 9526 109414 9590
rect 15102 9118 15166 9182
rect 16870 8982 16934 9046
rect 124718 8982 124782 9046
rect 1230 8846 1294 8910
rect 137502 8710 137566 8774
rect 124174 8574 124238 8638
rect 550 7622 614 7686
rect 15238 7622 15302 7686
rect 1230 6942 1294 7006
rect 137502 7078 137566 7142
rect 1230 5446 1294 5510
rect 137502 5446 137566 5510
rect 1230 3814 1294 3878
rect 16870 3814 16934 3878
rect 36726 3678 36790 3742
rect 137502 3814 137566 3878
rect 16598 2862 16662 2926
rect 17686 2862 17750 2926
rect 18774 2862 18838 2926
rect 20134 2862 20198 2926
rect 21086 2862 21150 2926
rect 22310 2862 22374 2926
rect 23670 2862 23734 2926
rect 24758 2862 24822 2926
rect 25982 2862 26046 2926
rect 27070 2862 27134 2926
rect 28158 2862 28222 2926
rect 29246 2862 29310 2926
rect 30606 2862 30670 2926
rect 31830 2862 31894 2926
rect 32918 2862 32982 2926
rect 34006 2862 34070 2926
rect 35094 2862 35158 2926
rect 36454 2862 36518 2926
rect 37542 2862 37606 2926
rect 38630 2862 38694 2926
rect 39990 2862 40054 2926
rect 41214 2862 41278 2926
rect 42302 2862 42366 2926
rect 43390 2862 43454 2926
rect 44478 2862 44542 2926
rect 45838 2862 45902 2926
rect 46926 2862 46990 2926
rect 48150 2862 48214 2926
rect 49238 2862 49302 2926
rect 50326 2862 50390 2926
rect 51686 2862 51750 2926
rect 52774 2862 52838 2926
rect 53862 2862 53926 2926
rect 54950 2862 55014 2926
rect 56310 2862 56374 2926
rect 57534 2862 57598 2926
rect 58622 2862 58686 2926
rect 59710 2862 59774 2926
rect 19318 2318 19382 2382
rect 2046 1638 2110 1702
rect 3814 1696 3870 1702
rect 3870 1696 3878 1702
rect 3814 1638 3878 1696
rect 5446 1696 5494 1702
rect 5494 1696 5510 1702
rect 5446 1638 5510 1696
rect 7214 1696 7230 1702
rect 7230 1696 7278 1702
rect 7214 1638 7278 1696
rect 8710 1638 8774 1702
rect 10478 1696 10534 1702
rect 10534 1696 10542 1702
rect 10478 1638 10542 1696
rect 12110 1638 12174 1702
rect 13878 1696 13894 1702
rect 13894 1696 13942 1702
rect 13878 1638 13942 1696
rect 15646 1638 15710 1702
rect 17142 1638 17206 1702
rect 19046 1638 19110 1702
rect 20542 1638 20606 1702
rect 22174 1638 22238 1702
rect 23942 1696 23974 1702
rect 23974 1696 24006 1702
rect 23942 1638 24006 1696
rect 25710 1638 25774 1702
rect 27206 1638 27270 1702
rect 28838 1638 28902 1702
rect 30470 1638 30534 1702
rect 32238 1638 32302 1702
rect 36726 1774 36790 1838
rect 34278 1638 34342 1702
rect 35638 1638 35702 1702
rect 37270 1638 37334 1702
rect 39038 1696 39094 1702
rect 39094 1696 39102 1702
rect 39038 1638 39102 1696
rect 40670 1638 40734 1702
rect 42438 1696 42454 1702
rect 42454 1696 42502 1702
rect 42438 1638 42502 1696
rect 44070 1638 44134 1702
rect 45702 1638 45766 1702
rect 47470 1696 47494 1702
rect 47494 1696 47534 1702
rect 47470 1638 47534 1696
rect 48966 1638 49030 1702
rect 50734 1638 50798 1702
rect 52502 1696 52534 1702
rect 52534 1696 52566 1702
rect 52502 1638 52566 1696
rect 54134 1638 54198 1702
rect 55902 1696 55950 1702
rect 55950 1696 55966 1702
rect 55902 1638 55966 1696
rect 57398 1638 57462 1702
rect 59166 1638 59230 1702
rect 60934 1696 60990 1702
rect 60990 1696 60998 1702
rect 60934 1638 60998 1696
rect 62702 1638 62766 1702
rect 64198 1638 64262 1702
rect 65830 1638 65894 1702
rect 67598 1696 67654 1702
rect 67654 1696 67662 1702
rect 67598 1638 67662 1696
rect 69230 1638 69294 1702
rect 71134 1638 71198 1702
rect 72630 1638 72694 1702
rect 74262 1638 74326 1702
rect 76030 1696 76054 1702
rect 76054 1696 76094 1702
rect 76030 1638 76094 1696
rect 77662 1638 77726 1702
rect 79294 1638 79358 1702
rect 81198 1638 81262 1702
rect 82694 1638 82758 1702
rect 84598 1638 84662 1702
rect 86094 1696 86134 1702
rect 86134 1696 86158 1702
rect 86094 1638 86158 1696
rect 87726 1638 87790 1702
rect 89358 1638 89422 1702
rect 91126 1696 91174 1702
rect 91174 1696 91190 1702
rect 91126 1638 91190 1696
rect 92894 1696 92910 1702
rect 92910 1696 92958 1702
rect 92894 1638 92958 1696
rect 94662 1638 94726 1702
rect 96158 1696 96214 1702
rect 96214 1696 96222 1702
rect 96158 1638 96222 1696
rect 97926 1696 97950 1702
rect 97950 1696 97990 1702
rect 97926 1638 97990 1696
rect 99694 1638 99758 1702
rect 101190 1638 101254 1702
rect 102958 1696 102990 1702
rect 102990 1696 103022 1702
rect 102958 1638 103022 1696
rect 104590 1696 104614 1702
rect 104614 1696 104654 1702
rect 104590 1638 104654 1696
rect 106222 1638 106286 1702
rect 107854 1638 107918 1702
rect 109622 1696 109654 1702
rect 109654 1696 109686 1702
rect 109622 1638 109686 1696
rect 111390 1638 111454 1702
rect 112886 1638 112950 1702
rect 114654 1696 114694 1702
rect 114694 1696 114718 1702
rect 114654 1638 114718 1696
rect 116286 1638 116350 1702
rect 118054 1696 118110 1702
rect 118110 1696 118118 1702
rect 118054 1638 118118 1696
rect 119686 1696 119734 1702
rect 119734 1696 119750 1702
rect 119686 1638 119750 1696
rect 121454 1696 121470 1702
rect 121470 1696 121518 1702
rect 121454 1638 121518 1696
rect 122950 1638 123014 1702
rect 125126 1638 125190 1702
rect 126350 1638 126414 1702
rect 128118 1696 128134 1702
rect 128134 1696 128182 1702
rect 128118 1638 128182 1696
rect 129886 1638 129950 1702
rect 131382 1638 131446 1702
rect 133150 1696 133174 1702
rect 133174 1696 133214 1702
rect 133150 1638 133214 1696
rect 134782 1638 134846 1702
rect 136550 1696 136590 1702
rect 136590 1696 136614 1702
rect 136550 1638 136614 1696
rect 958 1230 1022 1294
rect 1094 1230 1158 1294
rect 1230 1230 1294 1294
rect 2046 1230 2110 1294
rect 3814 1230 3878 1294
rect 5446 1230 5510 1294
rect 7214 1230 7278 1294
rect 8710 1230 8774 1294
rect 10478 1230 10542 1294
rect 12110 1230 12174 1294
rect 13878 1230 13942 1294
rect 15646 1230 15710 1294
rect 17142 1230 17206 1294
rect 19046 1230 19110 1294
rect 20542 1230 20606 1294
rect 22174 1230 22238 1294
rect 23942 1230 24006 1294
rect 25710 1230 25774 1294
rect 27206 1230 27270 1294
rect 28838 1230 28902 1294
rect 30470 1230 30534 1294
rect 32238 1230 32302 1294
rect 34278 1230 34342 1294
rect 35638 1230 35702 1294
rect 37270 1230 37334 1294
rect 39038 1230 39102 1294
rect 40670 1230 40734 1294
rect 42438 1230 42502 1294
rect 44070 1230 44134 1294
rect 45702 1230 45766 1294
rect 47470 1230 47534 1294
rect 48966 1230 49030 1294
rect 50734 1230 50798 1294
rect 52502 1230 52566 1294
rect 54134 1230 54198 1294
rect 55902 1230 55966 1294
rect 57398 1230 57462 1294
rect 59166 1230 59230 1294
rect 60934 1230 60998 1294
rect 62702 1230 62766 1294
rect 64198 1230 64262 1294
rect 65830 1230 65894 1294
rect 67598 1230 67662 1294
rect 69230 1230 69294 1294
rect 71134 1230 71198 1294
rect 72630 1230 72694 1294
rect 74262 1230 74326 1294
rect 76030 1230 76094 1294
rect 77662 1230 77726 1294
rect 79294 1230 79358 1294
rect 81198 1230 81262 1294
rect 82694 1230 82758 1294
rect 84598 1230 84662 1294
rect 86094 1230 86158 1294
rect 87726 1230 87790 1294
rect 89358 1230 89422 1294
rect 91126 1230 91190 1294
rect 92894 1230 92958 1294
rect 94662 1230 94726 1294
rect 96158 1230 96222 1294
rect 97926 1230 97990 1294
rect 99694 1230 99758 1294
rect 101190 1230 101254 1294
rect 102958 1230 103022 1294
rect 104590 1230 104654 1294
rect 106222 1230 106286 1294
rect 107854 1230 107918 1294
rect 109622 1230 109686 1294
rect 111390 1230 111454 1294
rect 112886 1230 112950 1294
rect 114654 1230 114718 1294
rect 116286 1230 116350 1294
rect 118054 1230 118118 1294
rect 119686 1230 119750 1294
rect 121454 1230 121518 1294
rect 122950 1230 123014 1294
rect 125126 1230 125190 1294
rect 126350 1230 126414 1294
rect 128118 1230 128182 1294
rect 129886 1230 129950 1294
rect 131382 1230 131446 1294
rect 133150 1230 133214 1294
rect 134782 1230 134846 1294
rect 136550 1230 136614 1294
rect 137502 1230 137566 1294
rect 137638 1230 137702 1294
rect 137774 1230 137838 1294
rect 958 1094 1022 1158
rect 1094 1094 1158 1158
rect 1230 1094 1294 1158
rect 137502 1094 137566 1158
rect 137638 1094 137702 1158
rect 137774 1094 137838 1158
rect 958 958 1022 1022
rect 1094 958 1158 1022
rect 1230 958 1294 1022
rect 137502 958 137566 1022
rect 137638 958 137702 1022
rect 137774 958 137838 1022
rect 278 550 342 614
rect 414 550 478 614
rect 550 550 614 614
rect 19318 550 19382 614
rect 138182 550 138246 614
rect 138318 550 138382 614
rect 138454 550 138518 614
rect 278 414 342 478
rect 414 414 478 478
rect 550 414 614 478
rect 138182 414 138246 478
rect 138318 414 138382 478
rect 138454 414 138518 478
rect 278 278 342 342
rect 414 278 478 342
rect 550 278 614 342
rect 138182 278 138246 342
rect 138318 278 138382 342
rect 138454 278 138518 342
<< metal4 >>
rect 272 133486 620 133492
rect 272 133422 278 133486
rect 342 133422 414 133486
rect 478 133422 550 133486
rect 614 133422 620 133486
rect 272 133350 620 133422
rect 272 133286 278 133350
rect 342 133286 414 133350
rect 478 133286 550 133350
rect 614 133286 620 133350
rect 272 133214 620 133286
rect 272 133150 278 133214
rect 342 133150 414 133214
rect 478 133150 550 133214
rect 614 133150 620 133214
rect 272 25910 620 133150
rect 272 25846 550 25910
rect 614 25846 620 25910
rect 272 20334 620 25846
rect 272 20270 550 20334
rect 614 20270 620 20334
rect 272 14758 620 20270
rect 272 14694 550 14758
rect 614 14694 620 14758
rect 272 10270 620 14694
rect 272 10206 550 10270
rect 614 10206 620 10270
rect 272 7686 620 10206
rect 272 7622 550 7686
rect 614 7622 620 7686
rect 272 614 620 7622
rect 952 132806 1300 132812
rect 952 132742 958 132806
rect 1022 132742 1094 132806
rect 1158 132742 1230 132806
rect 1294 132742 1300 132806
rect 952 132670 1300 132742
rect 952 132606 958 132670
rect 1022 132606 1094 132670
rect 1158 132606 1230 132670
rect 1294 132606 1300 132670
rect 952 132534 1300 132606
rect 952 132470 958 132534
rect 1022 132470 1094 132534
rect 1158 132470 1230 132534
rect 1294 132470 1300 132534
rect 952 129814 1300 132470
rect 2176 132534 2252 132540
rect 2176 132470 2182 132534
rect 2246 132470 2252 132534
rect 2176 132126 2252 132470
rect 2176 132094 2182 132126
rect 2181 132062 2182 132094
rect 2246 132094 2252 132126
rect 3672 132534 3748 132540
rect 3672 132470 3678 132534
rect 3742 132470 3748 132534
rect 3672 132126 3748 132470
rect 3672 132094 3678 132126
rect 2246 132062 2247 132094
rect 2181 132061 2247 132062
rect 3677 132062 3678 132094
rect 3742 132094 3748 132126
rect 5440 132534 5516 132540
rect 5440 132470 5446 132534
rect 5510 132470 5516 132534
rect 5440 132126 5516 132470
rect 5440 132094 5446 132126
rect 3742 132062 3743 132094
rect 3677 132061 3743 132062
rect 5445 132062 5446 132094
rect 5510 132094 5516 132126
rect 7208 132534 7284 132540
rect 7208 132470 7214 132534
rect 7278 132470 7284 132534
rect 7208 132126 7284 132470
rect 7208 132094 7214 132126
rect 5510 132062 5511 132094
rect 5445 132061 5511 132062
rect 7213 132062 7214 132094
rect 7278 132094 7284 132126
rect 8976 132534 9052 132540
rect 8976 132470 8982 132534
rect 9046 132470 9052 132534
rect 8976 132126 9052 132470
rect 8976 132094 8982 132126
rect 7278 132062 7279 132094
rect 7213 132061 7279 132062
rect 8981 132062 8982 132094
rect 9046 132094 9052 132126
rect 10472 132534 10548 132540
rect 10472 132470 10478 132534
rect 10542 132470 10548 132534
rect 10472 132126 10548 132470
rect 10472 132094 10478 132126
rect 9046 132062 9047 132094
rect 8981 132061 9047 132062
rect 10477 132062 10478 132094
rect 10542 132094 10548 132126
rect 12104 132534 12180 132540
rect 12104 132470 12110 132534
rect 12174 132470 12180 132534
rect 12104 132126 12180 132470
rect 12104 132094 12110 132126
rect 10542 132062 10543 132094
rect 10477 132061 10543 132062
rect 12109 132062 12110 132094
rect 12174 132094 12180 132126
rect 13872 132534 13948 132540
rect 13872 132470 13878 132534
rect 13942 132470 13948 132534
rect 13872 132126 13948 132470
rect 13872 132094 13878 132126
rect 12174 132062 12175 132094
rect 12109 132061 12175 132062
rect 13877 132062 13878 132094
rect 13942 132094 13948 132126
rect 15640 132534 15716 132540
rect 15640 132470 15646 132534
rect 15710 132470 15716 132534
rect 15640 132126 15716 132470
rect 15640 132094 15646 132126
rect 13942 132062 13943 132094
rect 13877 132061 13943 132062
rect 15645 132062 15646 132094
rect 15710 132094 15716 132126
rect 17136 132534 17212 132540
rect 17136 132470 17142 132534
rect 17206 132470 17212 132534
rect 17136 132126 17212 132470
rect 17136 132094 17142 132126
rect 15710 132062 15711 132094
rect 15645 132061 15711 132062
rect 17141 132062 17142 132094
rect 17206 132094 17212 132126
rect 18904 132534 18980 132540
rect 18904 132470 18910 132534
rect 18974 132470 18980 132534
rect 18904 132126 18980 132470
rect 18904 132094 18910 132126
rect 17206 132062 17207 132094
rect 17141 132061 17207 132062
rect 18909 132062 18910 132094
rect 18974 132094 18980 132126
rect 20672 132534 20748 132540
rect 20672 132470 20678 132534
rect 20742 132470 20748 132534
rect 20672 132126 20748 132470
rect 20672 132094 20678 132126
rect 18974 132062 18975 132094
rect 18909 132061 18975 132062
rect 20677 132062 20678 132094
rect 20742 132094 20748 132126
rect 22168 132534 22244 132540
rect 22168 132470 22174 132534
rect 22238 132470 22244 132534
rect 22168 132126 22244 132470
rect 22168 132094 22174 132126
rect 20742 132062 20743 132094
rect 20677 132061 20743 132062
rect 22173 132062 22174 132094
rect 22238 132094 22244 132126
rect 23936 132534 24012 132540
rect 23936 132470 23942 132534
rect 24006 132470 24012 132534
rect 23936 132126 24012 132470
rect 23936 132094 23942 132126
rect 22238 132062 22239 132094
rect 22173 132061 22239 132062
rect 23941 132062 23942 132094
rect 24006 132094 24012 132126
rect 25704 132534 25780 132540
rect 25704 132470 25710 132534
rect 25774 132470 25780 132534
rect 25704 132126 25780 132470
rect 25704 132094 25710 132126
rect 24006 132062 24007 132094
rect 23941 132061 24007 132062
rect 25709 132062 25710 132094
rect 25774 132094 25780 132126
rect 27200 132534 27276 132540
rect 27200 132470 27206 132534
rect 27270 132470 27276 132534
rect 27200 132126 27276 132470
rect 27200 132094 27206 132126
rect 25774 132062 25775 132094
rect 25709 132061 25775 132062
rect 27205 132062 27206 132094
rect 27270 132094 27276 132126
rect 28968 132534 29044 132540
rect 28968 132470 28974 132534
rect 29038 132470 29044 132534
rect 28968 132126 29044 132470
rect 28968 132094 28974 132126
rect 27270 132062 27271 132094
rect 27205 132061 27271 132062
rect 28973 132062 28974 132094
rect 29038 132094 29044 132126
rect 29038 132062 29039 132094
rect 28973 132061 29039 132062
rect 2040 131990 2116 131996
rect 2040 131926 2046 131990
rect 2110 131926 2116 131990
rect 2040 131582 2116 131926
rect 2040 131550 2046 131582
rect 2045 131518 2046 131550
rect 2110 131550 2116 131582
rect 2110 131518 2111 131550
rect 2045 131517 2111 131518
rect 952 129750 1230 129814
rect 1294 129750 1300 129814
rect 952 128182 1300 129750
rect 952 128118 1230 128182
rect 1294 128118 1300 128182
rect 952 126414 1300 128118
rect 29648 127638 29724 133764
rect 30736 132534 30812 132540
rect 30736 132470 30742 132534
rect 30806 132470 30812 132534
rect 30736 132126 30812 132470
rect 30736 132094 30742 132126
rect 30741 132062 30742 132094
rect 30806 132094 30812 132126
rect 30806 132062 30807 132094
rect 30741 132061 30807 132062
rect 29648 127606 29654 127638
rect 29653 127574 29654 127606
rect 29718 127606 29724 127638
rect 31960 127638 32036 133764
rect 32232 132534 32308 132540
rect 32232 132470 32238 132534
rect 32302 132470 32308 132534
rect 32232 132126 32308 132470
rect 32232 132094 32238 132126
rect 32237 132062 32238 132094
rect 32302 132094 32308 132126
rect 34136 132534 34212 132540
rect 34136 132470 34142 132534
rect 34206 132470 34212 132534
rect 34136 132126 34212 132470
rect 34136 132094 34142 132126
rect 32302 132062 32303 132094
rect 32237 132061 32303 132062
rect 34141 132062 34142 132094
rect 34206 132094 34212 132126
rect 34206 132062 34207 132094
rect 34141 132061 34207 132062
rect 31960 127606 31966 127638
rect 29718 127574 29719 127606
rect 29653 127573 29719 127574
rect 31965 127574 31966 127606
rect 32030 127606 32036 127638
rect 34544 127638 34620 133764
rect 35632 132534 35708 132540
rect 35632 132470 35638 132534
rect 35702 132470 35708 132534
rect 35632 132126 35708 132470
rect 35632 132094 35638 132126
rect 35637 132062 35638 132094
rect 35702 132094 35708 132126
rect 35702 132062 35703 132094
rect 35637 132061 35703 132062
rect 34544 127606 34550 127638
rect 32030 127574 32031 127606
rect 31965 127573 32031 127574
rect 34549 127574 34550 127606
rect 34614 127606 34620 127638
rect 36992 127638 37068 133764
rect 37400 132534 37476 132540
rect 37400 132470 37406 132534
rect 37470 132470 37476 132534
rect 37400 132126 37476 132470
rect 37400 132094 37406 132126
rect 37405 132062 37406 132094
rect 37470 132094 37476 132126
rect 39168 132534 39244 132540
rect 39168 132470 39174 132534
rect 39238 132470 39244 132534
rect 39168 132126 39244 132470
rect 39168 132094 39174 132126
rect 37470 132062 37471 132094
rect 37405 132061 37471 132062
rect 39173 132062 39174 132094
rect 39238 132094 39244 132126
rect 39238 132062 39239 132094
rect 39173 132061 39239 132062
rect 36992 127606 36998 127638
rect 34614 127574 34615 127606
rect 34549 127573 34615 127574
rect 36997 127574 36998 127606
rect 37062 127606 37068 127638
rect 39576 127638 39652 133764
rect 40664 132534 40740 132540
rect 40664 132470 40670 132534
rect 40734 132470 40740 132534
rect 40664 132126 40740 132470
rect 40664 132094 40670 132126
rect 40669 132062 40670 132094
rect 40734 132094 40740 132126
rect 40734 132062 40735 132094
rect 40669 132061 40735 132062
rect 39576 127606 39582 127638
rect 37062 127574 37063 127606
rect 36997 127573 37063 127574
rect 39581 127574 39582 127606
rect 39646 127606 39652 127638
rect 42024 127638 42100 133764
rect 42432 132534 42508 132540
rect 42432 132470 42438 132534
rect 42502 132470 42508 132534
rect 42432 132126 42508 132470
rect 42432 132094 42438 132126
rect 42437 132062 42438 132094
rect 42502 132094 42508 132126
rect 44200 132534 44276 132540
rect 44200 132470 44206 132534
rect 44270 132470 44276 132534
rect 44200 132126 44276 132470
rect 44200 132094 44206 132126
rect 42502 132062 42503 132094
rect 42437 132061 42503 132062
rect 44205 132062 44206 132094
rect 44270 132094 44276 132126
rect 44270 132062 44271 132094
rect 44205 132061 44271 132062
rect 42024 127606 42030 127638
rect 39646 127574 39647 127606
rect 39581 127573 39647 127574
rect 42029 127574 42030 127606
rect 42094 127606 42100 127638
rect 44608 127638 44684 133764
rect 45696 132534 45772 132540
rect 45696 132470 45702 132534
rect 45766 132470 45772 132534
rect 45696 132126 45772 132470
rect 45696 132094 45702 132126
rect 45701 132062 45702 132094
rect 45766 132094 45772 132126
rect 45766 132062 45767 132094
rect 45701 132061 45767 132062
rect 44608 127606 44614 127638
rect 42094 127574 42095 127606
rect 42029 127573 42095 127574
rect 44613 127574 44614 127606
rect 44678 127606 44684 127638
rect 47056 127638 47132 133764
rect 47464 132534 47540 132540
rect 47464 132470 47470 132534
rect 47534 132470 47540 132534
rect 47464 132126 47540 132470
rect 47464 132094 47470 132126
rect 47469 132062 47470 132094
rect 47534 132094 47540 132126
rect 49096 132534 49172 132540
rect 49096 132470 49102 132534
rect 49166 132470 49172 132534
rect 49096 132126 49172 132470
rect 49096 132094 49102 132126
rect 47534 132062 47535 132094
rect 47469 132061 47535 132062
rect 49101 132062 49102 132094
rect 49166 132094 49172 132126
rect 49166 132062 49167 132094
rect 49101 132061 49167 132062
rect 47056 127606 47062 127638
rect 44678 127574 44679 127606
rect 44613 127573 44679 127574
rect 47061 127574 47062 127606
rect 47126 127606 47132 127638
rect 49504 127638 49580 133764
rect 50728 132534 50804 132540
rect 50728 132470 50734 132534
rect 50798 132470 50804 132534
rect 50728 132126 50804 132470
rect 50728 132094 50734 132126
rect 50733 132062 50734 132094
rect 50798 132094 50804 132126
rect 50798 132062 50799 132094
rect 50733 132061 50799 132062
rect 49504 127606 49510 127638
rect 47126 127574 47127 127606
rect 47061 127573 47127 127574
rect 49509 127574 49510 127606
rect 49574 127606 49580 127638
rect 51952 127638 52028 133764
rect 52632 132534 52708 132540
rect 52632 132470 52638 132534
rect 52702 132470 52708 132534
rect 52632 132126 52708 132470
rect 52632 132094 52638 132126
rect 52637 132062 52638 132094
rect 52702 132094 52708 132126
rect 54128 132534 54204 132540
rect 54128 132470 54134 132534
rect 54198 132470 54204 132534
rect 54128 132126 54204 132470
rect 54128 132094 54134 132126
rect 52702 132062 52703 132094
rect 52637 132061 52703 132062
rect 54133 132062 54134 132094
rect 54198 132094 54204 132126
rect 54198 132062 54199 132094
rect 54133 132061 54199 132062
rect 51952 127606 51958 127638
rect 49574 127574 49575 127606
rect 49509 127573 49575 127574
rect 51957 127574 51958 127606
rect 52022 127606 52028 127638
rect 54400 127638 54476 133764
rect 55896 132534 55972 132540
rect 55896 132470 55902 132534
rect 55966 132470 55972 132534
rect 55896 132126 55972 132470
rect 55896 132094 55902 132126
rect 55901 132062 55902 132094
rect 55966 132094 55972 132126
rect 55966 132062 55967 132094
rect 55901 132061 55967 132062
rect 54400 127606 54406 127638
rect 52022 127574 52023 127606
rect 51957 127573 52023 127574
rect 54405 127574 54406 127606
rect 54470 127606 54476 127638
rect 56984 127638 57060 133764
rect 57664 132534 57740 132540
rect 57664 132470 57670 132534
rect 57734 132470 57740 132534
rect 57664 132126 57740 132470
rect 57664 132094 57670 132126
rect 57669 132062 57670 132094
rect 57734 132094 57740 132126
rect 59160 132534 59236 132540
rect 59160 132470 59166 132534
rect 59230 132470 59236 132534
rect 59160 132126 59236 132470
rect 59160 132094 59166 132126
rect 57734 132062 57735 132094
rect 57669 132061 57735 132062
rect 59165 132062 59166 132094
rect 59230 132094 59236 132126
rect 59230 132062 59231 132094
rect 59165 132061 59231 132062
rect 56984 127606 56990 127638
rect 54470 127574 54471 127606
rect 54405 127573 54471 127574
rect 56989 127574 56990 127606
rect 57054 127606 57060 127638
rect 59568 127638 59644 133764
rect 61064 132534 61140 132540
rect 61064 132470 61070 132534
rect 61134 132470 61140 132534
rect 61064 132126 61140 132470
rect 61064 132094 61070 132126
rect 61069 132062 61070 132094
rect 61134 132094 61140 132126
rect 61134 132062 61135 132094
rect 61069 132061 61135 132062
rect 59568 127606 59574 127638
rect 57054 127574 57055 127606
rect 56989 127573 57055 127574
rect 59573 127574 59574 127606
rect 59638 127606 59644 127638
rect 62016 127638 62092 133764
rect 62696 132534 62772 132540
rect 62696 132470 62702 132534
rect 62766 132470 62772 132534
rect 62696 132126 62772 132470
rect 62696 132094 62702 132126
rect 62701 132062 62702 132094
rect 62766 132094 62772 132126
rect 64192 132534 64268 132540
rect 64192 132470 64198 132534
rect 64262 132470 64268 132534
rect 64192 132126 64268 132470
rect 64192 132094 64198 132126
rect 62766 132062 62767 132094
rect 62701 132061 62767 132062
rect 64197 132062 64198 132094
rect 64262 132094 64268 132126
rect 64262 132062 64263 132094
rect 64197 132061 64263 132062
rect 62016 127606 62022 127638
rect 59638 127574 59639 127606
rect 59573 127573 59639 127574
rect 62021 127574 62022 127606
rect 62086 127606 62092 127638
rect 64600 127638 64676 133764
rect 66096 132534 66172 132540
rect 66096 132470 66102 132534
rect 66166 132470 66172 132534
rect 66096 132126 66172 132470
rect 66096 132094 66102 132126
rect 66101 132062 66102 132094
rect 66166 132094 66172 132126
rect 66166 132062 66167 132094
rect 66101 132061 66167 132062
rect 64600 127606 64606 127638
rect 62086 127574 62087 127606
rect 62021 127573 62087 127574
rect 64605 127574 64606 127606
rect 64670 127606 64676 127638
rect 67048 127638 67124 133764
rect 67728 132534 67804 132540
rect 67728 132470 67734 132534
rect 67798 132470 67804 132534
rect 67728 132126 67804 132470
rect 67728 132094 67734 132126
rect 67733 132062 67734 132094
rect 67798 132094 67804 132126
rect 69224 132534 69300 132540
rect 69224 132470 69230 132534
rect 69294 132470 69300 132534
rect 69224 132126 69300 132470
rect 69224 132094 69230 132126
rect 67798 132062 67799 132094
rect 67733 132061 67799 132062
rect 69229 132062 69230 132094
rect 69294 132094 69300 132126
rect 69294 132062 69295 132094
rect 69229 132061 69295 132062
rect 67048 127606 67054 127638
rect 64670 127574 64671 127606
rect 64605 127573 64671 127574
rect 67053 127574 67054 127606
rect 67118 127606 67124 127638
rect 69360 127638 69436 133764
rect 71128 132534 71204 132540
rect 71128 132470 71134 132534
rect 71198 132470 71204 132534
rect 71128 132126 71204 132470
rect 71128 132094 71134 132126
rect 71133 132062 71134 132094
rect 71198 132094 71204 132126
rect 71198 132062 71199 132094
rect 71133 132061 71199 132062
rect 69360 127606 69366 127638
rect 67118 127574 67119 127606
rect 67053 127573 67119 127574
rect 69365 127574 69366 127606
rect 69430 127606 69436 127638
rect 72080 127638 72156 133764
rect 72624 132534 72700 132540
rect 72624 132470 72630 132534
rect 72694 132470 72700 132534
rect 72624 132126 72700 132470
rect 72624 132094 72630 132126
rect 72629 132062 72630 132094
rect 72694 132094 72700 132126
rect 74256 132534 74332 132540
rect 74256 132470 74262 132534
rect 74326 132470 74332 132534
rect 74256 132126 74332 132470
rect 74256 132094 74262 132126
rect 72694 132062 72695 132094
rect 72629 132061 72695 132062
rect 74261 132062 74262 132094
rect 74326 132094 74332 132126
rect 74326 132062 74327 132094
rect 74261 132061 74327 132062
rect 72080 127606 72086 127638
rect 69430 127574 69431 127606
rect 69365 127573 69431 127574
rect 72085 127574 72086 127606
rect 72150 127606 72156 127638
rect 74392 127638 74468 133764
rect 76160 132534 76236 132540
rect 76160 132470 76166 132534
rect 76230 132470 76236 132534
rect 76160 132126 76236 132470
rect 76160 132094 76166 132126
rect 76165 132062 76166 132094
rect 76230 132094 76236 132126
rect 76230 132062 76231 132094
rect 76165 132061 76231 132062
rect 74392 127606 74398 127638
rect 72150 127574 72151 127606
rect 72085 127573 72151 127574
rect 74397 127574 74398 127606
rect 74462 127606 74468 127638
rect 76976 127638 77052 133764
rect 77656 132534 77732 132540
rect 77656 132470 77662 132534
rect 77726 132470 77732 132534
rect 77656 132126 77732 132470
rect 77656 132094 77662 132126
rect 77661 132062 77662 132094
rect 77726 132094 77732 132126
rect 79288 132534 79364 132540
rect 79288 132470 79294 132534
rect 79358 132470 79364 132534
rect 79288 132126 79364 132470
rect 79288 132094 79294 132126
rect 77726 132062 77727 132094
rect 77661 132061 77727 132062
rect 79293 132062 79294 132094
rect 79358 132094 79364 132126
rect 79358 132062 79359 132094
rect 79293 132061 79359 132062
rect 76976 127606 76982 127638
rect 74462 127574 74463 127606
rect 74397 127573 74463 127574
rect 76981 127574 76982 127606
rect 77046 127606 77052 127638
rect 79424 127638 79500 133764
rect 81192 132534 81268 132540
rect 81192 132470 81198 132534
rect 81262 132470 81268 132534
rect 81192 132126 81268 132470
rect 81192 132094 81198 132126
rect 81197 132062 81198 132094
rect 81262 132094 81268 132126
rect 81262 132062 81263 132094
rect 81197 132061 81263 132062
rect 79424 127606 79430 127638
rect 77046 127574 77047 127606
rect 76981 127573 77047 127574
rect 79429 127574 79430 127606
rect 79494 127606 79500 127638
rect 82008 127638 82084 133764
rect 82688 132534 82764 132540
rect 82688 132470 82694 132534
rect 82758 132470 82764 132534
rect 82688 132126 82764 132470
rect 82688 132094 82694 132126
rect 82693 132062 82694 132094
rect 82758 132094 82764 132126
rect 84320 132534 84396 132540
rect 84320 132470 84326 132534
rect 84390 132470 84396 132534
rect 84320 132126 84396 132470
rect 84320 132094 84326 132126
rect 82758 132062 82759 132094
rect 82693 132061 82759 132062
rect 84325 132062 84326 132094
rect 84390 132094 84396 132126
rect 84390 132062 84391 132094
rect 84325 132061 84391 132062
rect 82008 127606 82014 127638
rect 79494 127574 79495 127606
rect 79429 127573 79495 127574
rect 82013 127574 82014 127606
rect 82078 127606 82084 127638
rect 84456 127638 84532 133764
rect 86088 132534 86164 132540
rect 86088 132470 86094 132534
rect 86158 132470 86164 132534
rect 86088 132126 86164 132470
rect 86088 132094 86094 132126
rect 86093 132062 86094 132094
rect 86158 132094 86164 132126
rect 86158 132062 86159 132094
rect 86093 132061 86159 132062
rect 84456 127606 84462 127638
rect 82078 127574 82079 127606
rect 82013 127573 82079 127574
rect 84461 127574 84462 127606
rect 84526 127606 84532 127638
rect 87040 127638 87116 133764
rect 87720 132534 87796 132540
rect 87720 132470 87726 132534
rect 87790 132470 87796 132534
rect 87720 132126 87796 132470
rect 87720 132094 87726 132126
rect 87725 132062 87726 132094
rect 87790 132094 87796 132126
rect 87790 132062 87791 132094
rect 87725 132061 87791 132062
rect 87040 127606 87046 127638
rect 84526 127574 84527 127606
rect 84461 127573 84527 127574
rect 87045 127574 87046 127606
rect 87110 127606 87116 127638
rect 89488 127638 89564 133764
rect 89760 132534 89836 132540
rect 89760 132470 89766 132534
rect 89830 132470 89836 132534
rect 89760 132126 89836 132470
rect 89760 132094 89766 132126
rect 89765 132062 89766 132094
rect 89830 132094 89836 132126
rect 91120 132534 91196 132540
rect 91120 132470 91126 132534
rect 91190 132470 91196 132534
rect 91120 132126 91196 132470
rect 91120 132094 91126 132126
rect 89830 132062 89831 132094
rect 89765 132061 89831 132062
rect 91125 132062 91126 132094
rect 91190 132094 91196 132126
rect 91190 132062 91191 132094
rect 91125 132061 91191 132062
rect 89488 127606 89494 127638
rect 87110 127574 87111 127606
rect 87045 127573 87111 127574
rect 89493 127574 89494 127606
rect 89558 127606 89564 127638
rect 91936 127638 92012 133764
rect 92888 132534 92964 132540
rect 92888 132470 92894 132534
rect 92958 132470 92964 132534
rect 92888 132126 92964 132470
rect 92888 132094 92894 132126
rect 92893 132062 92894 132094
rect 92958 132094 92964 132126
rect 92958 132062 92959 132094
rect 92893 132061 92959 132062
rect 91936 127606 91942 127638
rect 89558 127574 89559 127606
rect 89493 127573 89559 127574
rect 91941 127574 91942 127606
rect 92006 127606 92012 127638
rect 94384 127638 94460 133764
rect 94656 132534 94732 132540
rect 94656 132470 94662 132534
rect 94726 132470 94732 132534
rect 94656 132126 94732 132470
rect 94656 132094 94662 132126
rect 94661 132062 94662 132094
rect 94726 132094 94732 132126
rect 96152 132534 96228 132540
rect 96152 132470 96158 132534
rect 96222 132470 96228 132534
rect 96152 132126 96228 132470
rect 96152 132094 96158 132126
rect 94726 132062 94727 132094
rect 94661 132061 94727 132062
rect 96157 132062 96158 132094
rect 96222 132094 96228 132126
rect 96222 132062 96223 132094
rect 96157 132061 96223 132062
rect 94384 127606 94390 127638
rect 92006 127574 92007 127606
rect 91941 127573 92007 127574
rect 94389 127574 94390 127606
rect 94454 127606 94460 127638
rect 96832 127638 96908 133764
rect 97920 132534 97996 132540
rect 97920 132470 97926 132534
rect 97990 132470 97996 132534
rect 97920 132126 97996 132470
rect 97920 132094 97926 132126
rect 97925 132062 97926 132094
rect 97990 132094 97996 132126
rect 97990 132062 97991 132094
rect 97925 132061 97991 132062
rect 96832 127606 96838 127638
rect 94454 127574 94455 127606
rect 94389 127573 94455 127574
rect 96837 127574 96838 127606
rect 96902 127606 96908 127638
rect 99416 127638 99492 133764
rect 99688 132534 99764 132540
rect 99688 132470 99694 132534
rect 99758 132470 99764 132534
rect 99688 132126 99764 132470
rect 99688 132094 99694 132126
rect 99693 132062 99694 132094
rect 99758 132094 99764 132126
rect 101184 132534 101260 132540
rect 101184 132470 101190 132534
rect 101254 132470 101260 132534
rect 101184 132126 101260 132470
rect 101184 132094 101190 132126
rect 99758 132062 99759 132094
rect 99693 132061 99759 132062
rect 101189 132062 101190 132094
rect 101254 132094 101260 132126
rect 101254 132062 101255 132094
rect 101189 132061 101255 132062
rect 99416 127606 99422 127638
rect 96902 127574 96903 127606
rect 96837 127573 96903 127574
rect 99421 127574 99422 127606
rect 99486 127606 99492 127638
rect 102000 127638 102076 133764
rect 102952 132534 103028 132540
rect 102952 132470 102958 132534
rect 103022 132470 103028 132534
rect 102952 132126 103028 132470
rect 102952 132094 102958 132126
rect 102957 132062 102958 132094
rect 103022 132094 103028 132126
rect 103022 132062 103023 132094
rect 102957 132061 103023 132062
rect 102000 127606 102006 127638
rect 99486 127574 99487 127606
rect 99421 127573 99487 127574
rect 102005 127574 102006 127606
rect 102070 127606 102076 127638
rect 104448 127638 104524 133764
rect 104720 132534 104796 132540
rect 104720 132470 104726 132534
rect 104790 132470 104796 132534
rect 104720 132126 104796 132470
rect 104720 132094 104726 132126
rect 104725 132062 104726 132094
rect 104790 132094 104796 132126
rect 106216 132534 106292 132540
rect 106216 132470 106222 132534
rect 106286 132470 106292 132534
rect 106216 132126 106292 132470
rect 106216 132094 106222 132126
rect 104790 132062 104791 132094
rect 104725 132061 104791 132062
rect 106221 132062 106222 132094
rect 106286 132094 106292 132126
rect 106286 132062 106287 132094
rect 106221 132061 106287 132062
rect 104448 127606 104454 127638
rect 102070 127574 102071 127606
rect 102005 127573 102071 127574
rect 104453 127574 104454 127606
rect 104518 127606 104524 127638
rect 107032 127638 107108 133764
rect 107848 132534 107924 132540
rect 107848 132470 107854 132534
rect 107918 132470 107924 132534
rect 107848 132126 107924 132470
rect 107848 132094 107854 132126
rect 107853 132062 107854 132094
rect 107918 132094 107924 132126
rect 109616 132534 109692 132540
rect 109616 132470 109622 132534
rect 109686 132470 109692 132534
rect 109616 132126 109692 132470
rect 109616 132094 109622 132126
rect 107918 132062 107919 132094
rect 107853 132061 107919 132062
rect 109621 132062 109622 132094
rect 109686 132094 109692 132126
rect 111384 132534 111460 132540
rect 111384 132470 111390 132534
rect 111454 132470 111460 132534
rect 111384 132126 111460 132470
rect 111384 132094 111390 132126
rect 109686 132062 109687 132094
rect 109621 132061 109687 132062
rect 111389 132062 111390 132094
rect 111454 132094 111460 132126
rect 112880 132534 112956 132540
rect 112880 132470 112886 132534
rect 112950 132470 112956 132534
rect 112880 132126 112956 132470
rect 112880 132094 112886 132126
rect 111454 132062 111455 132094
rect 111389 132061 111455 132062
rect 112885 132062 112886 132094
rect 112950 132094 112956 132126
rect 114648 132534 114724 132540
rect 114648 132470 114654 132534
rect 114718 132470 114724 132534
rect 114648 132126 114724 132470
rect 114648 132094 114654 132126
rect 112950 132062 112951 132094
rect 112885 132061 112951 132062
rect 114653 132062 114654 132094
rect 114718 132094 114724 132126
rect 116416 132534 116492 132540
rect 116416 132470 116422 132534
rect 116486 132470 116492 132534
rect 116416 132126 116492 132470
rect 116416 132094 116422 132126
rect 114718 132062 114719 132094
rect 114653 132061 114719 132062
rect 116421 132062 116422 132094
rect 116486 132094 116492 132126
rect 117912 132534 117988 132540
rect 117912 132470 117918 132534
rect 117982 132470 117988 132534
rect 117912 132126 117988 132470
rect 117912 132094 117918 132126
rect 116486 132062 116487 132094
rect 116421 132061 116487 132062
rect 117917 132062 117918 132094
rect 117982 132094 117988 132126
rect 119680 132534 119756 132540
rect 119680 132470 119686 132534
rect 119750 132470 119756 132534
rect 119680 132126 119756 132470
rect 119680 132094 119686 132126
rect 117982 132062 117983 132094
rect 117917 132061 117983 132062
rect 119685 132062 119686 132094
rect 119750 132094 119756 132126
rect 119750 132062 119751 132094
rect 119685 132061 119751 132062
rect 119680 131990 119756 131996
rect 119680 131926 119686 131990
rect 119750 131926 119756 131990
rect 119544 131310 119620 131316
rect 119544 131246 119550 131310
rect 119614 131246 119620 131310
rect 119408 129950 119484 129956
rect 119408 129886 119414 129950
rect 119478 129886 119484 129950
rect 117509 129134 117575 129135
rect 117509 129102 117510 129134
rect 117504 129070 117510 129102
rect 117574 129102 117575 129134
rect 117574 129070 117580 129102
rect 107032 127606 107038 127638
rect 104518 127574 104519 127606
rect 104453 127573 104519 127574
rect 107037 127574 107038 127606
rect 107102 127606 107108 127638
rect 117368 127774 117444 127780
rect 117368 127710 117374 127774
rect 117438 127710 117444 127774
rect 107102 127574 107103 127606
rect 107037 127573 107103 127574
rect 29925 127502 29991 127503
rect 29925 127470 29926 127502
rect 29920 127438 29926 127470
rect 29990 127470 29991 127502
rect 32509 127502 32575 127503
rect 32509 127470 32510 127502
rect 29990 127438 29996 127470
rect 29784 127230 29860 127236
rect 29784 127166 29790 127230
rect 29854 127166 29860 127230
rect 29784 126550 29860 127166
rect 29784 126518 29790 126550
rect 29789 126486 29790 126518
rect 29854 126518 29860 126550
rect 29854 126486 29855 126518
rect 29789 126485 29855 126486
rect 952 126350 1230 126414
rect 1294 126350 1300 126414
rect 952 124646 1300 126350
rect 29920 125734 29996 127438
rect 32504 127438 32510 127470
rect 32574 127470 32575 127502
rect 34957 127502 35023 127503
rect 34957 127470 34958 127502
rect 32574 127438 32580 127470
rect 32101 127230 32167 127231
rect 32101 127198 32102 127230
rect 32096 127166 32102 127198
rect 32166 127198 32167 127230
rect 32368 127230 32444 127236
rect 32166 127166 32172 127198
rect 32096 126550 32172 127166
rect 32096 126486 32102 126550
rect 32166 126486 32172 126550
rect 32368 127166 32374 127230
rect 32438 127166 32444 127230
rect 32368 126550 32444 127166
rect 32368 126518 32374 126550
rect 32096 126480 32172 126486
rect 32373 126486 32374 126518
rect 32438 126518 32444 126550
rect 32438 126486 32439 126518
rect 32373 126485 32439 126486
rect 29920 125670 29926 125734
rect 29990 125670 29996 125734
rect 30061 125734 30127 125735
rect 30061 125702 30062 125734
rect 29920 125664 29996 125670
rect 30056 125670 30062 125702
rect 30126 125702 30127 125734
rect 32504 125734 32580 127438
rect 34952 127438 34958 127470
rect 35022 127470 35023 127502
rect 37269 127502 37335 127503
rect 37269 127470 37270 127502
rect 35022 127438 35028 127470
rect 34816 127230 34892 127236
rect 34816 127166 34822 127230
rect 34886 127166 34892 127230
rect 34816 126550 34892 127166
rect 34816 126518 34822 126550
rect 34821 126486 34822 126518
rect 34886 126518 34892 126550
rect 34886 126486 34887 126518
rect 34821 126485 34887 126486
rect 30126 125670 30132 125702
rect 952 124582 1230 124646
rect 1294 124582 1300 124646
rect 952 123150 1300 124582
rect 30056 123830 30132 125670
rect 32504 125670 32510 125734
rect 32574 125670 32580 125734
rect 32645 125734 32711 125735
rect 32645 125702 32646 125734
rect 32504 125664 32580 125670
rect 32640 125670 32646 125702
rect 32710 125702 32711 125734
rect 34952 125734 35028 127438
rect 37264 127438 37270 127470
rect 37334 127470 37335 127502
rect 39989 127502 40055 127503
rect 39989 127470 39990 127502
rect 37334 127438 37340 127470
rect 37128 127230 37204 127236
rect 37128 127166 37134 127230
rect 37198 127166 37204 127230
rect 37128 126550 37204 127166
rect 37128 126518 37134 126550
rect 37133 126486 37134 126518
rect 37198 126518 37204 126550
rect 37198 126486 37199 126518
rect 37133 126485 37199 126486
rect 32710 125670 32716 125702
rect 30056 123766 30062 123830
rect 30126 123766 30132 123830
rect 30056 123760 30132 123766
rect 32640 123830 32716 125670
rect 34952 125670 34958 125734
rect 35022 125670 35028 125734
rect 35093 125734 35159 125735
rect 35093 125702 35094 125734
rect 34952 125664 35028 125670
rect 35088 125670 35094 125702
rect 35158 125702 35159 125734
rect 37264 125734 37340 127438
rect 39984 127438 39990 127470
rect 40054 127470 40055 127502
rect 42437 127502 42503 127503
rect 42437 127470 42438 127502
rect 40054 127438 40060 127470
rect 37400 127230 37476 127236
rect 37400 127166 37406 127230
rect 37470 127166 37476 127230
rect 37400 126550 37476 127166
rect 37400 126518 37406 126550
rect 37405 126486 37406 126518
rect 37470 126518 37476 126550
rect 39848 127230 39924 127236
rect 39848 127166 39854 127230
rect 39918 127166 39924 127230
rect 39848 126550 39924 127166
rect 39848 126518 39854 126550
rect 37470 126486 37471 126518
rect 37405 126485 37471 126486
rect 39853 126486 39854 126518
rect 39918 126518 39924 126550
rect 39918 126486 39919 126518
rect 39853 126485 39919 126486
rect 35158 125670 35164 125702
rect 32640 123766 32646 123830
rect 32710 123766 32716 123830
rect 32640 123760 32716 123766
rect 35088 123830 35164 125670
rect 37264 125670 37270 125734
rect 37334 125670 37340 125734
rect 37405 125734 37471 125735
rect 37405 125702 37406 125734
rect 37264 125664 37340 125670
rect 37400 125670 37406 125702
rect 37470 125702 37471 125734
rect 39984 125734 40060 127438
rect 42432 127438 42438 127470
rect 42502 127470 42503 127502
rect 44885 127502 44951 127503
rect 44885 127470 44886 127502
rect 42502 127438 42508 127470
rect 42160 127230 42236 127236
rect 42160 127166 42166 127230
rect 42230 127166 42236 127230
rect 42160 126550 42236 127166
rect 42160 126518 42166 126550
rect 42165 126486 42166 126518
rect 42230 126518 42236 126550
rect 42230 126486 42231 126518
rect 42165 126485 42231 126486
rect 37470 125670 37476 125702
rect 35088 123766 35094 123830
rect 35158 123766 35164 123830
rect 35088 123760 35164 123766
rect 37400 123830 37476 125670
rect 39984 125670 39990 125734
rect 40054 125670 40060 125734
rect 40125 125734 40191 125735
rect 40125 125702 40126 125734
rect 39984 125664 40060 125670
rect 40120 125670 40126 125702
rect 40190 125702 40191 125734
rect 42432 125734 42508 127438
rect 44880 127438 44886 127470
rect 44950 127470 44951 127502
rect 47333 127502 47399 127503
rect 47333 127470 47334 127502
rect 44950 127438 44956 127470
rect 44880 127372 44956 127438
rect 44744 127296 44956 127372
rect 47328 127438 47334 127470
rect 47398 127470 47399 127502
rect 49917 127502 49983 127503
rect 49917 127470 49918 127502
rect 47398 127438 47404 127470
rect 40190 125670 40196 125702
rect 37400 123766 37406 123830
rect 37470 123766 37476 123830
rect 37400 123760 37476 123766
rect 40120 123830 40196 125670
rect 42432 125670 42438 125734
rect 42502 125670 42508 125734
rect 42573 125734 42639 125735
rect 42573 125702 42574 125734
rect 42432 125664 42508 125670
rect 42568 125670 42574 125702
rect 42638 125702 42639 125734
rect 44744 125734 44820 127296
rect 44880 127230 44956 127236
rect 44880 127166 44886 127230
rect 44950 127166 44956 127230
rect 44880 126550 44956 127166
rect 44880 126518 44886 126550
rect 44885 126486 44886 126518
rect 44950 126518 44956 126550
rect 47192 127230 47268 127236
rect 47192 127166 47198 127230
rect 47262 127166 47268 127230
rect 47192 126550 47268 127166
rect 47192 126518 47198 126550
rect 44950 126486 44951 126518
rect 44885 126485 44951 126486
rect 47197 126486 47198 126518
rect 47262 126518 47268 126550
rect 47262 126486 47263 126518
rect 47197 126485 47263 126486
rect 42638 125670 42644 125702
rect 40120 123766 40126 123830
rect 40190 123766 40196 123830
rect 40120 123760 40196 123766
rect 42568 123830 42644 125670
rect 44744 125670 44750 125734
rect 44814 125670 44820 125734
rect 44885 125734 44951 125735
rect 44885 125702 44886 125734
rect 44744 125664 44820 125670
rect 44880 125670 44886 125702
rect 44950 125702 44951 125734
rect 47328 125734 47404 127438
rect 49912 127438 49918 127470
rect 49982 127470 49983 127502
rect 52365 127502 52431 127503
rect 52365 127470 52366 127502
rect 49982 127438 49988 127470
rect 49509 127230 49575 127231
rect 49509 127198 49510 127230
rect 49504 127166 49510 127198
rect 49574 127198 49575 127230
rect 49776 127230 49852 127236
rect 49574 127166 49580 127198
rect 49504 126550 49580 127166
rect 49504 126486 49510 126550
rect 49574 126486 49580 126550
rect 49776 127166 49782 127230
rect 49846 127166 49852 127230
rect 49776 126550 49852 127166
rect 49776 126518 49782 126550
rect 49504 126480 49580 126486
rect 49781 126486 49782 126518
rect 49846 126518 49852 126550
rect 49846 126486 49847 126518
rect 49781 126485 49847 126486
rect 44950 125670 44956 125702
rect 42568 123766 42574 123830
rect 42638 123766 42644 123830
rect 42568 123760 42644 123766
rect 44880 123830 44956 125670
rect 47328 125670 47334 125734
rect 47398 125670 47404 125734
rect 47469 125734 47535 125735
rect 47469 125702 47470 125734
rect 47328 125664 47404 125670
rect 47464 125670 47470 125702
rect 47534 125702 47535 125734
rect 49912 125734 49988 127438
rect 52360 127438 52366 127470
rect 52430 127470 52431 127502
rect 54949 127502 55015 127503
rect 54949 127470 54950 127502
rect 52430 127438 52436 127470
rect 52224 127230 52300 127236
rect 52224 127166 52230 127230
rect 52294 127166 52300 127230
rect 52224 126550 52300 127166
rect 52224 126518 52230 126550
rect 52229 126486 52230 126518
rect 52294 126518 52300 126550
rect 52294 126486 52295 126518
rect 52229 126485 52295 126486
rect 47534 125670 47540 125702
rect 44880 123766 44886 123830
rect 44950 123766 44956 123830
rect 44880 123760 44956 123766
rect 47464 123830 47540 125670
rect 49912 125670 49918 125734
rect 49982 125670 49988 125734
rect 50053 125734 50119 125735
rect 50053 125702 50054 125734
rect 49912 125664 49988 125670
rect 50048 125670 50054 125702
rect 50118 125702 50119 125734
rect 52360 125734 52436 127438
rect 54944 127438 54950 127470
rect 55014 127470 55015 127502
rect 57397 127502 57463 127503
rect 57397 127470 57398 127502
rect 55014 127438 55020 127470
rect 54808 127230 54884 127236
rect 54808 127166 54814 127230
rect 54878 127166 54884 127230
rect 54808 126550 54884 127166
rect 54808 126518 54814 126550
rect 54813 126486 54814 126518
rect 54878 126518 54884 126550
rect 54878 126486 54879 126518
rect 54813 126485 54879 126486
rect 50118 125670 50124 125702
rect 47464 123766 47470 123830
rect 47534 123766 47540 123830
rect 47464 123760 47540 123766
rect 50048 123830 50124 125670
rect 52360 125670 52366 125734
rect 52430 125670 52436 125734
rect 52501 125734 52567 125735
rect 52501 125702 52502 125734
rect 52360 125664 52436 125670
rect 52496 125670 52502 125702
rect 52566 125702 52567 125734
rect 54944 125734 55020 127438
rect 57392 127438 57398 127470
rect 57462 127470 57463 127502
rect 59845 127502 59911 127503
rect 59845 127470 59846 127502
rect 57462 127438 57468 127470
rect 56984 127230 57060 127236
rect 56984 127166 56990 127230
rect 57054 127166 57060 127230
rect 56984 126550 57060 127166
rect 56984 126518 56990 126550
rect 56989 126486 56990 126518
rect 57054 126518 57060 126550
rect 57256 127230 57332 127236
rect 57256 127166 57262 127230
rect 57326 127166 57332 127230
rect 57256 126550 57332 127166
rect 57256 126518 57262 126550
rect 57054 126486 57055 126518
rect 56989 126485 57055 126486
rect 57261 126486 57262 126518
rect 57326 126518 57332 126550
rect 57326 126486 57327 126518
rect 57261 126485 57327 126486
rect 52566 125670 52572 125702
rect 50048 123766 50054 123830
rect 50118 123766 50124 123830
rect 50048 123760 50124 123766
rect 52496 123830 52572 125670
rect 54944 125670 54950 125734
rect 55014 125670 55020 125734
rect 55085 125734 55151 125735
rect 55085 125702 55086 125734
rect 54944 125664 55020 125670
rect 55080 125670 55086 125702
rect 55150 125702 55151 125734
rect 57392 125734 57468 127438
rect 59840 127438 59846 127470
rect 59910 127470 59911 127502
rect 62429 127502 62495 127503
rect 62429 127470 62430 127502
rect 59910 127438 59916 127470
rect 59840 127372 59916 127438
rect 59704 127296 59916 127372
rect 62424 127438 62430 127470
rect 62494 127470 62495 127502
rect 64741 127502 64807 127503
rect 64741 127470 64742 127502
rect 62494 127438 62500 127470
rect 59568 127230 59644 127236
rect 59568 127166 59574 127230
rect 59638 127166 59644 127230
rect 59568 126550 59644 127166
rect 59568 126518 59574 126550
rect 59573 126486 59574 126518
rect 59638 126518 59644 126550
rect 59638 126486 59639 126518
rect 59573 126485 59639 126486
rect 55150 125670 55156 125702
rect 52496 123766 52502 123830
rect 52566 123766 52572 123830
rect 52496 123760 52572 123766
rect 55080 123830 55156 125670
rect 57392 125670 57398 125734
rect 57462 125670 57468 125734
rect 57533 125734 57599 125735
rect 57533 125702 57534 125734
rect 57392 125664 57468 125670
rect 57528 125670 57534 125702
rect 57598 125702 57599 125734
rect 59704 125734 59780 127296
rect 59840 127230 59916 127236
rect 59840 127166 59846 127230
rect 59910 127166 59916 127230
rect 59840 126550 59916 127166
rect 59840 126518 59846 126550
rect 59845 126486 59846 126518
rect 59910 126518 59916 126550
rect 62288 127230 62364 127236
rect 62288 127166 62294 127230
rect 62358 127166 62364 127230
rect 62288 126550 62364 127166
rect 62288 126518 62294 126550
rect 59910 126486 59911 126518
rect 59845 126485 59911 126486
rect 62293 126486 62294 126518
rect 62358 126518 62364 126550
rect 62358 126486 62359 126518
rect 62293 126485 62359 126486
rect 57598 125670 57604 125702
rect 55080 123766 55086 123830
rect 55150 123766 55156 123830
rect 55080 123760 55156 123766
rect 57528 123830 57604 125670
rect 59704 125670 59710 125734
rect 59774 125670 59780 125734
rect 59981 125734 60047 125735
rect 59981 125702 59982 125734
rect 59704 125664 59780 125670
rect 59976 125670 59982 125702
rect 60046 125702 60047 125734
rect 62424 125734 62500 127438
rect 64736 127438 64742 127470
rect 64806 127470 64807 127502
rect 67325 127502 67391 127503
rect 67325 127470 67326 127502
rect 64806 127438 64812 127470
rect 60046 125670 60052 125702
rect 57528 123766 57534 123830
rect 57598 123766 57604 123830
rect 57528 123760 57604 123766
rect 59976 123830 60052 125670
rect 62424 125670 62430 125734
rect 62494 125670 62500 125734
rect 62565 125734 62631 125735
rect 62565 125702 62566 125734
rect 62424 125664 62500 125670
rect 62560 125670 62566 125702
rect 62630 125702 62631 125734
rect 64736 125734 64812 127438
rect 67320 127438 67326 127470
rect 67390 127470 67391 127502
rect 69773 127502 69839 127503
rect 69773 127470 69774 127502
rect 67390 127438 67396 127470
rect 64872 127230 64948 127236
rect 64872 127166 64878 127230
rect 64942 127166 64948 127230
rect 67053 127230 67119 127231
rect 67053 127198 67054 127230
rect 64872 126550 64948 127166
rect 64872 126518 64878 126550
rect 64877 126486 64878 126518
rect 64942 126518 64948 126550
rect 67048 127166 67054 127198
rect 67118 127198 67119 127230
rect 67184 127230 67260 127236
rect 67118 127166 67124 127198
rect 67048 126550 67124 127166
rect 64942 126486 64943 126518
rect 64877 126485 64943 126486
rect 67048 126486 67054 126550
rect 67118 126486 67124 126550
rect 67184 127166 67190 127230
rect 67254 127166 67260 127230
rect 67184 126550 67260 127166
rect 67184 126518 67190 126550
rect 67048 126480 67124 126486
rect 67189 126486 67190 126518
rect 67254 126518 67260 126550
rect 67254 126486 67255 126518
rect 67189 126485 67255 126486
rect 62630 125670 62636 125702
rect 59976 123766 59982 123830
rect 60046 123766 60052 123830
rect 59976 123760 60052 123766
rect 62560 123830 62636 125670
rect 64736 125670 64742 125734
rect 64806 125670 64812 125734
rect 64877 125734 64943 125735
rect 64877 125702 64878 125734
rect 64736 125664 64812 125670
rect 64872 125670 64878 125702
rect 64942 125702 64943 125734
rect 67320 125734 67396 127438
rect 69768 127438 69774 127470
rect 69838 127470 69839 127502
rect 72357 127502 72423 127503
rect 72357 127470 72358 127502
rect 69838 127438 69844 127470
rect 69632 127230 69708 127236
rect 69632 127166 69638 127230
rect 69702 127166 69708 127230
rect 69632 126550 69708 127166
rect 69632 126518 69638 126550
rect 69637 126486 69638 126518
rect 69702 126518 69708 126550
rect 69702 126486 69703 126518
rect 69637 126485 69703 126486
rect 64942 125670 64948 125702
rect 62560 123766 62566 123830
rect 62630 123766 62636 123830
rect 62560 123760 62636 123766
rect 64872 123830 64948 125670
rect 67320 125670 67326 125734
rect 67390 125670 67396 125734
rect 67461 125734 67527 125735
rect 67461 125702 67462 125734
rect 67320 125664 67396 125670
rect 67456 125670 67462 125702
rect 67526 125702 67527 125734
rect 69768 125734 69844 127438
rect 72352 127438 72358 127470
rect 72422 127470 72423 127502
rect 74941 127502 75007 127503
rect 74941 127470 74942 127502
rect 72422 127438 72428 127470
rect 72216 127230 72292 127236
rect 72216 127166 72222 127230
rect 72286 127166 72292 127230
rect 72216 126550 72292 127166
rect 72216 126518 72222 126550
rect 72221 126486 72222 126518
rect 72286 126518 72292 126550
rect 72286 126486 72287 126518
rect 72221 126485 72287 126486
rect 67526 125670 67532 125702
rect 64872 123766 64878 123830
rect 64942 123766 64948 123830
rect 64872 123760 64948 123766
rect 67456 123830 67532 125670
rect 69768 125670 69774 125734
rect 69838 125670 69844 125734
rect 69909 125734 69975 125735
rect 69909 125702 69910 125734
rect 69768 125664 69844 125670
rect 69904 125670 69910 125702
rect 69974 125702 69975 125734
rect 72352 125734 72428 127438
rect 74936 127438 74942 127470
rect 75006 127470 75007 127502
rect 77389 127502 77455 127503
rect 77389 127470 77390 127502
rect 75006 127438 75012 127470
rect 74533 127230 74599 127231
rect 74533 127198 74534 127230
rect 74528 127166 74534 127198
rect 74598 127198 74599 127230
rect 74800 127230 74876 127236
rect 74598 127166 74604 127198
rect 74528 126550 74604 127166
rect 74528 126486 74534 126550
rect 74598 126486 74604 126550
rect 74800 127166 74806 127230
rect 74870 127166 74876 127230
rect 74800 126550 74876 127166
rect 74800 126518 74806 126550
rect 74528 126480 74604 126486
rect 74805 126486 74806 126518
rect 74870 126518 74876 126550
rect 74870 126486 74871 126518
rect 74805 126485 74871 126486
rect 69974 125670 69980 125702
rect 67456 123766 67462 123830
rect 67526 123766 67532 123830
rect 67456 123760 67532 123766
rect 69904 123830 69980 125670
rect 72352 125670 72358 125734
rect 72422 125670 72428 125734
rect 72493 125734 72559 125735
rect 72493 125702 72494 125734
rect 72352 125664 72428 125670
rect 72488 125670 72494 125702
rect 72558 125702 72559 125734
rect 74936 125734 75012 127438
rect 77384 127438 77390 127470
rect 77454 127470 77455 127502
rect 79837 127502 79903 127503
rect 79837 127470 79838 127502
rect 77454 127438 77460 127470
rect 77248 127230 77324 127236
rect 77248 127166 77254 127230
rect 77318 127166 77324 127230
rect 77248 126550 77324 127166
rect 77248 126518 77254 126550
rect 77253 126486 77254 126518
rect 77318 126518 77324 126550
rect 77318 126486 77319 126518
rect 77253 126485 77319 126486
rect 72558 125670 72564 125702
rect 69904 123766 69910 123830
rect 69974 123766 69980 123830
rect 69904 123760 69980 123766
rect 72488 123830 72564 125670
rect 74936 125670 74942 125734
rect 75006 125670 75012 125734
rect 75077 125734 75143 125735
rect 75077 125702 75078 125734
rect 74936 125664 75012 125670
rect 75072 125670 75078 125702
rect 75142 125702 75143 125734
rect 77384 125734 77460 127438
rect 79832 127438 79838 127470
rect 79902 127470 79903 127502
rect 82421 127502 82487 127503
rect 82421 127470 82422 127502
rect 79902 127438 79908 127470
rect 79832 127372 79908 127438
rect 79696 127296 79908 127372
rect 82416 127438 82422 127470
rect 82486 127470 82487 127502
rect 84869 127502 84935 127503
rect 84869 127470 84870 127502
rect 82486 127438 82492 127470
rect 79560 127230 79636 127236
rect 79560 127166 79566 127230
rect 79630 127166 79636 127230
rect 79560 126550 79636 127166
rect 79560 126518 79566 126550
rect 79565 126486 79566 126518
rect 79630 126518 79636 126550
rect 79630 126486 79631 126518
rect 79565 126485 79631 126486
rect 75142 125670 75148 125702
rect 72488 123766 72494 123830
rect 72558 123766 72564 123830
rect 72488 123760 72564 123766
rect 75072 123830 75148 125670
rect 77384 125670 77390 125734
rect 77454 125670 77460 125734
rect 77525 125734 77591 125735
rect 77525 125702 77526 125734
rect 77384 125664 77460 125670
rect 77520 125670 77526 125702
rect 77590 125702 77591 125734
rect 79696 125734 79772 127296
rect 79832 127230 79908 127236
rect 79832 127166 79838 127230
rect 79902 127166 79908 127230
rect 79832 126550 79908 127166
rect 79832 126518 79838 126550
rect 79837 126486 79838 126518
rect 79902 126518 79908 126550
rect 82008 127230 82084 127236
rect 82008 127166 82014 127230
rect 82078 127166 82084 127230
rect 82008 126550 82084 127166
rect 82008 126518 82014 126550
rect 79902 126486 79903 126518
rect 79837 126485 79903 126486
rect 82013 126486 82014 126518
rect 82078 126518 82084 126550
rect 82280 127230 82356 127236
rect 82280 127166 82286 127230
rect 82350 127166 82356 127230
rect 82280 126550 82356 127166
rect 82280 126518 82286 126550
rect 82078 126486 82079 126518
rect 82013 126485 82079 126486
rect 82285 126486 82286 126518
rect 82350 126518 82356 126550
rect 82350 126486 82351 126518
rect 82285 126485 82351 126486
rect 77590 125670 77596 125702
rect 75072 123766 75078 123830
rect 75142 123766 75148 123830
rect 75072 123760 75148 123766
rect 77520 123830 77596 125670
rect 79696 125670 79702 125734
rect 79766 125670 79772 125734
rect 79837 125734 79903 125735
rect 79837 125702 79838 125734
rect 79696 125664 79772 125670
rect 79832 125670 79838 125702
rect 79902 125702 79903 125734
rect 82416 125734 82492 127438
rect 84864 127438 84870 127470
rect 84934 127470 84935 127502
rect 87317 127502 87383 127503
rect 87317 127470 87318 127502
rect 84934 127438 84940 127470
rect 84456 127230 84532 127236
rect 84456 127166 84462 127230
rect 84526 127166 84532 127230
rect 84456 126550 84532 127166
rect 84456 126518 84462 126550
rect 84461 126486 84462 126518
rect 84526 126518 84532 126550
rect 84592 127230 84668 127236
rect 84592 127166 84598 127230
rect 84662 127166 84668 127230
rect 84592 126550 84668 127166
rect 84592 126518 84598 126550
rect 84526 126486 84527 126518
rect 84461 126485 84527 126486
rect 84597 126486 84598 126518
rect 84662 126518 84668 126550
rect 84662 126486 84663 126518
rect 84597 126485 84663 126486
rect 79902 125670 79908 125702
rect 77520 123766 77526 123830
rect 77590 123766 77596 123830
rect 77520 123760 77596 123766
rect 79832 123830 79908 125670
rect 82416 125670 82422 125734
rect 82486 125670 82492 125734
rect 82557 125734 82623 125735
rect 82557 125702 82558 125734
rect 82416 125664 82492 125670
rect 82552 125670 82558 125702
rect 82622 125702 82623 125734
rect 84864 125734 84940 127438
rect 87312 127438 87318 127470
rect 87382 127470 87383 127502
rect 89765 127502 89831 127503
rect 89765 127470 89766 127502
rect 87382 127438 87388 127470
rect 87312 127372 87388 127438
rect 87176 127296 87388 127372
rect 89760 127438 89766 127470
rect 89830 127470 89831 127502
rect 92349 127502 92415 127503
rect 92349 127470 92350 127502
rect 89830 127438 89836 127470
rect 82622 125670 82628 125702
rect 79832 123766 79838 123830
rect 79902 123766 79908 123830
rect 79832 123760 79908 123766
rect 82552 123830 82628 125670
rect 84864 125670 84870 125734
rect 84934 125670 84940 125734
rect 85005 125734 85071 125735
rect 85005 125702 85006 125734
rect 84864 125664 84940 125670
rect 85000 125670 85006 125702
rect 85070 125702 85071 125734
rect 87176 125734 87252 127296
rect 87312 127230 87388 127236
rect 87312 127166 87318 127230
rect 87382 127166 87388 127230
rect 87312 126550 87388 127166
rect 87312 126518 87318 126550
rect 87317 126486 87318 126518
rect 87382 126518 87388 126550
rect 89624 127230 89700 127236
rect 89624 127166 89630 127230
rect 89694 127166 89700 127230
rect 89624 126550 89700 127166
rect 89624 126518 89630 126550
rect 87382 126486 87383 126518
rect 87317 126485 87383 126486
rect 89629 126486 89630 126518
rect 89694 126518 89700 126550
rect 89694 126486 89695 126518
rect 89629 126485 89695 126486
rect 87861 126414 87927 126415
rect 87861 126382 87862 126414
rect 87856 126350 87862 126382
rect 87926 126382 87927 126414
rect 87926 126350 87932 126382
rect 85070 125670 85076 125702
rect 82552 123766 82558 123830
rect 82622 123766 82628 123830
rect 82552 123760 82628 123766
rect 85000 123830 85076 125670
rect 87176 125670 87182 125734
rect 87246 125670 87252 125734
rect 87317 125734 87383 125735
rect 87317 125702 87318 125734
rect 87176 125664 87252 125670
rect 87312 125670 87318 125702
rect 87382 125702 87383 125734
rect 87382 125670 87388 125702
rect 85000 123766 85006 123830
rect 85070 123766 85076 123830
rect 85000 123760 85076 123766
rect 87312 123830 87388 125670
rect 87312 123766 87318 123830
rect 87382 123766 87388 123830
rect 87312 123760 87388 123766
rect 952 123086 1230 123150
rect 1294 123086 1300 123150
rect 952 121518 1300 123086
rect 29920 123558 29996 123564
rect 29920 123494 29926 123558
rect 29990 123494 29996 123558
rect 29653 122062 29719 122063
rect 29653 122030 29654 122062
rect 29648 121998 29654 122030
rect 29718 122030 29719 122062
rect 29718 121998 29724 122030
rect 29648 121654 29724 121998
rect 29648 121590 29654 121654
rect 29718 121590 29724 121654
rect 29648 121584 29724 121590
rect 952 121454 1230 121518
rect 1294 121454 1300 121518
rect 952 119750 1300 121454
rect 29920 121110 29996 123494
rect 87856 122198 87932 126350
rect 89760 125734 89836 127438
rect 92344 127438 92350 127470
rect 92414 127470 92415 127502
rect 94797 127502 94863 127503
rect 94797 127470 94798 127502
rect 92414 127438 92420 127470
rect 92208 127230 92284 127236
rect 92208 127166 92214 127230
rect 92278 127166 92284 127230
rect 92208 126550 92284 127166
rect 92208 126518 92214 126550
rect 92213 126486 92214 126518
rect 92278 126518 92284 126550
rect 92278 126486 92279 126518
rect 92213 126485 92279 126486
rect 89760 125670 89766 125734
rect 89830 125670 89836 125734
rect 89901 125734 89967 125735
rect 89901 125702 89902 125734
rect 89760 125664 89836 125670
rect 89896 125670 89902 125702
rect 89966 125702 89967 125734
rect 92344 125734 92420 127438
rect 94792 127438 94798 127470
rect 94862 127470 94863 127502
rect 97381 127502 97447 127503
rect 97381 127470 97382 127502
rect 94862 127438 94868 127470
rect 94656 127230 94732 127236
rect 94656 127166 94662 127230
rect 94726 127166 94732 127230
rect 94656 126550 94732 127166
rect 94656 126518 94662 126550
rect 94661 126486 94662 126518
rect 94726 126518 94732 126550
rect 94726 126486 94727 126518
rect 94661 126485 94727 126486
rect 89966 125670 89972 125702
rect 89896 123830 89972 125670
rect 92344 125670 92350 125734
rect 92414 125670 92420 125734
rect 92485 125734 92551 125735
rect 92485 125702 92486 125734
rect 92344 125664 92420 125670
rect 92480 125670 92486 125702
rect 92550 125702 92551 125734
rect 94792 125734 94868 127438
rect 97376 127438 97382 127470
rect 97446 127470 97447 127502
rect 99829 127502 99895 127503
rect 99829 127470 99830 127502
rect 97446 127438 97452 127470
rect 97240 127230 97316 127236
rect 97240 127166 97246 127230
rect 97310 127166 97316 127230
rect 97240 126550 97316 127166
rect 97240 126518 97246 126550
rect 97245 126486 97246 126518
rect 97310 126518 97316 126550
rect 97310 126486 97311 126518
rect 97245 126485 97311 126486
rect 92550 125670 92556 125702
rect 89896 123766 89902 123830
rect 89966 123766 89972 123830
rect 89896 123760 89972 123766
rect 92480 123830 92556 125670
rect 94792 125670 94798 125734
rect 94862 125670 94868 125734
rect 94933 125734 94999 125735
rect 94933 125702 94934 125734
rect 94792 125664 94868 125670
rect 94928 125670 94934 125702
rect 94998 125702 94999 125734
rect 97376 125734 97452 127438
rect 99824 127438 99830 127470
rect 99894 127470 99895 127502
rect 102277 127502 102343 127503
rect 102277 127470 102278 127502
rect 99894 127438 99900 127470
rect 99416 127230 99492 127236
rect 99416 127166 99422 127230
rect 99486 127166 99492 127230
rect 99416 126550 99492 127166
rect 99416 126518 99422 126550
rect 99421 126486 99422 126518
rect 99486 126518 99492 126550
rect 99688 127230 99764 127236
rect 99688 127166 99694 127230
rect 99758 127166 99764 127230
rect 99688 126550 99764 127166
rect 99688 126518 99694 126550
rect 99486 126486 99487 126518
rect 99421 126485 99487 126486
rect 99693 126486 99694 126518
rect 99758 126518 99764 126550
rect 99758 126486 99759 126518
rect 99693 126485 99759 126486
rect 94998 125670 95004 125702
rect 92480 123766 92486 123830
rect 92550 123766 92556 123830
rect 92480 123760 92556 123766
rect 94928 123830 95004 125670
rect 97376 125670 97382 125734
rect 97446 125670 97452 125734
rect 97517 125734 97583 125735
rect 97517 125702 97518 125734
rect 97376 125664 97452 125670
rect 97512 125670 97518 125702
rect 97582 125702 97583 125734
rect 99824 125734 99900 127438
rect 102272 127438 102278 127470
rect 102342 127470 102343 127502
rect 104861 127502 104927 127503
rect 104861 127470 104862 127502
rect 102342 127438 102348 127470
rect 102272 127372 102348 127438
rect 102136 127296 102348 127372
rect 104856 127438 104862 127470
rect 104926 127470 104927 127502
rect 107309 127502 107375 127503
rect 107309 127470 107310 127502
rect 104926 127438 104932 127470
rect 97582 125670 97588 125702
rect 94928 123766 94934 123830
rect 94998 123766 95004 123830
rect 94928 123760 95004 123766
rect 97512 123830 97588 125670
rect 99824 125670 99830 125734
rect 99894 125670 99900 125734
rect 99965 125734 100031 125735
rect 99965 125702 99966 125734
rect 99824 125664 99900 125670
rect 99960 125670 99966 125702
rect 100030 125702 100031 125734
rect 102136 125734 102212 127296
rect 102272 127230 102348 127236
rect 102272 127166 102278 127230
rect 102342 127166 102348 127230
rect 102272 126550 102348 127166
rect 102272 126518 102278 126550
rect 102277 126486 102278 126518
rect 102342 126518 102348 126550
rect 104720 127230 104796 127236
rect 104720 127166 104726 127230
rect 104790 127166 104796 127230
rect 104720 126550 104796 127166
rect 104720 126518 104726 126550
rect 102342 126486 102343 126518
rect 102277 126485 102343 126486
rect 104725 126486 104726 126518
rect 104790 126518 104796 126550
rect 104790 126486 104791 126518
rect 104725 126485 104791 126486
rect 100030 125670 100036 125702
rect 97512 123766 97518 123830
rect 97582 123766 97588 123830
rect 97512 123760 97588 123766
rect 99960 123830 100036 125670
rect 102136 125670 102142 125734
rect 102206 125670 102212 125734
rect 102413 125734 102479 125735
rect 102413 125702 102414 125734
rect 102136 125664 102212 125670
rect 102408 125670 102414 125702
rect 102478 125702 102479 125734
rect 104856 125734 104932 127438
rect 107304 127438 107310 127470
rect 107374 127470 107375 127502
rect 107374 127438 107380 127470
rect 107168 127230 107244 127236
rect 107168 127166 107174 127230
rect 107238 127166 107244 127230
rect 107168 126550 107244 127166
rect 107168 126518 107174 126550
rect 107173 126486 107174 126518
rect 107238 126518 107244 126550
rect 107238 126486 107239 126518
rect 107173 126485 107239 126486
rect 102478 125670 102484 125702
rect 99960 123766 99966 123830
rect 100030 123766 100036 123830
rect 99960 123760 100036 123766
rect 102408 123830 102484 125670
rect 104856 125670 104862 125734
rect 104926 125670 104932 125734
rect 104997 125734 105063 125735
rect 104997 125702 104998 125734
rect 104856 125664 104932 125670
rect 104992 125670 104998 125702
rect 105062 125702 105063 125734
rect 107304 125734 107380 127438
rect 117237 126278 117303 126279
rect 117237 126246 117238 126278
rect 117232 126214 117238 126246
rect 117302 126246 117303 126278
rect 117302 126214 117308 126246
rect 105062 125670 105068 125702
rect 102408 123766 102414 123830
rect 102478 123766 102484 123830
rect 102408 123760 102484 123766
rect 104992 123830 105068 125670
rect 107304 125670 107310 125734
rect 107374 125670 107380 125734
rect 107445 125734 107511 125735
rect 107445 125702 107446 125734
rect 107304 125664 107380 125670
rect 107440 125670 107446 125702
rect 107510 125702 107511 125734
rect 107510 125670 107516 125702
rect 104992 123766 104998 123830
rect 105062 123766 105068 123830
rect 104992 123760 105068 123766
rect 107440 123830 107516 125670
rect 107440 123766 107446 123830
rect 107510 123766 107516 123830
rect 107440 123760 107516 123766
rect 116280 124918 116356 124924
rect 116280 124854 116286 124918
rect 116350 124854 116356 124918
rect 110165 123558 110231 123559
rect 110165 123526 110166 123558
rect 87856 122134 87862 122198
rect 87926 122134 87932 122198
rect 87856 122128 87932 122134
rect 110160 123494 110166 123526
rect 110230 123526 110231 123558
rect 110230 123494 110236 123526
rect 30333 122062 30399 122063
rect 30333 122030 30334 122062
rect 30328 121998 30334 122030
rect 30398 122030 30399 122062
rect 30464 122062 30540 122068
rect 30398 121998 30404 122030
rect 30328 121654 30404 121998
rect 30328 121590 30334 121654
rect 30398 121590 30404 121654
rect 30464 121998 30470 122062
rect 30534 121998 30540 122062
rect 30464 121654 30540 121998
rect 30464 121622 30470 121654
rect 30328 121584 30404 121590
rect 30469 121590 30470 121622
rect 30534 121622 30540 121654
rect 31688 122062 31764 122068
rect 31688 121998 31694 122062
rect 31758 121998 31764 122062
rect 32781 122062 32847 122063
rect 32781 122030 32782 122062
rect 31688 121654 31764 121998
rect 31688 121622 31694 121654
rect 30534 121590 30535 121622
rect 30469 121589 30535 121590
rect 31693 121590 31694 121622
rect 31758 121622 31764 121654
rect 32776 121998 32782 122030
rect 32846 122030 32847 122062
rect 33461 122062 33527 122063
rect 33461 122030 33462 122062
rect 32846 121998 32852 122030
rect 32776 121654 32852 121998
rect 31758 121590 31759 121622
rect 31693 121589 31759 121590
rect 32776 121590 32782 121654
rect 32846 121590 32852 121654
rect 32776 121584 32852 121590
rect 33456 121998 33462 122030
rect 33526 122030 33527 122062
rect 34136 122062 34212 122068
rect 33526 121998 33532 122030
rect 33456 121654 33532 121998
rect 33456 121590 33462 121654
rect 33526 121590 33532 121654
rect 34136 121998 34142 122062
rect 34206 121998 34212 122062
rect 34685 122062 34751 122063
rect 34685 122030 34686 122062
rect 34136 121654 34212 121998
rect 34136 121622 34142 121654
rect 33456 121584 33532 121590
rect 34141 121590 34142 121622
rect 34206 121622 34212 121654
rect 34680 121998 34686 122030
rect 34750 122030 34751 122062
rect 35360 122062 35436 122068
rect 34750 121998 34756 122030
rect 34680 121654 34756 121998
rect 34206 121590 34207 121622
rect 34141 121589 34207 121590
rect 34680 121590 34686 121654
rect 34750 121590 34756 121654
rect 35360 121998 35366 122062
rect 35430 121998 35436 122062
rect 35909 122062 35975 122063
rect 35909 122030 35910 122062
rect 35360 121654 35436 121998
rect 35360 121622 35366 121654
rect 34680 121584 34756 121590
rect 35365 121590 35366 121622
rect 35430 121622 35436 121654
rect 35904 121998 35910 122030
rect 35974 122030 35975 122062
rect 37133 122062 37199 122063
rect 37133 122030 37134 122062
rect 35974 121998 35980 122030
rect 35904 121654 35980 121998
rect 35430 121590 35431 121622
rect 35365 121589 35431 121590
rect 35904 121590 35910 121654
rect 35974 121590 35980 121654
rect 35904 121584 35980 121590
rect 37128 121998 37134 122030
rect 37198 122030 37199 122062
rect 38493 122062 38559 122063
rect 38493 122030 38494 122062
rect 37198 121998 37204 122030
rect 37128 121654 37204 121998
rect 37128 121590 37134 121654
rect 37198 121590 37204 121654
rect 37128 121584 37204 121590
rect 38488 121998 38494 122030
rect 38558 122030 38559 122062
rect 39168 122062 39244 122068
rect 38558 121998 38564 122030
rect 38488 121654 38564 121998
rect 38488 121590 38494 121654
rect 38558 121590 38564 121654
rect 39168 121998 39174 122062
rect 39238 121998 39244 122062
rect 39581 122062 39647 122063
rect 39581 122030 39582 122062
rect 39168 121654 39244 121998
rect 39168 121622 39174 121654
rect 38488 121584 38564 121590
rect 39173 121590 39174 121622
rect 39238 121622 39244 121654
rect 39576 121998 39582 122030
rect 39646 122030 39647 122062
rect 40392 122062 40468 122068
rect 39646 121998 39652 122030
rect 39576 121654 39652 121998
rect 39238 121590 39239 121622
rect 39173 121589 39239 121590
rect 39576 121590 39582 121654
rect 39646 121590 39652 121654
rect 40392 121998 40398 122062
rect 40462 121998 40468 122062
rect 40941 122062 41007 122063
rect 40941 122030 40942 122062
rect 40392 121654 40468 121998
rect 40392 121622 40398 121654
rect 39576 121584 39652 121590
rect 40397 121590 40398 121622
rect 40462 121622 40468 121654
rect 40936 121998 40942 122030
rect 41006 122030 41007 122062
rect 42165 122062 42231 122063
rect 42165 122030 42166 122062
rect 41006 121998 41012 122030
rect 40936 121654 41012 121998
rect 40462 121590 40463 121622
rect 40397 121589 40463 121590
rect 40936 121590 40942 121654
rect 41006 121590 41012 121654
rect 40936 121584 41012 121590
rect 42160 121998 42166 122030
rect 42230 122030 42231 122062
rect 42840 122062 42916 122068
rect 42230 121998 42236 122030
rect 42160 121654 42236 121998
rect 42160 121590 42166 121654
rect 42230 121590 42236 121654
rect 42840 121998 42846 122062
rect 42910 121998 42916 122062
rect 43389 122062 43455 122063
rect 43389 122030 43390 122062
rect 42840 121654 42916 121998
rect 42840 121622 42846 121654
rect 42160 121584 42236 121590
rect 42845 121590 42846 121622
rect 42910 121622 42916 121654
rect 43384 121998 43390 122030
rect 43454 122030 43455 122062
rect 43928 122062 44004 122068
rect 43454 121998 43460 122030
rect 43384 121654 43460 121998
rect 42910 121590 42911 121622
rect 42845 121589 42911 121590
rect 43384 121590 43390 121654
rect 43454 121590 43460 121654
rect 43928 121998 43934 122062
rect 43998 121998 44004 122062
rect 43928 121654 44004 121998
rect 43928 121622 43934 121654
rect 43384 121584 43460 121590
rect 43933 121590 43934 121622
rect 43998 121622 44004 121654
rect 44064 122062 44140 122068
rect 44064 121998 44070 122062
rect 44134 121998 44140 122062
rect 44613 122062 44679 122063
rect 44613 122030 44614 122062
rect 44064 121654 44140 121998
rect 44064 121622 44070 121654
rect 43998 121590 43999 121622
rect 43933 121589 43999 121590
rect 44069 121590 44070 121622
rect 44134 121622 44140 121654
rect 44608 121998 44614 122030
rect 44678 122030 44679 122062
rect 45696 122062 45772 122068
rect 44678 121998 44684 122030
rect 44608 121654 44684 121998
rect 44134 121590 44135 121622
rect 44069 121589 44135 121590
rect 44608 121590 44614 121654
rect 44678 121590 44684 121654
rect 45696 121998 45702 122062
rect 45766 121998 45772 122062
rect 45696 121654 45772 121998
rect 45696 121622 45702 121654
rect 44608 121584 44684 121590
rect 45701 121590 45702 121622
rect 45766 121622 45772 121654
rect 46648 122062 46724 122068
rect 46648 121998 46654 122062
rect 46718 121998 46724 122062
rect 46648 121654 46724 121998
rect 46648 121622 46654 121654
rect 45766 121590 45767 121622
rect 45701 121589 45767 121590
rect 46653 121590 46654 121622
rect 46718 121622 46724 121654
rect 47872 122062 47948 122068
rect 47872 121998 47878 122062
rect 47942 121998 47948 122062
rect 48421 122062 48487 122063
rect 48421 122030 48422 122062
rect 47872 121654 47948 121998
rect 47872 121622 47878 121654
rect 46718 121590 46719 121622
rect 46653 121589 46719 121590
rect 47877 121590 47878 121622
rect 47942 121622 47948 121654
rect 48416 121998 48422 122030
rect 48486 122030 48487 122062
rect 49096 122062 49172 122068
rect 48486 121998 48492 122030
rect 48416 121654 48492 121998
rect 47942 121590 47943 121622
rect 47877 121589 47943 121590
rect 48416 121590 48422 121654
rect 48486 121590 48492 121654
rect 49096 121998 49102 122062
rect 49166 121998 49172 122062
rect 49237 122062 49303 122063
rect 49237 122030 49238 122062
rect 49096 121654 49172 121998
rect 49096 121622 49102 121654
rect 48416 121584 48492 121590
rect 49101 121590 49102 121622
rect 49166 121622 49172 121654
rect 49232 121998 49238 122030
rect 49302 122030 49303 122062
rect 50320 122062 50396 122068
rect 49302 121998 49308 122030
rect 49232 121654 49308 121998
rect 49166 121590 49167 121622
rect 49101 121589 49167 121590
rect 49232 121590 49238 121654
rect 49302 121590 49308 121654
rect 50320 121998 50326 122062
rect 50390 121998 50396 122062
rect 50869 122062 50935 122063
rect 50869 122030 50870 122062
rect 50320 121654 50396 121998
rect 50320 121622 50326 121654
rect 49232 121584 49308 121590
rect 50325 121590 50326 121622
rect 50390 121622 50396 121654
rect 50864 121998 50870 122030
rect 50934 122030 50935 122062
rect 52229 122062 52295 122063
rect 52229 122030 52230 122062
rect 50934 121998 50940 122030
rect 50864 121654 50940 121998
rect 50390 121590 50391 121622
rect 50325 121589 50391 121590
rect 50864 121590 50870 121654
rect 50934 121590 50940 121654
rect 50864 121584 50940 121590
rect 52224 121998 52230 122030
rect 52294 122030 52295 122062
rect 52904 122062 52980 122068
rect 52294 121998 52300 122030
rect 52224 121654 52300 121998
rect 52224 121590 52230 121654
rect 52294 121590 52300 121654
rect 52904 121998 52910 122062
rect 52974 121998 52980 122062
rect 53317 122062 53383 122063
rect 53317 122030 53318 122062
rect 52904 121654 52980 121998
rect 52904 121622 52910 121654
rect 52224 121584 52300 121590
rect 52909 121590 52910 121622
rect 52974 121622 52980 121654
rect 53312 121998 53318 122030
rect 53382 122030 53383 122062
rect 54128 122062 54204 122068
rect 53382 121998 53388 122030
rect 53312 121654 53388 121998
rect 52974 121590 52975 121622
rect 52909 121589 52975 121590
rect 53312 121590 53318 121654
rect 53382 121590 53388 121654
rect 54128 121998 54134 122062
rect 54198 121998 54204 122062
rect 54677 122062 54743 122063
rect 54677 122030 54678 122062
rect 54128 121654 54204 121998
rect 54128 121622 54134 121654
rect 53312 121584 53388 121590
rect 54133 121590 54134 121622
rect 54198 121622 54204 121654
rect 54672 121998 54678 122030
rect 54742 122030 54743 122062
rect 55352 122062 55428 122068
rect 54742 121998 54748 122030
rect 54672 121654 54748 121998
rect 54198 121590 54199 121622
rect 54133 121589 54199 121590
rect 54672 121590 54678 121654
rect 54742 121590 54748 121654
rect 55352 121998 55358 122062
rect 55422 121998 55428 122062
rect 55352 121654 55428 121998
rect 55352 121622 55358 121654
rect 54672 121584 54748 121590
rect 55357 121590 55358 121622
rect 55422 121622 55428 121654
rect 56712 122062 56788 122068
rect 56712 121998 56718 122062
rect 56782 121998 56788 122062
rect 57125 122062 57191 122063
rect 57125 122030 57126 122062
rect 56712 121654 56788 121998
rect 56712 121622 56718 121654
rect 55422 121590 55423 121622
rect 55357 121589 55423 121590
rect 56717 121590 56718 121622
rect 56782 121622 56788 121654
rect 57120 121998 57126 122030
rect 57190 122030 57191 122062
rect 58077 122062 58143 122063
rect 58077 122030 58078 122062
rect 57190 121998 57196 122030
rect 57120 121654 57196 121998
rect 56782 121590 56783 121622
rect 56717 121589 56783 121590
rect 57120 121590 57126 121654
rect 57190 121590 57196 121654
rect 57120 121584 57196 121590
rect 58072 121998 58078 122030
rect 58142 122030 58143 122062
rect 59160 122062 59236 122068
rect 58142 121998 58148 122030
rect 58072 121654 58148 121998
rect 58072 121590 58078 121654
rect 58142 121590 58148 121654
rect 59160 121998 59166 122062
rect 59230 121998 59236 122062
rect 60933 122062 60999 122063
rect 60933 122030 60934 122062
rect 59160 121654 59236 121998
rect 59160 121622 59166 121654
rect 58072 121584 58148 121590
rect 59165 121590 59166 121622
rect 59230 121622 59236 121654
rect 60928 121998 60934 122030
rect 60998 122030 60999 122062
rect 61608 122062 61684 122068
rect 60998 121998 61004 122030
rect 60928 121654 61004 121998
rect 59230 121590 59231 121622
rect 59165 121589 59231 121590
rect 60928 121590 60934 121654
rect 60998 121590 61004 121654
rect 61608 121998 61614 122062
rect 61678 121998 61684 122062
rect 62157 122062 62223 122063
rect 62157 122030 62158 122062
rect 61608 121654 61684 121998
rect 61608 121622 61614 121654
rect 60928 121584 61004 121590
rect 61613 121590 61614 121622
rect 61678 121622 61684 121654
rect 62152 121998 62158 122030
rect 62222 122030 62223 122062
rect 62832 122062 62908 122068
rect 62222 121998 62228 122030
rect 62152 121654 62228 121998
rect 61678 121590 61679 121622
rect 61613 121589 61679 121590
rect 62152 121590 62158 121654
rect 62222 121590 62228 121654
rect 62832 121998 62838 122062
rect 62902 121998 62908 122062
rect 63381 122062 63447 122063
rect 63381 122030 63382 122062
rect 62832 121654 62908 121998
rect 62832 121622 62838 121654
rect 62152 121584 62228 121590
rect 62837 121590 62838 121622
rect 62902 121622 62908 121654
rect 63376 121998 63382 122030
rect 63446 122030 63447 122062
rect 64056 122062 64132 122068
rect 63446 121998 63452 122030
rect 63376 121654 63452 121998
rect 62902 121590 62903 121622
rect 62837 121589 62903 121590
rect 63376 121590 63382 121654
rect 63446 121590 63452 121654
rect 64056 121998 64062 122062
rect 64126 121998 64132 122062
rect 64605 122062 64671 122063
rect 64605 122030 64606 122062
rect 64056 121654 64132 121998
rect 64056 121622 64062 121654
rect 63376 121584 63452 121590
rect 64061 121590 64062 121622
rect 64126 121622 64132 121654
rect 64600 121998 64606 122030
rect 64670 122030 64671 122062
rect 65688 122062 65764 122068
rect 64670 121998 64676 122030
rect 64600 121654 64676 121998
rect 64126 121590 64127 121622
rect 64061 121589 64127 121590
rect 64600 121590 64606 121654
rect 64670 121590 64676 121654
rect 65688 121998 65694 122062
rect 65758 121998 65764 122062
rect 67189 122062 67255 122063
rect 67189 122030 67190 122062
rect 65688 121654 65764 121998
rect 65688 121622 65694 121654
rect 64600 121584 64676 121590
rect 65693 121590 65694 121622
rect 65758 121622 65764 121654
rect 67184 121998 67190 122030
rect 67254 122030 67255 122062
rect 67864 122062 67940 122068
rect 67254 121998 67260 122030
rect 67184 121654 67260 121998
rect 65758 121590 65759 121622
rect 65693 121589 65759 121590
rect 67184 121590 67190 121654
rect 67254 121590 67260 121654
rect 67864 121998 67870 122062
rect 67934 121998 67940 122062
rect 68413 122062 68479 122063
rect 68413 122030 68414 122062
rect 67864 121654 67940 121998
rect 67864 121622 67870 121654
rect 67184 121584 67260 121590
rect 67869 121590 67870 121622
rect 67934 121622 67940 121654
rect 68408 121998 68414 122030
rect 68478 122030 68479 122062
rect 69088 122062 69164 122068
rect 68478 121998 68484 122030
rect 68408 121654 68484 121998
rect 67934 121590 67935 121622
rect 67869 121589 67935 121590
rect 68408 121590 68414 121654
rect 68478 121590 68484 121654
rect 69088 121998 69094 122062
rect 69158 121998 69164 122062
rect 69637 122062 69703 122063
rect 69637 122030 69638 122062
rect 69088 121654 69164 121998
rect 69088 121622 69094 121654
rect 68408 121584 68484 121590
rect 69093 121590 69094 121622
rect 69158 121622 69164 121654
rect 69632 121998 69638 122030
rect 69702 122030 69703 122062
rect 70312 122062 70388 122068
rect 69702 121998 69708 122030
rect 69632 121654 69708 121998
rect 69158 121590 69159 121622
rect 69093 121589 69159 121590
rect 69632 121590 69638 121654
rect 69702 121590 69708 121654
rect 70312 121998 70318 122062
rect 70382 121998 70388 122062
rect 70861 122062 70927 122063
rect 70861 122030 70862 122062
rect 70312 121654 70388 121998
rect 70312 121622 70318 121654
rect 69632 121584 69708 121590
rect 70317 121590 70318 121622
rect 70382 121622 70388 121654
rect 70856 121998 70862 122030
rect 70926 122030 70927 122062
rect 72085 122062 72151 122063
rect 72085 122030 72086 122062
rect 70926 121998 70932 122030
rect 70856 121654 70932 121998
rect 70382 121590 70383 121622
rect 70317 121589 70383 121590
rect 70856 121590 70862 121654
rect 70926 121590 70932 121654
rect 70856 121584 70932 121590
rect 72080 121998 72086 122030
rect 72150 122030 72151 122062
rect 72765 122062 72831 122063
rect 72765 122030 72766 122062
rect 72150 121998 72156 122030
rect 72080 121654 72156 121998
rect 72080 121590 72086 121654
rect 72150 121590 72156 121654
rect 72080 121584 72156 121590
rect 72760 121998 72766 122030
rect 72830 122030 72831 122062
rect 72896 122062 72972 122068
rect 72830 121998 72836 122030
rect 72760 121654 72836 121998
rect 72760 121590 72766 121654
rect 72830 121590 72836 121654
rect 72896 121998 72902 122062
rect 72966 121998 72972 122062
rect 73309 122062 73375 122063
rect 73309 122030 73310 122062
rect 72896 121654 72972 121998
rect 72896 121622 72902 121654
rect 72760 121584 72836 121590
rect 72901 121590 72902 121622
rect 72966 121622 72972 121654
rect 73304 121998 73310 122030
rect 73374 122030 73375 122062
rect 74120 122062 74196 122068
rect 73374 121998 73380 122030
rect 73304 121654 73380 121998
rect 72966 121590 72967 121622
rect 72901 121589 72967 121590
rect 73304 121590 73310 121654
rect 73374 121590 73380 121654
rect 74120 121998 74126 122062
rect 74190 121998 74196 122062
rect 75213 122062 75279 122063
rect 75213 122030 75214 122062
rect 74120 121654 74196 121998
rect 74120 121622 74126 121654
rect 73304 121584 73380 121590
rect 74125 121590 74126 121622
rect 74190 121622 74196 121654
rect 75208 121998 75214 122030
rect 75278 122030 75279 122062
rect 75344 122062 75420 122068
rect 75278 121998 75284 122030
rect 75208 121654 75284 121998
rect 74190 121590 74191 121622
rect 74125 121589 74191 121590
rect 75208 121590 75214 121654
rect 75278 121590 75284 121654
rect 75344 121998 75350 122062
rect 75414 121998 75420 122062
rect 75893 122062 75959 122063
rect 75893 122030 75894 122062
rect 75344 121654 75420 121998
rect 75344 121622 75350 121654
rect 75208 121584 75284 121590
rect 75349 121590 75350 121622
rect 75414 121622 75420 121654
rect 75888 121998 75894 122030
rect 75958 122030 75959 122062
rect 76568 122062 76644 122068
rect 75958 121998 75964 122030
rect 75888 121654 75964 121998
rect 75414 121590 75415 121622
rect 75349 121589 75415 121590
rect 75888 121590 75894 121654
rect 75958 121590 75964 121654
rect 76568 121998 76574 122062
rect 76638 121998 76644 122062
rect 77117 122062 77183 122063
rect 77117 122030 77118 122062
rect 76568 121654 76644 121998
rect 76568 121622 76574 121654
rect 75888 121584 75964 121590
rect 76573 121590 76574 121622
rect 76638 121622 76644 121654
rect 77112 121998 77118 122030
rect 77182 122030 77183 122062
rect 77792 122062 77868 122068
rect 77182 121998 77188 122030
rect 77112 121654 77188 121998
rect 76638 121590 76639 121622
rect 76573 121589 76639 121590
rect 77112 121590 77118 121654
rect 77182 121590 77188 121654
rect 77792 121998 77798 122062
rect 77862 121998 77868 122062
rect 78341 122062 78407 122063
rect 78341 122030 78342 122062
rect 77792 121654 77868 121998
rect 77792 121622 77798 121654
rect 77112 121584 77188 121590
rect 77797 121590 77798 121622
rect 77862 121622 77868 121654
rect 78336 121998 78342 122030
rect 78406 122030 78407 122062
rect 79565 122062 79631 122063
rect 79565 122030 79566 122062
rect 78406 121998 78412 122030
rect 78336 121654 78412 121998
rect 77862 121590 77863 121622
rect 77797 121589 77863 121590
rect 78336 121590 78342 121654
rect 78406 121590 78412 121654
rect 78336 121584 78412 121590
rect 79560 121998 79566 122030
rect 79630 122030 79631 122062
rect 80517 122062 80583 122063
rect 80517 122030 80518 122062
rect 79630 121998 79636 122030
rect 79560 121654 79636 121998
rect 79560 121590 79566 121654
rect 79630 121590 79636 121654
rect 79560 121584 79636 121590
rect 80512 121998 80518 122030
rect 80582 122030 80583 122062
rect 81469 122062 81535 122063
rect 81469 122030 81470 122062
rect 80582 121998 80588 122030
rect 80512 121518 80588 121998
rect 81464 121998 81470 122030
rect 81534 122030 81535 122062
rect 81600 122062 81676 122068
rect 81534 121998 81540 122030
rect 81464 121654 81540 121998
rect 81464 121590 81470 121654
rect 81534 121590 81540 121654
rect 81600 121998 81606 122062
rect 81670 121998 81676 122062
rect 81600 121654 81676 121998
rect 81600 121622 81606 121654
rect 81464 121584 81540 121590
rect 81605 121590 81606 121622
rect 81670 121622 81676 121654
rect 82824 122062 82900 122068
rect 82824 121998 82830 122062
rect 82894 121998 82900 122062
rect 83373 122062 83439 122063
rect 83373 122030 83374 122062
rect 82824 121654 82900 121998
rect 82824 121622 82830 121654
rect 81670 121590 81671 121622
rect 81605 121589 81671 121590
rect 82829 121590 82830 121622
rect 82894 121622 82900 121654
rect 83368 121998 83374 122030
rect 83438 122030 83439 122062
rect 84048 122062 84124 122068
rect 83438 121998 83444 122030
rect 83368 121654 83444 121998
rect 82894 121590 82895 121622
rect 82829 121589 82895 121590
rect 83368 121590 83374 121654
rect 83438 121590 83444 121654
rect 84048 121998 84054 122062
rect 84118 121998 84124 122062
rect 84597 122062 84663 122063
rect 84597 122030 84598 122062
rect 84048 121654 84124 121998
rect 84048 121622 84054 121654
rect 83368 121584 83444 121590
rect 84053 121590 84054 121622
rect 84118 121622 84124 121654
rect 84592 121998 84598 122030
rect 84662 122030 84663 122062
rect 85408 122062 85484 122068
rect 84662 121998 84668 122030
rect 84592 121654 84668 121998
rect 84118 121590 84119 121622
rect 84053 121589 84119 121590
rect 84592 121590 84598 121654
rect 84662 121590 84668 121654
rect 85408 121998 85414 122062
rect 85478 121998 85484 122062
rect 85821 122062 85887 122063
rect 85821 122030 85822 122062
rect 85408 121654 85484 121998
rect 85408 121622 85414 121654
rect 84592 121584 84668 121590
rect 85413 121590 85414 121622
rect 85478 121622 85484 121654
rect 85816 121998 85822 122030
rect 85886 122030 85887 122062
rect 86496 122062 86572 122068
rect 85886 121998 85892 122030
rect 85816 121654 85892 121998
rect 85478 121590 85479 121622
rect 85413 121589 85479 121590
rect 85816 121590 85822 121654
rect 85886 121590 85892 121654
rect 86496 121998 86502 122062
rect 86566 121998 86572 122062
rect 87045 122062 87111 122063
rect 87045 122030 87046 122062
rect 86496 121654 86572 121998
rect 86496 121622 86502 121654
rect 85816 121584 85892 121590
rect 86501 121590 86502 121622
rect 86566 121622 86572 121654
rect 87040 121998 87046 122030
rect 87110 122030 87111 122062
rect 88405 122062 88471 122063
rect 88405 122030 88406 122062
rect 87110 121998 87116 122030
rect 87040 121654 87116 121998
rect 86566 121590 86567 121622
rect 86501 121589 86567 121590
rect 87040 121590 87046 121654
rect 87110 121590 87116 121654
rect 87040 121584 87116 121590
rect 88400 121998 88406 122030
rect 88470 122030 88471 122062
rect 89080 122062 89156 122068
rect 88470 121998 88476 122030
rect 88400 121654 88476 121998
rect 88400 121590 88406 121654
rect 88470 121590 88476 121654
rect 89080 121998 89086 122062
rect 89150 121998 89156 122062
rect 89221 122062 89287 122063
rect 89221 122030 89222 122062
rect 89080 121654 89156 121998
rect 89080 121622 89086 121654
rect 88400 121584 88476 121590
rect 89085 121590 89086 121622
rect 89150 121622 89156 121654
rect 89216 121998 89222 122030
rect 89286 122030 89287 122062
rect 90304 122062 90380 122068
rect 89286 121998 89292 122030
rect 89216 121654 89292 121998
rect 89150 121590 89151 121622
rect 89085 121589 89151 121590
rect 89216 121590 89222 121654
rect 89286 121590 89292 121654
rect 90304 121998 90310 122062
rect 90374 121998 90380 122062
rect 90853 122062 90919 122063
rect 90853 122030 90854 122062
rect 90304 121654 90380 121998
rect 90304 121622 90310 121654
rect 89216 121584 89292 121590
rect 90309 121590 90310 121622
rect 90374 121622 90380 121654
rect 90848 121998 90854 122030
rect 90918 122030 90919 122062
rect 91528 122062 91604 122068
rect 90918 121998 90924 122030
rect 90848 121654 90924 121998
rect 90374 121590 90375 121622
rect 90309 121589 90375 121590
rect 90848 121590 90854 121654
rect 90918 121590 90924 121654
rect 91528 121998 91534 122062
rect 91598 121998 91604 122062
rect 91528 121654 91604 121998
rect 91528 121622 91534 121654
rect 90848 121584 90924 121590
rect 91533 121590 91534 121622
rect 91598 121622 91604 121654
rect 92752 122062 92828 122068
rect 92752 121998 92758 122062
rect 92822 121998 92828 122062
rect 93301 122062 93367 122063
rect 93301 122030 93302 122062
rect 92752 121654 92828 121998
rect 92752 121622 92758 121654
rect 91598 121590 91599 121622
rect 91533 121589 91599 121590
rect 92757 121590 92758 121622
rect 92822 121622 92828 121654
rect 93296 121998 93302 122030
rect 93366 122030 93367 122062
rect 94253 122062 94319 122063
rect 94253 122030 94254 122062
rect 93366 121998 93372 122030
rect 93296 121654 93372 121998
rect 92822 121590 92823 121622
rect 92757 121589 92823 121590
rect 93296 121590 93302 121654
rect 93366 121590 93372 121654
rect 93296 121584 93372 121590
rect 94248 121998 94254 122030
rect 94318 122030 94319 122062
rect 95477 122062 95543 122063
rect 95477 122030 95478 122062
rect 94318 121998 94324 122030
rect 94248 121654 94324 121998
rect 94248 121590 94254 121654
rect 94318 121590 94324 121654
rect 94248 121584 94324 121590
rect 95472 121998 95478 122030
rect 95542 122030 95543 122062
rect 97109 122062 97175 122063
rect 97109 122030 97110 122062
rect 95542 121998 95548 122030
rect 80512 121454 80518 121518
rect 80582 121454 80588 121518
rect 80512 121448 80588 121454
rect 95472 121518 95548 121998
rect 97104 121998 97110 122030
rect 97174 122030 97175 122062
rect 97784 122062 97860 122068
rect 97174 121998 97180 122030
rect 97104 121654 97180 121998
rect 97104 121590 97110 121654
rect 97174 121590 97180 121654
rect 97784 121998 97790 122062
rect 97854 121998 97860 122062
rect 98333 122062 98399 122063
rect 98333 122030 98334 122062
rect 97784 121654 97860 121998
rect 97784 121622 97790 121654
rect 97104 121584 97180 121590
rect 97789 121590 97790 121622
rect 97854 121622 97860 121654
rect 98328 121998 98334 122030
rect 98398 122030 98399 122062
rect 99008 122062 99084 122068
rect 98398 121998 98404 122030
rect 98328 121654 98404 121998
rect 97854 121590 97855 121622
rect 97789 121589 97855 121590
rect 98328 121590 98334 121654
rect 98398 121590 98404 121654
rect 99008 121998 99014 122062
rect 99078 121998 99084 122062
rect 99557 122062 99623 122063
rect 99557 122030 99558 122062
rect 99008 121654 99084 121998
rect 99008 121622 99014 121654
rect 98328 121584 98404 121590
rect 99013 121590 99014 121622
rect 99078 121622 99084 121654
rect 99552 121998 99558 122030
rect 99622 122030 99623 122062
rect 100781 122062 100847 122063
rect 100781 122030 100782 122062
rect 99622 121998 99628 122030
rect 99552 121654 99628 121998
rect 99078 121590 99079 121622
rect 99013 121589 99079 121590
rect 99552 121590 99558 121654
rect 99622 121590 99628 121654
rect 99552 121584 99628 121590
rect 100776 121998 100782 122030
rect 100846 122030 100847 122062
rect 101592 122062 101668 122068
rect 100846 121998 100852 122030
rect 100776 121654 100852 121998
rect 100776 121590 100782 121654
rect 100846 121590 100852 121654
rect 101592 121998 101598 122062
rect 101662 121998 101668 122062
rect 102005 122062 102071 122063
rect 102005 122030 102006 122062
rect 101592 121654 101668 121998
rect 101592 121622 101598 121654
rect 100776 121584 100852 121590
rect 101597 121590 101598 121622
rect 101662 121622 101668 121654
rect 102000 121998 102006 122030
rect 102070 122030 102071 122062
rect 103365 122062 103431 122063
rect 103365 122030 103366 122062
rect 102070 121998 102076 122030
rect 102000 121654 102076 121998
rect 101662 121590 101663 121622
rect 101597 121589 101663 121590
rect 102000 121590 102006 121654
rect 102070 121590 102076 121654
rect 102000 121584 102076 121590
rect 103360 121998 103366 122030
rect 103430 122030 103431 122062
rect 103909 122062 103975 122063
rect 103909 122030 103910 122062
rect 103430 121998 103436 122030
rect 103360 121654 103436 121998
rect 103360 121590 103366 121654
rect 103430 121590 103436 121654
rect 103360 121584 103436 121590
rect 103904 121998 103910 122030
rect 103974 122030 103975 122062
rect 104040 122062 104116 122068
rect 103974 121998 103980 122030
rect 103904 121654 103980 121998
rect 103904 121590 103910 121654
rect 103974 121590 103980 121654
rect 104040 121998 104046 122062
rect 104110 121998 104116 122062
rect 104589 122062 104655 122063
rect 104589 122030 104590 122062
rect 104040 121654 104116 121998
rect 104040 121622 104046 121654
rect 103904 121584 103980 121590
rect 104045 121590 104046 121622
rect 104110 121622 104116 121654
rect 104584 121998 104590 122030
rect 104654 122030 104655 122062
rect 105813 122062 105879 122063
rect 105813 122030 105814 122062
rect 104654 121998 104660 122030
rect 104584 121654 104660 121998
rect 104110 121590 104111 121622
rect 104045 121589 104111 121590
rect 104584 121590 104590 121654
rect 104654 121590 104660 121654
rect 104584 121584 104660 121590
rect 105808 121998 105814 122030
rect 105878 122030 105879 122062
rect 107037 122062 107103 122063
rect 107037 122030 107038 122062
rect 105878 121998 105884 122030
rect 105808 121654 105884 121998
rect 105808 121590 105814 121654
rect 105878 121590 105884 121654
rect 105808 121584 105884 121590
rect 107032 121998 107038 122030
rect 107102 122030 107103 122062
rect 108120 122062 108196 122068
rect 107102 121998 107108 122030
rect 107032 121654 107108 121998
rect 107032 121590 107038 121654
rect 107102 121590 107108 121654
rect 108120 121998 108126 122062
rect 108190 121998 108196 122062
rect 109485 122062 109551 122063
rect 109485 122030 109486 122062
rect 108120 121654 108196 121998
rect 108120 121622 108126 121654
rect 107032 121584 107108 121590
rect 108125 121590 108126 121622
rect 108190 121622 108196 121654
rect 109480 121998 109486 122030
rect 109550 122030 109551 122062
rect 109550 121998 109556 122030
rect 109480 121654 109556 121998
rect 108190 121590 108191 121622
rect 108125 121589 108191 121590
rect 109480 121590 109486 121654
rect 109550 121590 109556 121654
rect 109480 121584 109556 121590
rect 95472 121454 95478 121518
rect 95542 121454 95548 121518
rect 95472 121448 95548 121454
rect 29920 121078 29926 121110
rect 29925 121046 29926 121078
rect 29990 121078 29996 121110
rect 110160 121110 110236 123494
rect 111661 121518 111727 121519
rect 111661 121486 111662 121518
rect 111656 121454 111662 121486
rect 111726 121486 111727 121518
rect 111726 121454 111732 121486
rect 111656 121246 111732 121454
rect 111656 121182 111662 121246
rect 111726 121182 111732 121246
rect 116280 121246 116356 124854
rect 117232 123700 117308 126214
rect 117368 125054 117444 127710
rect 117504 126414 117580 129070
rect 119408 127910 119484 129886
rect 119544 129270 119620 131246
rect 119680 130086 119756 131926
rect 119952 130902 120028 133764
rect 120632 133214 120708 133220
rect 120632 133150 120638 133214
rect 120702 133150 120708 133214
rect 120632 131446 120708 133150
rect 120632 131414 120638 131446
rect 120637 131382 120638 131414
rect 120702 131414 120708 131446
rect 120702 131382 120703 131414
rect 120637 131381 120703 131382
rect 119952 130870 119958 130902
rect 119957 130838 119958 130870
rect 120022 130870 120028 130902
rect 121176 130902 121252 133764
rect 123624 133214 123700 133220
rect 123624 133150 123630 133214
rect 123694 133150 123700 133214
rect 121448 132534 121524 132540
rect 121448 132470 121454 132534
rect 121518 132470 121524 132534
rect 121448 132126 121524 132470
rect 121448 132094 121454 132126
rect 121453 132062 121454 132094
rect 121518 132094 121524 132126
rect 123080 132534 123156 132540
rect 123080 132470 123086 132534
rect 123150 132470 123156 132534
rect 123080 132126 123156 132470
rect 123080 132094 123086 132126
rect 121518 132062 121519 132094
rect 121453 132061 121519 132062
rect 123085 132062 123086 132094
rect 123150 132094 123156 132126
rect 123150 132062 123151 132094
rect 123085 132061 123151 132062
rect 121176 130870 121182 130902
rect 120022 130838 120023 130870
rect 119957 130837 120023 130838
rect 121181 130838 121182 130870
rect 121246 130870 121252 130902
rect 121246 130838 121247 130870
rect 121181 130837 121247 130838
rect 123624 130494 123700 133150
rect 124712 132534 124788 132540
rect 124712 132470 124718 132534
rect 124782 132470 124788 132534
rect 124712 132126 124788 132470
rect 124712 132094 124718 132126
rect 124717 132062 124718 132094
rect 124782 132094 124788 132126
rect 126344 132534 126420 132540
rect 126344 132470 126350 132534
rect 126414 132470 126420 132534
rect 126344 132126 126420 132470
rect 126344 132094 126350 132126
rect 124782 132062 124783 132094
rect 124717 132061 124783 132062
rect 126349 132062 126350 132094
rect 126414 132094 126420 132126
rect 128112 132534 128188 132540
rect 128112 132470 128118 132534
rect 128182 132470 128188 132534
rect 128112 132126 128188 132470
rect 128112 132094 128118 132126
rect 126414 132062 126415 132094
rect 126349 132061 126415 132062
rect 128117 132062 128118 132094
rect 128182 132094 128188 132126
rect 129880 132534 129956 132540
rect 129880 132470 129886 132534
rect 129950 132470 129956 132534
rect 129880 132126 129956 132470
rect 129880 132094 129886 132126
rect 128182 132062 128183 132094
rect 128117 132061 128183 132062
rect 129885 132062 129886 132094
rect 129950 132094 129956 132126
rect 131376 132534 131452 132540
rect 131376 132470 131382 132534
rect 131446 132470 131452 132534
rect 131376 132126 131452 132470
rect 131376 132094 131382 132126
rect 129950 132062 129951 132094
rect 129885 132061 129951 132062
rect 131381 132062 131382 132094
rect 131446 132094 131452 132126
rect 131446 132062 131447 132094
rect 131381 132061 131447 132062
rect 123624 130462 123630 130494
rect 123629 130430 123630 130462
rect 123694 130462 123700 130494
rect 123694 130430 123695 130462
rect 123629 130429 123695 130430
rect 119680 130054 119686 130086
rect 119685 130022 119686 130054
rect 119750 130054 119756 130086
rect 123760 130358 123836 130364
rect 123760 130294 123766 130358
rect 123830 130294 123836 130358
rect 119750 130022 119751 130054
rect 119685 130021 119751 130022
rect 123629 129950 123695 129951
rect 123629 129918 123630 129950
rect 119544 129238 119550 129270
rect 119549 129206 119550 129238
rect 119614 129238 119620 129270
rect 123624 129886 123630 129918
rect 123694 129918 123695 129950
rect 123694 129886 123700 129918
rect 119614 129206 119615 129238
rect 119549 129205 119615 129206
rect 123624 128998 123700 129886
rect 123624 128934 123630 128998
rect 123694 128934 123700 128998
rect 123624 128928 123700 128934
rect 123629 128862 123695 128863
rect 123629 128830 123630 128862
rect 119408 127878 119414 127910
rect 119413 127846 119414 127878
rect 119478 127878 119484 127910
rect 123624 128798 123630 128830
rect 123694 128830 123695 128862
rect 123694 128798 123700 128830
rect 119478 127846 119479 127878
rect 119413 127845 119479 127846
rect 117504 126350 117510 126414
rect 117574 126350 117580 126414
rect 117504 126344 117580 126350
rect 123624 126278 123700 128798
rect 123760 127638 123836 130294
rect 132736 129814 132812 133764
rect 138176 133486 138524 133492
rect 138176 133422 138182 133486
rect 138246 133422 138318 133486
rect 138382 133422 138454 133486
rect 138518 133422 138524 133486
rect 138176 133350 138524 133422
rect 138176 133286 138182 133350
rect 138246 133286 138318 133350
rect 138382 133286 138454 133350
rect 138518 133286 138524 133350
rect 138176 133214 138524 133286
rect 138176 133150 138182 133214
rect 138246 133150 138318 133214
rect 138382 133150 138454 133214
rect 138518 133150 138524 133214
rect 137496 132806 137844 132812
rect 137496 132742 137502 132806
rect 137566 132742 137638 132806
rect 137702 132742 137774 132806
rect 137838 132742 137844 132806
rect 137496 132670 137844 132742
rect 137496 132606 137502 132670
rect 137566 132606 137638 132670
rect 137702 132606 137774 132670
rect 137838 132606 137844 132670
rect 133144 132534 133220 132540
rect 133144 132470 133150 132534
rect 133214 132470 133220 132534
rect 133144 132126 133220 132470
rect 133144 132094 133150 132126
rect 133149 132062 133150 132094
rect 133214 132094 133220 132126
rect 134912 132534 134988 132540
rect 134912 132470 134918 132534
rect 134982 132470 134988 132534
rect 134912 132126 134988 132470
rect 134912 132094 134918 132126
rect 133214 132062 133215 132094
rect 133149 132061 133215 132062
rect 134917 132062 134918 132094
rect 134982 132094 134988 132126
rect 136408 132534 136484 132540
rect 136408 132470 136414 132534
rect 136478 132470 136484 132534
rect 136408 132126 136484 132470
rect 136408 132094 136414 132126
rect 134982 132062 134983 132094
rect 134917 132061 134983 132062
rect 136413 132062 136414 132094
rect 136478 132094 136484 132126
rect 137496 132534 137844 132606
rect 137496 132470 137502 132534
rect 137566 132470 137638 132534
rect 137702 132470 137774 132534
rect 137838 132470 137844 132534
rect 136478 132062 136479 132094
rect 136413 132061 136479 132062
rect 136821 131990 136887 131991
rect 136821 131958 136822 131990
rect 136816 131926 136822 131958
rect 136886 131958 136887 131990
rect 136886 131926 136892 131958
rect 136816 131582 136892 131926
rect 136816 131518 136822 131582
rect 136886 131518 136892 131582
rect 136816 131512 136892 131518
rect 132736 129782 132742 129814
rect 132741 129750 132742 129782
rect 132806 129782 132812 129814
rect 137496 129814 137844 132470
rect 132806 129750 132807 129782
rect 132741 129749 132807 129750
rect 137496 129750 137502 129814
rect 137566 129750 137844 129814
rect 136821 128862 136887 128863
rect 136821 128830 136822 128862
rect 136816 128798 136822 128830
rect 136886 128830 136887 128862
rect 136886 128798 136892 128830
rect 136816 128182 136892 128798
rect 136816 128118 136822 128182
rect 136886 128118 136892 128182
rect 136816 128112 136892 128118
rect 137496 128182 137844 129750
rect 137496 128118 137502 128182
rect 137566 128118 137844 128182
rect 123760 127606 123766 127638
rect 123765 127574 123766 127606
rect 123830 127606 123836 127638
rect 123830 127574 123831 127606
rect 123765 127573 123831 127574
rect 123624 126214 123630 126278
rect 123694 126214 123700 126278
rect 123624 126208 123700 126214
rect 123896 127502 123972 127508
rect 123896 127438 123902 127502
rect 123966 127438 123972 127502
rect 117368 125022 117374 125054
rect 117373 124990 117374 125022
rect 117438 125022 117444 125054
rect 123760 126142 123836 126148
rect 123760 126078 123766 126142
rect 123830 126078 123836 126142
rect 117438 124990 117439 125022
rect 117373 124989 117439 124990
rect 123624 124646 123700 124652
rect 123624 124582 123630 124646
rect 123694 124582 123700 124646
rect 117232 123694 117444 123700
rect 117232 123630 117374 123694
rect 117438 123630 117444 123694
rect 117232 123624 117444 123630
rect 116280 121214 116286 121246
rect 111656 121176 111732 121182
rect 116285 121182 116286 121214
rect 116350 121214 116356 121246
rect 117368 123422 117444 123428
rect 117368 123358 117374 123422
rect 117438 123358 117444 123422
rect 116350 121182 116351 121214
rect 116285 121181 116351 121182
rect 29990 121046 29991 121078
rect 29925 121045 29991 121046
rect 110160 121046 110166 121110
rect 110230 121046 110236 121110
rect 115333 121110 115399 121111
rect 115333 121078 115334 121110
rect 110160 121040 110236 121046
rect 115328 121046 115334 121078
rect 115398 121078 115399 121110
rect 115398 121046 115404 121078
rect 115328 120702 115404 121046
rect 115328 120638 115334 120702
rect 115398 120638 115404 120702
rect 117368 120702 117444 123358
rect 123624 121926 123700 124582
rect 123760 123422 123836 126078
rect 123896 124782 123972 127438
rect 123896 124750 123902 124782
rect 123901 124718 123902 124750
rect 123966 124750 123972 124782
rect 137496 126550 137844 128118
rect 137496 126486 137502 126550
rect 137566 126486 137844 126550
rect 137496 124782 137844 126486
rect 123966 124718 123967 124750
rect 123901 124717 123967 124718
rect 137496 124718 137502 124782
rect 137566 124718 137844 124782
rect 123760 123390 123766 123422
rect 123765 123358 123766 123390
rect 123830 123390 123836 123422
rect 123830 123358 123831 123390
rect 123765 123357 123831 123358
rect 134645 123286 134711 123287
rect 134645 123254 134646 123286
rect 123624 121894 123630 121926
rect 123629 121862 123630 121894
rect 123694 121894 123700 121926
rect 134640 123222 134646 123254
rect 134710 123254 134711 123286
rect 134710 123222 134716 123254
rect 123694 121862 123695 121894
rect 123629 121861 123695 121862
rect 117368 120670 117374 120702
rect 115328 120632 115404 120638
rect 117373 120638 117374 120670
rect 117438 120670 117444 120702
rect 117438 120638 117439 120670
rect 117373 120637 117439 120638
rect 21760 120566 21836 120572
rect 21760 120502 21766 120566
rect 21830 120502 21836 120566
rect 22309 120566 22375 120567
rect 22309 120534 22310 120566
rect 21760 120294 21836 120502
rect 21760 120262 21766 120294
rect 21765 120230 21766 120262
rect 21830 120262 21836 120294
rect 22304 120502 22310 120534
rect 22374 120534 22375 120566
rect 22576 120566 22652 120572
rect 22374 120502 22380 120534
rect 22304 120294 22380 120502
rect 21830 120230 21831 120262
rect 21765 120229 21831 120230
rect 22304 120230 22310 120294
rect 22374 120230 22380 120294
rect 22576 120502 22582 120566
rect 22646 120502 22652 120566
rect 22989 120566 23055 120567
rect 22989 120534 22990 120566
rect 22576 120294 22652 120502
rect 22576 120262 22582 120294
rect 22304 120224 22380 120230
rect 22581 120230 22582 120262
rect 22646 120262 22652 120294
rect 22984 120502 22990 120534
rect 23054 120534 23055 120566
rect 23397 120566 23463 120567
rect 23397 120534 23398 120566
rect 23054 120502 23060 120534
rect 22984 120294 23060 120502
rect 22646 120230 22647 120262
rect 22581 120229 22647 120230
rect 22984 120230 22990 120294
rect 23054 120230 23060 120294
rect 22984 120224 23060 120230
rect 23392 120502 23398 120534
rect 23462 120534 23463 120566
rect 115197 120566 115263 120567
rect 115197 120534 115198 120566
rect 23462 120502 23468 120534
rect 23392 120294 23468 120502
rect 23392 120230 23398 120294
rect 23462 120230 23468 120294
rect 23392 120224 23468 120230
rect 115192 120502 115198 120534
rect 115262 120534 115263 120566
rect 115736 120566 115812 120572
rect 115262 120502 115268 120534
rect 115192 120294 115268 120502
rect 115192 120230 115198 120294
rect 115262 120230 115268 120294
rect 115736 120502 115742 120566
rect 115806 120502 115812 120566
rect 115736 120294 115812 120502
rect 115736 120262 115742 120294
rect 115192 120224 115268 120230
rect 115741 120230 115742 120262
rect 115806 120262 115812 120294
rect 116008 120566 116084 120572
rect 116008 120502 116014 120566
rect 116078 120502 116084 120566
rect 116965 120566 117031 120567
rect 116965 120534 116966 120566
rect 116008 120294 116084 120502
rect 116008 120262 116014 120294
rect 115806 120230 115807 120262
rect 115741 120229 115807 120230
rect 116013 120230 116014 120262
rect 116078 120262 116084 120294
rect 116960 120502 116966 120534
rect 117030 120534 117031 120566
rect 134640 120566 134716 123222
rect 137496 123014 137844 124718
rect 137496 122950 137502 123014
rect 137566 122950 137844 123014
rect 136192 122918 136258 122919
rect 136192 122854 136193 122918
rect 136257 122854 136258 122918
rect 136192 122853 136258 122854
rect 117030 120502 117036 120534
rect 116960 120294 117036 120502
rect 134640 120502 134646 120566
rect 134710 120502 134716 120566
rect 134640 120496 134716 120502
rect 116078 120230 116079 120262
rect 116013 120229 116079 120230
rect 116960 120230 116966 120294
rect 117030 120230 117036 120294
rect 116960 120224 117036 120230
rect 134640 120430 134716 120436
rect 134640 120366 134646 120430
rect 134710 120366 134716 120430
rect 21760 120158 21836 120164
rect 21760 120094 21766 120158
rect 21830 120094 21836 120158
rect 22581 120158 22647 120159
rect 22581 120126 22582 120158
rect 21760 119886 21836 120094
rect 21760 119854 21766 119886
rect 21765 119822 21766 119854
rect 21830 119854 21836 119886
rect 22576 120094 22582 120126
rect 22646 120126 22647 120158
rect 23120 120158 23196 120164
rect 22646 120094 22652 120126
rect 22576 119886 22652 120094
rect 21830 119822 21831 119854
rect 21765 119821 21831 119822
rect 22576 119822 22582 119886
rect 22646 119822 22652 119886
rect 23120 120094 23126 120158
rect 23190 120094 23196 120158
rect 23120 119886 23196 120094
rect 23120 119854 23126 119886
rect 22576 119816 22652 119822
rect 23125 119822 23126 119854
rect 23190 119854 23196 119886
rect 23528 120158 23604 120164
rect 23528 120094 23534 120158
rect 23598 120094 23604 120158
rect 23528 119886 23604 120094
rect 23528 119854 23534 119886
rect 23190 119822 23191 119854
rect 23125 119821 23191 119822
rect 23533 119822 23534 119854
rect 23598 119854 23604 119886
rect 115328 120158 115404 120164
rect 115328 120094 115334 120158
rect 115398 120094 115404 120158
rect 115741 120158 115807 120159
rect 115741 120126 115742 120158
rect 115328 119886 115404 120094
rect 115328 119854 115334 119886
rect 23598 119822 23599 119854
rect 23533 119821 23599 119822
rect 115333 119822 115334 119854
rect 115398 119854 115404 119886
rect 115736 120094 115742 120126
rect 115806 120126 115807 120158
rect 116824 120158 116900 120164
rect 115806 120094 115812 120126
rect 115736 119886 115812 120094
rect 115398 119822 115399 119854
rect 115333 119821 115399 119822
rect 115736 119822 115742 119886
rect 115806 119822 115812 119886
rect 116824 120094 116830 120158
rect 116894 120094 116900 120158
rect 116824 119886 116900 120094
rect 116824 119854 116830 119886
rect 115736 119816 115812 119822
rect 116829 119822 116830 119854
rect 116894 119854 116900 119886
rect 116894 119822 116895 119854
rect 116829 119821 116895 119822
rect 952 119686 1230 119750
rect 1294 119686 1300 119750
rect 21901 119750 21967 119751
rect 21901 119718 21902 119750
rect 952 118118 1300 119686
rect 21896 119686 21902 119718
rect 21966 119718 21967 119750
rect 22989 119750 23055 119751
rect 22989 119718 22990 119750
rect 21966 119686 21972 119718
rect 21896 119478 21972 119686
rect 21896 119414 21902 119478
rect 21966 119414 21972 119478
rect 21896 119408 21972 119414
rect 22984 119686 22990 119718
rect 23054 119718 23055 119750
rect 23397 119750 23463 119751
rect 23397 119718 23398 119750
rect 23054 119686 23060 119718
rect 22984 119478 23060 119686
rect 22984 119414 22990 119478
rect 23054 119414 23060 119478
rect 22984 119408 23060 119414
rect 23392 119686 23398 119718
rect 23462 119718 23463 119750
rect 115197 119750 115263 119751
rect 115197 119718 115198 119750
rect 23462 119686 23468 119718
rect 23392 119478 23468 119686
rect 23392 119414 23398 119478
rect 23462 119414 23468 119478
rect 23392 119408 23468 119414
rect 115192 119686 115198 119718
rect 115262 119718 115263 119750
rect 115605 119750 115671 119751
rect 115605 119718 115606 119750
rect 115262 119686 115268 119718
rect 115192 119478 115268 119686
rect 115192 119414 115198 119478
rect 115262 119414 115268 119478
rect 115192 119408 115268 119414
rect 115600 119686 115606 119718
rect 115670 119718 115671 119750
rect 116557 119750 116623 119751
rect 116557 119718 116558 119750
rect 115670 119686 115676 119718
rect 115600 119478 115676 119686
rect 115600 119414 115606 119478
rect 115670 119414 115676 119478
rect 115600 119408 115676 119414
rect 116552 119686 116558 119718
rect 116622 119718 116623 119750
rect 116965 119750 117031 119751
rect 116965 119718 116966 119750
rect 116622 119686 116628 119718
rect 116552 119478 116628 119686
rect 116552 119414 116558 119478
rect 116622 119414 116628 119478
rect 116552 119408 116628 119414
rect 116960 119686 116966 119718
rect 117030 119718 117031 119750
rect 117030 119686 117036 119718
rect 116960 119478 117036 119686
rect 116960 119414 116966 119478
rect 117030 119414 117036 119478
rect 116960 119408 117036 119414
rect 21760 119342 21836 119348
rect 21760 119278 21766 119342
rect 21830 119278 21836 119342
rect 22309 119342 22375 119343
rect 22309 119310 22310 119342
rect 21760 119070 21836 119278
rect 21760 119038 21766 119070
rect 21765 119006 21766 119038
rect 21830 119038 21836 119070
rect 22304 119278 22310 119310
rect 22374 119310 22375 119342
rect 22445 119342 22511 119343
rect 22445 119310 22446 119342
rect 22374 119278 22380 119310
rect 22304 119070 22380 119278
rect 21830 119006 21831 119038
rect 21765 119005 21831 119006
rect 22304 119006 22310 119070
rect 22374 119006 22380 119070
rect 22304 119000 22380 119006
rect 22440 119278 22446 119310
rect 22510 119310 22511 119342
rect 23125 119342 23191 119343
rect 23125 119310 23126 119342
rect 22510 119278 22516 119310
rect 22440 119070 22516 119278
rect 22440 119006 22446 119070
rect 22510 119006 22516 119070
rect 22440 119000 22516 119006
rect 23120 119278 23126 119310
rect 23190 119310 23191 119342
rect 23397 119342 23463 119343
rect 23397 119310 23398 119342
rect 23190 119278 23196 119310
rect 23120 119070 23196 119278
rect 23120 119006 23126 119070
rect 23190 119006 23196 119070
rect 23120 119000 23196 119006
rect 23392 119278 23398 119310
rect 23462 119310 23463 119342
rect 115328 119342 115404 119348
rect 23462 119278 23468 119310
rect 23392 119070 23468 119278
rect 23392 119006 23398 119070
rect 23462 119006 23468 119070
rect 115328 119278 115334 119342
rect 115398 119278 115404 119342
rect 115328 119070 115404 119278
rect 115328 119038 115334 119070
rect 23392 119000 23468 119006
rect 115333 119006 115334 119038
rect 115398 119038 115404 119070
rect 115736 119342 115812 119348
rect 115736 119278 115742 119342
rect 115806 119278 115812 119342
rect 115736 119070 115812 119278
rect 115736 119038 115742 119070
rect 115398 119006 115399 119038
rect 115333 119005 115399 119006
rect 115741 119006 115742 119038
rect 115806 119038 115812 119070
rect 116008 119342 116084 119348
rect 116008 119278 116014 119342
rect 116078 119278 116084 119342
rect 116285 119342 116351 119343
rect 116285 119310 116286 119342
rect 116008 119070 116084 119278
rect 116008 119038 116014 119070
rect 115806 119006 115807 119038
rect 115741 119005 115807 119006
rect 116013 119006 116014 119038
rect 116078 119038 116084 119070
rect 116280 119278 116286 119310
rect 116350 119310 116351 119342
rect 116965 119342 117031 119343
rect 116965 119310 116966 119342
rect 116350 119278 116356 119310
rect 116280 119070 116356 119278
rect 116078 119006 116079 119038
rect 116013 119005 116079 119006
rect 116280 119006 116286 119070
rect 116350 119006 116356 119070
rect 116280 119000 116356 119006
rect 116960 119278 116966 119310
rect 117030 119310 117031 119342
rect 117030 119278 117036 119310
rect 116960 119070 117036 119278
rect 116960 119006 116966 119070
rect 117030 119006 117036 119070
rect 116960 119000 117036 119006
rect 22581 118934 22647 118935
rect 22581 118902 22582 118934
rect 22576 118870 22582 118902
rect 22646 118902 22647 118934
rect 22984 118934 23060 118940
rect 22646 118870 22652 118902
rect 22576 118662 22652 118870
rect 22576 118598 22582 118662
rect 22646 118598 22652 118662
rect 22984 118870 22990 118934
rect 23054 118870 23060 118934
rect 22984 118662 23060 118870
rect 22984 118630 22990 118662
rect 22576 118592 22652 118598
rect 22989 118598 22990 118630
rect 23054 118630 23060 118662
rect 23392 118934 23468 118940
rect 23392 118870 23398 118934
rect 23462 118870 23468 118934
rect 23392 118662 23468 118870
rect 115192 118934 115268 118940
rect 115192 118870 115198 118934
rect 115262 118870 115268 118934
rect 28565 118798 28631 118799
rect 28565 118766 28566 118798
rect 23392 118630 23398 118662
rect 23054 118598 23055 118630
rect 22989 118597 23055 118598
rect 23397 118598 23398 118630
rect 23462 118630 23468 118662
rect 28560 118734 28566 118766
rect 28630 118766 28631 118798
rect 110301 118798 110367 118799
rect 110301 118766 110302 118798
rect 28630 118734 28636 118766
rect 23462 118598 23463 118630
rect 23397 118597 23463 118598
rect 22989 118526 23055 118527
rect 22989 118494 22990 118526
rect 22984 118462 22990 118494
rect 23054 118494 23055 118526
rect 23397 118526 23463 118527
rect 23397 118494 23398 118526
rect 23054 118462 23060 118494
rect 22984 118254 23060 118462
rect 22984 118190 22990 118254
rect 23054 118190 23060 118254
rect 22984 118184 23060 118190
rect 23392 118462 23398 118494
rect 23462 118494 23463 118526
rect 28429 118526 28495 118527
rect 28429 118494 28430 118526
rect 23462 118462 23468 118494
rect 23392 118254 23468 118462
rect 23392 118190 23398 118254
rect 23462 118190 23468 118254
rect 23392 118184 23468 118190
rect 28424 118462 28430 118494
rect 28494 118494 28495 118526
rect 28560 118526 28636 118734
rect 28494 118462 28500 118494
rect 952 118054 1230 118118
rect 1294 118054 1300 118118
rect 22173 118118 22239 118119
rect 22173 118086 22174 118118
rect 952 116350 1300 118054
rect 22168 118054 22174 118086
rect 22238 118086 22239 118118
rect 28424 118118 28500 118462
rect 28560 118462 28566 118526
rect 28630 118462 28636 118526
rect 28560 118456 28636 118462
rect 110296 118734 110302 118766
rect 110366 118766 110367 118798
rect 110366 118734 110372 118766
rect 110296 118526 110372 118734
rect 115192 118662 115268 118870
rect 115192 118630 115198 118662
rect 115197 118598 115198 118630
rect 115262 118630 115268 118662
rect 115600 118934 115676 118940
rect 115600 118870 115606 118934
rect 115670 118870 115676 118934
rect 115600 118662 115676 118870
rect 115600 118630 115606 118662
rect 115262 118598 115263 118630
rect 115197 118597 115263 118598
rect 115605 118598 115606 118630
rect 115670 118630 115676 118662
rect 116280 118934 116356 118940
rect 116280 118870 116286 118934
rect 116350 118870 116356 118934
rect 116280 118662 116356 118870
rect 116280 118630 116286 118662
rect 115670 118598 115671 118630
rect 115605 118597 115671 118598
rect 116285 118598 116286 118630
rect 116350 118630 116356 118662
rect 116350 118598 116351 118630
rect 116285 118597 116351 118598
rect 110296 118462 110302 118526
rect 110366 118462 110372 118526
rect 115197 118526 115263 118527
rect 115197 118494 115198 118526
rect 110296 118456 110372 118462
rect 115192 118462 115198 118494
rect 115262 118494 115263 118526
rect 115600 118526 115676 118532
rect 115262 118462 115268 118494
rect 22238 118054 22244 118086
rect 21765 117846 21831 117847
rect 21765 117814 21766 117846
rect 21760 117782 21766 117814
rect 21830 117814 21831 117846
rect 22168 117846 22244 118054
rect 28424 118054 28430 118118
rect 28494 118054 28500 118118
rect 28424 118048 28500 118054
rect 110296 118254 110372 118260
rect 110296 118190 110302 118254
rect 110366 118190 110372 118254
rect 21830 117782 21836 117814
rect 21760 117574 21836 117782
rect 22168 117782 22174 117846
rect 22238 117782 22244 117846
rect 22168 117776 22244 117782
rect 28424 117982 28500 117988
rect 28424 117918 28430 117982
rect 28494 117918 28500 117982
rect 110296 117982 110372 118190
rect 115192 118254 115268 118462
rect 115192 118190 115198 118254
rect 115262 118190 115268 118254
rect 115600 118462 115606 118526
rect 115670 118462 115676 118526
rect 115600 118254 115676 118462
rect 115600 118222 115606 118254
rect 115192 118184 115268 118190
rect 115605 118190 115606 118222
rect 115670 118222 115676 118254
rect 115670 118190 115671 118222
rect 115605 118189 115671 118190
rect 116285 118118 116351 118119
rect 116285 118086 116286 118118
rect 116280 118054 116286 118086
rect 116350 118086 116351 118118
rect 116350 118054 116356 118086
rect 110296 117950 110302 117982
rect 28424 117710 28500 117918
rect 110301 117918 110302 117950
rect 110366 117950 110372 117982
rect 110432 117982 110508 117988
rect 110366 117918 110367 117950
rect 110301 117917 110367 117918
rect 110432 117918 110438 117982
rect 110502 117918 110508 117982
rect 28424 117678 28430 117710
rect 28429 117646 28430 117678
rect 28494 117678 28500 117710
rect 110432 117710 110508 117918
rect 116280 117846 116356 118054
rect 116280 117782 116286 117846
rect 116350 117782 116356 117846
rect 116829 117846 116895 117847
rect 116829 117814 116830 117846
rect 116280 117776 116356 117782
rect 116824 117782 116830 117814
rect 116894 117814 116895 117846
rect 116894 117782 116900 117814
rect 110432 117678 110438 117710
rect 28494 117646 28495 117678
rect 28429 117645 28495 117646
rect 110437 117646 110438 117678
rect 110502 117678 110508 117710
rect 110502 117646 110503 117678
rect 110437 117645 110503 117646
rect 21760 117510 21766 117574
rect 21830 117510 21836 117574
rect 21760 117504 21836 117510
rect 28560 117574 28636 117580
rect 28560 117510 28566 117574
rect 28630 117510 28636 117574
rect 110165 117574 110231 117575
rect 110165 117542 110166 117574
rect 21896 117438 21972 117444
rect 21896 117374 21902 117438
rect 21966 117374 21972 117438
rect 22445 117438 22511 117439
rect 22445 117406 22446 117438
rect 21896 117166 21972 117374
rect 21896 117134 21902 117166
rect 21901 117102 21902 117134
rect 21966 117134 21972 117166
rect 22440 117374 22446 117406
rect 22510 117406 22511 117438
rect 22510 117374 22516 117406
rect 22440 117166 22516 117374
rect 21966 117102 21967 117134
rect 21901 117101 21967 117102
rect 22440 117102 22446 117166
rect 22510 117102 22516 117166
rect 28429 117166 28495 117167
rect 28429 117134 28430 117166
rect 22440 117096 22516 117102
rect 28424 117102 28430 117134
rect 28494 117134 28495 117166
rect 28560 117166 28636 117510
rect 110160 117510 110166 117542
rect 110230 117542 110231 117574
rect 116824 117574 116900 117782
rect 134640 117710 134716 120366
rect 134640 117678 134646 117710
rect 134645 117646 134646 117678
rect 134710 117678 134716 117710
rect 134710 117646 134711 117678
rect 134645 117645 134711 117646
rect 110230 117510 110236 117542
rect 110160 117302 110236 117510
rect 116824 117510 116830 117574
rect 116894 117510 116900 117574
rect 116824 117504 116900 117510
rect 110160 117238 110166 117302
rect 110230 117238 110236 117302
rect 110160 117232 110236 117238
rect 116552 117438 116628 117444
rect 116552 117374 116558 117438
rect 116622 117374 116628 117438
rect 28560 117134 28566 117166
rect 28494 117102 28500 117134
rect 21760 117030 21836 117036
rect 21760 116966 21766 117030
rect 21830 116966 21836 117030
rect 22989 117030 23055 117031
rect 22989 116998 22990 117030
rect 21760 116758 21836 116966
rect 21760 116726 21766 116758
rect 21765 116694 21766 116726
rect 21830 116726 21836 116758
rect 22984 116966 22990 116998
rect 23054 116998 23055 117030
rect 23528 117030 23604 117036
rect 23054 116966 23060 116998
rect 22984 116758 23060 116966
rect 21830 116694 21831 116726
rect 21765 116693 21831 116694
rect 22984 116694 22990 116758
rect 23054 116694 23060 116758
rect 23528 116966 23534 117030
rect 23598 116966 23604 117030
rect 23528 116758 23604 116966
rect 28424 116894 28500 117102
rect 28565 117102 28566 117134
rect 28630 117134 28636 117166
rect 116552 117166 116628 117374
rect 116552 117134 116558 117166
rect 28630 117102 28631 117134
rect 28565 117101 28631 117102
rect 116557 117102 116558 117134
rect 116622 117134 116628 117166
rect 116960 117438 117036 117444
rect 116960 117374 116966 117438
rect 117030 117374 117036 117438
rect 116960 117166 117036 117374
rect 116960 117134 116966 117166
rect 116622 117102 116623 117134
rect 116557 117101 116623 117102
rect 116965 117102 116966 117134
rect 117030 117134 117036 117166
rect 117030 117102 117031 117134
rect 116965 117101 117031 117102
rect 28424 116830 28430 116894
rect 28494 116830 28500 116894
rect 28424 116824 28500 116830
rect 115328 117030 115404 117036
rect 115328 116966 115334 117030
rect 115398 116966 115404 117030
rect 23528 116726 23534 116758
rect 22984 116688 23060 116694
rect 23533 116694 23534 116726
rect 23598 116726 23604 116758
rect 28560 116758 28636 116764
rect 23598 116694 23599 116726
rect 23533 116693 23599 116694
rect 28560 116694 28566 116758
rect 28630 116694 28636 116758
rect 115328 116758 115404 116966
rect 115328 116726 115334 116758
rect 952 116286 1230 116350
rect 1294 116286 1300 116350
rect 21896 116622 21972 116628
rect 21896 116558 21902 116622
rect 21966 116558 21972 116622
rect 23125 116622 23191 116623
rect 23125 116590 23126 116622
rect 21896 116350 21972 116558
rect 21896 116318 21902 116350
rect 952 114718 1300 116286
rect 21901 116286 21902 116318
rect 21966 116318 21972 116350
rect 23120 116558 23126 116590
rect 23190 116590 23191 116622
rect 23392 116622 23468 116628
rect 23190 116558 23196 116590
rect 23120 116350 23196 116558
rect 21966 116286 21967 116318
rect 21901 116285 21967 116286
rect 23120 116286 23126 116350
rect 23190 116286 23196 116350
rect 23392 116558 23398 116622
rect 23462 116558 23468 116622
rect 23392 116350 23468 116558
rect 23392 116318 23398 116350
rect 23120 116280 23196 116286
rect 23397 116286 23398 116318
rect 23462 116318 23468 116350
rect 28560 116350 28636 116694
rect 115333 116694 115334 116726
rect 115398 116726 115404 116758
rect 115736 117030 115812 117036
rect 115736 116966 115742 117030
rect 115806 116966 115812 117030
rect 115736 116758 115812 116966
rect 115736 116726 115742 116758
rect 115398 116694 115399 116726
rect 115333 116693 115399 116694
rect 115741 116694 115742 116726
rect 115806 116726 115812 116758
rect 116824 117030 116900 117036
rect 116824 116966 116830 117030
rect 116894 116966 116900 117030
rect 116824 116758 116900 116966
rect 116824 116726 116830 116758
rect 115806 116694 115807 116726
rect 115741 116693 115807 116694
rect 116829 116694 116830 116726
rect 116894 116726 116900 116758
rect 116894 116694 116895 116726
rect 116829 116693 116895 116694
rect 28560 116318 28566 116350
rect 23462 116286 23463 116318
rect 23397 116285 23463 116286
rect 28565 116286 28566 116318
rect 28630 116318 28636 116350
rect 115192 116622 115268 116628
rect 115192 116558 115198 116622
rect 115262 116558 115268 116622
rect 115741 116622 115807 116623
rect 115741 116590 115742 116622
rect 115192 116350 115268 116558
rect 115192 116318 115198 116350
rect 28630 116286 28631 116318
rect 28565 116285 28631 116286
rect 115197 116286 115198 116318
rect 115262 116318 115268 116350
rect 115736 116558 115742 116590
rect 115806 116590 115807 116622
rect 116552 116622 116628 116628
rect 115806 116558 115812 116590
rect 115736 116350 115812 116558
rect 115262 116286 115263 116318
rect 115197 116285 115263 116286
rect 115736 116286 115742 116350
rect 115806 116286 115812 116350
rect 116552 116558 116558 116622
rect 116622 116558 116628 116622
rect 116552 116350 116628 116558
rect 116552 116318 116558 116350
rect 115736 116280 115812 116286
rect 116557 116286 116558 116318
rect 116622 116318 116628 116350
rect 116960 116622 117036 116628
rect 116960 116558 116966 116622
rect 117030 116558 117036 116622
rect 116960 116350 117036 116558
rect 116960 116318 116966 116350
rect 116622 116286 116623 116318
rect 116557 116285 116623 116286
rect 116965 116286 116966 116318
rect 117030 116318 117036 116350
rect 117030 116286 117031 116318
rect 116965 116285 117031 116286
rect 21901 116214 21967 116215
rect 21901 116182 21902 116214
rect 21896 116150 21902 116182
rect 21966 116182 21967 116214
rect 22440 116214 22516 116220
rect 21966 116150 21972 116182
rect 21896 115942 21972 116150
rect 21896 115878 21902 115942
rect 21966 115878 21972 115942
rect 22440 116150 22446 116214
rect 22510 116150 22516 116214
rect 22989 116214 23055 116215
rect 22989 116182 22990 116214
rect 22440 115942 22516 116150
rect 22440 115910 22446 115942
rect 21896 115872 21972 115878
rect 22445 115878 22446 115910
rect 22510 115910 22516 115942
rect 22984 116150 22990 116182
rect 23054 116182 23055 116214
rect 23397 116214 23463 116215
rect 23397 116182 23398 116214
rect 23054 116150 23060 116182
rect 22984 115942 23060 116150
rect 22510 115878 22511 115910
rect 22445 115877 22511 115878
rect 22984 115878 22990 115942
rect 23054 115878 23060 115942
rect 22984 115872 23060 115878
rect 23392 116150 23398 116182
rect 23462 116182 23463 116214
rect 115197 116214 115263 116215
rect 115197 116182 115198 116214
rect 23462 116150 23468 116182
rect 23392 115942 23468 116150
rect 23392 115878 23398 115942
rect 23462 115878 23468 115942
rect 23392 115872 23468 115878
rect 115192 116150 115198 116182
rect 115262 116182 115263 116214
rect 115736 116214 115812 116220
rect 115262 116150 115268 116182
rect 115192 115942 115268 116150
rect 115192 115878 115198 115942
rect 115262 115878 115268 115942
rect 115736 116150 115742 116214
rect 115806 116150 115812 116214
rect 115736 115942 115812 116150
rect 115736 115910 115742 115942
rect 115192 115872 115268 115878
rect 115741 115878 115742 115910
rect 115806 115910 115812 115942
rect 116008 116214 116084 116220
rect 116008 116150 116014 116214
rect 116078 116150 116084 116214
rect 116285 116214 116351 116215
rect 116285 116182 116286 116214
rect 116008 115942 116084 116150
rect 116008 115910 116014 115942
rect 115806 115878 115807 115910
rect 115741 115877 115807 115878
rect 116013 115878 116014 115910
rect 116078 115910 116084 115942
rect 116280 116150 116286 116182
rect 116350 116182 116351 116214
rect 116965 116214 117031 116215
rect 116965 116182 116966 116214
rect 116350 116150 116356 116182
rect 116280 115942 116356 116150
rect 116078 115878 116079 115910
rect 116013 115877 116079 115878
rect 116280 115878 116286 115942
rect 116350 115878 116356 115942
rect 116280 115872 116356 115878
rect 116960 116150 116966 116182
rect 117030 116182 117031 116214
rect 117030 116150 117036 116182
rect 116960 115942 117036 116150
rect 116960 115878 116966 115942
rect 117030 115878 117036 115942
rect 116960 115872 117036 115878
rect 21760 115806 21836 115812
rect 21760 115742 21766 115806
rect 21830 115742 21836 115806
rect 21760 115534 21836 115742
rect 21760 115502 21766 115534
rect 21765 115470 21766 115502
rect 21830 115502 21836 115534
rect 22168 115806 22244 115812
rect 22168 115742 22174 115806
rect 22238 115742 22244 115806
rect 22168 115534 22244 115742
rect 22168 115502 22174 115534
rect 21830 115470 21831 115502
rect 21765 115469 21831 115470
rect 22173 115470 22174 115502
rect 22238 115502 22244 115534
rect 22576 115806 22652 115812
rect 22576 115742 22582 115806
rect 22646 115742 22652 115806
rect 22576 115534 22652 115742
rect 22576 115502 22582 115534
rect 22238 115470 22239 115502
rect 22173 115469 22239 115470
rect 22581 115470 22582 115502
rect 22646 115502 22652 115534
rect 23120 115806 23196 115812
rect 23120 115742 23126 115806
rect 23190 115742 23196 115806
rect 23533 115806 23599 115807
rect 23533 115774 23534 115806
rect 23120 115534 23196 115742
rect 23120 115502 23126 115534
rect 22646 115470 22647 115502
rect 22581 115469 22647 115470
rect 23125 115470 23126 115502
rect 23190 115502 23196 115534
rect 23528 115742 23534 115774
rect 23598 115774 23599 115806
rect 115328 115806 115404 115812
rect 23598 115742 23604 115774
rect 23528 115534 23604 115742
rect 23190 115470 23191 115502
rect 23125 115469 23191 115470
rect 23528 115470 23534 115534
rect 23598 115470 23604 115534
rect 115328 115742 115334 115806
rect 115398 115742 115404 115806
rect 115741 115806 115807 115807
rect 115741 115774 115742 115806
rect 115328 115534 115404 115742
rect 115328 115502 115334 115534
rect 23528 115464 23604 115470
rect 115333 115470 115334 115502
rect 115398 115502 115404 115534
rect 115736 115742 115742 115774
rect 115806 115774 115807 115806
rect 116829 115806 116895 115807
rect 116829 115774 116830 115806
rect 115806 115742 115812 115774
rect 115736 115534 115812 115742
rect 115398 115470 115399 115502
rect 115333 115469 115399 115470
rect 115736 115470 115742 115534
rect 115806 115470 115812 115534
rect 115736 115464 115812 115470
rect 116824 115742 116830 115774
rect 116894 115774 116895 115806
rect 116894 115742 116900 115774
rect 116824 115534 116900 115742
rect 116824 115470 116830 115534
rect 116894 115470 116900 115534
rect 116824 115464 116900 115470
rect 21896 115398 21972 115404
rect 21896 115334 21902 115398
rect 21966 115334 21972 115398
rect 21896 115126 21972 115334
rect 21896 115094 21902 115126
rect 21901 115062 21902 115094
rect 21966 115094 21972 115126
rect 22712 115398 22788 115404
rect 22712 115334 22718 115398
rect 22782 115334 22788 115398
rect 22712 115126 22788 115334
rect 22712 115094 22718 115126
rect 21966 115062 21967 115094
rect 21901 115061 21967 115062
rect 22717 115062 22718 115094
rect 22782 115094 22788 115126
rect 23120 115398 23196 115404
rect 23120 115334 23126 115398
rect 23190 115334 23196 115398
rect 23120 115126 23196 115334
rect 23120 115094 23126 115126
rect 22782 115062 22783 115094
rect 22717 115061 22783 115062
rect 23125 115062 23126 115094
rect 23190 115094 23196 115126
rect 23392 115398 23468 115404
rect 23392 115334 23398 115398
rect 23462 115334 23468 115398
rect 115333 115398 115399 115399
rect 115333 115366 115334 115398
rect 23392 115126 23468 115334
rect 23392 115094 23398 115126
rect 23190 115062 23191 115094
rect 23125 115061 23191 115062
rect 23397 115062 23398 115094
rect 23462 115094 23468 115126
rect 115328 115334 115334 115366
rect 115398 115366 115399 115398
rect 115600 115398 115676 115404
rect 115398 115334 115404 115366
rect 115328 115126 115404 115334
rect 23462 115062 23463 115094
rect 23397 115061 23463 115062
rect 115328 115062 115334 115126
rect 115398 115062 115404 115126
rect 115600 115334 115606 115398
rect 115670 115334 115676 115398
rect 116557 115398 116623 115399
rect 116557 115366 116558 115398
rect 115600 115126 115676 115334
rect 115600 115094 115606 115126
rect 115328 115056 115404 115062
rect 115605 115062 115606 115094
rect 115670 115094 115676 115126
rect 116552 115334 116558 115366
rect 116622 115366 116623 115398
rect 116965 115398 117031 115399
rect 116965 115366 116966 115398
rect 116622 115334 116628 115366
rect 116552 115126 116628 115334
rect 115670 115062 115671 115094
rect 115605 115061 115671 115062
rect 116552 115062 116558 115126
rect 116622 115062 116628 115126
rect 116552 115056 116628 115062
rect 116960 115334 116966 115366
rect 117030 115366 117031 115398
rect 117030 115334 117036 115366
rect 116960 115126 117036 115334
rect 116960 115062 116966 115126
rect 117030 115062 117036 115126
rect 116960 115056 117036 115062
rect 23125 114990 23191 114991
rect 23125 114958 23126 114990
rect 952 114654 1230 114718
rect 1294 114654 1300 114718
rect 952 113086 1300 114654
rect 23120 114926 23126 114958
rect 23190 114958 23191 114990
rect 23528 114990 23604 114996
rect 23190 114926 23196 114958
rect 23120 114718 23196 114926
rect 23120 114654 23126 114718
rect 23190 114654 23196 114718
rect 23528 114926 23534 114990
rect 23598 114926 23604 114990
rect 23528 114718 23604 114926
rect 115328 114990 115404 114996
rect 115328 114926 115334 114990
rect 115398 114926 115404 114990
rect 110301 114854 110367 114855
rect 110301 114822 110302 114854
rect 23528 114686 23534 114718
rect 23120 114648 23196 114654
rect 23533 114654 23534 114686
rect 23598 114686 23604 114718
rect 110296 114790 110302 114822
rect 110366 114822 110367 114854
rect 110366 114790 110372 114822
rect 23598 114654 23599 114686
rect 23533 114653 23599 114654
rect 22984 114582 23060 114588
rect 22984 114518 22990 114582
rect 23054 114518 23060 114582
rect 22984 114310 23060 114518
rect 22984 114278 22990 114310
rect 22989 114246 22990 114278
rect 23054 114278 23060 114310
rect 23392 114582 23468 114588
rect 23392 114518 23398 114582
rect 23462 114518 23468 114582
rect 23392 114310 23468 114518
rect 110296 114582 110372 114790
rect 115328 114718 115404 114926
rect 115328 114686 115334 114718
rect 115333 114654 115334 114686
rect 115398 114686 115404 114718
rect 115736 114990 115812 114996
rect 115736 114926 115742 114990
rect 115806 114926 115812 114990
rect 116149 114990 116215 114991
rect 116149 114958 116150 114990
rect 115736 114718 115812 114926
rect 115736 114686 115742 114718
rect 115398 114654 115399 114686
rect 115333 114653 115399 114654
rect 115741 114654 115742 114686
rect 115806 114686 115812 114718
rect 116144 114926 116150 114958
rect 116214 114958 116215 114990
rect 116214 114926 116220 114958
rect 116144 114718 116220 114926
rect 115806 114654 115807 114686
rect 115741 114653 115807 114654
rect 116144 114654 116150 114718
rect 116214 114654 116220 114718
rect 116144 114648 116220 114654
rect 135320 114718 135396 114724
rect 135320 114654 135326 114718
rect 135390 114654 135396 114718
rect 110296 114518 110302 114582
rect 110366 114518 110372 114582
rect 110296 114512 110372 114518
rect 115192 114582 115268 114588
rect 115192 114518 115198 114582
rect 115262 114518 115268 114582
rect 115741 114582 115807 114583
rect 115741 114550 115742 114582
rect 23392 114278 23398 114310
rect 23054 114246 23055 114278
rect 22989 114245 23055 114246
rect 23397 114246 23398 114278
rect 23462 114278 23468 114310
rect 115192 114310 115268 114518
rect 115192 114278 115198 114310
rect 23462 114246 23463 114278
rect 23397 114245 23463 114246
rect 115197 114246 115198 114278
rect 115262 114278 115268 114310
rect 115736 114518 115742 114550
rect 115806 114550 115807 114582
rect 115806 114518 115812 114550
rect 115736 114310 115812 114518
rect 115262 114246 115263 114278
rect 115197 114245 115263 114246
rect 115736 114246 115742 114310
rect 115806 114246 115812 114310
rect 115736 114240 115812 114246
rect 22445 114174 22511 114175
rect 22445 114142 22446 114174
rect 22440 114110 22446 114142
rect 22510 114142 22511 114174
rect 23120 114174 23196 114180
rect 22510 114110 22516 114142
rect 21760 113902 21836 113908
rect 21760 113838 21766 113902
rect 21830 113838 21836 113902
rect 21760 113630 21836 113838
rect 22440 113902 22516 114110
rect 22440 113838 22446 113902
rect 22510 113838 22516 113902
rect 23120 114110 23126 114174
rect 23190 114110 23196 114174
rect 23120 113902 23196 114110
rect 23120 113870 23126 113902
rect 22440 113832 22516 113838
rect 23125 113838 23126 113870
rect 23190 113870 23196 113902
rect 23392 114174 23468 114180
rect 23392 114110 23398 114174
rect 23462 114110 23468 114174
rect 23392 113902 23468 114110
rect 115192 114174 115268 114180
rect 115192 114110 115198 114174
rect 115262 114110 115268 114174
rect 23392 113870 23398 113902
rect 23190 113838 23191 113870
rect 23125 113837 23191 113838
rect 23397 113838 23398 113870
rect 23462 113870 23468 113902
rect 28560 114038 28636 114044
rect 28560 113974 28566 114038
rect 28630 113974 28636 114038
rect 23462 113838 23463 113870
rect 23397 113837 23463 113838
rect 28293 113766 28359 113767
rect 28293 113734 28294 113766
rect 21760 113598 21766 113630
rect 21765 113566 21766 113598
rect 21830 113598 21836 113630
rect 28288 113702 28294 113734
rect 28358 113734 28359 113766
rect 28560 113766 28636 113974
rect 115192 113902 115268 114110
rect 115192 113870 115198 113902
rect 115197 113838 115198 113870
rect 115262 113870 115268 113902
rect 115600 114174 115676 114180
rect 115600 114110 115606 114174
rect 115670 114110 115676 114174
rect 116421 114174 116487 114175
rect 116421 114142 116422 114174
rect 115600 113902 115676 114110
rect 115600 113870 115606 113902
rect 115262 113838 115263 113870
rect 115197 113837 115263 113838
rect 115605 113838 115606 113870
rect 115670 113870 115676 113902
rect 116416 114110 116422 114142
rect 116486 114142 116487 114174
rect 116486 114110 116492 114142
rect 116416 113902 116492 114110
rect 115670 113838 115671 113870
rect 115605 113837 115671 113838
rect 116416 113838 116422 113902
rect 116486 113838 116492 113902
rect 116416 113832 116492 113838
rect 116824 113902 116900 113908
rect 116824 113838 116830 113902
rect 116894 113838 116900 113902
rect 28560 113734 28566 113766
rect 28358 113702 28364 113734
rect 21830 113566 21831 113598
rect 21765 113565 21831 113566
rect 21896 113494 21972 113500
rect 21896 113430 21902 113494
rect 21966 113430 21972 113494
rect 22173 113494 22239 113495
rect 22173 113462 22174 113494
rect 21896 113222 21972 113430
rect 21896 113190 21902 113222
rect 21901 113158 21902 113190
rect 21966 113190 21972 113222
rect 22168 113430 22174 113462
rect 22238 113462 22239 113494
rect 22440 113494 22516 113500
rect 22238 113430 22244 113462
rect 22168 113222 22244 113430
rect 21966 113158 21967 113190
rect 21901 113157 21967 113158
rect 22168 113158 22174 113222
rect 22238 113158 22244 113222
rect 22440 113430 22446 113494
rect 22510 113430 22516 113494
rect 22440 113222 22516 113430
rect 28288 113358 28364 113702
rect 28565 113702 28566 113734
rect 28630 113734 28636 113766
rect 28630 113702 28631 113734
rect 28565 113701 28631 113702
rect 28288 113294 28294 113358
rect 28358 113294 28364 113358
rect 110432 113630 110508 113636
rect 110432 113566 110438 113630
rect 110502 113566 110508 113630
rect 116824 113630 116900 113838
rect 116824 113598 116830 113630
rect 110432 113358 110508 113566
rect 116829 113566 116830 113598
rect 116894 113598 116900 113630
rect 116894 113566 116895 113598
rect 116829 113565 116895 113566
rect 116829 113494 116895 113495
rect 116829 113462 116830 113494
rect 110432 113326 110438 113358
rect 28288 113288 28364 113294
rect 110437 113294 110438 113326
rect 110502 113326 110508 113358
rect 116824 113430 116830 113462
rect 116894 113462 116895 113494
rect 116894 113430 116900 113462
rect 110502 113294 110503 113326
rect 110437 113293 110503 113294
rect 22440 113190 22446 113222
rect 22168 113152 22244 113158
rect 22445 113158 22446 113190
rect 22510 113190 22516 113222
rect 28288 113222 28364 113228
rect 22510 113158 22511 113190
rect 22445 113157 22511 113158
rect 28288 113158 28294 113222
rect 28358 113158 28364 113222
rect 952 113022 1230 113086
rect 1294 113022 1300 113086
rect 21901 113086 21967 113087
rect 21901 113054 21902 113086
rect 952 111318 1300 113022
rect 21896 113022 21902 113054
rect 21966 113054 21967 113086
rect 22989 113086 23055 113087
rect 22989 113054 22990 113086
rect 21966 113022 21972 113054
rect 21896 112814 21972 113022
rect 21896 112750 21902 112814
rect 21966 112750 21972 112814
rect 21896 112744 21972 112750
rect 22984 113022 22990 113054
rect 23054 113054 23055 113086
rect 23392 113086 23468 113092
rect 23054 113022 23060 113054
rect 22984 112814 23060 113022
rect 22984 112750 22990 112814
rect 23054 112750 23060 112814
rect 23392 113022 23398 113086
rect 23462 113022 23468 113086
rect 23392 112814 23468 113022
rect 28288 112950 28364 113158
rect 116824 113222 116900 113430
rect 116824 113158 116830 113222
rect 116894 113158 116900 113222
rect 116824 113152 116900 113158
rect 28288 112918 28294 112950
rect 28293 112886 28294 112918
rect 28358 112918 28364 112950
rect 115192 113086 115268 113092
rect 115192 113022 115198 113086
rect 115262 113022 115268 113086
rect 28358 112886 28359 112918
rect 28293 112885 28359 112886
rect 23392 112782 23398 112814
rect 22984 112744 23060 112750
rect 23397 112750 23398 112782
rect 23462 112782 23468 112814
rect 115192 112814 115268 113022
rect 115192 112782 115198 112814
rect 23462 112750 23463 112782
rect 23397 112749 23463 112750
rect 115197 112750 115198 112782
rect 115262 112782 115268 112814
rect 115600 113086 115676 113092
rect 115600 113022 115606 113086
rect 115670 113022 115676 113086
rect 116965 113086 117031 113087
rect 116965 113054 116966 113086
rect 115600 112814 115676 113022
rect 115600 112782 115606 112814
rect 115262 112750 115263 112782
rect 115197 112749 115263 112750
rect 115605 112750 115606 112782
rect 115670 112782 115676 112814
rect 116960 113022 116966 113054
rect 117030 113054 117031 113086
rect 117030 113022 117036 113054
rect 116960 112814 117036 113022
rect 115670 112750 115671 112782
rect 115605 112749 115671 112750
rect 116960 112750 116966 112814
rect 117030 112750 117036 112814
rect 116960 112744 117036 112750
rect 21760 112678 21836 112684
rect 21760 112614 21766 112678
rect 21830 112614 21836 112678
rect 22173 112678 22239 112679
rect 22173 112646 22174 112678
rect 21760 112406 21836 112614
rect 21760 112374 21766 112406
rect 21765 112342 21766 112374
rect 21830 112374 21836 112406
rect 22168 112614 22174 112646
rect 22238 112646 22239 112678
rect 23120 112678 23196 112684
rect 22238 112614 22244 112646
rect 22168 112406 22244 112614
rect 21830 112342 21831 112374
rect 21765 112341 21831 112342
rect 22168 112342 22174 112406
rect 22238 112342 22244 112406
rect 23120 112614 23126 112678
rect 23190 112614 23196 112678
rect 23533 112678 23599 112679
rect 23533 112646 23534 112678
rect 23120 112406 23196 112614
rect 23120 112374 23126 112406
rect 22168 112336 22244 112342
rect 23125 112342 23126 112374
rect 23190 112374 23196 112406
rect 23528 112614 23534 112646
rect 23598 112646 23599 112678
rect 115197 112678 115263 112679
rect 115197 112646 115198 112678
rect 23598 112614 23604 112646
rect 23528 112406 23604 112614
rect 115192 112614 115198 112646
rect 115262 112646 115263 112678
rect 115736 112678 115812 112684
rect 115262 112614 115268 112646
rect 23190 112342 23191 112374
rect 23125 112341 23191 112342
rect 23528 112342 23534 112406
rect 23598 112342 23604 112406
rect 28429 112406 28495 112407
rect 28429 112374 28430 112406
rect 23528 112336 23604 112342
rect 28424 112342 28430 112374
rect 28494 112374 28495 112406
rect 110301 112406 110367 112407
rect 110301 112374 110302 112406
rect 28494 112342 28500 112374
rect 21896 112270 21972 112276
rect 21896 112206 21902 112270
rect 21966 112206 21972 112270
rect 21896 111998 21972 112206
rect 21896 111966 21902 111998
rect 21901 111934 21902 111966
rect 21966 111966 21972 111998
rect 22304 112270 22380 112276
rect 22304 112206 22310 112270
rect 22374 112206 22380 112270
rect 23125 112270 23191 112271
rect 23125 112238 23126 112270
rect 22304 111998 22380 112206
rect 22304 111966 22310 111998
rect 21966 111934 21967 111966
rect 21901 111933 21967 111934
rect 22309 111934 22310 111966
rect 22374 111966 22380 111998
rect 23120 112206 23126 112238
rect 23190 112238 23191 112270
rect 23392 112270 23468 112276
rect 23190 112206 23196 112238
rect 23120 111998 23196 112206
rect 22374 111934 22375 111966
rect 22309 111933 22375 111934
rect 23120 111934 23126 111998
rect 23190 111934 23196 111998
rect 23392 112206 23398 112270
rect 23462 112206 23468 112270
rect 23392 111998 23468 112206
rect 28424 112134 28500 112342
rect 28424 112070 28430 112134
rect 28494 112070 28500 112134
rect 28424 112064 28500 112070
rect 110296 112342 110302 112374
rect 110366 112374 110367 112406
rect 115192 112406 115268 112614
rect 110366 112342 110372 112374
rect 110296 112134 110372 112342
rect 115192 112342 115198 112406
rect 115262 112342 115268 112406
rect 115736 112614 115742 112678
rect 115806 112614 115812 112678
rect 115736 112406 115812 112614
rect 115736 112374 115742 112406
rect 115192 112336 115268 112342
rect 115741 112342 115742 112374
rect 115806 112374 115812 112406
rect 116144 112678 116220 112684
rect 116144 112614 116150 112678
rect 116214 112614 116220 112678
rect 116144 112406 116220 112614
rect 116144 112374 116150 112406
rect 115806 112342 115807 112374
rect 115741 112341 115807 112342
rect 116149 112342 116150 112374
rect 116214 112374 116220 112406
rect 116824 112678 116900 112684
rect 116824 112614 116830 112678
rect 116894 112614 116900 112678
rect 116824 112406 116900 112614
rect 116824 112374 116830 112406
rect 116214 112342 116215 112374
rect 116149 112341 116215 112342
rect 116829 112342 116830 112374
rect 116894 112374 116900 112406
rect 116894 112342 116895 112374
rect 116829 112341 116895 112342
rect 110296 112070 110302 112134
rect 110366 112070 110372 112134
rect 110296 112064 110372 112070
rect 115192 112270 115268 112276
rect 115192 112206 115198 112270
rect 115262 112206 115268 112270
rect 115741 112270 115807 112271
rect 115741 112238 115742 112270
rect 23392 111966 23398 111998
rect 23120 111928 23196 111934
rect 23397 111934 23398 111966
rect 23462 111966 23468 111998
rect 115192 111998 115268 112206
rect 115192 111966 115198 111998
rect 23462 111934 23463 111966
rect 23397 111933 23463 111934
rect 115197 111934 115198 111966
rect 115262 111966 115268 111998
rect 115736 112206 115742 112238
rect 115806 112238 115807 112270
rect 116008 112270 116084 112276
rect 115806 112206 115812 112238
rect 115736 111998 115812 112206
rect 115262 111934 115263 111966
rect 115197 111933 115263 111934
rect 115736 111934 115742 111998
rect 115806 111934 115812 111998
rect 116008 112206 116014 112270
rect 116078 112206 116084 112270
rect 116421 112270 116487 112271
rect 116421 112238 116422 112270
rect 116008 111998 116084 112206
rect 116008 111966 116014 111998
rect 115736 111928 115812 111934
rect 116013 111934 116014 111966
rect 116078 111966 116084 111998
rect 116416 112206 116422 112238
rect 116486 112238 116487 112270
rect 116829 112270 116895 112271
rect 116829 112238 116830 112270
rect 116486 112206 116492 112238
rect 116416 111998 116492 112206
rect 116078 111934 116079 111966
rect 116013 111933 116079 111934
rect 116416 111934 116422 111998
rect 116486 111934 116492 111998
rect 116416 111928 116492 111934
rect 116824 112206 116830 112238
rect 116894 112238 116895 112270
rect 116894 112206 116900 112238
rect 116824 111998 116900 112206
rect 135320 112134 135396 114654
rect 136195 112684 136255 122853
rect 136821 121790 136887 121791
rect 136821 121758 136822 121790
rect 136816 121726 136822 121758
rect 136886 121758 136887 121790
rect 136886 121726 136892 121758
rect 136816 121518 136892 121726
rect 136816 121454 136822 121518
rect 136886 121454 136892 121518
rect 136816 121448 136892 121454
rect 137496 121518 137844 122950
rect 137496 121454 137502 121518
rect 137566 121454 137844 121518
rect 137496 119750 137844 121454
rect 137496 119686 137502 119750
rect 137566 119686 137844 119750
rect 136816 119614 136892 119620
rect 136816 119550 136822 119614
rect 136886 119550 136892 119614
rect 136816 119206 136892 119550
rect 136816 119174 136822 119206
rect 136821 119142 136822 119174
rect 136886 119174 136892 119206
rect 136886 119142 136887 119174
rect 136821 119141 136887 119142
rect 137496 118118 137844 119686
rect 137496 118054 137502 118118
rect 137566 118054 137844 118118
rect 137496 116214 137844 118054
rect 137496 116150 137502 116214
rect 137566 116150 137844 116214
rect 137496 114582 137844 116150
rect 137496 114518 137502 114582
rect 137566 114518 137844 114582
rect 136821 113358 136887 113359
rect 136821 113326 136822 113358
rect 136816 113294 136822 113326
rect 136886 113326 136887 113358
rect 136886 113294 136892 113326
rect 136816 113086 136892 113294
rect 136816 113022 136822 113086
rect 136886 113022 136892 113086
rect 136816 113016 136892 113022
rect 137496 112950 137844 114518
rect 137496 112886 137502 112950
rect 137566 112886 137844 112950
rect 136192 112683 136258 112684
rect 136192 112619 136193 112683
rect 136257 112619 136258 112683
rect 136192 112618 136258 112619
rect 135320 112102 135326 112134
rect 135325 112070 135326 112102
rect 135390 112102 135396 112134
rect 135390 112070 135391 112102
rect 135325 112069 135391 112070
rect 116824 111934 116830 111998
rect 116894 111934 116900 111998
rect 116824 111928 116900 111934
rect 21901 111862 21967 111863
rect 21901 111830 21902 111862
rect 21896 111798 21902 111830
rect 21966 111830 21967 111862
rect 22168 111862 22244 111868
rect 21966 111798 21972 111830
rect 21896 111590 21972 111798
rect 21896 111526 21902 111590
rect 21966 111526 21972 111590
rect 22168 111798 22174 111862
rect 22238 111798 22244 111862
rect 22717 111862 22783 111863
rect 22717 111830 22718 111862
rect 22168 111590 22244 111798
rect 22168 111558 22174 111590
rect 21896 111520 21972 111526
rect 22173 111526 22174 111558
rect 22238 111558 22244 111590
rect 22712 111798 22718 111830
rect 22782 111830 22783 111862
rect 22989 111862 23055 111863
rect 22989 111830 22990 111862
rect 22782 111798 22788 111830
rect 22712 111590 22788 111798
rect 22238 111526 22239 111558
rect 22173 111525 22239 111526
rect 22712 111526 22718 111590
rect 22782 111526 22788 111590
rect 22712 111520 22788 111526
rect 22984 111798 22990 111830
rect 23054 111830 23055 111862
rect 23397 111862 23463 111863
rect 23397 111830 23398 111862
rect 23054 111798 23060 111830
rect 22984 111590 23060 111798
rect 22984 111526 22990 111590
rect 23054 111526 23060 111590
rect 22984 111520 23060 111526
rect 23392 111798 23398 111830
rect 23462 111830 23463 111862
rect 115328 111862 115404 111868
rect 23462 111798 23468 111830
rect 23392 111590 23468 111798
rect 23392 111526 23398 111590
rect 23462 111526 23468 111590
rect 115328 111798 115334 111862
rect 115398 111798 115404 111862
rect 115605 111862 115671 111863
rect 115605 111830 115606 111862
rect 115328 111590 115404 111798
rect 115328 111558 115334 111590
rect 23392 111520 23468 111526
rect 115333 111526 115334 111558
rect 115398 111558 115404 111590
rect 115600 111798 115606 111830
rect 115670 111830 115671 111862
rect 116008 111862 116084 111868
rect 115670 111798 115676 111830
rect 115600 111590 115676 111798
rect 115398 111526 115399 111558
rect 115333 111525 115399 111526
rect 115600 111526 115606 111590
rect 115670 111526 115676 111590
rect 116008 111798 116014 111862
rect 116078 111798 116084 111862
rect 116965 111862 117031 111863
rect 116965 111830 116966 111862
rect 116008 111590 116084 111798
rect 116008 111558 116014 111590
rect 115600 111520 115676 111526
rect 116013 111526 116014 111558
rect 116078 111558 116084 111590
rect 116960 111798 116966 111830
rect 117030 111830 117031 111862
rect 117030 111798 117036 111830
rect 116960 111590 117036 111798
rect 116078 111526 116079 111558
rect 116013 111525 116079 111526
rect 116960 111526 116966 111590
rect 117030 111526 117036 111590
rect 116960 111520 117036 111526
rect 952 111254 1230 111318
rect 1294 111254 1300 111318
rect 952 109686 1300 111254
rect 21760 111454 21836 111460
rect 21760 111390 21766 111454
rect 21830 111390 21836 111454
rect 21760 111182 21836 111390
rect 21760 111150 21766 111182
rect 21765 111118 21766 111150
rect 21830 111150 21836 111182
rect 22576 111454 22652 111460
rect 22576 111390 22582 111454
rect 22646 111390 22652 111454
rect 22576 111182 22652 111390
rect 22576 111150 22582 111182
rect 21830 111118 21831 111150
rect 21765 111117 21831 111118
rect 22581 111118 22582 111150
rect 22646 111150 22652 111182
rect 23120 111454 23196 111460
rect 23120 111390 23126 111454
rect 23190 111390 23196 111454
rect 23533 111454 23599 111455
rect 23533 111422 23534 111454
rect 23120 111182 23196 111390
rect 23120 111150 23126 111182
rect 22646 111118 22647 111150
rect 22581 111117 22647 111118
rect 23125 111118 23126 111150
rect 23190 111150 23196 111182
rect 23528 111390 23534 111422
rect 23598 111422 23599 111454
rect 115333 111454 115399 111455
rect 115333 111422 115334 111454
rect 23598 111390 23604 111422
rect 23528 111182 23604 111390
rect 23190 111118 23191 111150
rect 23125 111117 23191 111118
rect 23528 111118 23534 111182
rect 23598 111118 23604 111182
rect 23528 111112 23604 111118
rect 115328 111390 115334 111422
rect 115398 111422 115399 111454
rect 115741 111454 115807 111455
rect 115741 111422 115742 111454
rect 115398 111390 115404 111422
rect 115328 111182 115404 111390
rect 115328 111118 115334 111182
rect 115398 111118 115404 111182
rect 115328 111112 115404 111118
rect 115736 111390 115742 111422
rect 115806 111422 115807 111454
rect 116421 111454 116487 111455
rect 116421 111422 116422 111454
rect 115806 111390 115812 111422
rect 115736 111182 115812 111390
rect 115736 111118 115742 111182
rect 115806 111118 115812 111182
rect 115736 111112 115812 111118
rect 116416 111390 116422 111422
rect 116486 111422 116487 111454
rect 116824 111454 116900 111460
rect 116486 111390 116492 111422
rect 116416 111182 116492 111390
rect 116416 111118 116422 111182
rect 116486 111118 116492 111182
rect 116824 111390 116830 111454
rect 116894 111390 116900 111454
rect 116824 111182 116900 111390
rect 116824 111150 116830 111182
rect 116416 111112 116492 111118
rect 116829 111118 116830 111150
rect 116894 111150 116900 111182
rect 137496 111318 137844 112886
rect 137496 111254 137502 111318
rect 137566 111254 137844 111318
rect 116894 111118 116895 111150
rect 116829 111117 116895 111118
rect 22309 111046 22375 111047
rect 22309 111014 22310 111046
rect 22304 110982 22310 111014
rect 22374 111014 22375 111046
rect 22445 111046 22511 111047
rect 22445 111014 22446 111046
rect 22374 110982 22380 111014
rect 22304 110774 22380 110982
rect 22304 110710 22310 110774
rect 22374 110710 22380 110774
rect 22304 110704 22380 110710
rect 22440 110982 22446 111014
rect 22510 111014 22511 111046
rect 23120 111046 23196 111052
rect 22510 110982 22516 111014
rect 22440 110774 22516 110982
rect 22440 110710 22446 110774
rect 22510 110710 22516 110774
rect 23120 110982 23126 111046
rect 23190 110982 23196 111046
rect 23120 110774 23196 110982
rect 23120 110742 23126 110774
rect 22440 110704 22516 110710
rect 23125 110710 23126 110742
rect 23190 110742 23196 110774
rect 23392 111046 23468 111052
rect 23392 110982 23398 111046
rect 23462 110982 23468 111046
rect 23392 110774 23468 110982
rect 115192 111046 115268 111052
rect 115192 110982 115198 111046
rect 115262 110982 115268 111046
rect 23392 110742 23398 110774
rect 23190 110710 23191 110742
rect 23125 110709 23191 110710
rect 23397 110710 23398 110742
rect 23462 110742 23468 110774
rect 28288 110910 28364 110916
rect 28288 110846 28294 110910
rect 28358 110846 28364 110910
rect 23462 110710 23463 110742
rect 23397 110709 23463 110710
rect 23125 110638 23191 110639
rect 23125 110606 23126 110638
rect 23120 110574 23126 110606
rect 23190 110606 23191 110638
rect 23397 110638 23463 110639
rect 23397 110606 23398 110638
rect 23190 110574 23196 110606
rect 23120 110366 23196 110574
rect 23120 110302 23126 110366
rect 23190 110302 23196 110366
rect 23120 110296 23196 110302
rect 23392 110574 23398 110606
rect 23462 110606 23463 110638
rect 28288 110638 28364 110846
rect 115192 110774 115268 110982
rect 115192 110742 115198 110774
rect 115197 110710 115198 110742
rect 115262 110742 115268 110774
rect 115600 111046 115676 111052
rect 115600 110982 115606 111046
rect 115670 110982 115676 111046
rect 115600 110774 115676 110982
rect 115600 110742 115606 110774
rect 115262 110710 115263 110742
rect 115197 110709 115263 110710
rect 115605 110710 115606 110742
rect 115670 110742 115676 110774
rect 116552 111046 116628 111052
rect 116552 110982 116558 111046
rect 116622 110982 116628 111046
rect 116552 110774 116628 110982
rect 116552 110742 116558 110774
rect 115670 110710 115671 110742
rect 115605 110709 115671 110710
rect 116557 110710 116558 110742
rect 116622 110742 116628 110774
rect 116622 110710 116623 110742
rect 116557 110709 116623 110710
rect 28288 110606 28294 110638
rect 23462 110574 23468 110606
rect 23392 110366 23468 110574
rect 28293 110574 28294 110606
rect 28358 110606 28364 110638
rect 115197 110638 115263 110639
rect 115197 110606 115198 110638
rect 28358 110574 28359 110606
rect 28293 110573 28359 110574
rect 115192 110574 115198 110606
rect 115262 110606 115263 110638
rect 115736 110638 115812 110644
rect 115262 110574 115268 110606
rect 23392 110302 23398 110366
rect 23462 110302 23468 110366
rect 23392 110296 23468 110302
rect 115192 110366 115268 110574
rect 115192 110302 115198 110366
rect 115262 110302 115268 110366
rect 115736 110574 115742 110638
rect 115806 110574 115812 110638
rect 115736 110366 115812 110574
rect 115736 110334 115742 110366
rect 115192 110296 115268 110302
rect 115741 110302 115742 110334
rect 115806 110334 115812 110366
rect 115806 110302 115807 110334
rect 115741 110301 115807 110302
rect 22440 110230 22516 110236
rect 22440 110166 22446 110230
rect 22510 110166 22516 110230
rect 21901 109958 21967 109959
rect 21901 109926 21902 109958
rect 952 109622 1230 109686
rect 1294 109622 1300 109686
rect 952 108054 1300 109622
rect 21896 109894 21902 109926
rect 21966 109926 21967 109958
rect 22440 109958 22516 110166
rect 22440 109926 22446 109958
rect 21966 109894 21972 109926
rect 21896 109686 21972 109894
rect 22445 109894 22446 109926
rect 22510 109926 22516 109958
rect 22984 110230 23060 110236
rect 22984 110166 22990 110230
rect 23054 110166 23060 110230
rect 23533 110230 23599 110231
rect 23533 110198 23534 110230
rect 22984 109958 23060 110166
rect 22984 109926 22990 109958
rect 22510 109894 22511 109926
rect 22445 109893 22511 109894
rect 22989 109894 22990 109926
rect 23054 109926 23060 109958
rect 23528 110166 23534 110198
rect 23598 110198 23599 110230
rect 115192 110230 115268 110236
rect 23598 110166 23604 110198
rect 23528 109958 23604 110166
rect 115192 110166 115198 110230
rect 115262 110166 115268 110230
rect 115741 110230 115807 110231
rect 115741 110198 115742 110230
rect 28565 110094 28631 110095
rect 28565 110062 28566 110094
rect 23054 109894 23055 109926
rect 22989 109893 23055 109894
rect 23528 109894 23534 109958
rect 23598 109894 23604 109958
rect 23528 109888 23604 109894
rect 28560 110030 28566 110062
rect 28630 110062 28631 110094
rect 110160 110094 110236 110100
rect 28630 110030 28636 110062
rect 22309 109822 22375 109823
rect 22309 109790 22310 109822
rect 21896 109622 21902 109686
rect 21966 109622 21972 109686
rect 21896 109616 21972 109622
rect 22304 109758 22310 109790
rect 22374 109790 22375 109822
rect 28560 109822 28636 110030
rect 22374 109758 22380 109790
rect 22304 109692 22380 109758
rect 28560 109758 28566 109822
rect 28630 109758 28636 109822
rect 110160 110030 110166 110094
rect 110230 110030 110236 110094
rect 110160 109822 110236 110030
rect 115192 109958 115268 110166
rect 115192 109926 115198 109958
rect 115197 109894 115198 109926
rect 115262 109926 115268 109958
rect 115736 110166 115742 110198
rect 115806 110198 115807 110230
rect 116008 110230 116084 110236
rect 115806 110166 115812 110198
rect 115736 109958 115812 110166
rect 115262 109894 115263 109926
rect 115197 109893 115263 109894
rect 115736 109894 115742 109958
rect 115806 109894 115812 109958
rect 116008 110166 116014 110230
rect 116078 110166 116084 110230
rect 116008 109958 116084 110166
rect 116008 109926 116014 109958
rect 115736 109888 115812 109894
rect 116013 109894 116014 109926
rect 116078 109926 116084 109958
rect 116965 109958 117031 109959
rect 116965 109926 116966 109958
rect 116078 109894 116079 109926
rect 116013 109893 116079 109894
rect 116960 109894 116966 109926
rect 117030 109926 117031 109958
rect 117030 109894 117036 109926
rect 110160 109790 110166 109822
rect 28560 109752 28636 109758
rect 110165 109758 110166 109790
rect 110230 109790 110236 109822
rect 110230 109758 110231 109790
rect 110165 109757 110231 109758
rect 22304 109686 22516 109692
rect 22304 109622 22446 109686
rect 22510 109622 22516 109686
rect 22304 109616 22516 109622
rect 28288 109686 28364 109692
rect 28288 109622 28294 109686
rect 28358 109622 28364 109686
rect 110165 109686 110231 109687
rect 110165 109654 110166 109686
rect 21760 109550 21836 109556
rect 21760 109486 21766 109550
rect 21830 109486 21836 109550
rect 22445 109550 22511 109551
rect 22445 109518 22446 109550
rect 21760 109278 21836 109486
rect 21760 109246 21766 109278
rect 21765 109214 21766 109246
rect 21830 109246 21836 109278
rect 22440 109486 22446 109518
rect 22510 109518 22511 109550
rect 22510 109486 22516 109518
rect 22440 109278 22516 109486
rect 28288 109414 28364 109622
rect 28288 109382 28294 109414
rect 28293 109350 28294 109382
rect 28358 109382 28364 109414
rect 110160 109622 110166 109654
rect 110230 109654 110231 109686
rect 110301 109686 110367 109687
rect 110301 109654 110302 109686
rect 110230 109622 110236 109654
rect 110160 109414 110236 109622
rect 28358 109350 28359 109382
rect 28293 109349 28359 109350
rect 110160 109350 110166 109414
rect 110230 109350 110236 109414
rect 110160 109344 110236 109350
rect 110296 109622 110302 109654
rect 110366 109654 110367 109686
rect 116960 109686 117036 109894
rect 110366 109622 110372 109654
rect 21830 109214 21831 109246
rect 21765 109213 21831 109214
rect 22440 109214 22446 109278
rect 22510 109214 22516 109278
rect 28293 109278 28359 109279
rect 28293 109246 28294 109278
rect 22440 109208 22516 109214
rect 28288 109214 28294 109246
rect 28358 109246 28359 109278
rect 110296 109278 110372 109622
rect 116960 109622 116966 109686
rect 117030 109622 117036 109686
rect 116960 109616 117036 109622
rect 137496 109686 137844 111254
rect 137496 109622 137502 109686
rect 137566 109622 137844 109686
rect 116149 109550 116215 109551
rect 116149 109518 116150 109550
rect 116144 109486 116150 109518
rect 116214 109518 116215 109550
rect 116285 109550 116351 109551
rect 116285 109518 116286 109550
rect 116214 109486 116220 109518
rect 28358 109214 28364 109246
rect 21896 109142 21972 109148
rect 21896 109078 21902 109142
rect 21966 109078 21972 109142
rect 21896 108870 21972 109078
rect 28288 109006 28364 109214
rect 110296 109214 110302 109278
rect 110366 109214 110372 109278
rect 110296 109208 110372 109214
rect 110432 109278 110508 109284
rect 110432 109214 110438 109278
rect 110502 109214 110508 109278
rect 28288 108942 28294 109006
rect 28358 108942 28364 109006
rect 110432 109006 110508 109214
rect 116144 109278 116220 109486
rect 116144 109214 116150 109278
rect 116214 109214 116220 109278
rect 116144 109208 116220 109214
rect 116280 109486 116286 109518
rect 116350 109518 116351 109550
rect 116965 109550 117031 109551
rect 116965 109518 116966 109550
rect 116350 109486 116356 109518
rect 116280 109278 116356 109486
rect 116280 109214 116286 109278
rect 116350 109214 116356 109278
rect 116280 109208 116356 109214
rect 116960 109486 116966 109518
rect 117030 109518 117031 109550
rect 117030 109486 117036 109518
rect 116960 109278 117036 109486
rect 116960 109214 116966 109278
rect 117030 109214 117036 109278
rect 116960 109208 117036 109214
rect 110432 108974 110438 109006
rect 28288 108936 28364 108942
rect 110437 108942 110438 108974
rect 110502 108974 110508 109006
rect 116960 109142 117036 109148
rect 116960 109078 116966 109142
rect 117030 109078 117036 109142
rect 110502 108942 110503 108974
rect 110437 108941 110503 108942
rect 21896 108838 21902 108870
rect 21901 108806 21902 108838
rect 21966 108838 21972 108870
rect 28429 108870 28495 108871
rect 28429 108838 28430 108870
rect 21966 108806 21967 108838
rect 21901 108805 21967 108806
rect 28424 108806 28430 108838
rect 28494 108838 28495 108870
rect 116960 108870 117036 109078
rect 116960 108838 116966 108870
rect 28494 108806 28500 108838
rect 21901 108734 21967 108735
rect 21901 108702 21902 108734
rect 21896 108670 21902 108702
rect 21966 108702 21967 108734
rect 22309 108734 22375 108735
rect 22309 108702 22310 108734
rect 21966 108670 21972 108702
rect 21896 108462 21972 108670
rect 21896 108398 21902 108462
rect 21966 108398 21972 108462
rect 21896 108392 21972 108398
rect 22304 108670 22310 108702
rect 22374 108702 22375 108734
rect 23120 108734 23196 108740
rect 22374 108670 22380 108702
rect 22304 108462 22380 108670
rect 22304 108398 22310 108462
rect 22374 108398 22380 108462
rect 23120 108670 23126 108734
rect 23190 108670 23196 108734
rect 23397 108734 23463 108735
rect 23397 108702 23398 108734
rect 23120 108462 23196 108670
rect 23120 108430 23126 108462
rect 22304 108392 22380 108398
rect 23125 108398 23126 108430
rect 23190 108430 23196 108462
rect 23392 108670 23398 108702
rect 23462 108702 23463 108734
rect 23462 108670 23468 108702
rect 23392 108462 23468 108670
rect 23190 108398 23191 108430
rect 23125 108397 23191 108398
rect 23392 108398 23398 108462
rect 23462 108398 23468 108462
rect 23392 108392 23468 108398
rect 28424 108462 28500 108806
rect 116965 108806 116966 108838
rect 117030 108838 117036 108870
rect 117030 108806 117031 108838
rect 116965 108805 117031 108806
rect 115192 108734 115268 108740
rect 115192 108670 115198 108734
rect 115262 108670 115268 108734
rect 115605 108734 115671 108735
rect 115605 108702 115606 108734
rect 28424 108398 28430 108462
rect 28494 108398 28500 108462
rect 28424 108392 28500 108398
rect 28560 108462 28636 108468
rect 28560 108398 28566 108462
rect 28630 108398 28636 108462
rect 115192 108462 115268 108670
rect 115192 108430 115198 108462
rect 952 107990 1230 108054
rect 1294 107990 1300 108054
rect 21760 108326 21836 108332
rect 21760 108262 21766 108326
rect 21830 108262 21836 108326
rect 22173 108326 22239 108327
rect 22173 108294 22174 108326
rect 21760 108054 21836 108262
rect 21760 108022 21766 108054
rect 952 106150 1300 107990
rect 21765 107990 21766 108022
rect 21830 108022 21836 108054
rect 22168 108262 22174 108294
rect 22238 108294 22239 108326
rect 22989 108326 23055 108327
rect 22989 108294 22990 108326
rect 22238 108262 22244 108294
rect 22168 108054 22244 108262
rect 21830 107990 21831 108022
rect 21765 107989 21831 107990
rect 22168 107990 22174 108054
rect 22238 107990 22244 108054
rect 22168 107984 22244 107990
rect 22984 108262 22990 108294
rect 23054 108294 23055 108326
rect 23533 108326 23599 108327
rect 23533 108294 23534 108326
rect 23054 108262 23060 108294
rect 22984 108054 23060 108262
rect 22984 107990 22990 108054
rect 23054 107990 23060 108054
rect 22984 107984 23060 107990
rect 23528 108262 23534 108294
rect 23598 108294 23599 108326
rect 23598 108262 23604 108294
rect 23528 108054 23604 108262
rect 28560 108190 28636 108398
rect 115197 108398 115198 108430
rect 115262 108430 115268 108462
rect 115600 108670 115606 108702
rect 115670 108702 115671 108734
rect 116013 108734 116079 108735
rect 116013 108702 116014 108734
rect 115670 108670 115676 108702
rect 115600 108462 115676 108670
rect 115262 108398 115263 108430
rect 115197 108397 115263 108398
rect 115600 108398 115606 108462
rect 115670 108398 115676 108462
rect 115600 108392 115676 108398
rect 116008 108670 116014 108702
rect 116078 108702 116079 108734
rect 116965 108734 117031 108735
rect 116965 108702 116966 108734
rect 116078 108670 116084 108702
rect 116008 108462 116084 108670
rect 116008 108398 116014 108462
rect 116078 108398 116084 108462
rect 116008 108392 116084 108398
rect 116960 108670 116966 108702
rect 117030 108702 117031 108734
rect 117030 108670 117036 108702
rect 116960 108462 117036 108670
rect 116960 108398 116966 108462
rect 117030 108398 117036 108462
rect 116960 108392 117036 108398
rect 28560 108158 28566 108190
rect 28565 108126 28566 108158
rect 28630 108158 28636 108190
rect 115328 108326 115404 108332
rect 115328 108262 115334 108326
rect 115398 108262 115404 108326
rect 115741 108326 115807 108327
rect 115741 108294 115742 108326
rect 28630 108126 28631 108158
rect 28565 108125 28631 108126
rect 23528 107990 23534 108054
rect 23598 107990 23604 108054
rect 115328 108054 115404 108262
rect 115328 108022 115334 108054
rect 23528 107984 23604 107990
rect 115333 107990 115334 108022
rect 115398 108022 115404 108054
rect 115736 108262 115742 108294
rect 115806 108294 115807 108326
rect 116285 108326 116351 108327
rect 116285 108294 116286 108326
rect 115806 108262 115812 108294
rect 115736 108054 115812 108262
rect 115398 107990 115399 108022
rect 115333 107989 115399 107990
rect 115736 107990 115742 108054
rect 115806 107990 115812 108054
rect 115736 107984 115812 107990
rect 116280 108262 116286 108294
rect 116350 108294 116351 108326
rect 116824 108326 116900 108332
rect 116350 108262 116356 108294
rect 116280 108054 116356 108262
rect 116280 107990 116286 108054
rect 116350 107990 116356 108054
rect 116824 108262 116830 108326
rect 116894 108262 116900 108326
rect 116824 108054 116900 108262
rect 116824 108022 116830 108054
rect 116280 107984 116356 107990
rect 116829 107990 116830 108022
rect 116894 108022 116900 108054
rect 137496 108054 137844 109622
rect 116894 107990 116895 108022
rect 116829 107989 116895 107990
rect 137496 107990 137502 108054
rect 137566 107990 137844 108054
rect 21896 107918 21972 107924
rect 21896 107854 21902 107918
rect 21966 107854 21972 107918
rect 21896 107646 21972 107854
rect 21896 107614 21902 107646
rect 21901 107582 21902 107614
rect 21966 107614 21972 107646
rect 22304 107918 22380 107924
rect 22304 107854 22310 107918
rect 22374 107854 22380 107918
rect 22581 107918 22647 107919
rect 22581 107886 22582 107918
rect 22304 107646 22380 107854
rect 22304 107614 22310 107646
rect 21966 107582 21967 107614
rect 21901 107581 21967 107582
rect 22309 107582 22310 107614
rect 22374 107614 22380 107646
rect 22576 107854 22582 107886
rect 22646 107886 22647 107918
rect 23125 107918 23191 107919
rect 23125 107886 23126 107918
rect 22646 107854 22652 107886
rect 22576 107646 22652 107854
rect 22374 107582 22375 107614
rect 22309 107581 22375 107582
rect 22576 107582 22582 107646
rect 22646 107582 22652 107646
rect 22576 107576 22652 107582
rect 23120 107854 23126 107886
rect 23190 107886 23191 107918
rect 23392 107918 23468 107924
rect 23190 107854 23196 107886
rect 23120 107646 23196 107854
rect 23120 107582 23126 107646
rect 23190 107582 23196 107646
rect 23392 107854 23398 107918
rect 23462 107854 23468 107918
rect 23392 107646 23468 107854
rect 23392 107614 23398 107646
rect 23120 107576 23196 107582
rect 23397 107582 23398 107614
rect 23462 107614 23468 107646
rect 115192 107918 115268 107924
rect 115192 107854 115198 107918
rect 115262 107854 115268 107918
rect 115192 107646 115268 107854
rect 115192 107614 115198 107646
rect 23462 107582 23463 107614
rect 23397 107581 23463 107582
rect 115197 107582 115198 107614
rect 115262 107614 115268 107646
rect 115600 107918 115676 107924
rect 115600 107854 115606 107918
rect 115670 107854 115676 107918
rect 116149 107918 116215 107919
rect 116149 107886 116150 107918
rect 115600 107646 115676 107854
rect 115600 107614 115606 107646
rect 115262 107582 115263 107614
rect 115197 107581 115263 107582
rect 115605 107582 115606 107614
rect 115670 107614 115676 107646
rect 116144 107854 116150 107886
rect 116214 107886 116215 107918
rect 116421 107918 116487 107919
rect 116421 107886 116422 107918
rect 116214 107854 116220 107886
rect 116144 107646 116220 107854
rect 115670 107582 115671 107614
rect 115605 107581 115671 107582
rect 116144 107582 116150 107646
rect 116214 107582 116220 107646
rect 116144 107576 116220 107582
rect 116416 107854 116422 107886
rect 116486 107886 116487 107918
rect 116960 107918 117036 107924
rect 116486 107854 116492 107886
rect 116416 107646 116492 107854
rect 116416 107582 116422 107646
rect 116486 107582 116492 107646
rect 116960 107854 116966 107918
rect 117030 107854 117036 107918
rect 116960 107646 117036 107854
rect 116960 107614 116966 107646
rect 116416 107576 116492 107582
rect 116965 107582 116966 107614
rect 117030 107614 117036 107646
rect 117030 107582 117031 107614
rect 116965 107581 117031 107582
rect 21901 107510 21967 107511
rect 21901 107478 21902 107510
rect 21896 107446 21902 107478
rect 21966 107478 21967 107510
rect 22440 107510 22516 107516
rect 21966 107446 21972 107478
rect 21896 107238 21972 107446
rect 21896 107174 21902 107238
rect 21966 107174 21972 107238
rect 22440 107446 22446 107510
rect 22510 107446 22516 107510
rect 22440 107238 22516 107446
rect 22440 107206 22446 107238
rect 21896 107168 21972 107174
rect 22445 107174 22446 107206
rect 22510 107206 22516 107238
rect 22576 107510 22652 107516
rect 22576 107446 22582 107510
rect 22646 107446 22652 107510
rect 22576 107238 22652 107446
rect 22576 107206 22582 107238
rect 22510 107174 22511 107206
rect 22445 107173 22511 107174
rect 22581 107174 22582 107206
rect 22646 107206 22652 107238
rect 22984 107510 23060 107516
rect 22984 107446 22990 107510
rect 23054 107446 23060 107510
rect 22984 107238 23060 107446
rect 22984 107206 22990 107238
rect 22646 107174 22647 107206
rect 22581 107173 22647 107174
rect 22989 107174 22990 107206
rect 23054 107206 23060 107238
rect 23528 107510 23604 107516
rect 23528 107446 23534 107510
rect 23598 107446 23604 107510
rect 115197 107510 115263 107511
rect 115197 107478 115198 107510
rect 23528 107238 23604 107446
rect 23528 107206 23534 107238
rect 23054 107174 23055 107206
rect 22989 107173 23055 107174
rect 23533 107174 23534 107206
rect 23598 107206 23604 107238
rect 115192 107446 115198 107478
rect 115262 107478 115263 107510
rect 115605 107510 115671 107511
rect 115605 107478 115606 107510
rect 115262 107446 115268 107478
rect 115192 107238 115268 107446
rect 23598 107174 23599 107206
rect 23533 107173 23599 107174
rect 115192 107174 115198 107238
rect 115262 107174 115268 107238
rect 115192 107168 115268 107174
rect 115600 107446 115606 107478
rect 115670 107478 115671 107510
rect 116008 107510 116084 107516
rect 115670 107446 115676 107478
rect 115600 107238 115676 107446
rect 115600 107174 115606 107238
rect 115670 107174 115676 107238
rect 116008 107446 116014 107510
rect 116078 107446 116084 107510
rect 116965 107510 117031 107511
rect 116965 107478 116966 107510
rect 116008 107238 116084 107446
rect 116008 107206 116014 107238
rect 115600 107168 115676 107174
rect 116013 107174 116014 107206
rect 116078 107206 116084 107238
rect 116960 107446 116966 107478
rect 117030 107478 117031 107510
rect 117030 107446 117036 107478
rect 116960 107238 117036 107446
rect 116078 107174 116079 107206
rect 116013 107173 116079 107174
rect 116960 107174 116966 107238
rect 117030 107174 117036 107238
rect 116960 107168 117036 107174
rect 22173 107102 22239 107103
rect 22173 107070 22174 107102
rect 22168 107038 22174 107070
rect 22238 107070 22239 107102
rect 22581 107102 22647 107103
rect 22581 107070 22582 107102
rect 22238 107038 22244 107070
rect 22168 106830 22244 107038
rect 22168 106766 22174 106830
rect 22238 106766 22244 106830
rect 22168 106760 22244 106766
rect 22576 107038 22582 107070
rect 22646 107070 22647 107102
rect 23120 107102 23196 107108
rect 22646 107038 22652 107070
rect 22576 106830 22652 107038
rect 22576 106766 22582 106830
rect 22646 106766 22652 106830
rect 23120 107038 23126 107102
rect 23190 107038 23196 107102
rect 23120 106830 23196 107038
rect 23120 106798 23126 106830
rect 22576 106760 22652 106766
rect 23125 106766 23126 106798
rect 23190 106798 23196 106830
rect 23528 107102 23604 107108
rect 23528 107038 23534 107102
rect 23598 107038 23604 107102
rect 23528 106830 23604 107038
rect 23528 106798 23534 106830
rect 23190 106766 23191 106798
rect 23125 106765 23191 106766
rect 23533 106766 23534 106798
rect 23598 106798 23604 106830
rect 115192 107102 115268 107108
rect 115192 107038 115198 107102
rect 115262 107038 115268 107102
rect 115741 107102 115807 107103
rect 115741 107070 115742 107102
rect 115192 106830 115268 107038
rect 115192 106798 115198 106830
rect 23598 106766 23599 106798
rect 23533 106765 23599 106766
rect 115197 106766 115198 106798
rect 115262 106798 115268 106830
rect 115736 107038 115742 107070
rect 115806 107070 115807 107102
rect 116013 107102 116079 107103
rect 116013 107070 116014 107102
rect 115806 107038 115812 107070
rect 115736 106830 115812 107038
rect 115262 106766 115263 106798
rect 115197 106765 115263 106766
rect 115736 106766 115742 106830
rect 115806 106766 115812 106830
rect 115736 106760 115812 106766
rect 116008 107038 116014 107070
rect 116078 107070 116079 107102
rect 116078 107038 116084 107070
rect 116008 106830 116084 107038
rect 116008 106766 116014 106830
rect 116078 106766 116084 106830
rect 116008 106760 116084 106766
rect 21901 106694 21967 106695
rect 21901 106662 21902 106694
rect 21896 106630 21902 106662
rect 21966 106662 21967 106694
rect 22712 106694 22788 106700
rect 21966 106630 21972 106662
rect 21896 106422 21972 106630
rect 21896 106358 21902 106422
rect 21966 106358 21972 106422
rect 22712 106630 22718 106694
rect 22782 106630 22788 106694
rect 22712 106422 22788 106630
rect 22712 106390 22718 106422
rect 21896 106352 21972 106358
rect 22717 106358 22718 106390
rect 22782 106390 22788 106422
rect 23120 106694 23196 106700
rect 23120 106630 23126 106694
rect 23190 106630 23196 106694
rect 23397 106694 23463 106695
rect 23397 106662 23398 106694
rect 23120 106422 23196 106630
rect 23120 106390 23126 106422
rect 22782 106358 22783 106390
rect 22717 106357 22783 106358
rect 23125 106358 23126 106390
rect 23190 106390 23196 106422
rect 23392 106630 23398 106662
rect 23462 106662 23463 106694
rect 115197 106694 115263 106695
rect 115197 106662 115198 106694
rect 23462 106630 23468 106662
rect 23392 106422 23468 106630
rect 23190 106358 23191 106390
rect 23125 106357 23191 106358
rect 23392 106358 23398 106422
rect 23462 106358 23468 106422
rect 23392 106352 23468 106358
rect 115192 106630 115198 106662
rect 115262 106662 115263 106694
rect 115600 106694 115676 106700
rect 115262 106630 115268 106662
rect 115192 106422 115268 106630
rect 115192 106358 115198 106422
rect 115262 106358 115268 106422
rect 115600 106630 115606 106694
rect 115670 106630 115676 106694
rect 115600 106422 115676 106630
rect 115600 106390 115606 106422
rect 115192 106352 115268 106358
rect 115605 106358 115606 106390
rect 115670 106390 115676 106422
rect 116552 106694 116628 106700
rect 116552 106630 116558 106694
rect 116622 106630 116628 106694
rect 116552 106422 116628 106630
rect 116552 106390 116558 106422
rect 115670 106358 115671 106390
rect 115605 106357 115671 106358
rect 116557 106358 116558 106390
rect 116622 106390 116628 106422
rect 116960 106694 117036 106700
rect 116960 106630 116966 106694
rect 117030 106630 117036 106694
rect 116960 106422 117036 106630
rect 116960 106390 116966 106422
rect 116622 106358 116623 106390
rect 116557 106357 116623 106358
rect 116965 106358 116966 106390
rect 117030 106390 117036 106422
rect 117030 106358 117031 106390
rect 116965 106357 117031 106358
rect 22445 106286 22511 106287
rect 22445 106254 22446 106286
rect 952 106086 1230 106150
rect 1294 106086 1300 106150
rect 952 104654 1300 106086
rect 22440 106222 22446 106254
rect 22510 106254 22511 106286
rect 23125 106286 23191 106287
rect 23125 106254 23126 106286
rect 22510 106222 22516 106254
rect 21760 106014 21836 106020
rect 21760 105950 21766 106014
rect 21830 105950 21836 106014
rect 21760 105742 21836 105950
rect 22440 106014 22516 106222
rect 22440 105950 22446 106014
rect 22510 105950 22516 106014
rect 22440 105944 22516 105950
rect 23120 106222 23126 106254
rect 23190 106254 23191 106286
rect 23528 106286 23604 106292
rect 23190 106222 23196 106254
rect 23120 106014 23196 106222
rect 23120 105950 23126 106014
rect 23190 105950 23196 106014
rect 23528 106222 23534 106286
rect 23598 106222 23604 106286
rect 23528 106014 23604 106222
rect 115328 106286 115404 106292
rect 115328 106222 115334 106286
rect 115398 106222 115404 106286
rect 110301 106150 110367 106151
rect 110301 106118 110302 106150
rect 23528 105982 23534 106014
rect 23120 105944 23196 105950
rect 23533 105950 23534 105982
rect 23598 105982 23604 106014
rect 110296 106086 110302 106118
rect 110366 106118 110367 106150
rect 110366 106086 110372 106118
rect 23598 105950 23599 105982
rect 23533 105949 23599 105950
rect 21760 105710 21766 105742
rect 21765 105678 21766 105710
rect 21830 105710 21836 105742
rect 22984 105878 23060 105884
rect 22984 105814 22990 105878
rect 23054 105814 23060 105878
rect 23533 105878 23599 105879
rect 23533 105846 23534 105878
rect 21830 105678 21831 105710
rect 21765 105677 21831 105678
rect 22984 105606 23060 105814
rect 22984 105574 22990 105606
rect 22989 105542 22990 105574
rect 23054 105574 23060 105606
rect 23528 105814 23534 105846
rect 23598 105846 23599 105878
rect 110296 105878 110372 106086
rect 115328 106014 115404 106222
rect 115328 105982 115334 106014
rect 115333 105950 115334 105982
rect 115398 105982 115404 106014
rect 115736 106286 115812 106292
rect 115736 106222 115742 106286
rect 115806 106222 115812 106286
rect 115736 106014 115812 106222
rect 137496 106286 137844 107990
rect 137496 106222 137502 106286
rect 137566 106222 137844 106286
rect 115736 105982 115742 106014
rect 115398 105950 115399 105982
rect 115333 105949 115399 105950
rect 115741 105950 115742 105982
rect 115806 105982 115812 106014
rect 116829 106014 116895 106015
rect 116829 105982 116830 106014
rect 115806 105950 115807 105982
rect 115741 105949 115807 105950
rect 116824 105950 116830 105982
rect 116894 105982 116895 106014
rect 116894 105950 116900 105982
rect 23598 105814 23604 105846
rect 23528 105606 23604 105814
rect 110296 105814 110302 105878
rect 110366 105814 110372 105878
rect 115333 105878 115399 105879
rect 115333 105846 115334 105878
rect 110296 105808 110372 105814
rect 115328 105814 115334 105846
rect 115398 105846 115399 105878
rect 115741 105878 115807 105879
rect 115741 105846 115742 105878
rect 115398 105814 115404 105846
rect 23054 105542 23055 105574
rect 22989 105541 23055 105542
rect 23528 105542 23534 105606
rect 23598 105542 23604 105606
rect 23528 105536 23604 105542
rect 115328 105606 115404 105814
rect 115328 105542 115334 105606
rect 115398 105542 115404 105606
rect 115328 105536 115404 105542
rect 115736 105814 115742 105846
rect 115806 105846 115807 105878
rect 115806 105814 115812 105846
rect 115736 105606 115812 105814
rect 116824 105742 116900 105950
rect 116824 105678 116830 105742
rect 116894 105678 116900 105742
rect 116824 105672 116900 105678
rect 115736 105542 115742 105606
rect 115806 105542 115812 105606
rect 115736 105536 115812 105542
rect 22309 105470 22375 105471
rect 22309 105438 22310 105470
rect 22304 105406 22310 105438
rect 22374 105438 22375 105470
rect 22445 105470 22511 105471
rect 22445 105438 22446 105470
rect 22374 105406 22380 105438
rect 21901 105198 21967 105199
rect 21901 105166 21902 105198
rect 21896 105134 21902 105166
rect 21966 105166 21967 105198
rect 22304 105198 22380 105406
rect 21966 105134 21972 105166
rect 21896 104926 21972 105134
rect 22304 105134 22310 105198
rect 22374 105134 22380 105198
rect 22304 105128 22380 105134
rect 22440 105406 22446 105438
rect 22510 105438 22511 105470
rect 116421 105470 116487 105471
rect 116421 105438 116422 105470
rect 22510 105406 22516 105438
rect 22440 105198 22516 105406
rect 22440 105134 22446 105198
rect 22510 105134 22516 105198
rect 22440 105128 22516 105134
rect 116416 105406 116422 105438
rect 116486 105438 116487 105470
rect 116486 105406 116492 105438
rect 116416 105198 116492 105406
rect 116416 105134 116422 105198
rect 116486 105134 116492 105198
rect 116965 105198 117031 105199
rect 116965 105166 116966 105198
rect 116416 105128 116492 105134
rect 116960 105134 116966 105166
rect 117030 105166 117031 105198
rect 117030 105134 117036 105166
rect 28293 105062 28359 105063
rect 28293 105030 28294 105062
rect 21896 104862 21902 104926
rect 21966 104862 21972 104926
rect 21896 104856 21972 104862
rect 28288 104998 28294 105030
rect 28358 105030 28359 105062
rect 28358 104998 28364 105030
rect 952 104590 1230 104654
rect 1294 104590 1300 104654
rect 952 102750 1300 104590
rect 21896 104790 21972 104796
rect 21896 104726 21902 104790
rect 21966 104726 21972 104790
rect 22581 104790 22647 104791
rect 22581 104758 22582 104790
rect 21896 104518 21972 104726
rect 21896 104486 21902 104518
rect 21901 104454 21902 104486
rect 21966 104486 21972 104518
rect 22576 104726 22582 104758
rect 22646 104758 22647 104790
rect 22984 104790 23060 104796
rect 22646 104726 22652 104758
rect 22576 104518 22652 104726
rect 21966 104454 21967 104486
rect 21901 104453 21967 104454
rect 22576 104454 22582 104518
rect 22646 104454 22652 104518
rect 22984 104726 22990 104790
rect 23054 104726 23060 104790
rect 23533 104790 23599 104791
rect 23533 104758 23534 104790
rect 22984 104518 23060 104726
rect 22984 104486 22990 104518
rect 22576 104448 22652 104454
rect 22989 104454 22990 104486
rect 23054 104486 23060 104518
rect 23528 104726 23534 104758
rect 23598 104758 23599 104790
rect 28288 104790 28364 104998
rect 23598 104726 23604 104758
rect 23528 104518 23604 104726
rect 28288 104726 28294 104790
rect 28358 104726 28364 104790
rect 28288 104720 28364 104726
rect 28560 104926 28636 104932
rect 28560 104862 28566 104926
rect 28630 104862 28636 104926
rect 23054 104454 23055 104486
rect 22989 104453 23055 104454
rect 23528 104454 23534 104518
rect 23598 104454 23604 104518
rect 28429 104518 28495 104519
rect 28429 104486 28430 104518
rect 23528 104448 23604 104454
rect 28424 104454 28430 104486
rect 28494 104486 28495 104518
rect 28560 104518 28636 104862
rect 116960 104926 117036 105134
rect 116960 104862 116966 104926
rect 117030 104862 117036 104926
rect 116960 104856 117036 104862
rect 28560 104486 28566 104518
rect 28494 104454 28500 104486
rect 21896 104382 21972 104388
rect 21896 104318 21902 104382
rect 21966 104318 21972 104382
rect 22989 104382 23055 104383
rect 22989 104350 22990 104382
rect 21896 104110 21972 104318
rect 21896 104078 21902 104110
rect 21901 104046 21902 104078
rect 21966 104078 21972 104110
rect 22984 104318 22990 104350
rect 23054 104350 23055 104382
rect 23397 104382 23463 104383
rect 23397 104350 23398 104382
rect 23054 104318 23060 104350
rect 22984 104110 23060 104318
rect 21966 104046 21967 104078
rect 21901 104045 21967 104046
rect 22984 104046 22990 104110
rect 23054 104046 23060 104110
rect 22984 104040 23060 104046
rect 23392 104318 23398 104350
rect 23462 104350 23463 104382
rect 23462 104318 23468 104350
rect 23392 104110 23468 104318
rect 28424 104246 28500 104454
rect 28565 104454 28566 104486
rect 28630 104486 28636 104518
rect 115192 104790 115268 104796
rect 115192 104726 115198 104790
rect 115262 104726 115268 104790
rect 115192 104518 115268 104726
rect 115192 104486 115198 104518
rect 28630 104454 28631 104486
rect 28565 104453 28631 104454
rect 115197 104454 115198 104486
rect 115262 104486 115268 104518
rect 115600 104790 115676 104796
rect 115600 104726 115606 104790
rect 115670 104726 115676 104790
rect 116013 104790 116079 104791
rect 116013 104758 116014 104790
rect 115600 104518 115676 104726
rect 115600 104486 115606 104518
rect 115262 104454 115263 104486
rect 115197 104453 115263 104454
rect 115605 104454 115606 104486
rect 115670 104486 115676 104518
rect 116008 104726 116014 104758
rect 116078 104758 116079 104790
rect 116960 104790 117036 104796
rect 116078 104726 116084 104758
rect 116008 104518 116084 104726
rect 115670 104454 115671 104486
rect 115605 104453 115671 104454
rect 116008 104454 116014 104518
rect 116078 104454 116084 104518
rect 116960 104726 116966 104790
rect 117030 104726 117036 104790
rect 116960 104518 117036 104726
rect 116960 104486 116966 104518
rect 116008 104448 116084 104454
rect 116965 104454 116966 104486
rect 117030 104486 117036 104518
rect 137496 104518 137844 106222
rect 117030 104454 117031 104486
rect 116965 104453 117031 104454
rect 137496 104454 137502 104518
rect 137566 104454 137844 104518
rect 28424 104182 28430 104246
rect 28494 104182 28500 104246
rect 28424 104176 28500 104182
rect 115192 104382 115268 104388
rect 115192 104318 115198 104382
rect 115262 104318 115268 104382
rect 115605 104382 115671 104383
rect 115605 104350 115606 104382
rect 23392 104046 23398 104110
rect 23462 104046 23468 104110
rect 115192 104110 115268 104318
rect 115192 104078 115198 104110
rect 23392 104040 23468 104046
rect 115197 104046 115198 104078
rect 115262 104078 115268 104110
rect 115600 104318 115606 104350
rect 115670 104350 115671 104382
rect 116144 104382 116220 104388
rect 115670 104318 115676 104350
rect 115600 104110 115676 104318
rect 115262 104046 115263 104078
rect 115197 104045 115263 104046
rect 115600 104046 115606 104110
rect 115670 104046 115676 104110
rect 116144 104318 116150 104382
rect 116214 104318 116220 104382
rect 116965 104382 117031 104383
rect 116965 104350 116966 104382
rect 116144 104110 116220 104318
rect 116144 104078 116150 104110
rect 115600 104040 115676 104046
rect 116149 104046 116150 104078
rect 116214 104078 116220 104110
rect 116960 104318 116966 104350
rect 117030 104350 117031 104382
rect 117030 104318 117036 104350
rect 116960 104110 117036 104318
rect 116214 104046 116215 104078
rect 116149 104045 116215 104046
rect 116960 104046 116966 104110
rect 117030 104046 117036 104110
rect 116960 104040 117036 104046
rect 21760 103974 21836 103980
rect 21760 103910 21766 103974
rect 21830 103910 21836 103974
rect 22173 103974 22239 103975
rect 22173 103942 22174 103974
rect 21760 103702 21836 103910
rect 21760 103670 21766 103702
rect 21765 103638 21766 103670
rect 21830 103670 21836 103702
rect 22168 103910 22174 103942
rect 22238 103942 22239 103974
rect 23120 103974 23196 103980
rect 22238 103910 22244 103942
rect 22168 103702 22244 103910
rect 21830 103638 21831 103670
rect 21765 103637 21831 103638
rect 22168 103638 22174 103702
rect 22238 103638 22244 103702
rect 23120 103910 23126 103974
rect 23190 103910 23196 103974
rect 23120 103702 23196 103910
rect 23120 103670 23126 103702
rect 22168 103632 22244 103638
rect 23125 103638 23126 103670
rect 23190 103670 23196 103702
rect 23528 103974 23604 103980
rect 23528 103910 23534 103974
rect 23598 103910 23604 103974
rect 23528 103702 23604 103910
rect 23528 103670 23534 103702
rect 23190 103638 23191 103670
rect 23125 103637 23191 103638
rect 23533 103638 23534 103670
rect 23598 103670 23604 103702
rect 115328 103974 115404 103980
rect 115328 103910 115334 103974
rect 115398 103910 115404 103974
rect 115741 103974 115807 103975
rect 115741 103942 115742 103974
rect 115328 103702 115404 103910
rect 115328 103670 115334 103702
rect 23598 103638 23599 103670
rect 23533 103637 23599 103638
rect 115333 103638 115334 103670
rect 115398 103670 115404 103702
rect 115736 103910 115742 103942
rect 115806 103942 115807 103974
rect 116013 103974 116079 103975
rect 116013 103942 116014 103974
rect 115806 103910 115812 103942
rect 115736 103702 115812 103910
rect 115398 103638 115399 103670
rect 115333 103637 115399 103638
rect 115736 103638 115742 103702
rect 115806 103638 115812 103702
rect 115736 103632 115812 103638
rect 116008 103910 116014 103942
rect 116078 103942 116079 103974
rect 116829 103974 116895 103975
rect 116829 103942 116830 103974
rect 116078 103910 116084 103942
rect 116008 103702 116084 103910
rect 116008 103638 116014 103702
rect 116078 103638 116084 103702
rect 116008 103632 116084 103638
rect 116824 103910 116830 103942
rect 116894 103942 116895 103974
rect 116894 103910 116900 103942
rect 116824 103702 116900 103910
rect 116824 103638 116830 103702
rect 116894 103638 116900 103702
rect 116824 103632 116900 103638
rect 21765 103566 21831 103567
rect 21765 103534 21766 103566
rect 21760 103502 21766 103534
rect 21830 103534 21831 103566
rect 22304 103566 22380 103572
rect 21830 103502 21836 103534
rect 21760 103294 21836 103502
rect 21760 103230 21766 103294
rect 21830 103230 21836 103294
rect 22304 103502 22310 103566
rect 22374 103502 22380 103566
rect 23125 103566 23191 103567
rect 23125 103534 23126 103566
rect 22304 103294 22380 103502
rect 22304 103262 22310 103294
rect 21760 103224 21836 103230
rect 22309 103230 22310 103262
rect 22374 103262 22380 103294
rect 23120 103502 23126 103534
rect 23190 103534 23191 103566
rect 23392 103566 23468 103572
rect 23190 103502 23196 103534
rect 23120 103294 23196 103502
rect 22374 103230 22375 103262
rect 22309 103229 22375 103230
rect 23120 103230 23126 103294
rect 23190 103230 23196 103294
rect 23392 103502 23398 103566
rect 23462 103502 23468 103566
rect 115333 103566 115399 103567
rect 115333 103534 115334 103566
rect 23392 103294 23468 103502
rect 23392 103262 23398 103294
rect 23120 103224 23196 103230
rect 23397 103230 23398 103262
rect 23462 103262 23468 103294
rect 115328 103502 115334 103534
rect 115398 103534 115399 103566
rect 115741 103566 115807 103567
rect 115741 103534 115742 103566
rect 115398 103502 115404 103534
rect 115328 103294 115404 103502
rect 23462 103230 23463 103262
rect 23397 103229 23463 103230
rect 115328 103230 115334 103294
rect 115398 103230 115404 103294
rect 115328 103224 115404 103230
rect 115736 103502 115742 103534
rect 115806 103534 115807 103566
rect 116285 103566 116351 103567
rect 116285 103534 116286 103566
rect 115806 103502 115812 103534
rect 115736 103294 115812 103502
rect 115736 103230 115742 103294
rect 115806 103230 115812 103294
rect 115736 103224 115812 103230
rect 116280 103502 116286 103534
rect 116350 103534 116351 103566
rect 116829 103566 116895 103567
rect 116829 103534 116830 103566
rect 116350 103502 116356 103534
rect 116280 103294 116356 103502
rect 116280 103230 116286 103294
rect 116350 103230 116356 103294
rect 116280 103224 116356 103230
rect 116824 103502 116830 103534
rect 116894 103534 116895 103566
rect 116894 103502 116900 103534
rect 116824 103294 116900 103502
rect 116824 103230 116830 103294
rect 116894 103230 116900 103294
rect 116824 103224 116900 103230
rect 21901 103158 21967 103159
rect 21901 103126 21902 103158
rect 21896 103094 21902 103126
rect 21966 103126 21967 103158
rect 22168 103158 22244 103164
rect 21966 103094 21972 103126
rect 21896 102886 21972 103094
rect 21896 102822 21902 102886
rect 21966 102822 21972 102886
rect 22168 103094 22174 103158
rect 22238 103094 22244 103158
rect 22445 103158 22511 103159
rect 22445 103126 22446 103158
rect 22168 102886 22244 103094
rect 22168 102854 22174 102886
rect 21896 102816 21972 102822
rect 22173 102822 22174 102854
rect 22238 102854 22244 102886
rect 22440 103094 22446 103126
rect 22510 103126 22511 103158
rect 22989 103158 23055 103159
rect 22989 103126 22990 103158
rect 22510 103094 22516 103126
rect 22440 102886 22516 103094
rect 22238 102822 22239 102854
rect 22173 102821 22239 102822
rect 22440 102822 22446 102886
rect 22510 102822 22516 102886
rect 22440 102816 22516 102822
rect 22984 103094 22990 103126
rect 23054 103126 23055 103158
rect 23397 103158 23463 103159
rect 23397 103126 23398 103158
rect 23054 103094 23060 103126
rect 22984 102886 23060 103094
rect 22984 102822 22990 102886
rect 23054 102822 23060 102886
rect 22984 102816 23060 102822
rect 23392 103094 23398 103126
rect 23462 103126 23463 103158
rect 115328 103158 115404 103164
rect 23462 103094 23468 103126
rect 23392 102886 23468 103094
rect 23392 102822 23398 102886
rect 23462 102822 23468 102886
rect 115328 103094 115334 103158
rect 115398 103094 115404 103158
rect 115328 102886 115404 103094
rect 115328 102854 115334 102886
rect 23392 102816 23468 102822
rect 115333 102822 115334 102854
rect 115398 102854 115404 102886
rect 115736 103158 115812 103164
rect 115736 103094 115742 103158
rect 115806 103094 115812 103158
rect 116965 103158 117031 103159
rect 116965 103126 116966 103158
rect 115736 102886 115812 103094
rect 115736 102854 115742 102886
rect 115398 102822 115399 102854
rect 115333 102821 115399 102822
rect 115741 102822 115742 102854
rect 115806 102854 115812 102886
rect 116960 103094 116966 103126
rect 117030 103126 117031 103158
rect 117030 103094 117036 103126
rect 116960 102886 117036 103094
rect 115806 102822 115807 102854
rect 115741 102821 115807 102822
rect 116960 102822 116966 102886
rect 117030 102822 117036 102886
rect 116960 102816 117036 102822
rect 137496 102886 137844 104454
rect 137496 102822 137502 102886
rect 137566 102822 137844 102886
rect 952 102686 1230 102750
rect 1294 102686 1300 102750
rect 952 101254 1300 102686
rect 21760 102750 21836 102756
rect 21760 102686 21766 102750
rect 21830 102686 21836 102750
rect 22581 102750 22647 102751
rect 22581 102718 22582 102750
rect 21760 102478 21836 102686
rect 21760 102446 21766 102478
rect 21765 102414 21766 102446
rect 21830 102446 21836 102478
rect 22576 102686 22582 102718
rect 22646 102718 22647 102750
rect 23120 102750 23196 102756
rect 22646 102686 22652 102718
rect 22576 102478 22652 102686
rect 21830 102414 21831 102446
rect 21765 102413 21831 102414
rect 22576 102414 22582 102478
rect 22646 102414 22652 102478
rect 23120 102686 23126 102750
rect 23190 102686 23196 102750
rect 23120 102478 23196 102686
rect 23120 102446 23126 102478
rect 22576 102408 22652 102414
rect 23125 102414 23126 102446
rect 23190 102446 23196 102478
rect 23528 102750 23604 102756
rect 23528 102686 23534 102750
rect 23598 102686 23604 102750
rect 23528 102478 23604 102686
rect 23528 102446 23534 102478
rect 23190 102414 23191 102446
rect 23125 102413 23191 102414
rect 23533 102414 23534 102446
rect 23598 102446 23604 102478
rect 115192 102750 115268 102756
rect 115192 102686 115198 102750
rect 115262 102686 115268 102750
rect 115741 102750 115807 102751
rect 115741 102718 115742 102750
rect 115192 102478 115268 102686
rect 115192 102446 115198 102478
rect 23598 102414 23599 102446
rect 23533 102413 23599 102414
rect 115197 102414 115198 102446
rect 115262 102446 115268 102478
rect 115736 102686 115742 102718
rect 115806 102718 115807 102750
rect 116144 102750 116220 102756
rect 115806 102686 115812 102718
rect 115736 102478 115812 102686
rect 115262 102414 115263 102446
rect 115197 102413 115263 102414
rect 115736 102414 115742 102478
rect 115806 102414 115812 102478
rect 116144 102686 116150 102750
rect 116214 102686 116220 102750
rect 116421 102750 116487 102751
rect 116421 102718 116422 102750
rect 116144 102478 116220 102686
rect 116144 102446 116150 102478
rect 115736 102408 115812 102414
rect 116149 102414 116150 102446
rect 116214 102446 116220 102478
rect 116416 102686 116422 102718
rect 116486 102718 116487 102750
rect 116824 102750 116900 102756
rect 116486 102686 116492 102718
rect 116416 102478 116492 102686
rect 116214 102414 116215 102446
rect 116149 102413 116215 102414
rect 116416 102414 116422 102478
rect 116486 102414 116492 102478
rect 116824 102686 116830 102750
rect 116894 102686 116900 102750
rect 116824 102478 116900 102686
rect 116824 102446 116830 102478
rect 116416 102408 116492 102414
rect 116829 102414 116830 102446
rect 116894 102446 116900 102478
rect 116894 102414 116895 102446
rect 116829 102413 116895 102414
rect 22309 102342 22375 102343
rect 22309 102310 22310 102342
rect 22304 102278 22310 102310
rect 22374 102310 22375 102342
rect 22712 102342 22788 102348
rect 22374 102278 22380 102310
rect 21760 102070 21836 102076
rect 21760 102006 21766 102070
rect 21830 102006 21836 102070
rect 21760 101798 21836 102006
rect 22304 102070 22380 102278
rect 22712 102278 22718 102342
rect 22782 102278 22788 102342
rect 22989 102342 23055 102343
rect 22989 102310 22990 102342
rect 22304 102006 22310 102070
rect 22374 102006 22380 102070
rect 22445 102070 22511 102071
rect 22445 102038 22446 102070
rect 22304 102000 22380 102006
rect 22440 102006 22446 102038
rect 22510 102038 22511 102070
rect 22712 102070 22788 102278
rect 22712 102038 22718 102070
rect 22510 102006 22516 102038
rect 21760 101766 21766 101798
rect 21765 101734 21766 101766
rect 21830 101766 21836 101798
rect 22440 101798 22516 102006
rect 22717 102006 22718 102038
rect 22782 102038 22788 102070
rect 22984 102278 22990 102310
rect 23054 102310 23055 102342
rect 23397 102342 23463 102343
rect 23397 102310 23398 102342
rect 23054 102278 23060 102310
rect 22984 102070 23060 102278
rect 22782 102006 22783 102038
rect 22717 102005 22783 102006
rect 22984 102006 22990 102070
rect 23054 102006 23060 102070
rect 22984 102000 23060 102006
rect 23392 102278 23398 102310
rect 23462 102310 23463 102342
rect 115192 102342 115268 102348
rect 23462 102278 23468 102310
rect 23392 102070 23468 102278
rect 23392 102006 23398 102070
rect 23462 102006 23468 102070
rect 115192 102278 115198 102342
rect 115262 102278 115268 102342
rect 115192 102070 115268 102278
rect 115192 102038 115198 102070
rect 23392 102000 23468 102006
rect 115197 102006 115198 102038
rect 115262 102038 115268 102070
rect 115600 102342 115676 102348
rect 115600 102278 115606 102342
rect 115670 102278 115676 102342
rect 115600 102070 115676 102278
rect 115600 102038 115606 102070
rect 115262 102006 115263 102038
rect 115197 102005 115263 102006
rect 115605 102006 115606 102038
rect 115670 102038 115676 102070
rect 116552 102342 116628 102348
rect 116552 102278 116558 102342
rect 116622 102278 116628 102342
rect 116552 102070 116628 102278
rect 116552 102038 116558 102070
rect 115670 102006 115671 102038
rect 115605 102005 115671 102006
rect 116557 102006 116558 102038
rect 116622 102038 116628 102070
rect 116960 102070 117036 102076
rect 116622 102006 116623 102038
rect 116557 102005 116623 102006
rect 116960 102006 116966 102070
rect 117030 102006 117036 102070
rect 23125 101934 23191 101935
rect 23125 101902 23126 101934
rect 21830 101734 21831 101766
rect 21765 101733 21831 101734
rect 22440 101734 22446 101798
rect 22510 101734 22516 101798
rect 22440 101728 22516 101734
rect 23120 101870 23126 101902
rect 23190 101902 23191 101934
rect 23528 101934 23604 101940
rect 23190 101870 23196 101902
rect 23120 101662 23196 101870
rect 23120 101598 23126 101662
rect 23190 101598 23196 101662
rect 23528 101870 23534 101934
rect 23598 101870 23604 101934
rect 115197 101934 115263 101935
rect 115197 101902 115198 101934
rect 23528 101662 23604 101870
rect 115192 101870 115198 101902
rect 115262 101902 115263 101934
rect 115605 101934 115671 101935
rect 115605 101902 115606 101934
rect 115262 101870 115268 101902
rect 23528 101630 23534 101662
rect 23120 101592 23196 101598
rect 23533 101598 23534 101630
rect 23598 101630 23604 101662
rect 28293 101662 28359 101663
rect 28293 101630 28294 101662
rect 23598 101598 23599 101630
rect 23533 101597 23599 101598
rect 28288 101598 28294 101630
rect 28358 101630 28359 101662
rect 115192 101662 115268 101870
rect 28358 101598 28364 101630
rect 22712 101526 22788 101532
rect 22712 101462 22718 101526
rect 22782 101462 22788 101526
rect 952 101190 1230 101254
rect 1294 101190 1300 101254
rect 21901 101254 21967 101255
rect 21901 101222 21902 101254
rect 952 99622 1300 101190
rect 21896 101190 21902 101222
rect 21966 101222 21967 101254
rect 22712 101254 22788 101462
rect 28288 101390 28364 101598
rect 115192 101598 115198 101662
rect 115262 101598 115268 101662
rect 115192 101592 115268 101598
rect 115600 101870 115606 101902
rect 115670 101902 115671 101934
rect 115670 101870 115676 101902
rect 115600 101662 115676 101870
rect 116960 101798 117036 102006
rect 116960 101766 116966 101798
rect 116965 101734 116966 101766
rect 117030 101766 117036 101798
rect 117030 101734 117031 101766
rect 116965 101733 117031 101734
rect 115600 101598 115606 101662
rect 115670 101598 115676 101662
rect 115600 101592 115676 101598
rect 116280 101526 116356 101532
rect 116280 101462 116286 101526
rect 116350 101462 116356 101526
rect 28288 101326 28294 101390
rect 28358 101326 28364 101390
rect 28565 101390 28631 101391
rect 28565 101358 28566 101390
rect 28288 101320 28364 101326
rect 28560 101326 28566 101358
rect 28630 101358 28631 101390
rect 110160 101390 110236 101396
rect 28630 101326 28636 101358
rect 22712 101222 22718 101254
rect 21966 101190 21972 101222
rect 21896 100982 21972 101190
rect 22717 101190 22718 101222
rect 22782 101222 22788 101254
rect 22782 101190 22783 101222
rect 22717 101189 22783 101190
rect 28560 101118 28636 101326
rect 28560 101054 28566 101118
rect 28630 101054 28636 101118
rect 110160 101326 110166 101390
rect 110230 101326 110236 101390
rect 110160 101118 110236 101326
rect 116280 101254 116356 101462
rect 116280 101222 116286 101254
rect 116285 101190 116286 101222
rect 116350 101222 116356 101254
rect 116960 101254 117036 101260
rect 116350 101190 116351 101222
rect 116285 101189 116351 101190
rect 116960 101190 116966 101254
rect 117030 101190 117036 101254
rect 110160 101086 110166 101118
rect 28560 101048 28636 101054
rect 110165 101054 110166 101086
rect 110230 101086 110236 101118
rect 110230 101054 110231 101086
rect 110165 101053 110231 101054
rect 21896 100918 21902 100982
rect 21966 100918 21972 100982
rect 21896 100912 21972 100918
rect 28288 100982 28364 100988
rect 28288 100918 28294 100982
rect 28358 100918 28364 100982
rect 21760 100846 21836 100852
rect 21760 100782 21766 100846
rect 21830 100782 21836 100846
rect 22445 100846 22511 100847
rect 22445 100814 22446 100846
rect 21760 100574 21836 100782
rect 21760 100542 21766 100574
rect 21765 100510 21766 100542
rect 21830 100542 21836 100574
rect 22440 100782 22446 100814
rect 22510 100814 22511 100846
rect 22510 100782 22516 100814
rect 22440 100574 22516 100782
rect 28288 100710 28364 100918
rect 28288 100678 28294 100710
rect 28293 100646 28294 100678
rect 28358 100678 28364 100710
rect 110296 100982 110372 100988
rect 110296 100918 110302 100982
rect 110366 100918 110372 100982
rect 116960 100982 117036 101190
rect 116960 100950 116966 100982
rect 110296 100710 110372 100918
rect 116965 100918 116966 100950
rect 117030 100950 117036 100982
rect 137496 101254 137844 102822
rect 137496 101190 137502 101254
rect 137566 101190 137844 101254
rect 117030 100918 117031 100950
rect 116965 100917 117031 100918
rect 116149 100846 116215 100847
rect 116149 100814 116150 100846
rect 110296 100678 110302 100710
rect 28358 100646 28359 100678
rect 28293 100645 28359 100646
rect 110301 100646 110302 100678
rect 110366 100678 110372 100710
rect 116144 100782 116150 100814
rect 116214 100814 116215 100846
rect 116416 100846 116492 100852
rect 116214 100782 116220 100814
rect 110366 100646 110367 100678
rect 110301 100645 110367 100646
rect 21830 100510 21831 100542
rect 21765 100509 21831 100510
rect 22440 100510 22446 100574
rect 22510 100510 22516 100574
rect 110301 100574 110367 100575
rect 110301 100542 110302 100574
rect 22440 100504 22516 100510
rect 110296 100510 110302 100542
rect 110366 100542 110367 100574
rect 116144 100574 116220 100782
rect 110366 100510 110372 100542
rect 21765 100438 21831 100439
rect 21765 100406 21766 100438
rect 21760 100374 21766 100406
rect 21830 100406 21831 100438
rect 22984 100438 23060 100444
rect 21830 100374 21836 100406
rect 21760 100166 21836 100374
rect 21760 100102 21766 100166
rect 21830 100102 21836 100166
rect 22984 100374 22990 100438
rect 23054 100374 23060 100438
rect 22984 100166 23060 100374
rect 22984 100134 22990 100166
rect 21760 100096 21836 100102
rect 22989 100102 22990 100134
rect 23054 100134 23060 100166
rect 23392 100438 23468 100444
rect 23392 100374 23398 100438
rect 23462 100374 23468 100438
rect 28429 100438 28495 100439
rect 28429 100406 28430 100438
rect 23392 100166 23468 100374
rect 23392 100134 23398 100166
rect 23054 100102 23055 100134
rect 22989 100101 23055 100102
rect 23397 100102 23398 100134
rect 23462 100134 23468 100166
rect 28424 100374 28430 100406
rect 28494 100406 28495 100438
rect 28494 100374 28500 100406
rect 23462 100102 23463 100134
rect 23397 100101 23463 100102
rect 21901 100030 21967 100031
rect 21901 99998 21902 100030
rect 21896 99966 21902 99998
rect 21966 99998 21967 100030
rect 22168 100030 22244 100036
rect 21966 99966 21972 99998
rect 21896 99758 21972 99966
rect 21896 99694 21902 99758
rect 21966 99694 21972 99758
rect 22168 99966 22174 100030
rect 22238 99966 22244 100030
rect 22989 100030 23055 100031
rect 22989 99998 22990 100030
rect 22168 99758 22244 99966
rect 22168 99726 22174 99758
rect 21896 99688 21972 99694
rect 22173 99694 22174 99726
rect 22238 99726 22244 99758
rect 22984 99966 22990 99998
rect 23054 99998 23055 100030
rect 23397 100030 23463 100031
rect 23397 99998 23398 100030
rect 23054 99966 23060 99998
rect 22984 99758 23060 99966
rect 22238 99694 22239 99726
rect 22173 99693 22239 99694
rect 22984 99694 22990 99758
rect 23054 99694 23060 99758
rect 22984 99688 23060 99694
rect 23392 99966 23398 99998
rect 23462 99998 23463 100030
rect 28424 100030 28500 100374
rect 110296 100302 110372 100510
rect 116144 100510 116150 100574
rect 116214 100510 116220 100574
rect 116416 100782 116422 100846
rect 116486 100782 116492 100846
rect 116965 100846 117031 100847
rect 116965 100814 116966 100846
rect 116416 100574 116492 100782
rect 116416 100542 116422 100574
rect 116144 100504 116220 100510
rect 116421 100510 116422 100542
rect 116486 100542 116492 100574
rect 116960 100782 116966 100814
rect 117030 100814 117031 100846
rect 117030 100782 117036 100814
rect 116960 100574 117036 100782
rect 116486 100510 116487 100542
rect 116421 100509 116487 100510
rect 116960 100510 116966 100574
rect 117030 100510 117036 100574
rect 116960 100504 117036 100510
rect 115333 100438 115399 100439
rect 115333 100406 115334 100438
rect 110296 100238 110302 100302
rect 110366 100238 110372 100302
rect 110296 100232 110372 100238
rect 115328 100374 115334 100406
rect 115398 100406 115399 100438
rect 115741 100438 115807 100439
rect 115741 100406 115742 100438
rect 115398 100374 115404 100406
rect 115328 100166 115404 100374
rect 115328 100102 115334 100166
rect 115398 100102 115404 100166
rect 115328 100096 115404 100102
rect 115736 100374 115742 100406
rect 115806 100406 115807 100438
rect 116960 100438 117036 100444
rect 115806 100374 115812 100406
rect 115736 100166 115812 100374
rect 115736 100102 115742 100166
rect 115806 100102 115812 100166
rect 116960 100374 116966 100438
rect 117030 100374 117036 100438
rect 116960 100166 117036 100374
rect 116960 100134 116966 100166
rect 115736 100096 115812 100102
rect 116965 100102 116966 100134
rect 117030 100134 117036 100166
rect 117030 100102 117031 100134
rect 116965 100101 117031 100102
rect 23462 99966 23468 99998
rect 23392 99758 23468 99966
rect 28424 99966 28430 100030
rect 28494 99966 28500 100030
rect 28424 99960 28500 99966
rect 115192 100030 115268 100036
rect 115192 99966 115198 100030
rect 115262 99966 115268 100030
rect 23392 99694 23398 99758
rect 23462 99694 23468 99758
rect 28565 99758 28631 99759
rect 28565 99726 28566 99758
rect 23392 99688 23468 99694
rect 28560 99694 28566 99726
rect 28630 99726 28631 99758
rect 115192 99758 115268 99966
rect 115192 99726 115198 99758
rect 28630 99694 28636 99726
rect 952 99558 1230 99622
rect 1294 99558 1300 99622
rect 952 97854 1300 99558
rect 21760 99622 21836 99628
rect 21760 99558 21766 99622
rect 21830 99558 21836 99622
rect 22173 99622 22239 99623
rect 22173 99590 22174 99622
rect 21760 99350 21836 99558
rect 21760 99318 21766 99350
rect 21765 99286 21766 99318
rect 21830 99318 21836 99350
rect 22168 99558 22174 99590
rect 22238 99590 22239 99622
rect 22445 99622 22511 99623
rect 22445 99590 22446 99622
rect 22238 99558 22244 99590
rect 22168 99350 22244 99558
rect 21830 99286 21831 99318
rect 21765 99285 21831 99286
rect 22168 99286 22174 99350
rect 22238 99286 22244 99350
rect 22168 99280 22244 99286
rect 22440 99558 22446 99590
rect 22510 99590 22511 99622
rect 22989 99622 23055 99623
rect 22989 99590 22990 99622
rect 22510 99558 22516 99590
rect 22440 99350 22516 99558
rect 22440 99286 22446 99350
rect 22510 99286 22516 99350
rect 22440 99280 22516 99286
rect 22984 99558 22990 99590
rect 23054 99590 23055 99622
rect 23528 99622 23604 99628
rect 23054 99558 23060 99590
rect 22984 99350 23060 99558
rect 22984 99286 22990 99350
rect 23054 99286 23060 99350
rect 23528 99558 23534 99622
rect 23598 99558 23604 99622
rect 23528 99350 23604 99558
rect 28560 99486 28636 99694
rect 115197 99694 115198 99726
rect 115262 99726 115268 99758
rect 115600 100030 115676 100036
rect 115600 99966 115606 100030
rect 115670 99966 115676 100030
rect 116013 100030 116079 100031
rect 116013 99998 116014 100030
rect 115600 99758 115676 99966
rect 115600 99726 115606 99758
rect 115262 99694 115263 99726
rect 115197 99693 115263 99694
rect 115605 99694 115606 99726
rect 115670 99726 115676 99758
rect 116008 99966 116014 99998
rect 116078 99998 116079 100030
rect 116824 100030 116900 100036
rect 116078 99966 116084 99998
rect 116008 99758 116084 99966
rect 115670 99694 115671 99726
rect 115605 99693 115671 99694
rect 116008 99694 116014 99758
rect 116078 99694 116084 99758
rect 116824 99966 116830 100030
rect 116894 99966 116900 100030
rect 116824 99758 116900 99966
rect 116824 99726 116830 99758
rect 116008 99688 116084 99694
rect 116829 99694 116830 99726
rect 116894 99726 116900 99758
rect 116894 99694 116895 99726
rect 116829 99693 116895 99694
rect 115197 99622 115263 99623
rect 115197 99590 115198 99622
rect 28560 99422 28566 99486
rect 28630 99422 28636 99486
rect 28560 99416 28636 99422
rect 115192 99558 115198 99590
rect 115262 99590 115263 99622
rect 115741 99622 115807 99623
rect 115741 99590 115742 99622
rect 115262 99558 115268 99590
rect 23528 99318 23534 99350
rect 22984 99280 23060 99286
rect 23533 99286 23534 99318
rect 23598 99318 23604 99350
rect 115192 99350 115268 99558
rect 23598 99286 23599 99318
rect 23533 99285 23599 99286
rect 115192 99286 115198 99350
rect 115262 99286 115268 99350
rect 115192 99280 115268 99286
rect 115736 99558 115742 99590
rect 115806 99590 115807 99622
rect 116285 99622 116351 99623
rect 116285 99590 116286 99622
rect 115806 99558 115812 99590
rect 115736 99350 115812 99558
rect 115736 99286 115742 99350
rect 115806 99286 115812 99350
rect 115736 99280 115812 99286
rect 116280 99558 116286 99590
rect 116350 99590 116351 99622
rect 116421 99622 116487 99623
rect 116421 99590 116422 99622
rect 116350 99558 116356 99590
rect 116280 99350 116356 99558
rect 116280 99286 116286 99350
rect 116350 99286 116356 99350
rect 116280 99280 116356 99286
rect 116416 99558 116422 99590
rect 116486 99590 116487 99622
rect 116829 99622 116895 99623
rect 116829 99590 116830 99622
rect 116486 99558 116492 99590
rect 116416 99350 116492 99558
rect 116416 99286 116422 99350
rect 116486 99286 116492 99350
rect 116416 99280 116492 99286
rect 116824 99558 116830 99590
rect 116894 99590 116895 99622
rect 137496 99622 137844 101190
rect 116894 99558 116900 99590
rect 116824 99350 116900 99558
rect 116824 99286 116830 99350
rect 116894 99286 116900 99350
rect 116824 99280 116900 99286
rect 137496 99558 137502 99622
rect 137566 99558 137844 99622
rect 21896 99214 21972 99220
rect 21896 99150 21902 99214
rect 21966 99150 21972 99214
rect 22581 99214 22647 99215
rect 22581 99182 22582 99214
rect 21896 98942 21972 99150
rect 21896 98910 21902 98942
rect 21901 98878 21902 98910
rect 21966 98910 21972 98942
rect 22576 99150 22582 99182
rect 22646 99182 22647 99214
rect 22984 99214 23060 99220
rect 22646 99150 22652 99182
rect 22576 98942 22652 99150
rect 21966 98878 21967 98910
rect 21901 98877 21967 98878
rect 22576 98878 22582 98942
rect 22646 98878 22652 98942
rect 22984 99150 22990 99214
rect 23054 99150 23060 99214
rect 22984 98942 23060 99150
rect 22984 98910 22990 98942
rect 22576 98872 22652 98878
rect 22989 98878 22990 98910
rect 23054 98910 23060 98942
rect 23392 99214 23468 99220
rect 23392 99150 23398 99214
rect 23462 99150 23468 99214
rect 23392 98942 23468 99150
rect 23392 98910 23398 98942
rect 23054 98878 23055 98910
rect 22989 98877 23055 98878
rect 23397 98878 23398 98910
rect 23462 98910 23468 98942
rect 115192 99214 115268 99220
rect 115192 99150 115198 99214
rect 115262 99150 115268 99214
rect 115192 98942 115268 99150
rect 115192 98910 115198 98942
rect 23462 98878 23463 98910
rect 23397 98877 23463 98878
rect 115197 98878 115198 98910
rect 115262 98910 115268 98942
rect 115600 99214 115676 99220
rect 115600 99150 115606 99214
rect 115670 99150 115676 99214
rect 116149 99214 116215 99215
rect 116149 99182 116150 99214
rect 115600 98942 115676 99150
rect 115600 98910 115606 98942
rect 115262 98878 115263 98910
rect 115197 98877 115263 98878
rect 115605 98878 115606 98910
rect 115670 98910 115676 98942
rect 116144 99150 116150 99182
rect 116214 99182 116215 99214
rect 116552 99214 116628 99220
rect 116214 99150 116220 99182
rect 116144 98942 116220 99150
rect 115670 98878 115671 98910
rect 115605 98877 115671 98878
rect 116144 98878 116150 98942
rect 116214 98878 116220 98942
rect 116552 99150 116558 99214
rect 116622 99150 116628 99214
rect 116552 98942 116628 99150
rect 116552 98910 116558 98942
rect 116144 98872 116220 98878
rect 116557 98878 116558 98910
rect 116622 98910 116628 98942
rect 116960 99214 117036 99220
rect 116960 99150 116966 99214
rect 117030 99150 117036 99214
rect 116960 98942 117036 99150
rect 116960 98910 116966 98942
rect 116622 98878 116623 98910
rect 116557 98877 116623 98878
rect 116965 98878 116966 98910
rect 117030 98910 117036 98942
rect 117030 98878 117031 98910
rect 116965 98877 117031 98878
rect 21901 98806 21967 98807
rect 21901 98774 21902 98806
rect 21896 98742 21902 98774
rect 21966 98774 21967 98806
rect 22168 98806 22244 98812
rect 21966 98742 21972 98774
rect 21896 98534 21972 98742
rect 21896 98470 21902 98534
rect 21966 98470 21972 98534
rect 22168 98742 22174 98806
rect 22238 98742 22244 98806
rect 23125 98806 23191 98807
rect 23125 98774 23126 98806
rect 22168 98534 22244 98742
rect 22168 98502 22174 98534
rect 21896 98464 21972 98470
rect 22173 98470 22174 98502
rect 22238 98502 22244 98534
rect 23120 98742 23126 98774
rect 23190 98774 23191 98806
rect 23397 98806 23463 98807
rect 23397 98774 23398 98806
rect 23190 98742 23196 98774
rect 23120 98534 23196 98742
rect 22238 98470 22239 98502
rect 22173 98469 22239 98470
rect 23120 98470 23126 98534
rect 23190 98470 23196 98534
rect 23120 98464 23196 98470
rect 23392 98742 23398 98774
rect 23462 98774 23463 98806
rect 115197 98806 115263 98807
rect 115197 98774 115198 98806
rect 23462 98742 23468 98774
rect 23392 98534 23468 98742
rect 23392 98470 23398 98534
rect 23462 98470 23468 98534
rect 23392 98464 23468 98470
rect 115192 98742 115198 98774
rect 115262 98774 115263 98806
rect 115605 98806 115671 98807
rect 115605 98774 115606 98806
rect 115262 98742 115268 98774
rect 115192 98534 115268 98742
rect 115192 98470 115198 98534
rect 115262 98470 115268 98534
rect 115192 98464 115268 98470
rect 115600 98742 115606 98774
rect 115670 98774 115671 98806
rect 116008 98806 116084 98812
rect 115670 98742 115676 98774
rect 115600 98534 115676 98742
rect 115600 98470 115606 98534
rect 115670 98470 115676 98534
rect 116008 98742 116014 98806
rect 116078 98742 116084 98806
rect 116965 98806 117031 98807
rect 116965 98774 116966 98806
rect 116008 98534 116084 98742
rect 116008 98502 116014 98534
rect 115600 98464 115676 98470
rect 116013 98470 116014 98502
rect 116078 98502 116084 98534
rect 116960 98742 116966 98774
rect 117030 98774 117031 98806
rect 117030 98742 117036 98774
rect 116960 98534 117036 98742
rect 116078 98470 116079 98502
rect 116013 98469 116079 98470
rect 116960 98470 116966 98534
rect 117030 98470 117036 98534
rect 116960 98464 117036 98470
rect 22173 98398 22239 98399
rect 22173 98366 22174 98398
rect 22168 98334 22174 98366
rect 22238 98366 22239 98398
rect 22581 98398 22647 98399
rect 22581 98366 22582 98398
rect 22238 98334 22244 98366
rect 22168 98126 22244 98334
rect 22168 98062 22174 98126
rect 22238 98062 22244 98126
rect 22168 98056 22244 98062
rect 22576 98334 22582 98366
rect 22646 98366 22647 98398
rect 22989 98398 23055 98399
rect 22989 98366 22990 98398
rect 22646 98334 22652 98366
rect 22576 98126 22652 98334
rect 22576 98062 22582 98126
rect 22646 98062 22652 98126
rect 22576 98056 22652 98062
rect 22984 98334 22990 98366
rect 23054 98366 23055 98398
rect 23533 98398 23599 98399
rect 23533 98366 23534 98398
rect 23054 98334 23060 98366
rect 22984 98126 23060 98334
rect 22984 98062 22990 98126
rect 23054 98062 23060 98126
rect 22984 98056 23060 98062
rect 23528 98334 23534 98366
rect 23598 98366 23599 98398
rect 115328 98398 115404 98404
rect 23598 98334 23604 98366
rect 23528 98126 23604 98334
rect 23528 98062 23534 98126
rect 23598 98062 23604 98126
rect 115328 98334 115334 98398
rect 115398 98334 115404 98398
rect 115328 98126 115404 98334
rect 115328 98094 115334 98126
rect 23528 98056 23604 98062
rect 115333 98062 115334 98094
rect 115398 98094 115404 98126
rect 115736 98398 115812 98404
rect 115736 98334 115742 98398
rect 115806 98334 115812 98398
rect 116013 98398 116079 98399
rect 116013 98366 116014 98398
rect 115736 98126 115812 98334
rect 115736 98094 115742 98126
rect 115398 98062 115399 98094
rect 115333 98061 115399 98062
rect 115741 98062 115742 98094
rect 115806 98094 115812 98126
rect 116008 98334 116014 98366
rect 116078 98366 116079 98398
rect 116421 98398 116487 98399
rect 116421 98366 116422 98398
rect 116078 98334 116084 98366
rect 116008 98126 116084 98334
rect 115806 98062 115807 98094
rect 115741 98061 115807 98062
rect 116008 98062 116014 98126
rect 116078 98062 116084 98126
rect 116008 98056 116084 98062
rect 116416 98334 116422 98366
rect 116486 98366 116487 98398
rect 116486 98334 116492 98366
rect 116416 98126 116492 98334
rect 116416 98062 116422 98126
rect 116486 98062 116492 98126
rect 116416 98056 116492 98062
rect 952 97790 1230 97854
rect 1294 97790 1300 97854
rect 952 96222 1300 97790
rect 23120 97990 23196 97996
rect 23120 97926 23126 97990
rect 23190 97926 23196 97990
rect 23120 97718 23196 97926
rect 23120 97686 23126 97718
rect 23125 97654 23126 97686
rect 23190 97686 23196 97718
rect 23392 97990 23468 97996
rect 23392 97926 23398 97990
rect 23462 97926 23468 97990
rect 28293 97990 28359 97991
rect 28293 97958 28294 97990
rect 23392 97718 23468 97926
rect 23392 97686 23398 97718
rect 23190 97654 23191 97686
rect 23125 97653 23191 97654
rect 23397 97654 23398 97686
rect 23462 97686 23468 97718
rect 28288 97926 28294 97958
rect 28358 97958 28359 97990
rect 115197 97990 115263 97991
rect 115197 97958 115198 97990
rect 28358 97926 28364 97958
rect 23462 97654 23463 97686
rect 23397 97653 23463 97654
rect 22576 97582 22652 97588
rect 22576 97518 22582 97582
rect 22646 97518 22652 97582
rect 23125 97582 23191 97583
rect 23125 97550 23126 97582
rect 21760 97310 21836 97316
rect 21760 97246 21766 97310
rect 21830 97246 21836 97310
rect 22576 97310 22652 97518
rect 22576 97278 22582 97310
rect 21760 97038 21836 97246
rect 22581 97246 22582 97278
rect 22646 97278 22652 97310
rect 23120 97518 23126 97550
rect 23190 97550 23191 97582
rect 23397 97582 23463 97583
rect 23397 97550 23398 97582
rect 23190 97518 23196 97550
rect 23120 97310 23196 97518
rect 22646 97246 22647 97278
rect 22581 97245 22647 97246
rect 23120 97246 23126 97310
rect 23190 97246 23196 97310
rect 23120 97240 23196 97246
rect 23392 97518 23398 97550
rect 23462 97550 23463 97582
rect 28288 97582 28364 97926
rect 115192 97926 115198 97958
rect 115262 97958 115263 97990
rect 115605 97990 115671 97991
rect 115605 97958 115606 97990
rect 115262 97926 115268 97958
rect 115192 97718 115268 97926
rect 115192 97654 115198 97718
rect 115262 97654 115268 97718
rect 115192 97648 115268 97654
rect 115600 97926 115606 97958
rect 115670 97958 115671 97990
rect 115670 97926 115676 97958
rect 115600 97718 115676 97926
rect 115600 97654 115606 97718
rect 115670 97654 115676 97718
rect 115600 97648 115676 97654
rect 137496 97854 137844 99558
rect 137496 97790 137502 97854
rect 137566 97790 137844 97854
rect 23462 97518 23468 97550
rect 23392 97310 23468 97518
rect 28288 97518 28294 97582
rect 28358 97518 28364 97582
rect 28288 97512 28364 97518
rect 115328 97582 115404 97588
rect 115328 97518 115334 97582
rect 115398 97518 115404 97582
rect 23392 97246 23398 97310
rect 23462 97246 23468 97310
rect 23392 97240 23468 97246
rect 110160 97446 110236 97452
rect 110160 97382 110166 97446
rect 110230 97382 110236 97446
rect 110160 97174 110236 97382
rect 115328 97310 115404 97518
rect 115328 97278 115334 97310
rect 115333 97246 115334 97278
rect 115398 97278 115404 97310
rect 115736 97582 115812 97588
rect 115736 97518 115742 97582
rect 115806 97518 115812 97582
rect 116285 97582 116351 97583
rect 116285 97550 116286 97582
rect 115736 97310 115812 97518
rect 115736 97278 115742 97310
rect 115398 97246 115399 97278
rect 115333 97245 115399 97246
rect 115741 97246 115742 97278
rect 115806 97278 115812 97310
rect 116280 97518 116286 97550
rect 116350 97550 116351 97582
rect 116350 97518 116356 97550
rect 116280 97310 116356 97518
rect 115806 97246 115807 97278
rect 115741 97245 115807 97246
rect 116280 97246 116286 97310
rect 116350 97246 116356 97310
rect 116280 97240 116356 97246
rect 116824 97310 116900 97316
rect 116824 97246 116830 97310
rect 116894 97246 116900 97310
rect 110160 97142 110166 97174
rect 110165 97110 110166 97142
rect 110230 97142 110236 97174
rect 110230 97110 110231 97142
rect 110165 97109 110231 97110
rect 21760 97006 21766 97038
rect 21765 96974 21766 97006
rect 21830 97006 21836 97038
rect 28424 97038 28500 97044
rect 21830 96974 21831 97006
rect 21765 96973 21831 96974
rect 28424 96974 28430 97038
rect 28494 96974 28500 97038
rect 110301 97038 110367 97039
rect 110301 97006 110302 97038
rect 21901 96902 21967 96903
rect 21901 96870 21902 96902
rect 21896 96838 21902 96870
rect 21966 96870 21967 96902
rect 22717 96902 22783 96903
rect 22717 96870 22718 96902
rect 21966 96838 21972 96870
rect 21896 96630 21972 96838
rect 21896 96566 21902 96630
rect 21966 96566 21972 96630
rect 21896 96560 21972 96566
rect 22712 96838 22718 96870
rect 22782 96870 22783 96902
rect 22782 96838 22788 96870
rect 22712 96630 22788 96838
rect 28424 96766 28500 96974
rect 28424 96734 28430 96766
rect 28429 96702 28430 96734
rect 28494 96734 28500 96766
rect 110296 96974 110302 97006
rect 110366 97006 110367 97038
rect 116824 97038 116900 97246
rect 116824 97006 116830 97038
rect 110366 96974 110372 97006
rect 110296 96766 110372 96974
rect 116829 96974 116830 97006
rect 116894 97006 116900 97038
rect 116894 96974 116895 97006
rect 116829 96973 116895 96974
rect 28494 96702 28495 96734
rect 28429 96701 28495 96702
rect 110296 96702 110302 96766
rect 110366 96702 110372 96766
rect 110296 96696 110372 96702
rect 116552 96902 116628 96908
rect 116552 96838 116558 96902
rect 116622 96838 116628 96902
rect 22712 96566 22718 96630
rect 22782 96566 22788 96630
rect 116552 96630 116628 96838
rect 116552 96598 116558 96630
rect 22712 96560 22788 96566
rect 116557 96566 116558 96598
rect 116622 96598 116628 96630
rect 116960 96902 117036 96908
rect 116960 96838 116966 96902
rect 117030 96838 117036 96902
rect 116960 96630 117036 96838
rect 116960 96598 116966 96630
rect 116622 96566 116623 96598
rect 116557 96565 116623 96566
rect 116965 96566 116966 96598
rect 117030 96598 117036 96630
rect 117030 96566 117031 96598
rect 116965 96565 117031 96566
rect 952 96158 1230 96222
rect 1294 96158 1300 96222
rect 21760 96494 21836 96500
rect 21760 96430 21766 96494
rect 21830 96430 21836 96494
rect 21760 96222 21836 96430
rect 21760 96190 21766 96222
rect 952 94590 1300 96158
rect 21765 96158 21766 96190
rect 21830 96190 21836 96222
rect 22984 96494 23060 96500
rect 22984 96430 22990 96494
rect 23054 96430 23060 96494
rect 22984 96222 23060 96430
rect 22984 96190 22990 96222
rect 21830 96158 21831 96190
rect 21765 96157 21831 96158
rect 22989 96158 22990 96190
rect 23054 96190 23060 96222
rect 23528 96494 23604 96500
rect 23528 96430 23534 96494
rect 23598 96430 23604 96494
rect 23528 96222 23604 96430
rect 23528 96190 23534 96222
rect 23054 96158 23055 96190
rect 22989 96157 23055 96158
rect 23533 96158 23534 96190
rect 23598 96190 23604 96222
rect 115328 96494 115404 96500
rect 115328 96430 115334 96494
rect 115398 96430 115404 96494
rect 115328 96222 115404 96430
rect 115328 96190 115334 96222
rect 23598 96158 23599 96190
rect 23533 96157 23599 96158
rect 115333 96158 115334 96190
rect 115398 96190 115404 96222
rect 115736 96494 115812 96500
rect 115736 96430 115742 96494
rect 115806 96430 115812 96494
rect 116285 96494 116351 96495
rect 116285 96462 116286 96494
rect 115736 96222 115812 96430
rect 115736 96190 115742 96222
rect 115398 96158 115399 96190
rect 115333 96157 115399 96158
rect 115741 96158 115742 96190
rect 115806 96190 115812 96222
rect 116280 96430 116286 96462
rect 116350 96462 116351 96494
rect 116965 96494 117031 96495
rect 116965 96462 116966 96494
rect 116350 96430 116356 96462
rect 116280 96222 116356 96430
rect 115806 96158 115807 96190
rect 115741 96157 115807 96158
rect 116280 96158 116286 96222
rect 116350 96158 116356 96222
rect 116280 96152 116356 96158
rect 116960 96430 116966 96462
rect 117030 96462 117031 96494
rect 117030 96430 117036 96462
rect 116960 96222 117036 96430
rect 116960 96158 116966 96222
rect 117030 96158 117036 96222
rect 116960 96152 117036 96158
rect 21896 96086 21972 96092
rect 21896 96022 21902 96086
rect 21966 96022 21972 96086
rect 22173 96086 22239 96087
rect 22173 96054 22174 96086
rect 21896 95814 21972 96022
rect 21896 95782 21902 95814
rect 21901 95750 21902 95782
rect 21966 95782 21972 95814
rect 22168 96022 22174 96054
rect 22238 96054 22239 96086
rect 22712 96086 22788 96092
rect 22238 96022 22244 96054
rect 22168 95814 22244 96022
rect 21966 95750 21967 95782
rect 21901 95749 21967 95750
rect 22168 95750 22174 95814
rect 22238 95750 22244 95814
rect 22712 96022 22718 96086
rect 22782 96022 22788 96086
rect 22989 96086 23055 96087
rect 22989 96054 22990 96086
rect 22712 95814 22788 96022
rect 22712 95782 22718 95814
rect 22168 95744 22244 95750
rect 22717 95750 22718 95782
rect 22782 95782 22788 95814
rect 22984 96022 22990 96054
rect 23054 96054 23055 96086
rect 23392 96086 23468 96092
rect 23054 96022 23060 96054
rect 22984 95814 23060 96022
rect 22782 95750 22783 95782
rect 22717 95749 22783 95750
rect 22984 95750 22990 95814
rect 23054 95750 23060 95814
rect 23392 96022 23398 96086
rect 23462 96022 23468 96086
rect 115333 96086 115399 96087
rect 115333 96054 115334 96086
rect 23392 95814 23468 96022
rect 115328 96022 115334 96054
rect 115398 96054 115399 96086
rect 115741 96086 115807 96087
rect 115741 96054 115742 96086
rect 115398 96022 115404 96054
rect 23392 95782 23398 95814
rect 22984 95744 23060 95750
rect 23397 95750 23398 95782
rect 23462 95782 23468 95814
rect 28429 95814 28495 95815
rect 28429 95782 28430 95814
rect 23462 95750 23463 95782
rect 23397 95749 23463 95750
rect 28424 95750 28430 95782
rect 28494 95782 28495 95814
rect 110165 95814 110231 95815
rect 110165 95782 110166 95814
rect 28494 95750 28500 95782
rect 21896 95678 21972 95684
rect 21896 95614 21902 95678
rect 21966 95614 21972 95678
rect 22989 95678 23055 95679
rect 22989 95646 22990 95678
rect 21896 95406 21972 95614
rect 21896 95374 21902 95406
rect 21901 95342 21902 95374
rect 21966 95374 21972 95406
rect 22984 95614 22990 95646
rect 23054 95646 23055 95678
rect 23397 95678 23463 95679
rect 23397 95646 23398 95678
rect 23054 95614 23060 95646
rect 22984 95406 23060 95614
rect 21966 95342 21967 95374
rect 21901 95341 21967 95342
rect 22984 95342 22990 95406
rect 23054 95342 23060 95406
rect 22984 95336 23060 95342
rect 23392 95614 23398 95646
rect 23462 95646 23463 95678
rect 23462 95614 23468 95646
rect 23392 95406 23468 95614
rect 28424 95542 28500 95750
rect 28424 95478 28430 95542
rect 28494 95478 28500 95542
rect 28424 95472 28500 95478
rect 110160 95750 110166 95782
rect 110230 95782 110231 95814
rect 115328 95814 115404 96022
rect 110230 95750 110236 95782
rect 110160 95542 110236 95750
rect 115328 95750 115334 95814
rect 115398 95750 115404 95814
rect 115328 95744 115404 95750
rect 115736 96022 115742 96054
rect 115806 96054 115807 96086
rect 116552 96086 116628 96092
rect 115806 96022 115812 96054
rect 115736 95814 115812 96022
rect 115736 95750 115742 95814
rect 115806 95750 115812 95814
rect 116552 96022 116558 96086
rect 116622 96022 116628 96086
rect 116552 95814 116628 96022
rect 116552 95782 116558 95814
rect 115736 95744 115812 95750
rect 116557 95750 116558 95782
rect 116622 95782 116628 95814
rect 116960 96086 117036 96092
rect 116960 96022 116966 96086
rect 117030 96022 117036 96086
rect 116960 95814 117036 96022
rect 116960 95782 116966 95814
rect 116622 95750 116623 95782
rect 116557 95749 116623 95750
rect 116965 95750 116966 95782
rect 117030 95782 117036 95814
rect 137496 96086 137844 97790
rect 137496 96022 137502 96086
rect 137566 96022 137844 96086
rect 117030 95750 117031 95782
rect 116965 95749 117031 95750
rect 115197 95678 115263 95679
rect 115197 95646 115198 95678
rect 110160 95478 110166 95542
rect 110230 95478 110236 95542
rect 110160 95472 110236 95478
rect 115192 95614 115198 95646
rect 115262 95646 115263 95678
rect 115600 95678 115676 95684
rect 115262 95614 115268 95646
rect 23392 95342 23398 95406
rect 23462 95342 23468 95406
rect 23392 95336 23468 95342
rect 115192 95406 115268 95614
rect 115192 95342 115198 95406
rect 115262 95342 115268 95406
rect 115600 95614 115606 95678
rect 115670 95614 115676 95678
rect 115600 95406 115676 95614
rect 115600 95374 115606 95406
rect 115192 95336 115268 95342
rect 115605 95342 115606 95374
rect 115670 95374 115676 95406
rect 116144 95678 116220 95684
rect 116144 95614 116150 95678
rect 116214 95614 116220 95678
rect 116965 95678 117031 95679
rect 116965 95646 116966 95678
rect 116144 95406 116220 95614
rect 116144 95374 116150 95406
rect 115670 95342 115671 95374
rect 115605 95341 115671 95342
rect 116149 95342 116150 95374
rect 116214 95374 116220 95406
rect 116960 95614 116966 95646
rect 117030 95646 117031 95678
rect 117030 95614 117036 95646
rect 116960 95406 117036 95614
rect 116214 95342 116215 95374
rect 116149 95341 116215 95342
rect 116960 95342 116966 95406
rect 117030 95342 117036 95406
rect 116960 95336 117036 95342
rect 21765 95270 21831 95271
rect 21765 95238 21766 95270
rect 21760 95206 21766 95238
rect 21830 95238 21831 95270
rect 22168 95270 22244 95276
rect 21830 95206 21836 95238
rect 21760 94998 21836 95206
rect 21760 94934 21766 94998
rect 21830 94934 21836 94998
rect 22168 95206 22174 95270
rect 22238 95206 22244 95270
rect 22581 95270 22647 95271
rect 22581 95238 22582 95270
rect 22168 94998 22244 95206
rect 22168 94966 22174 94998
rect 21760 94928 21836 94934
rect 22173 94934 22174 94966
rect 22238 94966 22244 94998
rect 22576 95206 22582 95238
rect 22646 95238 22647 95270
rect 23120 95270 23196 95276
rect 22646 95206 22652 95238
rect 22576 94998 22652 95206
rect 22238 94934 22239 94966
rect 22173 94933 22239 94934
rect 22576 94934 22582 94998
rect 22646 94934 22652 94998
rect 23120 95206 23126 95270
rect 23190 95206 23196 95270
rect 23120 94998 23196 95206
rect 23120 94966 23126 94998
rect 22576 94928 22652 94934
rect 23125 94934 23126 94966
rect 23190 94966 23196 94998
rect 23528 95270 23604 95276
rect 23528 95206 23534 95270
rect 23598 95206 23604 95270
rect 23528 94998 23604 95206
rect 23528 94966 23534 94998
rect 23190 94934 23191 94966
rect 23125 94933 23191 94934
rect 23533 94934 23534 94966
rect 23598 94966 23604 94998
rect 115328 95270 115404 95276
rect 115328 95206 115334 95270
rect 115398 95206 115404 95270
rect 115741 95270 115807 95271
rect 115741 95238 115742 95270
rect 115328 94998 115404 95206
rect 115328 94966 115334 94998
rect 23598 94934 23599 94966
rect 23533 94933 23599 94934
rect 115333 94934 115334 94966
rect 115398 94966 115404 94998
rect 115736 95206 115742 95238
rect 115806 95238 115807 95270
rect 116013 95270 116079 95271
rect 116013 95238 116014 95270
rect 115806 95206 115812 95238
rect 115736 94998 115812 95206
rect 115398 94934 115399 94966
rect 115333 94933 115399 94934
rect 115736 94934 115742 94998
rect 115806 94934 115812 94998
rect 115736 94928 115812 94934
rect 116008 95206 116014 95238
rect 116078 95238 116079 95270
rect 116421 95270 116487 95271
rect 116421 95238 116422 95270
rect 116078 95206 116084 95238
rect 116008 94998 116084 95206
rect 116008 94934 116014 94998
rect 116078 94934 116084 94998
rect 116008 94928 116084 94934
rect 116416 95206 116422 95238
rect 116486 95238 116487 95270
rect 116824 95270 116900 95276
rect 116486 95206 116492 95238
rect 116416 94998 116492 95206
rect 116416 94934 116422 94998
rect 116486 94934 116492 94998
rect 116824 95206 116830 95270
rect 116894 95206 116900 95270
rect 116824 94998 116900 95206
rect 116824 94966 116830 94998
rect 116416 94928 116492 94934
rect 116829 94934 116830 94966
rect 116894 94966 116900 94998
rect 116894 94934 116895 94966
rect 116829 94933 116895 94934
rect 952 94526 1230 94590
rect 1294 94526 1300 94590
rect 21896 94862 21972 94868
rect 21896 94798 21902 94862
rect 21966 94798 21972 94862
rect 21896 94590 21972 94798
rect 21896 94558 21902 94590
rect 952 92958 1300 94526
rect 21901 94526 21902 94558
rect 21966 94558 21972 94590
rect 22304 94862 22380 94868
rect 22304 94798 22310 94862
rect 22374 94798 22380 94862
rect 22304 94590 22380 94798
rect 22304 94558 22310 94590
rect 21966 94526 21967 94558
rect 21901 94525 21967 94526
rect 22309 94526 22310 94558
rect 22374 94558 22380 94590
rect 23120 94862 23196 94868
rect 23120 94798 23126 94862
rect 23190 94798 23196 94862
rect 23533 94862 23599 94863
rect 23533 94830 23534 94862
rect 23120 94590 23196 94798
rect 23120 94558 23126 94590
rect 22374 94526 22375 94558
rect 22309 94525 22375 94526
rect 23125 94526 23126 94558
rect 23190 94558 23196 94590
rect 23528 94798 23534 94830
rect 23598 94830 23599 94862
rect 115192 94862 115268 94868
rect 23598 94798 23604 94830
rect 23528 94590 23604 94798
rect 23190 94526 23191 94558
rect 23125 94525 23191 94526
rect 23528 94526 23534 94590
rect 23598 94526 23604 94590
rect 115192 94798 115198 94862
rect 115262 94798 115268 94862
rect 115192 94590 115268 94798
rect 115192 94558 115198 94590
rect 23528 94520 23604 94526
rect 115197 94526 115198 94558
rect 115262 94558 115268 94590
rect 115600 94862 115676 94868
rect 115600 94798 115606 94862
rect 115670 94798 115676 94862
rect 116829 94862 116895 94863
rect 116829 94830 116830 94862
rect 115600 94590 115676 94798
rect 115600 94558 115606 94590
rect 115262 94526 115263 94558
rect 115197 94525 115263 94526
rect 115605 94526 115606 94558
rect 115670 94558 115676 94590
rect 116824 94798 116830 94830
rect 116894 94830 116895 94862
rect 116894 94798 116900 94830
rect 116824 94590 116900 94798
rect 115670 94526 115671 94558
rect 115605 94525 115671 94526
rect 116824 94526 116830 94590
rect 116894 94526 116900 94590
rect 116824 94520 116900 94526
rect 22576 94454 22652 94460
rect 22576 94390 22582 94454
rect 22646 94390 22652 94454
rect 23125 94454 23191 94455
rect 23125 94422 23126 94454
rect 22576 94182 22652 94390
rect 22576 94150 22582 94182
rect 22581 94118 22582 94150
rect 22646 94150 22652 94182
rect 23120 94390 23126 94422
rect 23190 94422 23191 94454
rect 23397 94454 23463 94455
rect 23397 94422 23398 94454
rect 23190 94390 23196 94422
rect 23120 94182 23196 94390
rect 22646 94118 22647 94150
rect 22581 94117 22647 94118
rect 23120 94118 23126 94182
rect 23190 94118 23196 94182
rect 23120 94112 23196 94118
rect 23392 94390 23398 94422
rect 23462 94422 23463 94454
rect 115328 94454 115404 94460
rect 23462 94390 23468 94422
rect 23392 94182 23468 94390
rect 115328 94390 115334 94454
rect 115398 94390 115404 94454
rect 115605 94454 115671 94455
rect 115605 94422 115606 94454
rect 110165 94318 110231 94319
rect 110165 94286 110166 94318
rect 23392 94118 23398 94182
rect 23462 94118 23468 94182
rect 23392 94112 23468 94118
rect 110160 94254 110166 94286
rect 110230 94286 110231 94318
rect 110230 94254 110236 94286
rect 23120 94046 23196 94052
rect 23120 93982 23126 94046
rect 23190 93982 23196 94046
rect 23120 93774 23196 93982
rect 23120 93742 23126 93774
rect 23125 93710 23126 93742
rect 23190 93742 23196 93774
rect 23528 94046 23604 94052
rect 23528 93982 23534 94046
rect 23598 93982 23604 94046
rect 23528 93774 23604 93982
rect 110160 94046 110236 94254
rect 115328 94182 115404 94390
rect 115328 94150 115334 94182
rect 115333 94118 115334 94150
rect 115398 94150 115404 94182
rect 115600 94390 115606 94422
rect 115670 94422 115671 94454
rect 116013 94454 116079 94455
rect 116013 94422 116014 94454
rect 115670 94390 115676 94422
rect 115600 94182 115676 94390
rect 115398 94118 115399 94150
rect 115333 94117 115399 94118
rect 115600 94118 115606 94182
rect 115670 94118 115676 94182
rect 115600 94112 115676 94118
rect 116008 94390 116014 94422
rect 116078 94422 116079 94454
rect 116285 94454 116351 94455
rect 116285 94422 116286 94454
rect 116078 94390 116084 94422
rect 116008 94182 116084 94390
rect 116008 94118 116014 94182
rect 116078 94118 116084 94182
rect 116008 94112 116084 94118
rect 116280 94390 116286 94422
rect 116350 94422 116351 94454
rect 137496 94454 137844 96022
rect 116350 94390 116356 94422
rect 116280 94182 116356 94390
rect 116280 94118 116286 94182
rect 116350 94118 116356 94182
rect 116280 94112 116356 94118
rect 137496 94390 137502 94454
rect 137566 94390 137844 94454
rect 110160 93982 110166 94046
rect 110230 93982 110236 94046
rect 115333 94046 115399 94047
rect 115333 94014 115334 94046
rect 110160 93976 110236 93982
rect 115328 93982 115334 94014
rect 115398 94014 115399 94046
rect 115736 94046 115812 94052
rect 115398 93982 115404 94014
rect 23528 93742 23534 93774
rect 23190 93710 23191 93742
rect 23125 93709 23191 93710
rect 23533 93710 23534 93742
rect 23598 93742 23604 93774
rect 115328 93774 115404 93982
rect 23598 93710 23599 93742
rect 23533 93709 23599 93710
rect 115328 93710 115334 93774
rect 115398 93710 115404 93774
rect 115736 93982 115742 94046
rect 115806 93982 115812 94046
rect 115736 93774 115812 93982
rect 115736 93742 115742 93774
rect 115328 93704 115404 93710
rect 115741 93710 115742 93742
rect 115806 93742 115812 93774
rect 115806 93710 115807 93742
rect 115741 93709 115807 93710
rect 22440 93638 22516 93644
rect 22440 93574 22446 93638
rect 22510 93574 22516 93638
rect 22989 93638 23055 93639
rect 22989 93606 22990 93638
rect 21901 93366 21967 93367
rect 21901 93334 21902 93366
rect 21896 93302 21902 93334
rect 21966 93334 21967 93366
rect 22440 93366 22516 93574
rect 22440 93334 22446 93366
rect 21966 93302 21972 93334
rect 21896 93094 21972 93302
rect 22445 93302 22446 93334
rect 22510 93334 22516 93366
rect 22984 93574 22990 93606
rect 23054 93606 23055 93638
rect 23397 93638 23463 93639
rect 23397 93606 23398 93638
rect 23054 93574 23060 93606
rect 22984 93366 23060 93574
rect 22510 93302 22511 93334
rect 22445 93301 22511 93302
rect 22984 93302 22990 93366
rect 23054 93302 23060 93366
rect 22984 93296 23060 93302
rect 23392 93574 23398 93606
rect 23462 93606 23463 93638
rect 115197 93638 115263 93639
rect 115197 93606 115198 93638
rect 23462 93574 23468 93606
rect 23392 93366 23468 93574
rect 115192 93574 115198 93606
rect 115262 93606 115263 93638
rect 115600 93638 115676 93644
rect 115262 93574 115268 93606
rect 28565 93502 28631 93503
rect 28565 93470 28566 93502
rect 23392 93302 23398 93366
rect 23462 93302 23468 93366
rect 23392 93296 23468 93302
rect 28560 93438 28566 93470
rect 28630 93470 28631 93502
rect 28630 93438 28636 93470
rect 28560 93230 28636 93438
rect 115192 93366 115268 93574
rect 115192 93302 115198 93366
rect 115262 93302 115268 93366
rect 115600 93574 115606 93638
rect 115670 93574 115676 93638
rect 116421 93638 116487 93639
rect 116421 93606 116422 93638
rect 115600 93366 115676 93574
rect 115600 93334 115606 93366
rect 115192 93296 115268 93302
rect 115605 93302 115606 93334
rect 115670 93334 115676 93366
rect 116416 93574 116422 93606
rect 116486 93606 116487 93638
rect 116486 93574 116492 93606
rect 116416 93366 116492 93574
rect 115670 93302 115671 93334
rect 115605 93301 115671 93302
rect 116416 93302 116422 93366
rect 116486 93302 116492 93366
rect 116416 93296 116492 93302
rect 116824 93366 116900 93372
rect 116824 93302 116830 93366
rect 116894 93302 116900 93366
rect 28560 93166 28566 93230
rect 28630 93166 28636 93230
rect 28560 93160 28636 93166
rect 21896 93030 21902 93094
rect 21966 93030 21972 93094
rect 21896 93024 21972 93030
rect 28288 93094 28364 93100
rect 28288 93030 28294 93094
rect 28358 93030 28364 93094
rect 110301 93094 110367 93095
rect 110301 93062 110302 93094
rect 952 92894 1230 92958
rect 1294 92894 1300 92958
rect 952 91190 1300 92894
rect 21760 92958 21836 92964
rect 21760 92894 21766 92958
rect 21830 92894 21836 92958
rect 22581 92958 22647 92959
rect 22581 92926 22582 92958
rect 21760 92686 21836 92894
rect 21760 92654 21766 92686
rect 21765 92622 21766 92654
rect 21830 92654 21836 92686
rect 22576 92894 22582 92926
rect 22646 92926 22647 92958
rect 22646 92894 22652 92926
rect 22576 92686 22652 92894
rect 28288 92822 28364 93030
rect 28288 92790 28294 92822
rect 28293 92758 28294 92790
rect 28358 92790 28364 92822
rect 110296 93030 110302 93062
rect 110366 93062 110367 93094
rect 116824 93094 116900 93302
rect 116824 93062 116830 93094
rect 110366 93030 110372 93062
rect 110296 92822 110372 93030
rect 116829 93030 116830 93062
rect 116894 93062 116900 93094
rect 116894 93030 116895 93062
rect 116829 93029 116895 93030
rect 116421 92958 116487 92959
rect 116421 92926 116422 92958
rect 28358 92758 28359 92790
rect 28293 92757 28359 92758
rect 110296 92758 110302 92822
rect 110366 92758 110372 92822
rect 110296 92752 110372 92758
rect 116416 92894 116422 92926
rect 116486 92926 116487 92958
rect 116829 92958 116895 92959
rect 116829 92926 116830 92958
rect 116486 92894 116492 92926
rect 21830 92622 21831 92654
rect 21765 92621 21831 92622
rect 22576 92622 22582 92686
rect 22646 92622 22652 92686
rect 28565 92686 28631 92687
rect 28565 92654 28566 92686
rect 22576 92616 22652 92622
rect 28560 92622 28566 92654
rect 28630 92654 28631 92686
rect 110301 92686 110367 92687
rect 110301 92654 110302 92686
rect 28630 92622 28636 92654
rect 21901 92550 21967 92551
rect 21901 92518 21902 92550
rect 21896 92486 21902 92518
rect 21966 92518 21967 92550
rect 21966 92486 21972 92518
rect 21896 92278 21972 92486
rect 28429 92414 28495 92415
rect 28429 92382 28430 92414
rect 21896 92214 21902 92278
rect 21966 92214 21972 92278
rect 21896 92208 21972 92214
rect 28424 92350 28430 92382
rect 28494 92382 28495 92414
rect 28560 92414 28636 92622
rect 28494 92350 28500 92382
rect 21760 92142 21836 92148
rect 21760 92078 21766 92142
rect 21830 92078 21836 92142
rect 22445 92142 22511 92143
rect 22445 92110 22446 92142
rect 21760 91870 21836 92078
rect 21760 91838 21766 91870
rect 21765 91806 21766 91838
rect 21830 91838 21836 91870
rect 22440 92078 22446 92110
rect 22510 92110 22511 92142
rect 23125 92142 23191 92143
rect 23125 92110 23126 92142
rect 22510 92078 22516 92110
rect 22440 91870 22516 92078
rect 21830 91806 21831 91838
rect 21765 91805 21831 91806
rect 22440 91806 22446 91870
rect 22510 91806 22516 91870
rect 22440 91800 22516 91806
rect 23120 92078 23126 92110
rect 23190 92110 23191 92142
rect 23528 92142 23604 92148
rect 23190 92078 23196 92110
rect 23120 91870 23196 92078
rect 23120 91806 23126 91870
rect 23190 91806 23196 91870
rect 23528 92078 23534 92142
rect 23598 92078 23604 92142
rect 23528 91870 23604 92078
rect 28424 92142 28500 92350
rect 28560 92350 28566 92414
rect 28630 92350 28636 92414
rect 28560 92344 28636 92350
rect 110296 92622 110302 92654
rect 110366 92654 110367 92686
rect 116416 92686 116492 92894
rect 110366 92622 110372 92654
rect 110296 92414 110372 92622
rect 116416 92622 116422 92686
rect 116486 92622 116492 92686
rect 116416 92616 116492 92622
rect 116824 92894 116830 92926
rect 116894 92926 116895 92958
rect 137496 92958 137844 94390
rect 116894 92894 116900 92926
rect 116824 92686 116900 92894
rect 116824 92622 116830 92686
rect 116894 92622 116900 92686
rect 116824 92616 116900 92622
rect 137496 92894 137502 92958
rect 137566 92894 137844 92958
rect 110296 92350 110302 92414
rect 110366 92350 110372 92414
rect 110296 92344 110372 92350
rect 116960 92550 117036 92556
rect 116960 92486 116966 92550
rect 117030 92486 117036 92550
rect 116960 92278 117036 92486
rect 116960 92246 116966 92278
rect 116965 92214 116966 92246
rect 117030 92246 117036 92278
rect 117030 92214 117031 92246
rect 116965 92213 117031 92214
rect 28424 92078 28430 92142
rect 28494 92078 28500 92142
rect 28424 92072 28500 92078
rect 115328 92142 115404 92148
rect 115328 92078 115334 92142
rect 115398 92078 115404 92142
rect 115605 92142 115671 92143
rect 115605 92110 115606 92142
rect 23528 91838 23534 91870
rect 23120 91800 23196 91806
rect 23533 91806 23534 91838
rect 23598 91838 23604 91870
rect 110432 91870 110508 91876
rect 23598 91806 23599 91838
rect 23533 91805 23599 91806
rect 110432 91806 110438 91870
rect 110502 91806 110508 91870
rect 115328 91870 115404 92078
rect 115328 91838 115334 91870
rect 21765 91734 21831 91735
rect 21765 91702 21766 91734
rect 21760 91670 21766 91702
rect 21830 91702 21831 91734
rect 22304 91734 22380 91740
rect 21830 91670 21836 91702
rect 21760 91462 21836 91670
rect 21760 91398 21766 91462
rect 21830 91398 21836 91462
rect 22304 91670 22310 91734
rect 22374 91670 22380 91734
rect 22304 91462 22380 91670
rect 22304 91430 22310 91462
rect 21760 91392 21836 91398
rect 22309 91398 22310 91430
rect 22374 91430 22380 91462
rect 22712 91734 22788 91740
rect 22712 91670 22718 91734
rect 22782 91670 22788 91734
rect 22712 91462 22788 91670
rect 22712 91430 22718 91462
rect 22374 91398 22375 91430
rect 22309 91397 22375 91398
rect 22717 91398 22718 91430
rect 22782 91430 22788 91462
rect 22984 91734 23060 91740
rect 22984 91670 22990 91734
rect 23054 91670 23060 91734
rect 23533 91734 23599 91735
rect 23533 91702 23534 91734
rect 22984 91462 23060 91670
rect 22984 91430 22990 91462
rect 22782 91398 22783 91430
rect 22717 91397 22783 91398
rect 22989 91398 22990 91430
rect 23054 91430 23060 91462
rect 23528 91670 23534 91702
rect 23598 91702 23599 91734
rect 23598 91670 23604 91702
rect 23528 91462 23604 91670
rect 110432 91598 110508 91806
rect 115333 91806 115334 91838
rect 115398 91838 115404 91870
rect 115600 92078 115606 92110
rect 115670 92110 115671 92142
rect 116285 92142 116351 92143
rect 116285 92110 116286 92142
rect 115670 92078 115676 92110
rect 115600 91870 115676 92078
rect 115398 91806 115399 91838
rect 115333 91805 115399 91806
rect 115600 91806 115606 91870
rect 115670 91806 115676 91870
rect 115600 91800 115676 91806
rect 116280 92078 116286 92110
rect 116350 92110 116351 92142
rect 116965 92142 117031 92143
rect 116965 92110 116966 92142
rect 116350 92078 116356 92110
rect 116280 91870 116356 92078
rect 116280 91806 116286 91870
rect 116350 91806 116356 91870
rect 116280 91800 116356 91806
rect 116960 92078 116966 92110
rect 117030 92110 117031 92142
rect 117030 92078 117036 92110
rect 116960 91870 117036 92078
rect 116960 91806 116966 91870
rect 117030 91806 117036 91870
rect 116960 91800 117036 91806
rect 115333 91734 115399 91735
rect 115333 91702 115334 91734
rect 110432 91566 110438 91598
rect 110437 91534 110438 91566
rect 110502 91566 110508 91598
rect 115328 91670 115334 91702
rect 115398 91702 115399 91734
rect 115600 91734 115676 91740
rect 115398 91670 115404 91702
rect 110502 91534 110503 91566
rect 110437 91533 110503 91534
rect 23054 91398 23055 91430
rect 22989 91397 23055 91398
rect 23528 91398 23534 91462
rect 23598 91398 23604 91462
rect 23528 91392 23604 91398
rect 115328 91462 115404 91670
rect 115328 91398 115334 91462
rect 115398 91398 115404 91462
rect 115600 91670 115606 91734
rect 115670 91670 115676 91734
rect 116149 91734 116215 91735
rect 116149 91702 116150 91734
rect 115600 91462 115676 91670
rect 115600 91430 115606 91462
rect 115328 91392 115404 91398
rect 115605 91398 115606 91430
rect 115670 91430 115676 91462
rect 116144 91670 116150 91702
rect 116214 91702 116215 91734
rect 116960 91734 117036 91740
rect 116214 91670 116220 91702
rect 116144 91462 116220 91670
rect 115670 91398 115671 91430
rect 115605 91397 115671 91398
rect 116144 91398 116150 91462
rect 116214 91398 116220 91462
rect 116960 91670 116966 91734
rect 117030 91670 117036 91734
rect 116960 91462 117036 91670
rect 116960 91430 116966 91462
rect 116144 91392 116220 91398
rect 116965 91398 116966 91430
rect 117030 91430 117036 91462
rect 117030 91398 117031 91430
rect 116965 91397 117031 91398
rect 952 91126 1230 91190
rect 1294 91126 1300 91190
rect 952 89558 1300 91126
rect 21896 91326 21972 91332
rect 21896 91262 21902 91326
rect 21966 91262 21972 91326
rect 21896 91054 21972 91262
rect 21896 91022 21902 91054
rect 21901 90990 21902 91022
rect 21966 91022 21972 91054
rect 22168 91326 22244 91332
rect 22168 91262 22174 91326
rect 22238 91262 22244 91326
rect 22168 91054 22244 91262
rect 22168 91022 22174 91054
rect 21966 90990 21967 91022
rect 21901 90989 21967 90990
rect 22173 90990 22174 91022
rect 22238 91022 22244 91054
rect 22712 91326 22788 91332
rect 22712 91262 22718 91326
rect 22782 91262 22788 91326
rect 22989 91326 23055 91327
rect 22989 91294 22990 91326
rect 22712 91054 22788 91262
rect 22712 91022 22718 91054
rect 22238 90990 22239 91022
rect 22173 90989 22239 90990
rect 22717 90990 22718 91022
rect 22782 91022 22788 91054
rect 22984 91262 22990 91294
rect 23054 91294 23055 91326
rect 23397 91326 23463 91327
rect 23397 91294 23398 91326
rect 23054 91262 23060 91294
rect 22984 91054 23060 91262
rect 22782 90990 22783 91022
rect 22717 90989 22783 90990
rect 22984 90990 22990 91054
rect 23054 90990 23060 91054
rect 22984 90984 23060 90990
rect 23392 91262 23398 91294
rect 23462 91294 23463 91326
rect 115197 91326 115263 91327
rect 115197 91294 115198 91326
rect 23462 91262 23468 91294
rect 23392 91054 23468 91262
rect 23392 90990 23398 91054
rect 23462 90990 23468 91054
rect 23392 90984 23468 90990
rect 115192 91262 115198 91294
rect 115262 91294 115263 91326
rect 115605 91326 115671 91327
rect 115605 91294 115606 91326
rect 115262 91262 115268 91294
rect 115192 91054 115268 91262
rect 115192 90990 115198 91054
rect 115262 90990 115268 91054
rect 115192 90984 115268 90990
rect 115600 91262 115606 91294
rect 115670 91294 115671 91326
rect 116144 91326 116220 91332
rect 115670 91262 115676 91294
rect 115600 91054 115676 91262
rect 115600 90990 115606 91054
rect 115670 90990 115676 91054
rect 116144 91262 116150 91326
rect 116214 91262 116220 91326
rect 116965 91326 117031 91327
rect 116965 91294 116966 91326
rect 116144 91054 116220 91262
rect 116144 91022 116150 91054
rect 115600 90984 115676 90990
rect 116149 90990 116150 91022
rect 116214 91022 116220 91054
rect 116960 91262 116966 91294
rect 117030 91294 117031 91326
rect 117030 91262 117036 91294
rect 116960 91054 117036 91262
rect 116214 90990 116215 91022
rect 116149 90989 116215 90990
rect 116960 90990 116966 91054
rect 117030 90990 117036 91054
rect 116960 90984 117036 90990
rect 137496 91190 137844 92894
rect 137496 91126 137502 91190
rect 137566 91126 137844 91190
rect 21765 90918 21831 90919
rect 21765 90886 21766 90918
rect 21760 90854 21766 90886
rect 21830 90886 21831 90918
rect 22173 90918 22239 90919
rect 22173 90886 22174 90918
rect 21830 90854 21836 90886
rect 21760 90646 21836 90854
rect 21760 90582 21766 90646
rect 21830 90582 21836 90646
rect 21760 90576 21836 90582
rect 22168 90854 22174 90886
rect 22238 90886 22239 90918
rect 22581 90918 22647 90919
rect 22581 90886 22582 90918
rect 22238 90854 22244 90886
rect 22168 90646 22244 90854
rect 22168 90582 22174 90646
rect 22238 90582 22244 90646
rect 22168 90576 22244 90582
rect 22576 90854 22582 90886
rect 22646 90886 22647 90918
rect 22989 90918 23055 90919
rect 22989 90886 22990 90918
rect 22646 90854 22652 90886
rect 22576 90646 22652 90854
rect 22576 90582 22582 90646
rect 22646 90582 22652 90646
rect 22576 90576 22652 90582
rect 22984 90854 22990 90886
rect 23054 90886 23055 90918
rect 23528 90918 23604 90924
rect 23054 90854 23060 90886
rect 22984 90646 23060 90854
rect 22984 90582 22990 90646
rect 23054 90582 23060 90646
rect 23528 90854 23534 90918
rect 23598 90854 23604 90918
rect 115333 90918 115399 90919
rect 115333 90886 115334 90918
rect 23528 90646 23604 90854
rect 23528 90614 23534 90646
rect 22984 90576 23060 90582
rect 23533 90582 23534 90614
rect 23598 90614 23604 90646
rect 115328 90854 115334 90886
rect 115398 90886 115399 90918
rect 115736 90918 115812 90924
rect 115398 90854 115404 90886
rect 115328 90646 115404 90854
rect 23598 90582 23599 90614
rect 23533 90581 23599 90582
rect 115328 90582 115334 90646
rect 115398 90582 115404 90646
rect 115736 90854 115742 90918
rect 115806 90854 115812 90918
rect 116421 90918 116487 90919
rect 116421 90886 116422 90918
rect 115736 90646 115812 90854
rect 115736 90614 115742 90646
rect 115328 90576 115404 90582
rect 115741 90582 115742 90614
rect 115806 90614 115812 90646
rect 116416 90854 116422 90886
rect 116486 90886 116487 90918
rect 116824 90918 116900 90924
rect 116486 90854 116492 90886
rect 116416 90646 116492 90854
rect 115806 90582 115807 90614
rect 115741 90581 115807 90582
rect 116416 90582 116422 90646
rect 116486 90582 116492 90646
rect 116824 90854 116830 90918
rect 116894 90854 116900 90918
rect 116824 90646 116900 90854
rect 116824 90614 116830 90646
rect 116416 90576 116492 90582
rect 116829 90582 116830 90614
rect 116894 90614 116900 90646
rect 116894 90582 116895 90614
rect 116829 90581 116895 90582
rect 22440 90510 22516 90516
rect 22440 90446 22446 90510
rect 22510 90446 22516 90510
rect 23125 90510 23191 90511
rect 23125 90478 23126 90510
rect 22440 90238 22516 90446
rect 22440 90206 22446 90238
rect 22445 90174 22446 90206
rect 22510 90206 22516 90238
rect 23120 90446 23126 90478
rect 23190 90478 23191 90510
rect 23533 90510 23599 90511
rect 23533 90478 23534 90510
rect 23190 90446 23196 90478
rect 23120 90238 23196 90446
rect 22510 90174 22511 90206
rect 22445 90173 22511 90174
rect 23120 90174 23126 90238
rect 23190 90174 23196 90238
rect 23120 90168 23196 90174
rect 23528 90446 23534 90478
rect 23598 90478 23599 90510
rect 115333 90510 115399 90511
rect 115333 90478 115334 90510
rect 23598 90446 23604 90478
rect 23528 90238 23604 90446
rect 23528 90174 23534 90238
rect 23598 90174 23604 90238
rect 23528 90168 23604 90174
rect 115328 90446 115334 90478
rect 115398 90478 115399 90510
rect 115741 90510 115807 90511
rect 115741 90478 115742 90510
rect 115398 90446 115404 90478
rect 115328 90238 115404 90446
rect 115328 90174 115334 90238
rect 115398 90174 115404 90238
rect 115328 90168 115404 90174
rect 115736 90446 115742 90478
rect 115806 90478 115807 90510
rect 116149 90510 116215 90511
rect 116149 90478 116150 90510
rect 115806 90446 115812 90478
rect 115736 90238 115812 90446
rect 115736 90174 115742 90238
rect 115806 90174 115812 90238
rect 115736 90168 115812 90174
rect 116144 90446 116150 90478
rect 116214 90478 116215 90510
rect 116280 90510 116356 90516
rect 116214 90446 116220 90478
rect 116144 90238 116220 90446
rect 116144 90174 116150 90238
rect 116214 90174 116220 90238
rect 116280 90446 116286 90510
rect 116350 90446 116356 90510
rect 116280 90238 116356 90446
rect 116280 90206 116286 90238
rect 116144 90168 116220 90174
rect 116285 90174 116286 90206
rect 116350 90206 116356 90238
rect 116350 90174 116351 90206
rect 116285 90173 116351 90174
rect 21765 90102 21831 90103
rect 21765 90070 21766 90102
rect 21760 90038 21766 90070
rect 21830 90070 21831 90102
rect 22168 90102 22244 90108
rect 21830 90038 21836 90070
rect 21760 89830 21836 90038
rect 21760 89766 21766 89830
rect 21830 89766 21836 89830
rect 22168 90038 22174 90102
rect 22238 90038 22244 90102
rect 22168 89830 22244 90038
rect 22168 89798 22174 89830
rect 21760 89760 21836 89766
rect 22173 89766 22174 89798
rect 22238 89798 22244 89830
rect 22984 90102 23060 90108
rect 22984 90038 22990 90102
rect 23054 90038 23060 90102
rect 22984 89830 23060 90038
rect 22984 89798 22990 89830
rect 22238 89766 22239 89798
rect 22173 89765 22239 89766
rect 22989 89766 22990 89798
rect 23054 89798 23060 89830
rect 23528 90102 23604 90108
rect 23528 90038 23534 90102
rect 23598 90038 23604 90102
rect 115197 90102 115263 90103
rect 115197 90070 115198 90102
rect 23528 89830 23604 90038
rect 23528 89798 23534 89830
rect 23054 89766 23055 89798
rect 22989 89765 23055 89766
rect 23533 89766 23534 89798
rect 23598 89798 23604 89830
rect 115192 90038 115198 90070
rect 115262 90070 115263 90102
rect 115736 90102 115812 90108
rect 115262 90038 115268 90070
rect 115192 89830 115268 90038
rect 23598 89766 23599 89798
rect 23533 89765 23599 89766
rect 115192 89766 115198 89830
rect 115262 89766 115268 89830
rect 115736 90038 115742 90102
rect 115806 90038 115812 90102
rect 115736 89830 115812 90038
rect 115736 89798 115742 89830
rect 115192 89760 115268 89766
rect 115741 89766 115742 89798
rect 115806 89798 115812 89830
rect 116008 90102 116084 90108
rect 116008 90038 116014 90102
rect 116078 90038 116084 90102
rect 116285 90102 116351 90103
rect 116285 90070 116286 90102
rect 116008 89830 116084 90038
rect 116008 89798 116014 89830
rect 115806 89766 115807 89798
rect 115741 89765 115807 89766
rect 116013 89766 116014 89798
rect 116078 89798 116084 89830
rect 116280 90038 116286 90070
rect 116350 90070 116351 90102
rect 116824 90102 116900 90108
rect 116350 90038 116356 90070
rect 116280 89830 116356 90038
rect 116078 89766 116079 89798
rect 116013 89765 116079 89766
rect 116280 89766 116286 89830
rect 116350 89766 116356 89830
rect 116824 90038 116830 90102
rect 116894 90038 116900 90102
rect 116824 89830 116900 90038
rect 116824 89798 116830 89830
rect 116280 89760 116356 89766
rect 116829 89766 116830 89798
rect 116894 89798 116900 89830
rect 116894 89766 116895 89798
rect 116829 89765 116895 89766
rect 22581 89694 22647 89695
rect 22581 89662 22582 89694
rect 952 89494 1230 89558
rect 1294 89494 1300 89558
rect 952 87654 1300 89494
rect 22576 89630 22582 89662
rect 22646 89662 22647 89694
rect 22989 89694 23055 89695
rect 22989 89662 22990 89694
rect 22646 89630 22652 89662
rect 21765 89422 21831 89423
rect 21765 89390 21766 89422
rect 21760 89358 21766 89390
rect 21830 89390 21831 89422
rect 22576 89422 22652 89630
rect 21830 89358 21836 89390
rect 21760 89150 21836 89358
rect 22576 89358 22582 89422
rect 22646 89358 22652 89422
rect 22576 89352 22652 89358
rect 22984 89630 22990 89662
rect 23054 89662 23055 89694
rect 23533 89694 23599 89695
rect 23533 89662 23534 89694
rect 23054 89630 23060 89662
rect 22984 89422 23060 89630
rect 22984 89358 22990 89422
rect 23054 89358 23060 89422
rect 22984 89352 23060 89358
rect 23528 89630 23534 89662
rect 23598 89662 23599 89694
rect 115192 89694 115268 89700
rect 23598 89630 23604 89662
rect 23528 89422 23604 89630
rect 115192 89630 115198 89694
rect 115262 89630 115268 89694
rect 23528 89358 23534 89422
rect 23598 89358 23604 89422
rect 23528 89352 23604 89358
rect 28288 89558 28364 89564
rect 28288 89494 28294 89558
rect 28358 89494 28364 89558
rect 21760 89086 21766 89150
rect 21830 89086 21836 89150
rect 21760 89080 21836 89086
rect 22440 89286 22516 89292
rect 22440 89222 22446 89286
rect 22510 89222 22516 89286
rect 28288 89286 28364 89494
rect 115192 89422 115268 89630
rect 115192 89390 115198 89422
rect 115197 89358 115198 89390
rect 115262 89390 115268 89422
rect 115736 89694 115812 89700
rect 115736 89630 115742 89694
rect 115806 89630 115812 89694
rect 115736 89422 115812 89630
rect 137496 89558 137844 91126
rect 137496 89494 137502 89558
rect 137566 89494 137844 89558
rect 115736 89390 115742 89422
rect 115262 89358 115263 89390
rect 115197 89357 115263 89358
rect 115741 89358 115742 89390
rect 115806 89390 115812 89422
rect 116960 89422 117036 89428
rect 115806 89358 115807 89390
rect 115741 89357 115807 89358
rect 116960 89358 116966 89422
rect 117030 89358 117036 89422
rect 28288 89254 28294 89286
rect 21901 89014 21967 89015
rect 21901 88982 21902 89014
rect 21896 88950 21902 88982
rect 21966 88982 21967 89014
rect 22168 89014 22244 89020
rect 21966 88950 21972 88982
rect 21896 88742 21972 88950
rect 21896 88678 21902 88742
rect 21966 88678 21972 88742
rect 21896 88672 21972 88678
rect 22168 88950 22174 89014
rect 22238 88950 22244 89014
rect 22440 89014 22516 89222
rect 28293 89222 28294 89254
rect 28358 89254 28364 89286
rect 28358 89222 28359 89254
rect 28293 89221 28359 89222
rect 116960 89150 117036 89358
rect 116960 89118 116966 89150
rect 116965 89086 116966 89118
rect 117030 89118 117036 89150
rect 117030 89086 117031 89118
rect 116965 89085 117031 89086
rect 22440 88982 22446 89014
rect 21760 88606 21836 88612
rect 21760 88542 21766 88606
rect 21830 88542 21836 88606
rect 22168 88606 22244 88950
rect 22445 88950 22446 88982
rect 22510 88982 22516 89014
rect 110165 89014 110231 89015
rect 110165 88982 110166 89014
rect 22510 88950 22511 88982
rect 22445 88949 22511 88950
rect 110160 88950 110166 88982
rect 110230 88982 110231 89014
rect 116557 89014 116623 89015
rect 116557 88982 116558 89014
rect 110230 88950 110236 88982
rect 110160 88742 110236 88950
rect 116552 88950 116558 88982
rect 116622 88982 116623 89014
rect 116824 89014 116900 89020
rect 116622 88950 116628 88982
rect 110160 88678 110166 88742
rect 110230 88678 110236 88742
rect 110301 88742 110367 88743
rect 110301 88710 110302 88742
rect 110160 88672 110236 88678
rect 110296 88678 110302 88710
rect 110366 88710 110367 88742
rect 110366 88678 110372 88710
rect 22168 88574 22174 88606
rect 21760 88334 21836 88542
rect 22173 88542 22174 88574
rect 22238 88574 22244 88606
rect 22238 88542 22239 88574
rect 22173 88541 22239 88542
rect 110296 88470 110372 88678
rect 116552 88606 116628 88950
rect 116824 88950 116830 89014
rect 116894 88950 116900 89014
rect 116824 88742 116900 88950
rect 116824 88710 116830 88742
rect 116829 88678 116830 88710
rect 116894 88710 116900 88742
rect 116894 88678 116895 88710
rect 116829 88677 116895 88678
rect 116552 88542 116558 88606
rect 116622 88542 116628 88606
rect 116829 88606 116895 88607
rect 116829 88574 116830 88606
rect 116552 88536 116628 88542
rect 116824 88542 116830 88574
rect 116894 88574 116895 88606
rect 116894 88542 116900 88574
rect 110296 88406 110302 88470
rect 110366 88406 110372 88470
rect 110296 88400 110372 88406
rect 110432 88470 110508 88476
rect 110432 88406 110438 88470
rect 110502 88406 110508 88470
rect 21760 88302 21766 88334
rect 21765 88270 21766 88302
rect 21830 88302 21836 88334
rect 21830 88270 21831 88302
rect 21765 88269 21831 88270
rect 21896 88198 21972 88204
rect 21896 88134 21902 88198
rect 21966 88134 21972 88198
rect 21896 87926 21972 88134
rect 21896 87894 21902 87926
rect 21901 87862 21902 87894
rect 21966 87894 21972 87926
rect 22712 88198 22788 88204
rect 22712 88134 22718 88198
rect 22782 88134 22788 88198
rect 22712 87926 22788 88134
rect 22712 87894 22718 87926
rect 21966 87862 21967 87894
rect 21901 87861 21967 87862
rect 22717 87862 22718 87894
rect 22782 87894 22788 87926
rect 23120 88198 23196 88204
rect 23120 88134 23126 88198
rect 23190 88134 23196 88198
rect 23120 87926 23196 88134
rect 23120 87894 23126 87926
rect 22782 87862 22783 87894
rect 22717 87861 22783 87862
rect 23125 87862 23126 87894
rect 23190 87894 23196 87926
rect 23392 88198 23468 88204
rect 23392 88134 23398 88198
rect 23462 88134 23468 88198
rect 110432 88198 110508 88406
rect 116280 88470 116356 88476
rect 116280 88406 116286 88470
rect 116350 88406 116356 88470
rect 110432 88166 110438 88198
rect 23392 87926 23468 88134
rect 110437 88134 110438 88166
rect 110502 88166 110508 88198
rect 115192 88198 115268 88204
rect 110502 88134 110503 88166
rect 110437 88133 110503 88134
rect 115192 88134 115198 88198
rect 115262 88134 115268 88198
rect 115605 88198 115671 88199
rect 115605 88166 115606 88198
rect 23392 87894 23398 87926
rect 23190 87862 23191 87894
rect 23125 87861 23191 87862
rect 23397 87862 23398 87894
rect 23462 87894 23468 87926
rect 28288 87926 28364 87932
rect 23462 87862 23463 87894
rect 23397 87861 23463 87862
rect 28288 87862 28294 87926
rect 28358 87862 28364 87926
rect 115192 87926 115268 88134
rect 115192 87894 115198 87926
rect 952 87590 1230 87654
rect 1294 87590 1300 87654
rect 952 86158 1300 87590
rect 21760 87790 21836 87796
rect 21760 87726 21766 87790
rect 21830 87726 21836 87790
rect 23125 87790 23191 87791
rect 23125 87758 23126 87790
rect 21760 87518 21836 87726
rect 21760 87486 21766 87518
rect 21765 87454 21766 87486
rect 21830 87486 21836 87518
rect 23120 87726 23126 87758
rect 23190 87758 23191 87790
rect 23528 87790 23604 87796
rect 23190 87726 23196 87758
rect 23120 87518 23196 87726
rect 21830 87454 21831 87486
rect 21765 87453 21831 87454
rect 23120 87454 23126 87518
rect 23190 87454 23196 87518
rect 23528 87726 23534 87790
rect 23598 87726 23604 87790
rect 23528 87518 23604 87726
rect 28288 87654 28364 87862
rect 115197 87862 115198 87894
rect 115262 87894 115268 87926
rect 115600 88134 115606 88166
rect 115670 88166 115671 88198
rect 116280 88198 116356 88406
rect 116824 88334 116900 88542
rect 116824 88270 116830 88334
rect 116894 88270 116900 88334
rect 116824 88264 116900 88270
rect 116280 88166 116286 88198
rect 115670 88134 115676 88166
rect 115600 87926 115676 88134
rect 116285 88134 116286 88166
rect 116350 88166 116356 88198
rect 116552 88198 116628 88204
rect 116350 88134 116351 88166
rect 116285 88133 116351 88134
rect 116552 88134 116558 88198
rect 116622 88134 116628 88198
rect 115262 87862 115263 87894
rect 115197 87861 115263 87862
rect 115600 87862 115606 87926
rect 115670 87862 115676 87926
rect 116552 87926 116628 88134
rect 116552 87894 116558 87926
rect 115600 87856 115676 87862
rect 116557 87862 116558 87894
rect 116622 87894 116628 87926
rect 116960 88198 117036 88204
rect 116960 88134 116966 88198
rect 117030 88134 117036 88198
rect 116960 87926 117036 88134
rect 116960 87894 116966 87926
rect 116622 87862 116623 87894
rect 116557 87861 116623 87862
rect 116965 87862 116966 87894
rect 117030 87894 117036 87926
rect 117030 87862 117031 87894
rect 116965 87861 117031 87862
rect 28288 87622 28294 87654
rect 28293 87590 28294 87622
rect 28358 87622 28364 87654
rect 115328 87790 115404 87796
rect 115328 87726 115334 87790
rect 115398 87726 115404 87790
rect 28358 87590 28359 87622
rect 28293 87589 28359 87590
rect 23528 87486 23534 87518
rect 23120 87448 23196 87454
rect 23533 87454 23534 87486
rect 23598 87486 23604 87518
rect 115328 87518 115404 87726
rect 115328 87486 115334 87518
rect 23598 87454 23599 87486
rect 23533 87453 23599 87454
rect 115333 87454 115334 87486
rect 115398 87486 115404 87518
rect 115736 87790 115812 87796
rect 115736 87726 115742 87790
rect 115806 87726 115812 87790
rect 116149 87790 116215 87791
rect 116149 87758 116150 87790
rect 115736 87518 115812 87726
rect 115736 87486 115742 87518
rect 115398 87454 115399 87486
rect 115333 87453 115399 87454
rect 115741 87454 115742 87486
rect 115806 87486 115812 87518
rect 116144 87726 116150 87758
rect 116214 87758 116215 87790
rect 116280 87790 116356 87796
rect 116214 87726 116220 87758
rect 116144 87518 116220 87726
rect 115806 87454 115807 87486
rect 115741 87453 115807 87454
rect 116144 87454 116150 87518
rect 116214 87454 116220 87518
rect 116280 87726 116286 87790
rect 116350 87726 116356 87790
rect 116280 87518 116356 87726
rect 116280 87486 116286 87518
rect 116144 87448 116220 87454
rect 116285 87454 116286 87486
rect 116350 87486 116356 87518
rect 116416 87790 116492 87796
rect 116416 87726 116422 87790
rect 116486 87726 116492 87790
rect 116965 87790 117031 87791
rect 116965 87758 116966 87790
rect 116416 87518 116492 87726
rect 116416 87486 116422 87518
rect 116350 87454 116351 87486
rect 116285 87453 116351 87454
rect 116421 87454 116422 87486
rect 116486 87486 116492 87518
rect 116960 87726 116966 87758
rect 117030 87758 117031 87790
rect 137496 87790 137844 89494
rect 117030 87726 117036 87758
rect 116960 87518 117036 87726
rect 116486 87454 116487 87486
rect 116421 87453 116487 87454
rect 116960 87454 116966 87518
rect 117030 87454 117036 87518
rect 116960 87448 117036 87454
rect 137496 87726 137502 87790
rect 137566 87726 137844 87790
rect 21765 87382 21831 87383
rect 21765 87350 21766 87382
rect 21760 87318 21766 87350
rect 21830 87350 21831 87382
rect 22173 87382 22239 87383
rect 22173 87350 22174 87382
rect 21830 87318 21836 87350
rect 21760 87110 21836 87318
rect 21760 87046 21766 87110
rect 21830 87046 21836 87110
rect 21760 87040 21836 87046
rect 22168 87318 22174 87350
rect 22238 87350 22239 87382
rect 22581 87382 22647 87383
rect 22581 87350 22582 87382
rect 22238 87318 22244 87350
rect 22168 87110 22244 87318
rect 22168 87046 22174 87110
rect 22238 87046 22244 87110
rect 22168 87040 22244 87046
rect 22576 87318 22582 87350
rect 22646 87350 22647 87382
rect 22984 87382 23060 87388
rect 22646 87318 22652 87350
rect 22576 87110 22652 87318
rect 22576 87046 22582 87110
rect 22646 87046 22652 87110
rect 22984 87318 22990 87382
rect 23054 87318 23060 87382
rect 23533 87382 23599 87383
rect 23533 87350 23534 87382
rect 22984 87110 23060 87318
rect 22984 87078 22990 87110
rect 22576 87040 22652 87046
rect 22989 87046 22990 87078
rect 23054 87078 23060 87110
rect 23528 87318 23534 87350
rect 23598 87350 23599 87382
rect 115192 87382 115268 87388
rect 23598 87318 23604 87350
rect 23528 87110 23604 87318
rect 23054 87046 23055 87078
rect 22989 87045 23055 87046
rect 23528 87046 23534 87110
rect 23598 87046 23604 87110
rect 115192 87318 115198 87382
rect 115262 87318 115268 87382
rect 115741 87382 115807 87383
rect 115741 87350 115742 87382
rect 115192 87110 115268 87318
rect 115192 87078 115198 87110
rect 23528 87040 23604 87046
rect 115197 87046 115198 87078
rect 115262 87078 115268 87110
rect 115736 87318 115742 87350
rect 115806 87350 115807 87382
rect 116008 87382 116084 87388
rect 115806 87318 115812 87350
rect 115736 87110 115812 87318
rect 115262 87046 115263 87078
rect 115197 87045 115263 87046
rect 115736 87046 115742 87110
rect 115806 87046 115812 87110
rect 116008 87318 116014 87382
rect 116078 87318 116084 87382
rect 116285 87382 116351 87383
rect 116285 87350 116286 87382
rect 116008 87110 116084 87318
rect 116008 87078 116014 87110
rect 115736 87040 115812 87046
rect 116013 87046 116014 87078
rect 116078 87078 116084 87110
rect 116280 87318 116286 87350
rect 116350 87350 116351 87382
rect 116960 87382 117036 87388
rect 116350 87318 116356 87350
rect 116280 87110 116356 87318
rect 116078 87046 116079 87078
rect 116013 87045 116079 87046
rect 116280 87046 116286 87110
rect 116350 87046 116356 87110
rect 116960 87318 116966 87382
rect 117030 87318 117036 87382
rect 116960 87110 117036 87318
rect 116960 87078 116966 87110
rect 116280 87040 116356 87046
rect 116965 87046 116966 87078
rect 117030 87078 117036 87110
rect 117030 87046 117031 87078
rect 116965 87045 117031 87046
rect 21901 86974 21967 86975
rect 21901 86942 21902 86974
rect 21896 86910 21902 86942
rect 21966 86942 21967 86974
rect 23120 86974 23196 86980
rect 21966 86910 21972 86942
rect 21896 86702 21972 86910
rect 21896 86638 21902 86702
rect 21966 86638 21972 86702
rect 23120 86910 23126 86974
rect 23190 86910 23196 86974
rect 23120 86702 23196 86910
rect 23120 86670 23126 86702
rect 21896 86632 21972 86638
rect 23125 86638 23126 86670
rect 23190 86670 23196 86702
rect 23392 86974 23468 86980
rect 23392 86910 23398 86974
rect 23462 86910 23468 86974
rect 115197 86974 115263 86975
rect 115197 86942 115198 86974
rect 23392 86702 23468 86910
rect 23392 86670 23398 86702
rect 23190 86638 23191 86670
rect 23125 86637 23191 86638
rect 23397 86638 23398 86670
rect 23462 86670 23468 86702
rect 115192 86910 115198 86942
rect 115262 86942 115263 86974
rect 115600 86974 115676 86980
rect 115262 86910 115268 86942
rect 115192 86702 115268 86910
rect 23462 86638 23463 86670
rect 23397 86637 23463 86638
rect 115192 86638 115198 86702
rect 115262 86638 115268 86702
rect 115600 86910 115606 86974
rect 115670 86910 115676 86974
rect 115600 86702 115676 86910
rect 115600 86670 115606 86702
rect 115192 86632 115268 86638
rect 115605 86638 115606 86670
rect 115670 86670 115676 86702
rect 116144 86974 116220 86980
rect 116144 86910 116150 86974
rect 116214 86910 116220 86974
rect 116965 86974 117031 86975
rect 116965 86942 116966 86974
rect 116144 86702 116220 86910
rect 116144 86670 116150 86702
rect 115670 86638 115671 86670
rect 115605 86637 115671 86638
rect 116149 86638 116150 86670
rect 116214 86670 116220 86702
rect 116960 86910 116966 86942
rect 117030 86942 117031 86974
rect 117030 86910 117036 86942
rect 116960 86702 117036 86910
rect 116214 86638 116215 86670
rect 116149 86637 116215 86638
rect 116960 86638 116966 86702
rect 117030 86638 117036 86702
rect 116960 86632 117036 86638
rect 21760 86566 21836 86572
rect 21760 86502 21766 86566
rect 21830 86502 21836 86566
rect 22445 86566 22511 86567
rect 22445 86534 22446 86566
rect 21760 86294 21836 86502
rect 21760 86262 21766 86294
rect 21765 86230 21766 86262
rect 21830 86262 21836 86294
rect 22440 86502 22446 86534
rect 22510 86534 22511 86566
rect 22989 86566 23055 86567
rect 22989 86534 22990 86566
rect 22510 86502 22516 86534
rect 22440 86294 22516 86502
rect 21830 86230 21831 86262
rect 21765 86229 21831 86230
rect 22440 86230 22446 86294
rect 22510 86230 22516 86294
rect 22440 86224 22516 86230
rect 22984 86502 22990 86534
rect 23054 86534 23055 86566
rect 23528 86566 23604 86572
rect 23054 86502 23060 86534
rect 22984 86294 23060 86502
rect 22984 86230 22990 86294
rect 23054 86230 23060 86294
rect 23528 86502 23534 86566
rect 23598 86502 23604 86566
rect 23528 86294 23604 86502
rect 23528 86262 23534 86294
rect 22984 86224 23060 86230
rect 23533 86230 23534 86262
rect 23598 86262 23604 86294
rect 115328 86566 115404 86572
rect 115328 86502 115334 86566
rect 115398 86502 115404 86566
rect 115741 86566 115807 86567
rect 115741 86534 115742 86566
rect 115328 86294 115404 86502
rect 115328 86262 115334 86294
rect 23598 86230 23599 86262
rect 23533 86229 23599 86230
rect 115333 86230 115334 86262
rect 115398 86262 115404 86294
rect 115736 86502 115742 86534
rect 115806 86534 115807 86566
rect 116013 86566 116079 86567
rect 116013 86534 116014 86566
rect 115806 86502 115812 86534
rect 115736 86294 115812 86502
rect 115398 86230 115399 86262
rect 115333 86229 115399 86230
rect 115736 86230 115742 86294
rect 115806 86230 115812 86294
rect 115736 86224 115812 86230
rect 116008 86502 116014 86534
rect 116078 86534 116079 86566
rect 116421 86566 116487 86567
rect 116421 86534 116422 86566
rect 116078 86502 116084 86534
rect 116008 86294 116084 86502
rect 116008 86230 116014 86294
rect 116078 86230 116084 86294
rect 116008 86224 116084 86230
rect 116416 86502 116422 86534
rect 116486 86534 116487 86566
rect 116824 86566 116900 86572
rect 116486 86502 116492 86534
rect 116416 86294 116492 86502
rect 116416 86230 116422 86294
rect 116486 86230 116492 86294
rect 116824 86502 116830 86566
rect 116894 86502 116900 86566
rect 116824 86294 116900 86502
rect 116824 86262 116830 86294
rect 116416 86224 116492 86230
rect 116829 86230 116830 86262
rect 116894 86262 116900 86294
rect 116894 86230 116895 86262
rect 116829 86229 116895 86230
rect 952 86094 1230 86158
rect 1294 86094 1300 86158
rect 21765 86158 21831 86159
rect 21765 86126 21766 86158
rect 952 84390 1300 86094
rect 21760 86094 21766 86126
rect 21830 86126 21831 86158
rect 22304 86158 22380 86164
rect 21830 86094 21836 86126
rect 21760 85886 21836 86094
rect 21760 85822 21766 85886
rect 21830 85822 21836 85886
rect 22304 86094 22310 86158
rect 22374 86094 22380 86158
rect 22304 85886 22380 86094
rect 22304 85854 22310 85886
rect 21760 85816 21836 85822
rect 22309 85822 22310 85854
rect 22374 85854 22380 85886
rect 22984 86158 23060 86164
rect 22984 86094 22990 86158
rect 23054 86094 23060 86158
rect 23533 86158 23599 86159
rect 23533 86126 23534 86158
rect 22984 85886 23060 86094
rect 22984 85854 22990 85886
rect 22374 85822 22375 85854
rect 22309 85821 22375 85822
rect 22989 85822 22990 85854
rect 23054 85854 23060 85886
rect 23528 86094 23534 86126
rect 23598 86126 23599 86158
rect 115333 86158 115399 86159
rect 115333 86126 115334 86158
rect 23598 86094 23604 86126
rect 23528 85886 23604 86094
rect 23054 85822 23055 85854
rect 22989 85821 23055 85822
rect 23528 85822 23534 85886
rect 23598 85822 23604 85886
rect 23528 85816 23604 85822
rect 115328 86094 115334 86126
rect 115398 86126 115399 86158
rect 115600 86158 115676 86164
rect 115398 86094 115404 86126
rect 115328 85886 115404 86094
rect 115328 85822 115334 85886
rect 115398 85822 115404 85886
rect 115600 86094 115606 86158
rect 115670 86094 115676 86158
rect 116829 86158 116895 86159
rect 116829 86126 116830 86158
rect 115600 85886 115676 86094
rect 115600 85854 115606 85886
rect 115328 85816 115404 85822
rect 115605 85822 115606 85854
rect 115670 85854 115676 85886
rect 116824 86094 116830 86126
rect 116894 86126 116895 86158
rect 116894 86094 116900 86126
rect 116824 85886 116900 86094
rect 115670 85822 115671 85854
rect 115605 85821 115671 85822
rect 116824 85822 116830 85886
rect 116894 85822 116900 85886
rect 116824 85816 116900 85822
rect 137496 86022 137844 87726
rect 137496 85958 137502 86022
rect 137566 85958 137844 86022
rect 22440 85750 22516 85756
rect 22440 85686 22446 85750
rect 22510 85686 22516 85750
rect 22717 85750 22783 85751
rect 22717 85718 22718 85750
rect 21765 85478 21831 85479
rect 21765 85446 21766 85478
rect 21760 85414 21766 85446
rect 21830 85446 21831 85478
rect 22440 85478 22516 85686
rect 22440 85446 22446 85478
rect 21830 85414 21836 85446
rect 21760 85206 21836 85414
rect 22445 85414 22446 85446
rect 22510 85446 22516 85478
rect 22712 85686 22718 85718
rect 22782 85718 22783 85750
rect 22984 85750 23060 85756
rect 22782 85686 22788 85718
rect 22712 85478 22788 85686
rect 22510 85414 22511 85446
rect 22445 85413 22511 85414
rect 22712 85414 22718 85478
rect 22782 85414 22788 85478
rect 22984 85686 22990 85750
rect 23054 85686 23060 85750
rect 22984 85478 23060 85686
rect 22984 85446 22990 85478
rect 22712 85408 22788 85414
rect 22989 85414 22990 85446
rect 23054 85446 23060 85478
rect 23528 85750 23604 85756
rect 23528 85686 23534 85750
rect 23598 85686 23604 85750
rect 23528 85478 23604 85686
rect 115328 85750 115404 85756
rect 115328 85686 115334 85750
rect 115398 85686 115404 85750
rect 115605 85750 115671 85751
rect 115605 85718 115606 85750
rect 110165 85614 110231 85615
rect 110165 85582 110166 85614
rect 23528 85446 23534 85478
rect 23054 85414 23055 85446
rect 22989 85413 23055 85414
rect 23533 85414 23534 85446
rect 23598 85446 23604 85478
rect 110160 85550 110166 85582
rect 110230 85582 110231 85614
rect 110230 85550 110236 85582
rect 23598 85414 23599 85446
rect 23533 85413 23599 85414
rect 22989 85342 23055 85343
rect 22989 85310 22990 85342
rect 21760 85142 21766 85206
rect 21830 85142 21836 85206
rect 21760 85136 21836 85142
rect 22984 85278 22990 85310
rect 23054 85310 23055 85342
rect 23528 85342 23604 85348
rect 23054 85278 23060 85310
rect 22984 85070 23060 85278
rect 22984 85006 22990 85070
rect 23054 85006 23060 85070
rect 23528 85278 23534 85342
rect 23598 85278 23604 85342
rect 23528 85070 23604 85278
rect 110160 85342 110236 85550
rect 115328 85478 115404 85686
rect 115328 85446 115334 85478
rect 115333 85414 115334 85446
rect 115398 85446 115404 85478
rect 115600 85686 115606 85718
rect 115670 85718 115671 85750
rect 116008 85750 116084 85756
rect 115670 85686 115676 85718
rect 115600 85478 115676 85686
rect 115398 85414 115399 85446
rect 115333 85413 115399 85414
rect 115600 85414 115606 85478
rect 115670 85414 115676 85478
rect 116008 85686 116014 85750
rect 116078 85686 116084 85750
rect 116008 85478 116084 85686
rect 116008 85446 116014 85478
rect 115600 85408 115676 85414
rect 116013 85414 116014 85446
rect 116078 85446 116084 85478
rect 116960 85478 117036 85484
rect 116078 85414 116079 85446
rect 116013 85413 116079 85414
rect 116960 85414 116966 85478
rect 117030 85414 117036 85478
rect 110160 85278 110166 85342
rect 110230 85278 110236 85342
rect 110160 85272 110236 85278
rect 115328 85342 115404 85348
rect 115328 85278 115334 85342
rect 115398 85278 115404 85342
rect 115741 85342 115807 85343
rect 115741 85310 115742 85342
rect 23528 85038 23534 85070
rect 22984 85000 23060 85006
rect 23533 85006 23534 85038
rect 23598 85038 23604 85070
rect 115328 85070 115404 85278
rect 115328 85038 115334 85070
rect 23598 85006 23599 85038
rect 23533 85005 23599 85006
rect 115333 85006 115334 85038
rect 115398 85038 115404 85070
rect 115736 85278 115742 85310
rect 115806 85310 115807 85342
rect 115806 85278 115812 85310
rect 115736 85070 115812 85278
rect 116960 85206 117036 85414
rect 116960 85174 116966 85206
rect 116965 85142 116966 85174
rect 117030 85174 117036 85206
rect 117030 85142 117031 85174
rect 116965 85141 117031 85142
rect 115398 85006 115399 85038
rect 115333 85005 115399 85006
rect 115736 85006 115742 85070
rect 115806 85006 115812 85070
rect 115736 85000 115812 85006
rect 22712 84934 22788 84940
rect 22712 84870 22718 84934
rect 22782 84870 22788 84934
rect 21901 84662 21967 84663
rect 21901 84630 21902 84662
rect 952 84326 1230 84390
rect 1294 84326 1300 84390
rect 952 82758 1300 84326
rect 21896 84598 21902 84630
rect 21966 84630 21967 84662
rect 22712 84662 22788 84870
rect 116552 84934 116628 84940
rect 116552 84870 116558 84934
rect 116622 84870 116628 84934
rect 28565 84798 28631 84799
rect 28565 84766 28566 84798
rect 22712 84630 22718 84662
rect 21966 84598 21972 84630
rect 21896 84390 21972 84598
rect 22717 84598 22718 84630
rect 22782 84630 22788 84662
rect 28560 84734 28566 84766
rect 28630 84766 28631 84798
rect 28630 84734 28636 84766
rect 22782 84598 22783 84630
rect 22717 84597 22783 84598
rect 28560 84526 28636 84734
rect 116552 84662 116628 84870
rect 116552 84630 116558 84662
rect 116557 84598 116558 84630
rect 116622 84630 116628 84662
rect 116965 84662 117031 84663
rect 116965 84630 116966 84662
rect 116622 84598 116623 84630
rect 116557 84597 116623 84598
rect 116960 84598 116966 84630
rect 117030 84630 117031 84662
rect 117030 84598 117036 84630
rect 28560 84462 28566 84526
rect 28630 84462 28636 84526
rect 28560 84456 28636 84462
rect 21896 84326 21902 84390
rect 21966 84326 21972 84390
rect 28429 84390 28495 84391
rect 28429 84358 28430 84390
rect 21896 84320 21972 84326
rect 28424 84326 28430 84358
rect 28494 84358 28495 84390
rect 110160 84390 110236 84396
rect 28494 84326 28500 84358
rect 21760 84254 21836 84260
rect 21760 84190 21766 84254
rect 21830 84190 21836 84254
rect 21760 83982 21836 84190
rect 21760 83950 21766 83982
rect 21765 83918 21766 83950
rect 21830 83950 21836 83982
rect 22576 84254 22652 84260
rect 22576 84190 22582 84254
rect 22646 84190 22652 84254
rect 22576 83982 22652 84190
rect 28424 84118 28500 84326
rect 28424 84054 28430 84118
rect 28494 84054 28500 84118
rect 110160 84326 110166 84390
rect 110230 84326 110236 84390
rect 110160 84118 110236 84326
rect 116960 84390 117036 84598
rect 116960 84326 116966 84390
rect 117030 84326 117036 84390
rect 116960 84320 117036 84326
rect 137496 84526 137844 85958
rect 137496 84462 137502 84526
rect 137566 84462 137844 84526
rect 116829 84254 116895 84255
rect 116829 84222 116830 84254
rect 110160 84086 110166 84118
rect 28424 84048 28500 84054
rect 110165 84054 110166 84086
rect 110230 84086 110236 84118
rect 116824 84190 116830 84222
rect 116894 84222 116895 84254
rect 116894 84190 116900 84222
rect 110230 84054 110231 84086
rect 110165 84053 110231 84054
rect 22576 83950 22582 83982
rect 21830 83918 21831 83950
rect 21765 83917 21831 83918
rect 22581 83918 22582 83950
rect 22646 83950 22652 83982
rect 28424 83982 28500 83988
rect 22646 83918 22647 83950
rect 22581 83917 22647 83918
rect 28424 83918 28430 83982
rect 28494 83918 28500 83982
rect 21901 83846 21967 83847
rect 21901 83814 21902 83846
rect 21896 83782 21902 83814
rect 21966 83814 21967 83846
rect 23120 83846 23196 83852
rect 21966 83782 21972 83814
rect 21896 83574 21972 83782
rect 21896 83510 21902 83574
rect 21966 83510 21972 83574
rect 23120 83782 23126 83846
rect 23190 83782 23196 83846
rect 23397 83846 23463 83847
rect 23397 83814 23398 83846
rect 23120 83574 23196 83782
rect 23120 83542 23126 83574
rect 21896 83504 21972 83510
rect 23125 83510 23126 83542
rect 23190 83542 23196 83574
rect 23392 83782 23398 83814
rect 23462 83814 23463 83846
rect 23462 83782 23468 83814
rect 23392 83574 23468 83782
rect 28424 83710 28500 83918
rect 116824 83982 116900 84190
rect 116824 83918 116830 83982
rect 116894 83918 116900 83982
rect 116824 83912 116900 83918
rect 115197 83846 115263 83847
rect 115197 83814 115198 83846
rect 28424 83678 28430 83710
rect 28429 83646 28430 83678
rect 28494 83678 28500 83710
rect 115192 83782 115198 83814
rect 115262 83814 115263 83846
rect 115605 83846 115671 83847
rect 115605 83814 115606 83846
rect 115262 83782 115268 83814
rect 28494 83646 28495 83678
rect 28429 83645 28495 83646
rect 23190 83510 23191 83542
rect 23125 83509 23191 83510
rect 23392 83510 23398 83574
rect 23462 83510 23468 83574
rect 23392 83504 23468 83510
rect 115192 83574 115268 83782
rect 115192 83510 115198 83574
rect 115262 83510 115268 83574
rect 115192 83504 115268 83510
rect 115600 83782 115606 83814
rect 115670 83814 115671 83846
rect 116960 83846 117036 83852
rect 115670 83782 115676 83814
rect 115600 83574 115676 83782
rect 115600 83510 115606 83574
rect 115670 83510 115676 83574
rect 116960 83782 116966 83846
rect 117030 83782 117036 83846
rect 116960 83574 117036 83782
rect 116960 83542 116966 83574
rect 115600 83504 115676 83510
rect 116965 83510 116966 83542
rect 117030 83542 117036 83574
rect 117030 83510 117031 83542
rect 116965 83509 117031 83510
rect 21760 83438 21836 83444
rect 21760 83374 21766 83438
rect 21830 83374 21836 83438
rect 22309 83438 22375 83439
rect 22309 83406 22310 83438
rect 21760 83166 21836 83374
rect 21760 83134 21766 83166
rect 21765 83102 21766 83134
rect 21830 83134 21836 83166
rect 22304 83374 22310 83406
rect 22374 83406 22375 83438
rect 22984 83438 23060 83444
rect 22374 83374 22380 83406
rect 22304 83166 22380 83374
rect 21830 83102 21831 83134
rect 21765 83101 21831 83102
rect 22304 83102 22310 83166
rect 22374 83102 22380 83166
rect 22984 83374 22990 83438
rect 23054 83374 23060 83438
rect 23397 83438 23463 83439
rect 23397 83406 23398 83438
rect 22984 83166 23060 83374
rect 22984 83134 22990 83166
rect 22304 83096 22380 83102
rect 22989 83102 22990 83134
rect 23054 83134 23060 83166
rect 23392 83374 23398 83406
rect 23462 83406 23463 83438
rect 115197 83438 115263 83439
rect 115197 83406 115198 83438
rect 23462 83374 23468 83406
rect 23392 83166 23468 83374
rect 23054 83102 23055 83134
rect 22989 83101 23055 83102
rect 23392 83102 23398 83166
rect 23462 83102 23468 83166
rect 23392 83096 23468 83102
rect 115192 83374 115198 83406
rect 115262 83406 115263 83438
rect 115736 83438 115812 83444
rect 115262 83374 115268 83406
rect 115192 83166 115268 83374
rect 115192 83102 115198 83166
rect 115262 83102 115268 83166
rect 115736 83374 115742 83438
rect 115806 83374 115812 83438
rect 115736 83166 115812 83374
rect 115736 83134 115742 83166
rect 115192 83096 115268 83102
rect 115741 83102 115742 83134
rect 115806 83134 115812 83166
rect 116008 83438 116084 83444
rect 116008 83374 116014 83438
rect 116078 83374 116084 83438
rect 116008 83166 116084 83374
rect 116008 83134 116014 83166
rect 115806 83102 115807 83134
rect 115741 83101 115807 83102
rect 116013 83102 116014 83134
rect 116078 83134 116084 83166
rect 116416 83438 116492 83444
rect 116416 83374 116422 83438
rect 116486 83374 116492 83438
rect 116965 83438 117031 83439
rect 116965 83406 116966 83438
rect 116416 83166 116492 83374
rect 116416 83134 116422 83166
rect 116078 83102 116079 83134
rect 116013 83101 116079 83102
rect 116421 83102 116422 83134
rect 116486 83134 116492 83166
rect 116960 83374 116966 83406
rect 117030 83406 117031 83438
rect 117030 83374 117036 83406
rect 116960 83166 117036 83374
rect 116486 83102 116487 83134
rect 116421 83101 116487 83102
rect 116960 83102 116966 83166
rect 117030 83102 117036 83166
rect 116960 83096 117036 83102
rect 21765 83030 21831 83031
rect 21765 82998 21766 83030
rect 952 82694 1230 82758
rect 1294 82694 1300 82758
rect 952 81126 1300 82694
rect 21760 82966 21766 82998
rect 21830 82998 21831 83030
rect 22173 83030 22239 83031
rect 22173 82998 22174 83030
rect 21830 82966 21836 82998
rect 21760 82758 21836 82966
rect 21760 82694 21766 82758
rect 21830 82694 21836 82758
rect 21760 82688 21836 82694
rect 22168 82966 22174 82998
rect 22238 82998 22239 83030
rect 22581 83030 22647 83031
rect 22581 82998 22582 83030
rect 22238 82966 22244 82998
rect 22168 82758 22244 82966
rect 22168 82694 22174 82758
rect 22238 82694 22244 82758
rect 22168 82688 22244 82694
rect 22576 82966 22582 82998
rect 22646 82998 22647 83030
rect 22984 83030 23060 83036
rect 22646 82966 22652 82998
rect 22576 82758 22652 82966
rect 22576 82694 22582 82758
rect 22646 82694 22652 82758
rect 22984 82966 22990 83030
rect 23054 82966 23060 83030
rect 22984 82758 23060 82966
rect 22984 82726 22990 82758
rect 22576 82688 22652 82694
rect 22989 82694 22990 82726
rect 23054 82726 23060 82758
rect 23392 83030 23468 83036
rect 23392 82966 23398 83030
rect 23462 82966 23468 83030
rect 23392 82758 23468 82966
rect 23392 82726 23398 82758
rect 23054 82694 23055 82726
rect 22989 82693 23055 82694
rect 23397 82694 23398 82726
rect 23462 82726 23468 82758
rect 115192 83030 115268 83036
rect 115192 82966 115198 83030
rect 115262 82966 115268 83030
rect 115741 83030 115807 83031
rect 115741 82998 115742 83030
rect 115192 82758 115268 82966
rect 115192 82726 115198 82758
rect 23462 82694 23463 82726
rect 23397 82693 23463 82694
rect 115197 82694 115198 82726
rect 115262 82726 115268 82758
rect 115736 82966 115742 82998
rect 115806 82998 115807 83030
rect 116008 83030 116084 83036
rect 115806 82966 115812 82998
rect 115736 82758 115812 82966
rect 115262 82694 115263 82726
rect 115197 82693 115263 82694
rect 115736 82694 115742 82758
rect 115806 82694 115812 82758
rect 116008 82966 116014 83030
rect 116078 82966 116084 83030
rect 116829 83030 116895 83031
rect 116829 82998 116830 83030
rect 116008 82758 116084 82966
rect 116008 82726 116014 82758
rect 115736 82688 115812 82694
rect 116013 82694 116014 82726
rect 116078 82726 116084 82758
rect 116824 82966 116830 82998
rect 116894 82998 116895 83030
rect 116894 82966 116900 82998
rect 116824 82758 116900 82966
rect 116078 82694 116079 82726
rect 116013 82693 116079 82694
rect 116824 82694 116830 82758
rect 116894 82694 116900 82758
rect 116824 82688 116900 82694
rect 137496 82758 137844 84462
rect 137496 82694 137502 82758
rect 137566 82694 137844 82758
rect 21896 82622 21972 82628
rect 21896 82558 21902 82622
rect 21966 82558 21972 82622
rect 21896 82350 21972 82558
rect 21896 82318 21902 82350
rect 21901 82286 21902 82318
rect 21966 82318 21972 82350
rect 22440 82622 22516 82628
rect 22440 82558 22446 82622
rect 22510 82558 22516 82622
rect 22440 82350 22516 82558
rect 22440 82318 22446 82350
rect 21966 82286 21967 82318
rect 21901 82285 21967 82286
rect 22445 82286 22446 82318
rect 22510 82318 22516 82350
rect 23120 82622 23196 82628
rect 23120 82558 23126 82622
rect 23190 82558 23196 82622
rect 23397 82622 23463 82623
rect 23397 82590 23398 82622
rect 23120 82350 23196 82558
rect 23120 82318 23126 82350
rect 22510 82286 22511 82318
rect 22445 82285 22511 82286
rect 23125 82286 23126 82318
rect 23190 82318 23196 82350
rect 23392 82558 23398 82590
rect 23462 82590 23463 82622
rect 115197 82622 115263 82623
rect 115197 82590 115198 82622
rect 23462 82558 23468 82590
rect 23392 82350 23468 82558
rect 23190 82286 23191 82318
rect 23125 82285 23191 82286
rect 23392 82286 23398 82350
rect 23462 82286 23468 82350
rect 23392 82280 23468 82286
rect 115192 82558 115198 82590
rect 115262 82590 115263 82622
rect 115600 82622 115676 82628
rect 115262 82558 115268 82590
rect 115192 82350 115268 82558
rect 115192 82286 115198 82350
rect 115262 82286 115268 82350
rect 115600 82558 115606 82622
rect 115670 82558 115676 82622
rect 116013 82622 116079 82623
rect 116013 82590 116014 82622
rect 115600 82350 115676 82558
rect 115600 82318 115606 82350
rect 115192 82280 115268 82286
rect 115605 82286 115606 82318
rect 115670 82318 115676 82350
rect 116008 82558 116014 82590
rect 116078 82590 116079 82622
rect 116965 82622 117031 82623
rect 116965 82590 116966 82622
rect 116078 82558 116084 82590
rect 116008 82350 116084 82558
rect 115670 82286 115671 82318
rect 115605 82285 115671 82286
rect 116008 82286 116014 82350
rect 116078 82286 116084 82350
rect 116008 82280 116084 82286
rect 116960 82558 116966 82590
rect 117030 82590 117031 82622
rect 117030 82558 117036 82590
rect 116960 82350 117036 82558
rect 116960 82286 116966 82350
rect 117030 82286 117036 82350
rect 116960 82280 117036 82286
rect 21765 82214 21831 82215
rect 21765 82182 21766 82214
rect 21760 82150 21766 82182
rect 21830 82182 21831 82214
rect 22576 82214 22652 82220
rect 21830 82150 21836 82182
rect 21760 81942 21836 82150
rect 21760 81878 21766 81942
rect 21830 81878 21836 81942
rect 22576 82150 22582 82214
rect 22646 82150 22652 82214
rect 22576 81942 22652 82150
rect 22576 81910 22582 81942
rect 21760 81872 21836 81878
rect 22581 81878 22582 81910
rect 22646 81910 22652 81942
rect 23120 82214 23196 82220
rect 23120 82150 23126 82214
rect 23190 82150 23196 82214
rect 23120 81942 23196 82150
rect 23120 81910 23126 81942
rect 22646 81878 22647 81910
rect 22581 81877 22647 81878
rect 23125 81878 23126 81910
rect 23190 81910 23196 81942
rect 23528 82214 23604 82220
rect 23528 82150 23534 82214
rect 23598 82150 23604 82214
rect 23528 81942 23604 82150
rect 23528 81910 23534 81942
rect 23190 81878 23191 81910
rect 23125 81877 23191 81878
rect 23533 81878 23534 81910
rect 23598 81910 23604 81942
rect 115328 82214 115404 82220
rect 115328 82150 115334 82214
rect 115398 82150 115404 82214
rect 115741 82214 115807 82215
rect 115741 82182 115742 82214
rect 115328 81942 115404 82150
rect 115328 81910 115334 81942
rect 23598 81878 23599 81910
rect 23533 81877 23599 81878
rect 115333 81878 115334 81910
rect 115398 81910 115404 81942
rect 115736 82150 115742 82182
rect 115806 82182 115807 82214
rect 116013 82214 116079 82215
rect 116013 82182 116014 82214
rect 115806 82150 115812 82182
rect 115736 81942 115812 82150
rect 115398 81878 115399 81910
rect 115333 81877 115399 81878
rect 115736 81878 115742 81942
rect 115806 81878 115812 81942
rect 115736 81872 115812 81878
rect 116008 82150 116014 82182
rect 116078 82182 116079 82214
rect 116421 82214 116487 82215
rect 116421 82182 116422 82214
rect 116078 82150 116084 82182
rect 116008 81942 116084 82150
rect 116008 81878 116014 81942
rect 116078 81878 116084 81942
rect 116008 81872 116084 81878
rect 116416 82150 116422 82182
rect 116486 82182 116487 82214
rect 116829 82214 116895 82215
rect 116829 82182 116830 82214
rect 116486 82150 116492 82182
rect 116416 81942 116492 82150
rect 116416 81878 116422 81942
rect 116486 81878 116492 81942
rect 116416 81872 116492 81878
rect 116824 82150 116830 82182
rect 116894 82182 116895 82214
rect 116894 82150 116900 82182
rect 116824 81942 116900 82150
rect 116824 81878 116830 81942
rect 116894 81878 116900 81942
rect 116824 81872 116900 81878
rect 22304 81806 22380 81812
rect 22304 81742 22310 81806
rect 22374 81742 22380 81806
rect 22581 81806 22647 81807
rect 22581 81774 22582 81806
rect 22304 81534 22380 81742
rect 22304 81502 22310 81534
rect 22309 81470 22310 81502
rect 22374 81502 22380 81534
rect 22576 81742 22582 81774
rect 22646 81774 22647 81806
rect 23125 81806 23191 81807
rect 23125 81774 23126 81806
rect 22646 81742 22652 81774
rect 22576 81534 22652 81742
rect 22374 81470 22375 81502
rect 22309 81469 22375 81470
rect 22576 81470 22582 81534
rect 22646 81470 22652 81534
rect 22576 81464 22652 81470
rect 23120 81742 23126 81774
rect 23190 81774 23191 81806
rect 23533 81806 23599 81807
rect 23533 81774 23534 81806
rect 23190 81742 23196 81774
rect 23120 81534 23196 81742
rect 23120 81470 23126 81534
rect 23190 81470 23196 81534
rect 23120 81464 23196 81470
rect 23528 81742 23534 81774
rect 23598 81774 23599 81806
rect 115192 81806 115268 81812
rect 23598 81742 23604 81774
rect 23528 81534 23604 81742
rect 23528 81470 23534 81534
rect 23598 81470 23604 81534
rect 115192 81742 115198 81806
rect 115262 81742 115268 81806
rect 115192 81534 115268 81742
rect 115192 81502 115198 81534
rect 23528 81464 23604 81470
rect 115197 81470 115198 81502
rect 115262 81502 115268 81534
rect 115600 81806 115676 81812
rect 115600 81742 115606 81806
rect 115670 81742 115676 81806
rect 116285 81806 116351 81807
rect 116285 81774 116286 81806
rect 115600 81534 115676 81742
rect 115600 81502 115606 81534
rect 115262 81470 115263 81502
rect 115197 81469 115263 81470
rect 115605 81470 115606 81502
rect 115670 81502 115676 81534
rect 116280 81742 116286 81774
rect 116350 81774 116351 81806
rect 116350 81742 116356 81774
rect 116280 81534 116356 81742
rect 115670 81470 115671 81502
rect 115605 81469 115671 81470
rect 116280 81470 116286 81534
rect 116350 81470 116356 81534
rect 116280 81464 116356 81470
rect 952 81062 1230 81126
rect 1294 81062 1300 81126
rect 22984 81398 23060 81404
rect 22984 81334 22990 81398
rect 23054 81334 23060 81398
rect 22984 81126 23060 81334
rect 22984 81094 22990 81126
rect 952 79494 1300 81062
rect 22989 81062 22990 81094
rect 23054 81094 23060 81126
rect 23528 81398 23604 81404
rect 23528 81334 23534 81398
rect 23598 81334 23604 81398
rect 115197 81398 115263 81399
rect 115197 81366 115198 81398
rect 23528 81126 23604 81334
rect 115192 81334 115198 81366
rect 115262 81366 115263 81398
rect 115605 81398 115671 81399
rect 115605 81366 115606 81398
rect 115262 81334 115268 81366
rect 23528 81094 23534 81126
rect 23054 81062 23055 81094
rect 22989 81061 23055 81062
rect 23533 81062 23534 81094
rect 23598 81094 23604 81126
rect 28288 81126 28364 81132
rect 23598 81062 23599 81094
rect 23533 81061 23599 81062
rect 28288 81062 28294 81126
rect 28358 81062 28364 81126
rect 22168 80990 22244 80996
rect 22168 80926 22174 80990
rect 22238 80926 22244 80990
rect 21896 80718 21972 80724
rect 21896 80654 21902 80718
rect 21966 80654 21972 80718
rect 22168 80718 22244 80926
rect 28288 80854 28364 81062
rect 115192 81126 115268 81334
rect 115192 81062 115198 81126
rect 115262 81062 115268 81126
rect 115192 81056 115268 81062
rect 115600 81334 115606 81366
rect 115670 81366 115671 81398
rect 115670 81334 115676 81366
rect 115600 81126 115676 81334
rect 115600 81062 115606 81126
rect 115670 81062 115676 81126
rect 115600 81056 115676 81062
rect 137496 81126 137844 82694
rect 137496 81062 137502 81126
rect 137566 81062 137844 81126
rect 116144 80990 116220 80996
rect 116144 80926 116150 80990
rect 116214 80926 116220 80990
rect 28288 80822 28294 80854
rect 28293 80790 28294 80822
rect 28358 80822 28364 80854
rect 28565 80854 28631 80855
rect 28565 80822 28566 80854
rect 28358 80790 28359 80822
rect 28293 80789 28359 80790
rect 28560 80790 28566 80822
rect 28630 80822 28631 80854
rect 28630 80790 28636 80822
rect 22168 80686 22174 80718
rect 21896 80446 21972 80654
rect 22173 80654 22174 80686
rect 22238 80686 22244 80718
rect 22238 80654 22239 80686
rect 22173 80653 22239 80654
rect 21896 80414 21902 80446
rect 21901 80382 21902 80414
rect 21966 80414 21972 80446
rect 22440 80582 22516 80588
rect 22440 80518 22446 80582
rect 22510 80518 22516 80582
rect 21966 80382 21967 80414
rect 21901 80381 21967 80382
rect 21901 80310 21967 80311
rect 21901 80278 21902 80310
rect 21896 80246 21902 80278
rect 21966 80278 21967 80310
rect 22440 80310 22516 80518
rect 28560 80582 28636 80790
rect 116144 80718 116220 80926
rect 116144 80686 116150 80718
rect 116149 80654 116150 80686
rect 116214 80686 116220 80718
rect 116829 80718 116895 80719
rect 116829 80686 116830 80718
rect 116214 80654 116215 80686
rect 116149 80653 116215 80654
rect 116824 80654 116830 80686
rect 116894 80686 116895 80718
rect 116894 80654 116900 80686
rect 28560 80518 28566 80582
rect 28630 80518 28636 80582
rect 28560 80512 28636 80518
rect 28288 80446 28364 80452
rect 28288 80382 28294 80446
rect 28358 80382 28364 80446
rect 22440 80278 22446 80310
rect 21966 80246 21972 80278
rect 21896 80038 21972 80246
rect 22445 80246 22446 80278
rect 22510 80278 22516 80310
rect 22717 80310 22783 80311
rect 22717 80278 22718 80310
rect 22510 80246 22511 80278
rect 22445 80245 22511 80246
rect 22712 80246 22718 80278
rect 22782 80278 22783 80310
rect 22782 80246 22788 80278
rect 21896 79974 21902 80038
rect 21966 79974 21972 80038
rect 21896 79968 21972 79974
rect 22712 80038 22788 80246
rect 28288 80174 28364 80382
rect 28288 80142 28294 80174
rect 28293 80110 28294 80142
rect 28358 80142 28364 80174
rect 110432 80446 110508 80452
rect 110432 80382 110438 80446
rect 110502 80382 110508 80446
rect 110432 80174 110508 80382
rect 116824 80446 116900 80654
rect 116824 80382 116830 80446
rect 116894 80382 116900 80446
rect 116824 80376 116900 80382
rect 116013 80310 116079 80311
rect 116013 80278 116014 80310
rect 110432 80142 110438 80174
rect 28358 80110 28359 80142
rect 28293 80109 28359 80110
rect 110437 80110 110438 80142
rect 110502 80142 110508 80174
rect 116008 80246 116014 80278
rect 116078 80278 116079 80310
rect 116285 80310 116351 80311
rect 116285 80278 116286 80310
rect 116078 80246 116084 80278
rect 110502 80110 110503 80142
rect 110437 80109 110503 80110
rect 22712 79974 22718 80038
rect 22782 79974 22788 80038
rect 22712 79968 22788 79974
rect 110160 80038 110236 80044
rect 110160 79974 110166 80038
rect 110230 79974 110236 80038
rect 21760 79902 21836 79908
rect 21760 79838 21766 79902
rect 21830 79838 21836 79902
rect 22989 79902 23055 79903
rect 22989 79870 22990 79902
rect 21760 79630 21836 79838
rect 21760 79598 21766 79630
rect 21765 79566 21766 79598
rect 21830 79598 21836 79630
rect 22984 79838 22990 79870
rect 23054 79870 23055 79902
rect 23528 79902 23604 79908
rect 23054 79838 23060 79870
rect 22984 79630 23060 79838
rect 21830 79566 21831 79598
rect 21765 79565 21831 79566
rect 22984 79566 22990 79630
rect 23054 79566 23060 79630
rect 23528 79838 23534 79902
rect 23598 79838 23604 79902
rect 23528 79630 23604 79838
rect 110160 79766 110236 79974
rect 116008 80038 116084 80246
rect 116008 79974 116014 80038
rect 116078 79974 116084 80038
rect 116008 79968 116084 79974
rect 116280 80246 116286 80278
rect 116350 80278 116351 80310
rect 116824 80310 116900 80316
rect 116350 80246 116356 80278
rect 116280 80038 116356 80246
rect 116280 79974 116286 80038
rect 116350 79974 116356 80038
rect 116824 80246 116830 80310
rect 116894 80246 116900 80310
rect 116824 80038 116900 80246
rect 116824 80006 116830 80038
rect 116280 79968 116356 79974
rect 116829 79974 116830 80006
rect 116894 80006 116900 80038
rect 116894 79974 116895 80006
rect 116829 79973 116895 79974
rect 115333 79902 115399 79903
rect 115333 79870 115334 79902
rect 110160 79734 110166 79766
rect 110165 79702 110166 79734
rect 110230 79734 110236 79766
rect 115328 79838 115334 79870
rect 115398 79870 115399 79902
rect 115741 79902 115807 79903
rect 115741 79870 115742 79902
rect 115398 79838 115404 79870
rect 110230 79702 110231 79734
rect 110165 79701 110231 79702
rect 23528 79598 23534 79630
rect 22984 79560 23060 79566
rect 23533 79566 23534 79598
rect 23598 79598 23604 79630
rect 115328 79630 115404 79838
rect 23598 79566 23599 79598
rect 23533 79565 23599 79566
rect 115328 79566 115334 79630
rect 115398 79566 115404 79630
rect 115328 79560 115404 79566
rect 115736 79838 115742 79870
rect 115806 79870 115807 79902
rect 116824 79902 116900 79908
rect 115806 79838 115812 79870
rect 115736 79630 115812 79838
rect 116824 79838 116830 79902
rect 116894 79838 116900 79902
rect 115736 79566 115742 79630
rect 115806 79566 115812 79630
rect 115736 79560 115812 79566
rect 116280 79766 116356 79772
rect 116280 79702 116286 79766
rect 116350 79702 116356 79766
rect 952 79430 1230 79494
rect 1294 79430 1300 79494
rect 21901 79494 21967 79495
rect 21901 79462 21902 79494
rect 952 77726 1300 79430
rect 21896 79430 21902 79462
rect 21966 79462 21967 79494
rect 22712 79494 22788 79500
rect 21966 79430 21972 79462
rect 21896 79222 21972 79430
rect 21896 79158 21902 79222
rect 21966 79158 21972 79222
rect 22712 79430 22718 79494
rect 22782 79430 22788 79494
rect 22712 79222 22788 79430
rect 22712 79190 22718 79222
rect 21896 79152 21972 79158
rect 22717 79158 22718 79190
rect 22782 79190 22788 79222
rect 23120 79494 23196 79500
rect 23120 79430 23126 79494
rect 23190 79430 23196 79494
rect 23120 79222 23196 79430
rect 23120 79190 23126 79222
rect 22782 79158 22783 79190
rect 22717 79157 22783 79158
rect 23125 79158 23126 79190
rect 23190 79190 23196 79222
rect 23392 79494 23468 79500
rect 23392 79430 23398 79494
rect 23462 79430 23468 79494
rect 23392 79222 23468 79430
rect 115192 79494 115268 79500
rect 115192 79430 115198 79494
rect 115262 79430 115268 79494
rect 23392 79190 23398 79222
rect 23190 79158 23191 79190
rect 23125 79157 23191 79158
rect 23397 79158 23398 79190
rect 23462 79190 23468 79222
rect 28288 79222 28364 79228
rect 23462 79158 23463 79190
rect 23397 79157 23463 79158
rect 28288 79158 28294 79222
rect 28358 79158 28364 79222
rect 115192 79222 115268 79430
rect 115192 79190 115198 79222
rect 21760 79086 21836 79092
rect 21760 79022 21766 79086
rect 21830 79022 21836 79086
rect 23125 79086 23191 79087
rect 23125 79054 23126 79086
rect 21760 78814 21836 79022
rect 21760 78782 21766 78814
rect 21765 78750 21766 78782
rect 21830 78782 21836 78814
rect 23120 79022 23126 79054
rect 23190 79054 23191 79086
rect 23397 79086 23463 79087
rect 23397 79054 23398 79086
rect 23190 79022 23196 79054
rect 23120 78814 23196 79022
rect 21830 78750 21831 78782
rect 21765 78749 21831 78750
rect 23120 78750 23126 78814
rect 23190 78750 23196 78814
rect 23120 78744 23196 78750
rect 23392 79022 23398 79054
rect 23462 79054 23463 79086
rect 23462 79022 23468 79054
rect 23392 78814 23468 79022
rect 28288 78950 28364 79158
rect 115197 79158 115198 79190
rect 115262 79190 115268 79222
rect 115600 79494 115676 79500
rect 115600 79430 115606 79494
rect 115670 79430 115676 79494
rect 116280 79494 116356 79702
rect 116824 79630 116900 79838
rect 116824 79598 116830 79630
rect 116829 79566 116830 79598
rect 116894 79598 116900 79630
rect 116894 79566 116895 79598
rect 116829 79565 116895 79566
rect 116280 79462 116286 79494
rect 115600 79222 115676 79430
rect 116285 79430 116286 79462
rect 116350 79462 116356 79494
rect 116552 79494 116628 79500
rect 116350 79430 116351 79462
rect 116285 79429 116351 79430
rect 116552 79430 116558 79494
rect 116622 79430 116628 79494
rect 116965 79494 117031 79495
rect 116965 79462 116966 79494
rect 115600 79190 115606 79222
rect 115262 79158 115263 79190
rect 115197 79157 115263 79158
rect 115605 79158 115606 79190
rect 115670 79190 115676 79222
rect 116552 79222 116628 79430
rect 116552 79190 116558 79222
rect 115670 79158 115671 79190
rect 115605 79157 115671 79158
rect 116557 79158 116558 79190
rect 116622 79190 116628 79222
rect 116960 79430 116966 79462
rect 117030 79462 117031 79494
rect 137496 79494 137844 81062
rect 117030 79430 117036 79462
rect 116960 79222 117036 79430
rect 116622 79158 116623 79190
rect 116557 79157 116623 79158
rect 116960 79158 116966 79222
rect 117030 79158 117036 79222
rect 116960 79152 117036 79158
rect 137496 79430 137502 79494
rect 137566 79430 137844 79494
rect 115197 79086 115263 79087
rect 115197 79054 115198 79086
rect 28288 78918 28294 78950
rect 28293 78886 28294 78918
rect 28358 78918 28364 78950
rect 115192 79022 115198 79054
rect 115262 79054 115263 79086
rect 115736 79086 115812 79092
rect 115262 79022 115268 79054
rect 28358 78886 28359 78918
rect 28293 78885 28359 78886
rect 23392 78750 23398 78814
rect 23462 78750 23468 78814
rect 23392 78744 23468 78750
rect 115192 78814 115268 79022
rect 115192 78750 115198 78814
rect 115262 78750 115268 78814
rect 115736 79022 115742 79086
rect 115806 79022 115812 79086
rect 115736 78814 115812 79022
rect 115736 78782 115742 78814
rect 115192 78744 115268 78750
rect 115741 78750 115742 78782
rect 115806 78782 115812 78814
rect 116008 79086 116084 79092
rect 116008 79022 116014 79086
rect 116078 79022 116084 79086
rect 116965 79086 117031 79087
rect 116965 79054 116966 79086
rect 116008 78814 116084 79022
rect 116008 78782 116014 78814
rect 115806 78750 115807 78782
rect 115741 78749 115807 78750
rect 116013 78750 116014 78782
rect 116078 78782 116084 78814
rect 116960 79022 116966 79054
rect 117030 79054 117031 79086
rect 117030 79022 117036 79054
rect 116960 78814 117036 79022
rect 116078 78750 116079 78782
rect 116013 78749 116079 78750
rect 116960 78750 116966 78814
rect 117030 78750 117036 78814
rect 116960 78744 117036 78750
rect 21896 78678 21972 78684
rect 21896 78614 21902 78678
rect 21966 78614 21972 78678
rect 21896 78406 21972 78614
rect 21896 78374 21902 78406
rect 21901 78342 21902 78374
rect 21966 78374 21972 78406
rect 22304 78678 22380 78684
rect 22304 78614 22310 78678
rect 22374 78614 22380 78678
rect 22581 78678 22647 78679
rect 22581 78646 22582 78678
rect 22304 78406 22380 78614
rect 22304 78374 22310 78406
rect 21966 78342 21967 78374
rect 21901 78341 21967 78342
rect 22309 78342 22310 78374
rect 22374 78374 22380 78406
rect 22576 78614 22582 78646
rect 22646 78646 22647 78678
rect 22984 78678 23060 78684
rect 22646 78614 22652 78646
rect 22576 78406 22652 78614
rect 22374 78342 22375 78374
rect 22309 78341 22375 78342
rect 22576 78342 22582 78406
rect 22646 78342 22652 78406
rect 22984 78614 22990 78678
rect 23054 78614 23060 78678
rect 22984 78406 23060 78614
rect 22984 78374 22990 78406
rect 22576 78336 22652 78342
rect 22989 78342 22990 78374
rect 23054 78374 23060 78406
rect 23392 78678 23468 78684
rect 23392 78614 23398 78678
rect 23462 78614 23468 78678
rect 115333 78678 115399 78679
rect 115333 78646 115334 78678
rect 23392 78406 23468 78614
rect 23392 78374 23398 78406
rect 23054 78342 23055 78374
rect 22989 78341 23055 78342
rect 23397 78342 23398 78374
rect 23462 78374 23468 78406
rect 115328 78614 115334 78646
rect 115398 78646 115399 78678
rect 115741 78678 115807 78679
rect 115741 78646 115742 78678
rect 115398 78614 115404 78646
rect 115328 78406 115404 78614
rect 23462 78342 23463 78374
rect 23397 78341 23463 78342
rect 115328 78342 115334 78406
rect 115398 78342 115404 78406
rect 115328 78336 115404 78342
rect 115736 78614 115742 78646
rect 115806 78646 115807 78678
rect 116008 78678 116084 78684
rect 115806 78614 115812 78646
rect 115736 78406 115812 78614
rect 115736 78342 115742 78406
rect 115806 78342 115812 78406
rect 116008 78614 116014 78678
rect 116078 78614 116084 78678
rect 116008 78406 116084 78614
rect 116008 78374 116014 78406
rect 115736 78336 115812 78342
rect 116013 78342 116014 78374
rect 116078 78374 116084 78406
rect 116960 78678 117036 78684
rect 116960 78614 116966 78678
rect 117030 78614 117036 78678
rect 116960 78406 117036 78614
rect 116960 78374 116966 78406
rect 116078 78342 116079 78374
rect 116013 78341 116079 78342
rect 116965 78342 116966 78374
rect 117030 78374 117036 78406
rect 117030 78342 117031 78374
rect 116965 78341 117031 78342
rect 21901 78270 21967 78271
rect 21901 78238 21902 78270
rect 21896 78206 21902 78238
rect 21966 78238 21967 78270
rect 22309 78270 22375 78271
rect 22309 78238 22310 78270
rect 21966 78206 21972 78238
rect 21896 77998 21972 78206
rect 21896 77934 21902 77998
rect 21966 77934 21972 77998
rect 21896 77928 21972 77934
rect 22304 78206 22310 78238
rect 22374 78238 22375 78270
rect 22989 78270 23055 78271
rect 22989 78238 22990 78270
rect 22374 78206 22380 78238
rect 22304 77998 22380 78206
rect 22304 77934 22310 77998
rect 22374 77934 22380 77998
rect 22304 77928 22380 77934
rect 22984 78206 22990 78238
rect 23054 78238 23055 78270
rect 23397 78270 23463 78271
rect 23397 78238 23398 78270
rect 23054 78206 23060 78238
rect 22984 77998 23060 78206
rect 22984 77934 22990 77998
rect 23054 77934 23060 77998
rect 22984 77928 23060 77934
rect 23392 78206 23398 78238
rect 23462 78238 23463 78270
rect 115328 78270 115404 78276
rect 23462 78206 23468 78238
rect 23392 77998 23468 78206
rect 23392 77934 23398 77998
rect 23462 77934 23468 77998
rect 115328 78206 115334 78270
rect 115398 78206 115404 78270
rect 115328 77998 115404 78206
rect 115328 77966 115334 77998
rect 23392 77928 23468 77934
rect 115333 77934 115334 77966
rect 115398 77966 115404 77998
rect 115600 78270 115676 78276
rect 115600 78206 115606 78270
rect 115670 78206 115676 78270
rect 116013 78270 116079 78271
rect 116013 78238 116014 78270
rect 115600 77998 115676 78206
rect 115600 77966 115606 77998
rect 115398 77934 115399 77966
rect 115333 77933 115399 77934
rect 115605 77934 115606 77966
rect 115670 77966 115676 77998
rect 116008 78206 116014 78238
rect 116078 78238 116079 78270
rect 116960 78270 117036 78276
rect 116078 78206 116084 78238
rect 116008 77998 116084 78206
rect 115670 77934 115671 77966
rect 115605 77933 115671 77934
rect 116008 77934 116014 77998
rect 116078 77934 116084 77998
rect 116960 78206 116966 78270
rect 117030 78206 117036 78270
rect 116960 77998 117036 78206
rect 116960 77966 116966 77998
rect 116008 77928 116084 77934
rect 116965 77934 116966 77966
rect 117030 77966 117036 77998
rect 117030 77934 117031 77966
rect 116965 77933 117031 77934
rect 22445 77862 22511 77863
rect 22445 77830 22446 77862
rect 952 77662 1230 77726
rect 1294 77662 1300 77726
rect 952 75958 1300 77662
rect 22440 77798 22446 77830
rect 22510 77830 22511 77862
rect 23120 77862 23196 77868
rect 22510 77798 22516 77830
rect 22440 77590 22516 77798
rect 22440 77526 22446 77590
rect 22510 77526 22516 77590
rect 23120 77798 23126 77862
rect 23190 77798 23196 77862
rect 23120 77590 23196 77798
rect 23120 77558 23126 77590
rect 22440 77520 22516 77526
rect 23125 77526 23126 77558
rect 23190 77558 23196 77590
rect 23528 77862 23604 77868
rect 23528 77798 23534 77862
rect 23598 77798 23604 77862
rect 115333 77862 115399 77863
rect 115333 77830 115334 77862
rect 23528 77590 23604 77798
rect 115328 77798 115334 77830
rect 115398 77830 115399 77862
rect 115741 77862 115807 77863
rect 115741 77830 115742 77862
rect 115398 77798 115404 77830
rect 23528 77558 23534 77590
rect 23190 77526 23191 77558
rect 23125 77525 23191 77526
rect 23533 77526 23534 77558
rect 23598 77558 23604 77590
rect 28288 77726 28364 77732
rect 28288 77662 28294 77726
rect 28358 77662 28364 77726
rect 23598 77526 23599 77558
rect 23533 77525 23599 77526
rect 22984 77454 23060 77460
rect 22984 77390 22990 77454
rect 23054 77390 23060 77454
rect 22984 77182 23060 77390
rect 22984 77150 22990 77182
rect 22989 77118 22990 77150
rect 23054 77150 23060 77182
rect 23392 77454 23468 77460
rect 23392 77390 23398 77454
rect 23462 77390 23468 77454
rect 28288 77454 28364 77662
rect 28288 77422 28294 77454
rect 23392 77182 23468 77390
rect 28293 77390 28294 77422
rect 28358 77422 28364 77454
rect 110432 77726 110508 77732
rect 110432 77662 110438 77726
rect 110502 77662 110508 77726
rect 110432 77454 110508 77662
rect 115328 77590 115404 77798
rect 115328 77526 115334 77590
rect 115398 77526 115404 77590
rect 115328 77520 115404 77526
rect 115736 77798 115742 77830
rect 115806 77830 115807 77862
rect 116285 77862 116351 77863
rect 116285 77830 116286 77862
rect 115806 77798 115812 77830
rect 115736 77590 115812 77798
rect 115736 77526 115742 77590
rect 115806 77526 115812 77590
rect 115736 77520 115812 77526
rect 116280 77798 116286 77830
rect 116350 77830 116351 77862
rect 116350 77798 116356 77830
rect 116280 77590 116356 77798
rect 116280 77526 116286 77590
rect 116350 77526 116356 77590
rect 116280 77520 116356 77526
rect 137496 77590 137844 79430
rect 137496 77526 137502 77590
rect 137566 77526 137844 77590
rect 110432 77422 110438 77454
rect 28358 77390 28359 77422
rect 28293 77389 28359 77390
rect 110437 77390 110438 77422
rect 110502 77422 110508 77454
rect 115333 77454 115399 77455
rect 115333 77422 115334 77454
rect 110502 77390 110503 77422
rect 110437 77389 110503 77390
rect 115328 77390 115334 77422
rect 115398 77422 115399 77454
rect 115600 77454 115676 77460
rect 115398 77390 115404 77422
rect 23392 77150 23398 77182
rect 23054 77118 23055 77150
rect 22989 77117 23055 77118
rect 23397 77118 23398 77150
rect 23462 77150 23468 77182
rect 115328 77182 115404 77390
rect 23462 77118 23463 77150
rect 23397 77117 23463 77118
rect 115328 77118 115334 77182
rect 115398 77118 115404 77182
rect 115600 77390 115606 77454
rect 115670 77390 115676 77454
rect 115600 77182 115676 77390
rect 115600 77150 115606 77182
rect 115328 77112 115404 77118
rect 115605 77118 115606 77150
rect 115670 77150 115676 77182
rect 115670 77118 115671 77150
rect 115605 77117 115671 77118
rect 22576 77046 22652 77052
rect 22576 76982 22582 77046
rect 22646 76982 22652 77046
rect 21760 76774 21836 76780
rect 21760 76710 21766 76774
rect 21830 76710 21836 76774
rect 22576 76774 22652 76982
rect 22576 76742 22582 76774
rect 21760 76502 21836 76710
rect 22581 76710 22582 76742
rect 22646 76742 22652 76774
rect 22984 77046 23060 77052
rect 22984 76982 22990 77046
rect 23054 76982 23060 77046
rect 22984 76774 23060 76982
rect 22984 76742 22990 76774
rect 22646 76710 22647 76742
rect 22581 76709 22647 76710
rect 22989 76710 22990 76742
rect 23054 76742 23060 76774
rect 23528 77046 23604 77052
rect 23528 76982 23534 77046
rect 23598 76982 23604 77046
rect 23528 76774 23604 76982
rect 115328 77046 115404 77052
rect 115328 76982 115334 77046
rect 115398 76982 115404 77046
rect 23528 76742 23534 76774
rect 23054 76710 23055 76742
rect 22989 76709 23055 76710
rect 23533 76710 23534 76742
rect 23598 76742 23604 76774
rect 110432 76910 110508 76916
rect 110432 76846 110438 76910
rect 110502 76846 110508 76910
rect 23598 76710 23599 76742
rect 23533 76709 23599 76710
rect 110432 76638 110508 76846
rect 115328 76774 115404 76982
rect 115328 76742 115334 76774
rect 115333 76710 115334 76742
rect 115398 76742 115404 76774
rect 115736 77046 115812 77052
rect 115736 76982 115742 77046
rect 115806 76982 115812 77046
rect 115736 76774 115812 76982
rect 115736 76742 115742 76774
rect 115398 76710 115399 76742
rect 115333 76709 115399 76710
rect 115741 76710 115742 76742
rect 115806 76742 115812 76774
rect 116008 77046 116084 77052
rect 116008 76982 116014 77046
rect 116078 76982 116084 77046
rect 116008 76774 116084 76982
rect 116008 76742 116014 76774
rect 115806 76710 115807 76742
rect 115741 76709 115807 76710
rect 116013 76710 116014 76742
rect 116078 76742 116084 76774
rect 116824 76774 116900 76780
rect 116078 76710 116079 76742
rect 116013 76709 116079 76710
rect 116824 76710 116830 76774
rect 116894 76710 116900 76774
rect 110432 76606 110438 76638
rect 110437 76574 110438 76606
rect 110502 76606 110508 76638
rect 110502 76574 110503 76606
rect 110437 76573 110503 76574
rect 21760 76470 21766 76502
rect 21765 76438 21766 76470
rect 21830 76470 21836 76502
rect 28288 76502 28364 76508
rect 21830 76438 21831 76470
rect 21765 76437 21831 76438
rect 28288 76438 28294 76502
rect 28358 76438 28364 76502
rect 110301 76502 110367 76503
rect 110301 76470 110302 76502
rect 21896 76366 21972 76372
rect 21896 76302 21902 76366
rect 21966 76302 21972 76366
rect 22581 76366 22647 76367
rect 22581 76334 22582 76366
rect 21896 76094 21972 76302
rect 21896 76062 21902 76094
rect 21901 76030 21902 76062
rect 21966 76062 21972 76094
rect 22576 76302 22582 76334
rect 22646 76334 22647 76366
rect 22646 76302 22652 76334
rect 22576 76094 22652 76302
rect 28288 76230 28364 76438
rect 28288 76198 28294 76230
rect 28293 76166 28294 76198
rect 28358 76198 28364 76230
rect 110296 76438 110302 76470
rect 110366 76470 110367 76502
rect 116824 76502 116900 76710
rect 116824 76470 116830 76502
rect 110366 76438 110372 76470
rect 110296 76230 110372 76438
rect 116829 76438 116830 76470
rect 116894 76470 116900 76502
rect 116894 76438 116895 76470
rect 116829 76437 116895 76438
rect 116149 76366 116215 76367
rect 116149 76334 116150 76366
rect 28358 76166 28359 76198
rect 28293 76165 28359 76166
rect 110296 76166 110302 76230
rect 110366 76166 110372 76230
rect 110296 76160 110372 76166
rect 116144 76302 116150 76334
rect 116214 76334 116215 76366
rect 116552 76366 116628 76372
rect 116214 76302 116220 76334
rect 21966 76030 21967 76062
rect 21901 76029 21967 76030
rect 22576 76030 22582 76094
rect 22646 76030 22652 76094
rect 28565 76094 28631 76095
rect 28565 76062 28566 76094
rect 22576 76024 22652 76030
rect 28560 76030 28566 76062
rect 28630 76062 28631 76094
rect 116144 76094 116220 76302
rect 28630 76030 28636 76062
rect 952 75894 1230 75958
rect 1294 75894 1300 75958
rect 952 74190 1300 75894
rect 21760 75958 21836 75964
rect 21760 75894 21766 75958
rect 21830 75894 21836 75958
rect 21760 75686 21836 75894
rect 28560 75822 28636 76030
rect 116144 76030 116150 76094
rect 116214 76030 116220 76094
rect 116552 76302 116558 76366
rect 116622 76302 116628 76366
rect 116552 76094 116628 76302
rect 116552 76062 116558 76094
rect 116144 76024 116220 76030
rect 116557 76030 116558 76062
rect 116622 76062 116628 76094
rect 116960 76366 117036 76372
rect 116960 76302 116966 76366
rect 117030 76302 117036 76366
rect 116960 76094 117036 76302
rect 116960 76062 116966 76094
rect 116622 76030 116623 76062
rect 116557 76029 116623 76030
rect 116965 76030 116966 76062
rect 117030 76062 117036 76094
rect 117030 76030 117031 76062
rect 116965 76029 117031 76030
rect 28560 75758 28566 75822
rect 28630 75758 28636 75822
rect 28560 75752 28636 75758
rect 116824 75958 116900 75964
rect 116824 75894 116830 75958
rect 116894 75894 116900 75958
rect 21760 75654 21766 75686
rect 21765 75622 21766 75654
rect 21830 75654 21836 75686
rect 116824 75686 116900 75894
rect 116824 75654 116830 75686
rect 21830 75622 21831 75654
rect 21765 75621 21831 75622
rect 116829 75622 116830 75654
rect 116894 75654 116900 75686
rect 137496 75958 137844 77526
rect 137496 75894 137502 75958
rect 137566 75894 137844 75958
rect 116894 75622 116895 75654
rect 116829 75621 116895 75622
rect 21765 75550 21831 75551
rect 21765 75518 21766 75550
rect 21760 75486 21766 75518
rect 21830 75518 21831 75550
rect 22440 75550 22516 75556
rect 21830 75486 21836 75518
rect 21760 75278 21836 75486
rect 21760 75214 21766 75278
rect 21830 75214 21836 75278
rect 22440 75486 22446 75550
rect 22510 75486 22516 75550
rect 22989 75550 23055 75551
rect 22989 75518 22990 75550
rect 22440 75278 22516 75486
rect 22440 75246 22446 75278
rect 21760 75208 21836 75214
rect 22445 75214 22446 75246
rect 22510 75246 22516 75278
rect 22984 75486 22990 75518
rect 23054 75518 23055 75550
rect 23528 75550 23604 75556
rect 23054 75486 23060 75518
rect 22984 75278 23060 75486
rect 22510 75214 22511 75246
rect 22445 75213 22511 75214
rect 22984 75214 22990 75278
rect 23054 75214 23060 75278
rect 23528 75486 23534 75550
rect 23598 75486 23604 75550
rect 115333 75550 115399 75551
rect 115333 75518 115334 75550
rect 23528 75278 23604 75486
rect 115328 75486 115334 75518
rect 115398 75518 115399 75550
rect 115741 75550 115807 75551
rect 115741 75518 115742 75550
rect 115398 75486 115404 75518
rect 23528 75246 23534 75278
rect 22984 75208 23060 75214
rect 23533 75214 23534 75246
rect 23598 75246 23604 75278
rect 28424 75278 28500 75284
rect 23598 75214 23599 75246
rect 23533 75213 23599 75214
rect 28424 75214 28430 75278
rect 28494 75214 28500 75278
rect 21901 75142 21967 75143
rect 21901 75110 21902 75142
rect 21896 75078 21902 75110
rect 21966 75110 21967 75142
rect 22712 75142 22788 75148
rect 21966 75078 21972 75110
rect 21896 74870 21972 75078
rect 21896 74806 21902 74870
rect 21966 74806 21972 74870
rect 22712 75078 22718 75142
rect 22782 75078 22788 75142
rect 22712 74870 22788 75078
rect 22712 74838 22718 74870
rect 21896 74800 21972 74806
rect 22717 74806 22718 74838
rect 22782 74838 22788 74870
rect 23120 75142 23196 75148
rect 23120 75078 23126 75142
rect 23190 75078 23196 75142
rect 23120 74870 23196 75078
rect 23120 74838 23126 74870
rect 22782 74806 22783 74838
rect 22717 74805 22783 74806
rect 23125 74806 23126 74838
rect 23190 74838 23196 74870
rect 23392 75142 23468 75148
rect 23392 75078 23398 75142
rect 23462 75078 23468 75142
rect 23392 74870 23468 75078
rect 28424 75006 28500 75214
rect 115328 75278 115404 75486
rect 115328 75214 115334 75278
rect 115398 75214 115404 75278
rect 115328 75208 115404 75214
rect 115736 75486 115742 75518
rect 115806 75518 115807 75550
rect 116144 75550 116220 75556
rect 115806 75486 115812 75518
rect 115736 75278 115812 75486
rect 115736 75214 115742 75278
rect 115806 75214 115812 75278
rect 116144 75486 116150 75550
rect 116214 75486 116220 75550
rect 116421 75550 116487 75551
rect 116421 75518 116422 75550
rect 116144 75278 116220 75486
rect 116144 75246 116150 75278
rect 115736 75208 115812 75214
rect 116149 75214 116150 75246
rect 116214 75246 116220 75278
rect 116416 75486 116422 75518
rect 116486 75518 116487 75550
rect 116829 75550 116895 75551
rect 116829 75518 116830 75550
rect 116486 75486 116492 75518
rect 116416 75278 116492 75486
rect 116214 75214 116215 75246
rect 116149 75213 116215 75214
rect 116416 75214 116422 75278
rect 116486 75214 116492 75278
rect 116416 75208 116492 75214
rect 116824 75486 116830 75518
rect 116894 75518 116895 75550
rect 116894 75486 116900 75518
rect 116824 75278 116900 75486
rect 116824 75214 116830 75278
rect 116894 75214 116900 75278
rect 116824 75208 116900 75214
rect 28424 74974 28430 75006
rect 28429 74942 28430 74974
rect 28494 74974 28500 75006
rect 115192 75142 115268 75148
rect 115192 75078 115198 75142
rect 115262 75078 115268 75142
rect 28494 74942 28495 74974
rect 28429 74941 28495 74942
rect 23392 74838 23398 74870
rect 23190 74806 23191 74838
rect 23125 74805 23191 74806
rect 23397 74806 23398 74838
rect 23462 74838 23468 74870
rect 115192 74870 115268 75078
rect 115192 74838 115198 74870
rect 23462 74806 23463 74838
rect 23397 74805 23463 74806
rect 115197 74806 115198 74838
rect 115262 74838 115268 74870
rect 115600 75142 115676 75148
rect 115600 75078 115606 75142
rect 115670 75078 115676 75142
rect 115600 74870 115676 75078
rect 115600 74838 115606 74870
rect 115262 74806 115263 74838
rect 115197 74805 115263 74806
rect 115605 74806 115606 74838
rect 115670 74838 115676 74870
rect 116552 75142 116628 75148
rect 116552 75078 116558 75142
rect 116622 75078 116628 75142
rect 116552 74870 116628 75078
rect 116552 74838 116558 74870
rect 115670 74806 115671 74838
rect 115605 74805 115671 74806
rect 116557 74806 116558 74838
rect 116622 74838 116628 74870
rect 116960 75142 117036 75148
rect 116960 75078 116966 75142
rect 117030 75078 117036 75142
rect 116960 74870 117036 75078
rect 116960 74838 116966 74870
rect 116622 74806 116623 74838
rect 116557 74805 116623 74806
rect 116965 74806 116966 74838
rect 117030 74838 117036 74870
rect 117030 74806 117031 74838
rect 116965 74805 117031 74806
rect 21760 74734 21836 74740
rect 21760 74670 21766 74734
rect 21830 74670 21836 74734
rect 21760 74462 21836 74670
rect 21760 74430 21766 74462
rect 21765 74398 21766 74430
rect 21830 74430 21836 74462
rect 22168 74734 22244 74740
rect 22168 74670 22174 74734
rect 22238 74670 22244 74734
rect 22445 74734 22511 74735
rect 22445 74702 22446 74734
rect 22168 74462 22244 74670
rect 22168 74430 22174 74462
rect 21830 74398 21831 74430
rect 21765 74397 21831 74398
rect 22173 74398 22174 74430
rect 22238 74430 22244 74462
rect 22440 74670 22446 74702
rect 22510 74702 22511 74734
rect 23120 74734 23196 74740
rect 22510 74670 22516 74702
rect 22440 74462 22516 74670
rect 22238 74398 22239 74430
rect 22173 74397 22239 74398
rect 22440 74398 22446 74462
rect 22510 74398 22516 74462
rect 23120 74670 23126 74734
rect 23190 74670 23196 74734
rect 23397 74734 23463 74735
rect 23397 74702 23398 74734
rect 23120 74462 23196 74670
rect 23120 74430 23126 74462
rect 22440 74392 22516 74398
rect 23125 74398 23126 74430
rect 23190 74430 23196 74462
rect 23392 74670 23398 74702
rect 23462 74702 23463 74734
rect 115197 74734 115263 74735
rect 115197 74702 115198 74734
rect 23462 74670 23468 74702
rect 23392 74462 23468 74670
rect 23190 74398 23191 74430
rect 23125 74397 23191 74398
rect 23392 74398 23398 74462
rect 23462 74398 23468 74462
rect 23392 74392 23468 74398
rect 115192 74670 115198 74702
rect 115262 74702 115263 74734
rect 115605 74734 115671 74735
rect 115605 74702 115606 74734
rect 115262 74670 115268 74702
rect 115192 74462 115268 74670
rect 115192 74398 115198 74462
rect 115262 74398 115268 74462
rect 115192 74392 115268 74398
rect 115600 74670 115606 74702
rect 115670 74702 115671 74734
rect 116008 74734 116084 74740
rect 115670 74670 115676 74702
rect 115600 74462 115676 74670
rect 115600 74398 115606 74462
rect 115670 74398 115676 74462
rect 116008 74670 116014 74734
rect 116078 74670 116084 74734
rect 116965 74734 117031 74735
rect 116965 74702 116966 74734
rect 116008 74462 116084 74670
rect 116008 74430 116014 74462
rect 115600 74392 115676 74398
rect 116013 74398 116014 74430
rect 116078 74430 116084 74462
rect 116960 74670 116966 74702
rect 117030 74702 117031 74734
rect 117030 74670 117036 74702
rect 116960 74462 117036 74670
rect 116078 74398 116079 74430
rect 116013 74397 116079 74398
rect 116960 74398 116966 74462
rect 117030 74398 117036 74462
rect 116960 74392 117036 74398
rect 21765 74326 21831 74327
rect 21765 74294 21766 74326
rect 952 74126 1230 74190
rect 1294 74126 1300 74190
rect 952 72694 1300 74126
rect 21760 74262 21766 74294
rect 21830 74294 21831 74326
rect 22581 74326 22647 74327
rect 22581 74294 22582 74326
rect 21830 74262 21836 74294
rect 21760 74054 21836 74262
rect 21760 73990 21766 74054
rect 21830 73990 21836 74054
rect 21760 73984 21836 73990
rect 22576 74262 22582 74294
rect 22646 74294 22647 74326
rect 22984 74326 23060 74332
rect 22646 74262 22652 74294
rect 22576 74054 22652 74262
rect 22576 73990 22582 74054
rect 22646 73990 22652 74054
rect 22984 74262 22990 74326
rect 23054 74262 23060 74326
rect 22984 74054 23060 74262
rect 22984 74022 22990 74054
rect 22576 73984 22652 73990
rect 22989 73990 22990 74022
rect 23054 74022 23060 74054
rect 23392 74326 23468 74332
rect 23392 74262 23398 74326
rect 23462 74262 23468 74326
rect 23392 74054 23468 74262
rect 23392 74022 23398 74054
rect 23054 73990 23055 74022
rect 22989 73989 23055 73990
rect 23397 73990 23398 74022
rect 23462 74022 23468 74054
rect 115192 74326 115268 74332
rect 115192 74262 115198 74326
rect 115262 74262 115268 74326
rect 115192 74054 115268 74262
rect 115192 74022 115198 74054
rect 23462 73990 23463 74022
rect 23397 73989 23463 73990
rect 115197 73990 115198 74022
rect 115262 74022 115268 74054
rect 115600 74326 115676 74332
rect 115600 74262 115606 74326
rect 115670 74262 115676 74326
rect 116013 74326 116079 74327
rect 116013 74294 116014 74326
rect 115600 74054 115676 74262
rect 115600 74022 115606 74054
rect 115262 73990 115263 74022
rect 115197 73989 115263 73990
rect 115605 73990 115606 74022
rect 115670 74022 115676 74054
rect 116008 74262 116014 74294
rect 116078 74294 116079 74326
rect 116960 74326 117036 74332
rect 116078 74262 116084 74294
rect 116008 74054 116084 74262
rect 115670 73990 115671 74022
rect 115605 73989 115671 73990
rect 116008 73990 116014 74054
rect 116078 73990 116084 74054
rect 116960 74262 116966 74326
rect 117030 74262 117036 74326
rect 116960 74054 117036 74262
rect 116960 74022 116966 74054
rect 116008 73984 116084 73990
rect 116965 73990 116966 74022
rect 117030 74022 117036 74054
rect 137496 74326 137844 75894
rect 137496 74262 137502 74326
rect 137566 74262 137844 74326
rect 117030 73990 117031 74022
rect 116965 73989 117031 73990
rect 22712 73918 22788 73924
rect 22712 73854 22718 73918
rect 22782 73854 22788 73918
rect 22989 73918 23055 73919
rect 22989 73886 22990 73918
rect 22712 73646 22788 73854
rect 22712 73614 22718 73646
rect 22717 73582 22718 73614
rect 22782 73614 22788 73646
rect 22984 73854 22990 73886
rect 23054 73886 23055 73918
rect 23397 73918 23463 73919
rect 23397 73886 23398 73918
rect 23054 73854 23060 73886
rect 22984 73646 23060 73854
rect 22782 73582 22783 73614
rect 22717 73581 22783 73582
rect 22984 73582 22990 73646
rect 23054 73582 23060 73646
rect 22984 73576 23060 73582
rect 23392 73854 23398 73886
rect 23462 73886 23463 73918
rect 115192 73918 115268 73924
rect 23462 73854 23468 73886
rect 23392 73646 23468 73854
rect 23392 73582 23398 73646
rect 23462 73582 23468 73646
rect 115192 73854 115198 73918
rect 115262 73854 115268 73918
rect 115605 73918 115671 73919
rect 115605 73886 115606 73918
rect 115192 73646 115268 73854
rect 115192 73614 115198 73646
rect 23392 73576 23468 73582
rect 115197 73582 115198 73614
rect 115262 73614 115268 73646
rect 115600 73854 115606 73886
rect 115670 73886 115671 73918
rect 116144 73918 116220 73924
rect 115670 73854 115676 73886
rect 115600 73646 115676 73854
rect 115262 73582 115263 73614
rect 115197 73581 115263 73582
rect 115600 73582 115606 73646
rect 115670 73582 115676 73646
rect 116144 73854 116150 73918
rect 116214 73854 116220 73918
rect 116144 73646 116220 73854
rect 116144 73614 116150 73646
rect 115600 73576 115676 73582
rect 116149 73582 116150 73614
rect 116214 73614 116220 73646
rect 116214 73582 116215 73614
rect 116149 73581 116215 73582
rect 21901 73510 21967 73511
rect 21901 73478 21902 73510
rect 21896 73446 21902 73478
rect 21966 73478 21967 73510
rect 22168 73510 22244 73516
rect 21966 73446 21972 73478
rect 21896 73238 21972 73446
rect 21896 73174 21902 73238
rect 21966 73174 21972 73238
rect 22168 73446 22174 73510
rect 22238 73446 22244 73510
rect 22989 73510 23055 73511
rect 22989 73478 22990 73510
rect 22168 73238 22244 73446
rect 22168 73206 22174 73238
rect 21896 73168 21972 73174
rect 22173 73174 22174 73206
rect 22238 73206 22244 73238
rect 22984 73446 22990 73478
rect 23054 73478 23055 73510
rect 23533 73510 23599 73511
rect 23533 73478 23534 73510
rect 23054 73446 23060 73478
rect 22984 73238 23060 73446
rect 22238 73174 22239 73206
rect 22173 73173 22239 73174
rect 22984 73174 22990 73238
rect 23054 73174 23060 73238
rect 22984 73168 23060 73174
rect 23528 73446 23534 73478
rect 23598 73478 23599 73510
rect 115333 73510 115399 73511
rect 115333 73478 115334 73510
rect 23598 73446 23604 73478
rect 23528 73238 23604 73446
rect 23528 73174 23534 73238
rect 23598 73174 23604 73238
rect 23528 73168 23604 73174
rect 115328 73446 115334 73478
rect 115398 73478 115399 73510
rect 115736 73510 115812 73516
rect 115398 73446 115404 73478
rect 115328 73238 115404 73446
rect 115328 73174 115334 73238
rect 115398 73174 115404 73238
rect 115736 73446 115742 73510
rect 115806 73446 115812 73510
rect 116013 73510 116079 73511
rect 116013 73478 116014 73510
rect 115736 73238 115812 73446
rect 115736 73206 115742 73238
rect 115328 73168 115404 73174
rect 115741 73174 115742 73206
rect 115806 73206 115812 73238
rect 116008 73446 116014 73478
rect 116078 73478 116079 73510
rect 116824 73510 116900 73516
rect 116078 73446 116084 73478
rect 116008 73238 116084 73446
rect 115806 73174 115807 73206
rect 115741 73173 115807 73174
rect 116008 73174 116014 73238
rect 116078 73174 116084 73238
rect 116824 73446 116830 73510
rect 116894 73446 116900 73510
rect 116824 73238 116900 73446
rect 116824 73206 116830 73238
rect 116008 73168 116084 73174
rect 116829 73174 116830 73206
rect 116894 73206 116900 73238
rect 116894 73174 116895 73206
rect 116829 73173 116895 73174
rect 22440 73102 22516 73108
rect 22440 73038 22446 73102
rect 22510 73038 22516 73102
rect 952 72630 1230 72694
rect 1294 72630 1300 72694
rect 952 71062 1300 72630
rect 21896 72830 21972 72836
rect 21896 72766 21902 72830
rect 21966 72766 21972 72830
rect 22440 72830 22516 73038
rect 22440 72798 22446 72830
rect 21896 72558 21972 72766
rect 22445 72766 22446 72798
rect 22510 72798 22516 72830
rect 22984 73102 23060 73108
rect 22984 73038 22990 73102
rect 23054 73038 23060 73102
rect 22984 72830 23060 73038
rect 22984 72798 22990 72830
rect 22510 72766 22511 72798
rect 22445 72765 22511 72766
rect 22989 72766 22990 72798
rect 23054 72798 23060 72830
rect 23392 73102 23468 73108
rect 23392 73038 23398 73102
rect 23462 73038 23468 73102
rect 115333 73102 115399 73103
rect 115333 73070 115334 73102
rect 23392 72830 23468 73038
rect 115328 73038 115334 73070
rect 115398 73070 115399 73102
rect 115741 73102 115807 73103
rect 115741 73070 115742 73102
rect 115398 73038 115404 73070
rect 23392 72798 23398 72830
rect 23054 72766 23055 72798
rect 22989 72765 23055 72766
rect 23397 72766 23398 72798
rect 23462 72798 23468 72830
rect 28424 72966 28500 72972
rect 28424 72902 28430 72966
rect 28494 72902 28500 72966
rect 23462 72766 23463 72798
rect 23397 72765 23463 72766
rect 28424 72694 28500 72902
rect 115328 72830 115404 73038
rect 115328 72766 115334 72830
rect 115398 72766 115404 72830
rect 115328 72760 115404 72766
rect 115736 73038 115742 73070
rect 115806 73070 115807 73102
rect 116008 73102 116084 73108
rect 115806 73038 115812 73070
rect 115736 72830 115812 73038
rect 115736 72766 115742 72830
rect 115806 72766 115812 72830
rect 116008 73038 116014 73102
rect 116078 73038 116084 73102
rect 116421 73102 116487 73103
rect 116421 73070 116422 73102
rect 116008 72830 116084 73038
rect 116008 72798 116014 72830
rect 115736 72760 115812 72766
rect 116013 72766 116014 72798
rect 116078 72798 116084 72830
rect 116416 73038 116422 73070
rect 116486 73070 116487 73102
rect 116486 73038 116492 73070
rect 116416 72830 116492 73038
rect 116078 72766 116079 72798
rect 116013 72765 116079 72766
rect 116416 72766 116422 72830
rect 116486 72766 116492 72830
rect 116965 72830 117031 72831
rect 116965 72798 116966 72830
rect 116416 72760 116492 72766
rect 116960 72766 116966 72798
rect 117030 72798 117031 72830
rect 117030 72766 117036 72798
rect 28424 72662 28430 72694
rect 28429 72630 28430 72662
rect 28494 72662 28500 72694
rect 28494 72630 28495 72662
rect 28429 72629 28495 72630
rect 21896 72526 21902 72558
rect 21901 72494 21902 72526
rect 21966 72526 21972 72558
rect 28429 72558 28495 72559
rect 28429 72526 28430 72558
rect 21966 72494 21967 72526
rect 21901 72493 21967 72494
rect 28424 72494 28430 72526
rect 28494 72526 28495 72558
rect 110432 72558 110508 72564
rect 28494 72494 28500 72526
rect 21765 72422 21831 72423
rect 21765 72390 21766 72422
rect 21760 72358 21766 72390
rect 21830 72390 21831 72422
rect 22168 72422 22244 72428
rect 21830 72358 21836 72390
rect 21760 72150 21836 72358
rect 21760 72086 21766 72150
rect 21830 72086 21836 72150
rect 22168 72358 22174 72422
rect 22238 72358 22244 72422
rect 22168 72150 22244 72358
rect 22168 72118 22174 72150
rect 21760 72080 21836 72086
rect 22173 72086 22174 72118
rect 22238 72118 22244 72150
rect 22576 72422 22652 72428
rect 22576 72358 22582 72422
rect 22646 72358 22652 72422
rect 22576 72150 22652 72358
rect 28424 72286 28500 72494
rect 28424 72222 28430 72286
rect 28494 72222 28500 72286
rect 110432 72494 110438 72558
rect 110502 72494 110508 72558
rect 110432 72286 110508 72494
rect 116960 72558 117036 72766
rect 116960 72494 116966 72558
rect 117030 72494 117036 72558
rect 116960 72488 117036 72494
rect 137496 72694 137844 74262
rect 137496 72630 137502 72694
rect 137566 72630 137844 72694
rect 116013 72422 116079 72423
rect 116013 72390 116014 72422
rect 110432 72254 110438 72286
rect 28424 72216 28500 72222
rect 110437 72222 110438 72254
rect 110502 72254 110508 72286
rect 116008 72358 116014 72390
rect 116078 72390 116079 72422
rect 116829 72422 116895 72423
rect 116829 72390 116830 72422
rect 116078 72358 116084 72390
rect 110502 72222 110503 72254
rect 110437 72221 110503 72222
rect 22576 72118 22582 72150
rect 22238 72086 22239 72118
rect 22173 72085 22239 72086
rect 22581 72086 22582 72118
rect 22646 72118 22652 72150
rect 28293 72150 28359 72151
rect 28293 72118 28294 72150
rect 22646 72086 22647 72118
rect 22581 72085 22647 72086
rect 28288 72086 28294 72118
rect 28358 72118 28359 72150
rect 116008 72150 116084 72358
rect 28358 72086 28364 72118
rect 21896 72014 21972 72020
rect 21896 71950 21902 72014
rect 21966 71950 21972 72014
rect 21896 71742 21972 71950
rect 28288 71878 28364 72086
rect 116008 72086 116014 72150
rect 116078 72086 116084 72150
rect 116008 72080 116084 72086
rect 116824 72358 116830 72390
rect 116894 72390 116895 72422
rect 116894 72358 116900 72390
rect 116824 72150 116900 72358
rect 116824 72086 116830 72150
rect 116894 72086 116900 72150
rect 116824 72080 116900 72086
rect 116829 72014 116895 72015
rect 116829 71982 116830 72014
rect 28288 71814 28294 71878
rect 28358 71814 28364 71878
rect 28288 71808 28364 71814
rect 116824 71950 116830 71982
rect 116894 71982 116895 72014
rect 116894 71950 116900 71982
rect 21896 71710 21902 71742
rect 21901 71678 21902 71710
rect 21966 71710 21972 71742
rect 116824 71742 116900 71950
rect 21966 71678 21967 71710
rect 21901 71677 21967 71678
rect 116824 71678 116830 71742
rect 116894 71678 116900 71742
rect 116824 71672 116900 71678
rect 21901 71606 21967 71607
rect 21901 71574 21902 71606
rect 21896 71542 21902 71574
rect 21966 71574 21967 71606
rect 22440 71606 22516 71612
rect 21966 71542 21972 71574
rect 21896 71334 21972 71542
rect 21896 71270 21902 71334
rect 21966 71270 21972 71334
rect 22440 71542 22446 71606
rect 22510 71542 22516 71606
rect 22717 71606 22783 71607
rect 22717 71574 22718 71606
rect 22440 71334 22516 71542
rect 22440 71302 22446 71334
rect 21896 71264 21972 71270
rect 22445 71270 22446 71302
rect 22510 71302 22516 71334
rect 22712 71542 22718 71574
rect 22782 71574 22783 71606
rect 22984 71606 23060 71612
rect 22782 71542 22788 71574
rect 22712 71334 22788 71542
rect 22510 71270 22511 71302
rect 22445 71269 22511 71270
rect 22712 71270 22718 71334
rect 22782 71270 22788 71334
rect 22984 71542 22990 71606
rect 23054 71542 23060 71606
rect 22984 71334 23060 71542
rect 22984 71302 22990 71334
rect 22712 71264 22788 71270
rect 22989 71270 22990 71302
rect 23054 71302 23060 71334
rect 23528 71606 23604 71612
rect 23528 71542 23534 71606
rect 23598 71542 23604 71606
rect 115197 71606 115263 71607
rect 115197 71574 115198 71606
rect 23528 71334 23604 71542
rect 23528 71302 23534 71334
rect 23054 71270 23055 71302
rect 22989 71269 23055 71270
rect 23533 71270 23534 71302
rect 23598 71302 23604 71334
rect 115192 71542 115198 71574
rect 115262 71574 115263 71606
rect 115736 71606 115812 71612
rect 115262 71542 115268 71574
rect 115192 71334 115268 71542
rect 23598 71270 23599 71302
rect 23533 71269 23599 71270
rect 115192 71270 115198 71334
rect 115262 71270 115268 71334
rect 115736 71542 115742 71606
rect 115806 71542 115812 71606
rect 115736 71334 115812 71542
rect 115736 71302 115742 71334
rect 115192 71264 115268 71270
rect 115741 71270 115742 71302
rect 115806 71302 115812 71334
rect 116008 71606 116084 71612
rect 116008 71542 116014 71606
rect 116078 71542 116084 71606
rect 116285 71606 116351 71607
rect 116285 71574 116286 71606
rect 116008 71334 116084 71542
rect 116008 71302 116014 71334
rect 115806 71270 115807 71302
rect 115741 71269 115807 71270
rect 116013 71270 116014 71302
rect 116078 71302 116084 71334
rect 116280 71542 116286 71574
rect 116350 71574 116351 71606
rect 116824 71606 116900 71612
rect 116350 71542 116356 71574
rect 116280 71334 116356 71542
rect 116078 71270 116079 71302
rect 116013 71269 116079 71270
rect 116280 71270 116286 71334
rect 116350 71270 116356 71334
rect 116824 71542 116830 71606
rect 116894 71542 116900 71606
rect 116824 71334 116900 71542
rect 116824 71302 116830 71334
rect 116280 71264 116356 71270
rect 116829 71270 116830 71302
rect 116894 71302 116900 71334
rect 116894 71270 116895 71302
rect 116829 71269 116895 71270
rect 952 70998 1230 71062
rect 1294 70998 1300 71062
rect 952 69294 1300 70998
rect 21760 71198 21836 71204
rect 21760 71134 21766 71198
rect 21830 71134 21836 71198
rect 22173 71198 22239 71199
rect 22173 71166 22174 71198
rect 21760 70926 21836 71134
rect 21760 70894 21766 70926
rect 21765 70862 21766 70894
rect 21830 70894 21836 70926
rect 22168 71134 22174 71166
rect 22238 71166 22239 71198
rect 22576 71198 22652 71204
rect 22238 71134 22244 71166
rect 22168 70926 22244 71134
rect 21830 70862 21831 70894
rect 21765 70861 21831 70862
rect 22168 70862 22174 70926
rect 22238 70862 22244 70926
rect 22576 71134 22582 71198
rect 22646 71134 22652 71198
rect 22989 71198 23055 71199
rect 22989 71166 22990 71198
rect 22576 70926 22652 71134
rect 22576 70894 22582 70926
rect 22168 70856 22244 70862
rect 22581 70862 22582 70894
rect 22646 70894 22652 70926
rect 22984 71134 22990 71166
rect 23054 71166 23055 71198
rect 23528 71198 23604 71204
rect 23054 71134 23060 71166
rect 22984 70926 23060 71134
rect 22646 70862 22647 70894
rect 22581 70861 22647 70862
rect 22984 70862 22990 70926
rect 23054 70862 23060 70926
rect 23528 71134 23534 71198
rect 23598 71134 23604 71198
rect 115333 71198 115399 71199
rect 115333 71166 115334 71198
rect 23528 70926 23604 71134
rect 23528 70894 23534 70926
rect 22984 70856 23060 70862
rect 23533 70862 23534 70894
rect 23598 70894 23604 70926
rect 115328 71134 115334 71166
rect 115398 71166 115399 71198
rect 115741 71198 115807 71199
rect 115741 71166 115742 71198
rect 115398 71134 115404 71166
rect 115328 70926 115404 71134
rect 23598 70862 23599 70894
rect 23533 70861 23599 70862
rect 115328 70862 115334 70926
rect 115398 70862 115404 70926
rect 115328 70856 115404 70862
rect 115736 71134 115742 71166
rect 115806 71166 115807 71198
rect 116280 71198 116356 71204
rect 115806 71134 115812 71166
rect 115736 70926 115812 71134
rect 115736 70862 115742 70926
rect 115806 70862 115812 70926
rect 116280 71134 116286 71198
rect 116350 71134 116356 71198
rect 116829 71198 116895 71199
rect 116829 71166 116830 71198
rect 116280 70926 116356 71134
rect 116280 70894 116286 70926
rect 115736 70856 115812 70862
rect 116285 70862 116286 70894
rect 116350 70894 116356 70926
rect 116824 71134 116830 71166
rect 116894 71166 116895 71198
rect 116894 71134 116900 71166
rect 116824 70926 116900 71134
rect 116350 70862 116351 70894
rect 116285 70861 116351 70862
rect 116824 70862 116830 70926
rect 116894 70862 116900 70926
rect 116824 70856 116900 70862
rect 137496 71062 137844 72630
rect 137496 70998 137502 71062
rect 137566 70998 137844 71062
rect 21901 70790 21967 70791
rect 21901 70758 21902 70790
rect 21896 70726 21902 70758
rect 21966 70758 21967 70790
rect 22717 70790 22783 70791
rect 22717 70758 22718 70790
rect 21966 70726 21972 70758
rect 21896 70518 21972 70726
rect 21896 70454 21902 70518
rect 21966 70454 21972 70518
rect 21896 70448 21972 70454
rect 22712 70726 22718 70758
rect 22782 70758 22783 70790
rect 23120 70790 23196 70796
rect 22782 70726 22788 70758
rect 22712 70518 22788 70726
rect 22712 70454 22718 70518
rect 22782 70454 22788 70518
rect 23120 70726 23126 70790
rect 23190 70726 23196 70790
rect 23397 70790 23463 70791
rect 23397 70758 23398 70790
rect 23120 70518 23196 70726
rect 23120 70486 23126 70518
rect 22712 70448 22788 70454
rect 23125 70454 23126 70486
rect 23190 70486 23196 70518
rect 23392 70726 23398 70758
rect 23462 70758 23463 70790
rect 115192 70790 115268 70796
rect 23462 70726 23468 70758
rect 23392 70518 23468 70726
rect 23190 70454 23191 70486
rect 23125 70453 23191 70454
rect 23392 70454 23398 70518
rect 23462 70454 23468 70518
rect 115192 70726 115198 70790
rect 115262 70726 115268 70790
rect 115192 70518 115268 70726
rect 115192 70486 115198 70518
rect 23392 70448 23468 70454
rect 115197 70454 115198 70486
rect 115262 70486 115268 70518
rect 115600 70790 115676 70796
rect 115600 70726 115606 70790
rect 115670 70726 115676 70790
rect 115600 70518 115676 70726
rect 115600 70486 115606 70518
rect 115262 70454 115263 70486
rect 115197 70453 115263 70454
rect 115605 70454 115606 70486
rect 115670 70486 115676 70518
rect 116552 70790 116628 70796
rect 116552 70726 116558 70790
rect 116622 70726 116628 70790
rect 116965 70790 117031 70791
rect 116965 70758 116966 70790
rect 116552 70518 116628 70726
rect 116552 70486 116558 70518
rect 115670 70454 115671 70486
rect 115605 70453 115671 70454
rect 116557 70454 116558 70486
rect 116622 70486 116628 70518
rect 116960 70726 116966 70758
rect 117030 70758 117031 70790
rect 117030 70726 117036 70758
rect 116960 70518 117036 70726
rect 116622 70454 116623 70486
rect 116557 70453 116623 70454
rect 116960 70454 116966 70518
rect 117030 70454 117036 70518
rect 116960 70448 117036 70454
rect 21901 70382 21967 70383
rect 21901 70350 21902 70382
rect 21896 70318 21902 70350
rect 21966 70350 21967 70382
rect 22445 70382 22511 70383
rect 22445 70350 22446 70382
rect 21966 70318 21972 70350
rect 21896 70110 21972 70318
rect 21896 70046 21902 70110
rect 21966 70046 21972 70110
rect 21896 70040 21972 70046
rect 22440 70318 22446 70350
rect 22510 70350 22511 70382
rect 23125 70382 23191 70383
rect 23125 70350 23126 70382
rect 22510 70318 22516 70350
rect 22440 70110 22516 70318
rect 22440 70046 22446 70110
rect 22510 70046 22516 70110
rect 22440 70040 22516 70046
rect 23120 70318 23126 70350
rect 23190 70350 23191 70382
rect 23528 70382 23604 70388
rect 23190 70318 23196 70350
rect 23120 70110 23196 70318
rect 23120 70046 23126 70110
rect 23190 70046 23196 70110
rect 23528 70318 23534 70382
rect 23598 70318 23604 70382
rect 23528 70110 23604 70318
rect 23528 70078 23534 70110
rect 23120 70040 23196 70046
rect 23533 70046 23534 70078
rect 23598 70078 23604 70110
rect 24208 70382 24284 70388
rect 24208 70318 24214 70382
rect 24278 70318 24284 70382
rect 24208 70110 24284 70318
rect 24208 70078 24214 70110
rect 23598 70046 23599 70078
rect 23533 70045 23599 70046
rect 24213 70046 24214 70078
rect 24278 70078 24284 70110
rect 113288 70382 113364 70388
rect 113288 70318 113294 70382
rect 113358 70318 113364 70382
rect 115197 70382 115263 70383
rect 115197 70350 115198 70382
rect 24278 70046 24279 70078
rect 24213 70045 24279 70046
rect 22173 69974 22239 69975
rect 22173 69942 22174 69974
rect 22168 69910 22174 69942
rect 22238 69942 22239 69974
rect 22581 69974 22647 69975
rect 22581 69942 22582 69974
rect 22238 69910 22244 69942
rect 22168 69702 22244 69910
rect 22168 69638 22174 69702
rect 22238 69638 22244 69702
rect 22168 69632 22244 69638
rect 22576 69910 22582 69942
rect 22646 69942 22647 69974
rect 22984 69974 23060 69980
rect 22646 69910 22652 69942
rect 22576 69702 22652 69910
rect 22576 69638 22582 69702
rect 22646 69638 22652 69702
rect 22984 69910 22990 69974
rect 23054 69910 23060 69974
rect 22984 69702 23060 69910
rect 22984 69670 22990 69702
rect 22576 69632 22652 69638
rect 22989 69638 22990 69670
rect 23054 69670 23060 69702
rect 23392 69974 23468 69980
rect 23392 69910 23398 69974
rect 23462 69910 23468 69974
rect 23392 69702 23468 69910
rect 23392 69670 23398 69702
rect 23054 69638 23055 69670
rect 22989 69637 23055 69638
rect 23397 69638 23398 69670
rect 23462 69670 23468 69702
rect 113288 69702 113364 70318
rect 115192 70318 115198 70350
rect 115262 70350 115263 70382
rect 115736 70382 115812 70388
rect 115262 70318 115268 70350
rect 115192 70110 115268 70318
rect 115192 70046 115198 70110
rect 115262 70046 115268 70110
rect 115736 70318 115742 70382
rect 115806 70318 115812 70382
rect 116149 70382 116215 70383
rect 116149 70350 116150 70382
rect 115736 70110 115812 70318
rect 115736 70078 115742 70110
rect 115192 70040 115268 70046
rect 115741 70046 115742 70078
rect 115806 70078 115812 70110
rect 116144 70318 116150 70350
rect 116214 70350 116215 70382
rect 116965 70382 117031 70383
rect 116965 70350 116966 70382
rect 116214 70318 116220 70350
rect 116144 70110 116220 70318
rect 115806 70046 115807 70078
rect 115741 70045 115807 70046
rect 116144 70046 116150 70110
rect 116214 70046 116220 70110
rect 116144 70040 116220 70046
rect 116960 70318 116966 70350
rect 117030 70350 117031 70382
rect 117030 70318 117036 70350
rect 116960 70110 117036 70318
rect 116960 70046 116966 70110
rect 117030 70046 117036 70110
rect 116960 70040 117036 70046
rect 113288 69670 113294 69702
rect 23462 69638 23463 69670
rect 23397 69637 23463 69638
rect 113293 69638 113294 69670
rect 113358 69670 113364 69702
rect 115192 69974 115268 69980
rect 115192 69910 115198 69974
rect 115262 69910 115268 69974
rect 115192 69702 115268 69910
rect 115192 69670 115198 69702
rect 113358 69638 113359 69670
rect 113293 69637 113359 69638
rect 115197 69638 115198 69670
rect 115262 69670 115268 69702
rect 115600 69974 115676 69980
rect 115600 69910 115606 69974
rect 115670 69910 115676 69974
rect 115600 69702 115676 69910
rect 115600 69670 115606 69702
rect 115262 69638 115263 69670
rect 115197 69637 115263 69638
rect 115605 69638 115606 69670
rect 115670 69670 115676 69702
rect 116008 69974 116084 69980
rect 116008 69910 116014 69974
rect 116078 69910 116084 69974
rect 116008 69702 116084 69910
rect 116008 69670 116014 69702
rect 115670 69638 115671 69670
rect 115605 69637 115671 69638
rect 116013 69638 116014 69670
rect 116078 69670 116084 69702
rect 116552 69974 116628 69980
rect 116552 69910 116558 69974
rect 116622 69910 116628 69974
rect 116552 69702 116628 69910
rect 116552 69670 116558 69702
rect 116078 69638 116079 69670
rect 116013 69637 116079 69638
rect 116557 69638 116558 69670
rect 116622 69670 116628 69702
rect 116622 69638 116623 69670
rect 116557 69637 116623 69638
rect 952 69230 1230 69294
rect 1294 69230 1300 69294
rect 21896 69566 21972 69572
rect 21896 69502 21902 69566
rect 21966 69502 21972 69566
rect 21896 69294 21972 69502
rect 21896 69262 21902 69294
rect 952 67662 1300 69230
rect 21901 69230 21902 69262
rect 21966 69262 21972 69294
rect 22440 69566 22516 69572
rect 22440 69502 22446 69566
rect 22510 69502 22516 69566
rect 22989 69566 23055 69567
rect 22989 69534 22990 69566
rect 22440 69294 22516 69502
rect 22440 69262 22446 69294
rect 21966 69230 21967 69262
rect 21901 69229 21967 69230
rect 22445 69230 22446 69262
rect 22510 69262 22516 69294
rect 22984 69502 22990 69534
rect 23054 69534 23055 69566
rect 23397 69566 23463 69567
rect 23397 69534 23398 69566
rect 23054 69502 23060 69534
rect 22984 69294 23060 69502
rect 22510 69230 22511 69262
rect 22445 69229 22511 69230
rect 22984 69230 22990 69294
rect 23054 69230 23060 69294
rect 22984 69224 23060 69230
rect 23392 69502 23398 69534
rect 23462 69534 23463 69566
rect 115192 69566 115268 69572
rect 23462 69502 23468 69534
rect 23392 69294 23468 69502
rect 23392 69230 23398 69294
rect 23462 69230 23468 69294
rect 115192 69502 115198 69566
rect 115262 69502 115268 69566
rect 115605 69566 115671 69567
rect 115605 69534 115606 69566
rect 115192 69294 115268 69502
rect 115192 69262 115198 69294
rect 23392 69224 23468 69230
rect 115197 69230 115198 69262
rect 115262 69262 115268 69294
rect 115600 69502 115606 69534
rect 115670 69534 115671 69566
rect 116144 69566 116220 69572
rect 115670 69502 115676 69534
rect 115600 69294 115676 69502
rect 115262 69230 115263 69262
rect 115197 69229 115263 69230
rect 115600 69230 115606 69294
rect 115670 69230 115676 69294
rect 116144 69502 116150 69566
rect 116214 69502 116220 69566
rect 116829 69566 116895 69567
rect 116829 69534 116830 69566
rect 116144 69294 116220 69502
rect 116144 69262 116150 69294
rect 115600 69224 115676 69230
rect 116149 69230 116150 69262
rect 116214 69262 116220 69294
rect 116824 69502 116830 69534
rect 116894 69534 116895 69566
rect 116894 69502 116900 69534
rect 116824 69294 116900 69502
rect 116214 69230 116215 69262
rect 116149 69229 116215 69230
rect 116824 69230 116830 69294
rect 116894 69230 116900 69294
rect 116824 69224 116900 69230
rect 137496 69294 137844 70998
rect 137496 69230 137502 69294
rect 137566 69230 137844 69294
rect 22576 69158 22652 69164
rect 22576 69094 22582 69158
rect 22646 69094 22652 69158
rect 21896 68886 21972 68892
rect 21896 68822 21902 68886
rect 21966 68822 21972 68886
rect 22576 68886 22652 69094
rect 22576 68854 22582 68886
rect 21896 68614 21972 68822
rect 22581 68822 22582 68854
rect 22646 68854 22652 68886
rect 23120 69158 23196 69164
rect 23120 69094 23126 69158
rect 23190 69094 23196 69158
rect 23533 69158 23599 69159
rect 23533 69126 23534 69158
rect 23120 68886 23196 69094
rect 23120 68854 23126 68886
rect 22646 68822 22647 68854
rect 22581 68821 22647 68822
rect 23125 68822 23126 68854
rect 23190 68854 23196 68886
rect 23528 69094 23534 69126
rect 23598 69126 23599 69158
rect 115328 69158 115404 69164
rect 23598 69094 23604 69126
rect 23528 68886 23604 69094
rect 115328 69094 115334 69158
rect 115398 69094 115404 69158
rect 23190 68822 23191 68854
rect 23125 68821 23191 68822
rect 23528 68822 23534 68886
rect 23598 68822 23604 68886
rect 23528 68816 23604 68822
rect 28288 69022 28364 69028
rect 28288 68958 28294 69022
rect 28358 68958 28364 69022
rect 23125 68750 23191 68751
rect 23125 68718 23126 68750
rect 21896 68582 21902 68614
rect 21901 68550 21902 68582
rect 21966 68582 21972 68614
rect 23120 68686 23126 68718
rect 23190 68718 23191 68750
rect 23392 68750 23468 68756
rect 23190 68686 23196 68718
rect 21966 68550 21967 68582
rect 21901 68549 21967 68550
rect 23120 68478 23196 68686
rect 23120 68414 23126 68478
rect 23190 68414 23196 68478
rect 23392 68686 23398 68750
rect 23462 68686 23468 68750
rect 28288 68750 28364 68958
rect 110432 69022 110508 69028
rect 110432 68958 110438 69022
rect 110502 68958 110508 69022
rect 28288 68718 28294 68750
rect 23392 68478 23468 68686
rect 28293 68686 28294 68718
rect 28358 68718 28364 68750
rect 28424 68750 28500 68756
rect 28358 68686 28359 68718
rect 28293 68685 28359 68686
rect 28424 68686 28430 68750
rect 28494 68686 28500 68750
rect 110432 68750 110508 68958
rect 115328 68886 115404 69094
rect 115328 68854 115334 68886
rect 115333 68822 115334 68854
rect 115398 68854 115404 68886
rect 115736 69158 115812 69164
rect 115736 69094 115742 69158
rect 115806 69094 115812 69158
rect 116285 69158 116351 69159
rect 116285 69126 116286 69158
rect 115736 68886 115812 69094
rect 115736 68854 115742 68886
rect 115398 68822 115399 68854
rect 115333 68821 115399 68822
rect 115741 68822 115742 68854
rect 115806 68854 115812 68886
rect 116280 69094 116286 69126
rect 116350 69126 116351 69158
rect 116350 69094 116356 69126
rect 116280 68886 116356 69094
rect 115806 68822 115807 68854
rect 115741 68821 115807 68822
rect 116280 68822 116286 68886
rect 116350 68822 116356 68886
rect 116280 68816 116356 68822
rect 116960 68886 117036 68892
rect 116960 68822 116966 68886
rect 117030 68822 117036 68886
rect 110432 68718 110438 68750
rect 23392 68446 23398 68478
rect 23120 68408 23196 68414
rect 23397 68414 23398 68446
rect 23462 68446 23468 68478
rect 23462 68414 23463 68446
rect 23397 68413 23463 68414
rect 22173 68342 22239 68343
rect 22173 68310 22174 68342
rect 22168 68278 22174 68310
rect 22238 68310 22239 68342
rect 22581 68342 22647 68343
rect 22581 68310 22582 68342
rect 22238 68278 22244 68310
rect 21760 68070 21836 68076
rect 21760 68006 21766 68070
rect 21830 68006 21836 68070
rect 21760 67798 21836 68006
rect 22168 68070 22244 68278
rect 22168 68006 22174 68070
rect 22238 68006 22244 68070
rect 22168 68000 22244 68006
rect 22576 68278 22582 68310
rect 22646 68310 22647 68342
rect 28424 68342 28500 68686
rect 110437 68686 110438 68718
rect 110502 68718 110508 68750
rect 115333 68750 115399 68751
rect 115333 68718 115334 68750
rect 110502 68686 110503 68718
rect 110437 68685 110503 68686
rect 115328 68686 115334 68718
rect 115398 68718 115399 68750
rect 115741 68750 115807 68751
rect 115741 68718 115742 68750
rect 115398 68686 115404 68718
rect 115328 68478 115404 68686
rect 115328 68414 115334 68478
rect 115398 68414 115404 68478
rect 115328 68408 115404 68414
rect 115736 68686 115742 68718
rect 115806 68718 115807 68750
rect 115806 68686 115812 68718
rect 115736 68478 115812 68686
rect 116960 68614 117036 68822
rect 116960 68582 116966 68614
rect 116965 68550 116966 68582
rect 117030 68582 117036 68614
rect 117030 68550 117031 68582
rect 116965 68549 117031 68550
rect 115736 68414 115742 68478
rect 115806 68414 115812 68478
rect 115736 68408 115812 68414
rect 28424 68310 28430 68342
rect 22646 68278 22652 68310
rect 22576 68070 22652 68278
rect 28429 68278 28430 68310
rect 28494 68310 28500 68342
rect 116008 68342 116084 68348
rect 28494 68278 28495 68310
rect 28429 68277 28495 68278
rect 116008 68278 116014 68342
rect 116078 68278 116084 68342
rect 22576 68006 22582 68070
rect 22646 68006 22652 68070
rect 22576 68000 22652 68006
rect 110432 68206 110508 68212
rect 110432 68142 110438 68206
rect 110502 68142 110508 68206
rect 110432 67934 110508 68142
rect 116008 68070 116084 68278
rect 116008 68038 116014 68070
rect 116013 68006 116014 68038
rect 116078 68038 116084 68070
rect 116824 68070 116900 68076
rect 116078 68006 116079 68038
rect 116013 68005 116079 68006
rect 116824 68006 116830 68070
rect 116894 68006 116900 68070
rect 110432 67902 110438 67934
rect 110437 67870 110438 67902
rect 110502 67902 110508 67934
rect 110502 67870 110503 67902
rect 110437 67869 110503 67870
rect 21760 67766 21766 67798
rect 21765 67734 21766 67766
rect 21830 67766 21836 67798
rect 116824 67798 116900 68006
rect 116824 67766 116830 67798
rect 21830 67734 21831 67766
rect 21765 67733 21831 67734
rect 116829 67734 116830 67766
rect 116894 67766 116900 67798
rect 116894 67734 116895 67766
rect 116829 67733 116895 67734
rect 952 67598 1230 67662
rect 1294 67598 1300 67662
rect 21765 67662 21831 67663
rect 21765 67630 21766 67662
rect 952 65894 1300 67598
rect 21760 67598 21766 67630
rect 21830 67630 21831 67662
rect 22576 67662 22652 67668
rect 21830 67598 21836 67630
rect 21760 67390 21836 67598
rect 21760 67326 21766 67390
rect 21830 67326 21836 67390
rect 22576 67598 22582 67662
rect 22646 67598 22652 67662
rect 22576 67390 22652 67598
rect 116552 67662 116628 67668
rect 116552 67598 116558 67662
rect 116622 67598 116628 67662
rect 116829 67662 116895 67663
rect 116829 67630 116830 67662
rect 22576 67358 22582 67390
rect 21760 67320 21836 67326
rect 22581 67326 22582 67358
rect 22646 67358 22652 67390
rect 110301 67390 110367 67391
rect 110301 67358 110302 67390
rect 22646 67326 22647 67358
rect 22581 67325 22647 67326
rect 110296 67326 110302 67358
rect 110366 67358 110367 67390
rect 116552 67390 116628 67598
rect 116552 67358 116558 67390
rect 110366 67326 110372 67358
rect 21901 67254 21967 67255
rect 21901 67222 21902 67254
rect 21896 67190 21902 67222
rect 21966 67222 21967 67254
rect 22984 67254 23060 67260
rect 21966 67190 21972 67222
rect 21896 66982 21972 67190
rect 21896 66918 21902 66982
rect 21966 66918 21972 66982
rect 22984 67190 22990 67254
rect 23054 67190 23060 67254
rect 22984 66982 23060 67190
rect 22984 66950 22990 66982
rect 21896 66912 21972 66918
rect 22989 66918 22990 66950
rect 23054 66950 23060 66982
rect 23528 67254 23604 67260
rect 23528 67190 23534 67254
rect 23598 67190 23604 67254
rect 23528 66982 23604 67190
rect 110296 67118 110372 67326
rect 116557 67326 116558 67358
rect 116622 67358 116628 67390
rect 116824 67598 116830 67630
rect 116894 67630 116895 67662
rect 116894 67598 116900 67630
rect 116824 67390 116900 67598
rect 116622 67326 116623 67358
rect 116557 67325 116623 67326
rect 116824 67326 116830 67390
rect 116894 67326 116900 67390
rect 116824 67320 116900 67326
rect 137496 67526 137844 69230
rect 137496 67462 137502 67526
rect 137566 67462 137844 67526
rect 115197 67254 115263 67255
rect 115197 67222 115198 67254
rect 110296 67054 110302 67118
rect 110366 67054 110372 67118
rect 110296 67048 110372 67054
rect 115192 67190 115198 67222
rect 115262 67222 115263 67254
rect 115605 67254 115671 67255
rect 115605 67222 115606 67254
rect 115262 67190 115268 67222
rect 23528 66950 23534 66982
rect 23054 66918 23055 66950
rect 22989 66917 23055 66918
rect 23533 66918 23534 66950
rect 23598 66950 23604 66982
rect 115192 66982 115268 67190
rect 23598 66918 23599 66950
rect 23533 66917 23599 66918
rect 115192 66918 115198 66982
rect 115262 66918 115268 66982
rect 115192 66912 115268 66918
rect 115600 67190 115606 67222
rect 115670 67222 115671 67254
rect 116965 67254 117031 67255
rect 116965 67222 116966 67254
rect 115670 67190 115676 67222
rect 115600 66982 115676 67190
rect 115600 66918 115606 66982
rect 115670 66918 115676 66982
rect 115600 66912 115676 66918
rect 116960 67190 116966 67222
rect 117030 67222 117031 67254
rect 117030 67190 117036 67222
rect 116960 66982 117036 67190
rect 116960 66918 116966 66982
rect 117030 66918 117036 66982
rect 116960 66912 117036 66918
rect 21760 66846 21836 66852
rect 21760 66782 21766 66846
rect 21830 66782 21836 66846
rect 21760 66574 21836 66782
rect 21760 66542 21766 66574
rect 21765 66510 21766 66542
rect 21830 66542 21836 66574
rect 22576 66846 22652 66852
rect 22576 66782 22582 66846
rect 22646 66782 22652 66846
rect 22989 66846 23055 66847
rect 22989 66814 22990 66846
rect 22576 66574 22652 66782
rect 22576 66542 22582 66574
rect 21830 66510 21831 66542
rect 21765 66509 21831 66510
rect 22581 66510 22582 66542
rect 22646 66542 22652 66574
rect 22984 66782 22990 66814
rect 23054 66814 23055 66846
rect 23528 66846 23604 66852
rect 23054 66782 23060 66814
rect 22984 66574 23060 66782
rect 22646 66510 22647 66542
rect 22581 66509 22647 66510
rect 22984 66510 22990 66574
rect 23054 66510 23060 66574
rect 23528 66782 23534 66846
rect 23598 66782 23604 66846
rect 115333 66846 115399 66847
rect 115333 66814 115334 66846
rect 23528 66574 23604 66782
rect 23528 66542 23534 66574
rect 22984 66504 23060 66510
rect 23533 66510 23534 66542
rect 23598 66542 23604 66574
rect 115328 66782 115334 66814
rect 115398 66814 115399 66846
rect 115741 66846 115807 66847
rect 115741 66814 115742 66846
rect 115398 66782 115404 66814
rect 115328 66574 115404 66782
rect 23598 66510 23599 66542
rect 23533 66509 23599 66510
rect 115328 66510 115334 66574
rect 115398 66510 115404 66574
rect 115328 66504 115404 66510
rect 115736 66782 115742 66814
rect 115806 66814 115807 66846
rect 116280 66846 116356 66852
rect 115806 66782 115812 66814
rect 115736 66574 115812 66782
rect 115736 66510 115742 66574
rect 115806 66510 115812 66574
rect 116280 66782 116286 66846
rect 116350 66782 116356 66846
rect 116829 66846 116895 66847
rect 116829 66814 116830 66846
rect 116280 66574 116356 66782
rect 116280 66542 116286 66574
rect 115736 66504 115812 66510
rect 116285 66510 116286 66542
rect 116350 66542 116356 66574
rect 116824 66782 116830 66814
rect 116894 66814 116895 66846
rect 116894 66782 116900 66814
rect 116824 66574 116900 66782
rect 116350 66510 116351 66542
rect 116285 66509 116351 66510
rect 116824 66510 116830 66574
rect 116894 66510 116900 66574
rect 116824 66504 116900 66510
rect 21901 66438 21967 66439
rect 21901 66406 21902 66438
rect 21896 66374 21902 66406
rect 21966 66406 21967 66438
rect 22445 66438 22511 66439
rect 22445 66406 22446 66438
rect 21966 66374 21972 66406
rect 21896 66166 21972 66374
rect 21896 66102 21902 66166
rect 21966 66102 21972 66166
rect 21896 66096 21972 66102
rect 22440 66374 22446 66406
rect 22510 66406 22511 66438
rect 23120 66438 23196 66444
rect 22510 66374 22516 66406
rect 22440 66166 22516 66374
rect 22440 66102 22446 66166
rect 22510 66102 22516 66166
rect 23120 66374 23126 66438
rect 23190 66374 23196 66438
rect 23397 66438 23463 66439
rect 23397 66406 23398 66438
rect 23120 66166 23196 66374
rect 23120 66134 23126 66166
rect 22440 66096 22516 66102
rect 23125 66102 23126 66134
rect 23190 66134 23196 66166
rect 23392 66374 23398 66406
rect 23462 66406 23463 66438
rect 115192 66438 115268 66444
rect 23462 66374 23468 66406
rect 23392 66166 23468 66374
rect 23190 66102 23191 66134
rect 23125 66101 23191 66102
rect 23392 66102 23398 66166
rect 23462 66102 23468 66166
rect 115192 66374 115198 66438
rect 115262 66374 115268 66438
rect 115192 66166 115268 66374
rect 115192 66134 115198 66166
rect 23392 66096 23468 66102
rect 115197 66102 115198 66134
rect 115262 66134 115268 66166
rect 115600 66438 115676 66444
rect 115600 66374 115606 66438
rect 115670 66374 115676 66438
rect 115600 66166 115676 66374
rect 115600 66134 115606 66166
rect 115262 66102 115263 66134
rect 115197 66101 115263 66102
rect 115605 66102 115606 66134
rect 115670 66134 115676 66166
rect 116552 66438 116628 66444
rect 116552 66374 116558 66438
rect 116622 66374 116628 66438
rect 116552 66166 116628 66374
rect 116552 66134 116558 66166
rect 115670 66102 115671 66134
rect 115605 66101 115671 66102
rect 116557 66102 116558 66134
rect 116622 66134 116628 66166
rect 116960 66438 117036 66444
rect 116960 66374 116966 66438
rect 117030 66374 117036 66438
rect 116960 66166 117036 66374
rect 116960 66134 116966 66166
rect 116622 66102 116623 66134
rect 116557 66101 116623 66102
rect 116965 66102 116966 66134
rect 117030 66134 117036 66166
rect 117030 66102 117031 66134
rect 116965 66101 117031 66102
rect 952 65830 1230 65894
rect 1294 65830 1300 65894
rect 952 64398 1300 65830
rect 21760 66030 21836 66036
rect 21760 65966 21766 66030
rect 21830 65966 21836 66030
rect 22309 66030 22375 66031
rect 22309 65998 22310 66030
rect 21760 65758 21836 65966
rect 21760 65726 21766 65758
rect 21765 65694 21766 65726
rect 21830 65726 21836 65758
rect 22304 65966 22310 65998
rect 22374 65998 22375 66030
rect 23125 66030 23191 66031
rect 23125 65998 23126 66030
rect 22374 65966 22380 65998
rect 22304 65758 22380 65966
rect 21830 65694 21831 65726
rect 21765 65693 21831 65694
rect 22304 65694 22310 65758
rect 22374 65694 22380 65758
rect 22304 65688 22380 65694
rect 23120 65966 23126 65998
rect 23190 65998 23191 66030
rect 23528 66030 23604 66036
rect 23190 65966 23196 65998
rect 23120 65758 23196 65966
rect 23120 65694 23126 65758
rect 23190 65694 23196 65758
rect 23528 65966 23534 66030
rect 23598 65966 23604 66030
rect 115197 66030 115263 66031
rect 115197 65998 115198 66030
rect 23528 65758 23604 65966
rect 23528 65726 23534 65758
rect 23120 65688 23196 65694
rect 23533 65694 23534 65726
rect 23598 65726 23604 65758
rect 115192 65966 115198 65998
rect 115262 65998 115263 66030
rect 115605 66030 115671 66031
rect 115605 65998 115606 66030
rect 115262 65966 115268 65998
rect 115192 65758 115268 65966
rect 23598 65694 23599 65726
rect 23533 65693 23599 65694
rect 115192 65694 115198 65758
rect 115262 65694 115268 65758
rect 115192 65688 115268 65694
rect 115600 65966 115606 65998
rect 115670 65998 115671 66030
rect 116149 66030 116215 66031
rect 116149 65998 116150 66030
rect 115670 65966 115676 65998
rect 115600 65758 115676 65966
rect 115600 65694 115606 65758
rect 115670 65694 115676 65758
rect 115600 65688 115676 65694
rect 116144 65966 116150 65998
rect 116214 65998 116215 66030
rect 116416 66030 116492 66036
rect 116214 65966 116220 65998
rect 116144 65758 116220 65966
rect 116144 65694 116150 65758
rect 116214 65694 116220 65758
rect 116416 65966 116422 66030
rect 116486 65966 116492 66030
rect 116416 65758 116492 65966
rect 116416 65726 116422 65758
rect 116144 65688 116220 65694
rect 116421 65694 116422 65726
rect 116486 65726 116492 65758
rect 116824 66030 116900 66036
rect 116824 65966 116830 66030
rect 116894 65966 116900 66030
rect 116824 65758 116900 65966
rect 116824 65726 116830 65758
rect 116486 65694 116487 65726
rect 116421 65693 116487 65694
rect 116829 65694 116830 65726
rect 116894 65726 116900 65758
rect 137496 66030 137844 67462
rect 137496 65966 137502 66030
rect 137566 65966 137844 66030
rect 116894 65694 116895 65726
rect 116829 65693 116895 65694
rect 21896 65622 21972 65628
rect 21896 65558 21902 65622
rect 21966 65558 21972 65622
rect 22581 65622 22647 65623
rect 22581 65590 22582 65622
rect 21896 65350 21972 65558
rect 21896 65318 21902 65350
rect 21901 65286 21902 65318
rect 21966 65318 21972 65350
rect 22576 65558 22582 65590
rect 22646 65590 22647 65622
rect 22989 65622 23055 65623
rect 22989 65590 22990 65622
rect 22646 65558 22652 65590
rect 22576 65350 22652 65558
rect 21966 65286 21967 65318
rect 21901 65285 21967 65286
rect 22576 65286 22582 65350
rect 22646 65286 22652 65350
rect 22576 65280 22652 65286
rect 22984 65558 22990 65590
rect 23054 65590 23055 65622
rect 23533 65622 23599 65623
rect 23533 65590 23534 65622
rect 23054 65558 23060 65590
rect 22984 65350 23060 65558
rect 22984 65286 22990 65350
rect 23054 65286 23060 65350
rect 22984 65280 23060 65286
rect 23528 65558 23534 65590
rect 23598 65590 23599 65622
rect 115192 65622 115268 65628
rect 23598 65558 23604 65590
rect 23528 65350 23604 65558
rect 23528 65286 23534 65350
rect 23598 65286 23604 65350
rect 115192 65558 115198 65622
rect 115262 65558 115268 65622
rect 115192 65350 115268 65558
rect 115192 65318 115198 65350
rect 23528 65280 23604 65286
rect 115197 65286 115198 65318
rect 115262 65318 115268 65350
rect 115600 65622 115676 65628
rect 115600 65558 115606 65622
rect 115670 65558 115676 65622
rect 115600 65350 115676 65558
rect 115600 65318 115606 65350
rect 115262 65286 115263 65318
rect 115197 65285 115263 65286
rect 115605 65286 115606 65318
rect 115670 65318 115676 65350
rect 116008 65622 116084 65628
rect 116008 65558 116014 65622
rect 116078 65558 116084 65622
rect 116829 65622 116895 65623
rect 116829 65590 116830 65622
rect 116008 65350 116084 65558
rect 116008 65318 116014 65350
rect 115670 65286 115671 65318
rect 115605 65285 115671 65286
rect 116013 65286 116014 65318
rect 116078 65318 116084 65350
rect 116824 65558 116830 65590
rect 116894 65590 116895 65622
rect 116894 65558 116900 65590
rect 116824 65350 116900 65558
rect 116078 65286 116079 65318
rect 116013 65285 116079 65286
rect 116824 65286 116830 65350
rect 116894 65286 116900 65350
rect 116824 65280 116900 65286
rect 22309 65214 22375 65215
rect 22309 65182 22310 65214
rect 22304 65150 22310 65182
rect 22374 65182 22375 65214
rect 22445 65214 22511 65215
rect 22445 65182 22446 65214
rect 22374 65150 22380 65182
rect 22304 64942 22380 65150
rect 22304 64878 22310 64942
rect 22374 64878 22380 64942
rect 22304 64872 22380 64878
rect 22440 65150 22446 65182
rect 22510 65182 22511 65214
rect 23120 65214 23196 65220
rect 22510 65150 22516 65182
rect 22440 64942 22516 65150
rect 22440 64878 22446 64942
rect 22510 64878 22516 64942
rect 23120 65150 23126 65214
rect 23190 65150 23196 65214
rect 23120 64942 23196 65150
rect 23120 64910 23126 64942
rect 22440 64872 22516 64878
rect 23125 64878 23126 64910
rect 23190 64910 23196 64942
rect 23392 65214 23468 65220
rect 23392 65150 23398 65214
rect 23462 65150 23468 65214
rect 115197 65214 115263 65215
rect 115197 65182 115198 65214
rect 23392 64942 23468 65150
rect 23392 64910 23398 64942
rect 23190 64878 23191 64910
rect 23125 64877 23191 64878
rect 23397 64878 23398 64910
rect 23462 64910 23468 64942
rect 115192 65150 115198 65182
rect 115262 65182 115263 65214
rect 115600 65214 115676 65220
rect 115262 65150 115268 65182
rect 115192 64942 115268 65150
rect 23462 64878 23463 64910
rect 23397 64877 23463 64878
rect 115192 64878 115198 64942
rect 115262 64878 115268 64942
rect 115600 65150 115606 65214
rect 115670 65150 115676 65214
rect 115600 64942 115676 65150
rect 115600 64910 115606 64942
rect 115192 64872 115268 64878
rect 115605 64878 115606 64910
rect 115670 64910 115676 64942
rect 116144 65214 116220 65220
rect 116144 65150 116150 65214
rect 116214 65150 116220 65214
rect 116144 64942 116220 65150
rect 116144 64910 116150 64942
rect 115670 64878 115671 64910
rect 115605 64877 115671 64878
rect 116149 64878 116150 64910
rect 116214 64910 116220 64942
rect 116214 64878 116215 64910
rect 116149 64877 116215 64878
rect 22989 64806 23055 64807
rect 22989 64774 22990 64806
rect 22984 64742 22990 64774
rect 23054 64774 23055 64806
rect 23533 64806 23599 64807
rect 23533 64774 23534 64806
rect 23054 64742 23060 64774
rect 22984 64534 23060 64742
rect 22984 64470 22990 64534
rect 23054 64470 23060 64534
rect 22984 64464 23060 64470
rect 23528 64742 23534 64774
rect 23598 64774 23599 64806
rect 115328 64806 115404 64812
rect 23598 64742 23604 64774
rect 23528 64534 23604 64742
rect 23528 64470 23534 64534
rect 23598 64470 23604 64534
rect 115328 64742 115334 64806
rect 115398 64742 115404 64806
rect 115741 64806 115807 64807
rect 115741 64774 115742 64806
rect 115328 64534 115404 64742
rect 115328 64502 115334 64534
rect 23528 64464 23604 64470
rect 115333 64470 115334 64502
rect 115398 64502 115404 64534
rect 115736 64742 115742 64774
rect 115806 64774 115807 64806
rect 115806 64742 115812 64774
rect 115736 64534 115812 64742
rect 115398 64470 115399 64502
rect 115333 64469 115399 64470
rect 115736 64470 115742 64534
rect 115806 64470 115812 64534
rect 115736 64464 115812 64470
rect 952 64334 1230 64398
rect 1294 64334 1300 64398
rect 22173 64398 22239 64399
rect 22173 64366 22174 64398
rect 952 62630 1300 64334
rect 22168 64334 22174 64366
rect 22238 64366 22239 64398
rect 22581 64398 22647 64399
rect 22581 64366 22582 64398
rect 22238 64334 22244 64366
rect 21896 64126 21972 64132
rect 21896 64062 21902 64126
rect 21966 64062 21972 64126
rect 21896 63854 21972 64062
rect 22168 64126 22244 64334
rect 22168 64062 22174 64126
rect 22238 64062 22244 64126
rect 22168 64056 22244 64062
rect 22576 64334 22582 64366
rect 22646 64366 22647 64398
rect 116008 64398 116084 64404
rect 22646 64334 22652 64366
rect 22576 64126 22652 64334
rect 116008 64334 116014 64398
rect 116078 64334 116084 64398
rect 110165 64262 110231 64263
rect 110165 64230 110166 64262
rect 22576 64062 22582 64126
rect 22646 64062 22652 64126
rect 22576 64056 22652 64062
rect 110160 64198 110166 64230
rect 110230 64230 110231 64262
rect 110230 64198 110236 64230
rect 110160 63990 110236 64198
rect 116008 64126 116084 64334
rect 116008 64094 116014 64126
rect 116013 64062 116014 64094
rect 116078 64094 116084 64126
rect 116552 64398 116628 64404
rect 116552 64334 116558 64398
rect 116622 64334 116628 64398
rect 116552 64126 116628 64334
rect 137496 64262 137844 65966
rect 137496 64198 137502 64262
rect 137566 64198 137844 64262
rect 116552 64094 116558 64126
rect 116078 64062 116079 64094
rect 116013 64061 116079 64062
rect 116557 64062 116558 64094
rect 116622 64094 116628 64126
rect 116824 64126 116900 64132
rect 116622 64062 116623 64094
rect 116557 64061 116623 64062
rect 116824 64062 116830 64126
rect 116894 64062 116900 64126
rect 110160 63926 110166 63990
rect 110230 63926 110236 63990
rect 110160 63920 110236 63926
rect 21896 63822 21902 63854
rect 21901 63790 21902 63822
rect 21966 63822 21972 63854
rect 28560 63854 28636 63860
rect 21966 63790 21967 63822
rect 21901 63789 21967 63790
rect 28560 63790 28566 63854
rect 28630 63790 28636 63854
rect 21765 63718 21831 63719
rect 21765 63686 21766 63718
rect 21760 63654 21766 63686
rect 21830 63686 21831 63718
rect 22309 63718 22375 63719
rect 22309 63686 22310 63718
rect 21830 63654 21836 63686
rect 21760 63446 21836 63654
rect 21760 63382 21766 63446
rect 21830 63382 21836 63446
rect 21760 63376 21836 63382
rect 22304 63654 22310 63686
rect 22374 63686 22375 63718
rect 22374 63654 22380 63686
rect 22304 63446 22380 63654
rect 28560 63582 28636 63790
rect 28560 63550 28566 63582
rect 28565 63518 28566 63550
rect 28630 63550 28636 63582
rect 110432 63854 110508 63860
rect 110432 63790 110438 63854
rect 110502 63790 110508 63854
rect 116824 63854 116900 64062
rect 116824 63822 116830 63854
rect 110432 63582 110508 63790
rect 116829 63790 116830 63822
rect 116894 63822 116900 63854
rect 116894 63790 116895 63822
rect 116829 63789 116895 63790
rect 110432 63550 110438 63582
rect 28630 63518 28631 63550
rect 28565 63517 28631 63518
rect 110437 63518 110438 63550
rect 110502 63550 110508 63582
rect 116280 63718 116356 63724
rect 116280 63654 116286 63718
rect 116350 63654 116356 63718
rect 110502 63518 110503 63550
rect 110437 63517 110503 63518
rect 22304 63382 22310 63446
rect 22374 63382 22380 63446
rect 28293 63446 28359 63447
rect 28293 63414 28294 63446
rect 22304 63376 22380 63382
rect 28288 63382 28294 63414
rect 28358 63414 28359 63446
rect 116280 63446 116356 63654
rect 116280 63414 116286 63446
rect 28358 63382 28364 63414
rect 21896 63310 21972 63316
rect 21896 63246 21902 63310
rect 21966 63246 21972 63310
rect 23125 63310 23191 63311
rect 23125 63278 23126 63310
rect 21896 63038 21972 63246
rect 21896 63006 21902 63038
rect 21901 62974 21902 63006
rect 21966 63006 21972 63038
rect 23120 63246 23126 63278
rect 23190 63278 23191 63310
rect 23392 63310 23468 63316
rect 23190 63246 23196 63278
rect 23120 63038 23196 63246
rect 21966 62974 21967 63006
rect 21901 62973 21967 62974
rect 23120 62974 23126 63038
rect 23190 62974 23196 63038
rect 23392 63246 23398 63310
rect 23462 63246 23468 63310
rect 23392 63038 23468 63246
rect 28288 63174 28364 63382
rect 116285 63382 116286 63414
rect 116350 63414 116356 63446
rect 116824 63718 116900 63724
rect 116824 63654 116830 63718
rect 116894 63654 116900 63718
rect 116824 63446 116900 63654
rect 116824 63414 116830 63446
rect 116350 63382 116351 63414
rect 116285 63381 116351 63382
rect 116829 63382 116830 63414
rect 116894 63414 116900 63446
rect 116894 63382 116895 63414
rect 116829 63381 116895 63382
rect 28288 63110 28294 63174
rect 28358 63110 28364 63174
rect 28288 63104 28364 63110
rect 115192 63310 115268 63316
rect 115192 63246 115198 63310
rect 115262 63246 115268 63310
rect 23392 63006 23398 63038
rect 23120 62968 23196 62974
rect 23397 62974 23398 63006
rect 23462 63006 23468 63038
rect 115192 63038 115268 63246
rect 115192 63006 115198 63038
rect 23462 62974 23463 63006
rect 23397 62973 23463 62974
rect 115197 62974 115198 63006
rect 115262 63006 115268 63038
rect 115600 63310 115676 63316
rect 115600 63246 115606 63310
rect 115670 63246 115676 63310
rect 115600 63038 115676 63246
rect 115600 63006 115606 63038
rect 115262 62974 115263 63006
rect 115197 62973 115263 62974
rect 115605 62974 115606 63006
rect 115670 63006 115676 63038
rect 116960 63310 117036 63316
rect 116960 63246 116966 63310
rect 117030 63246 117036 63310
rect 116960 63038 117036 63246
rect 116960 63006 116966 63038
rect 115670 62974 115671 63006
rect 115605 62973 115671 62974
rect 116965 62974 116966 63006
rect 117030 63006 117036 63038
rect 117030 62974 117031 63006
rect 116965 62973 117031 62974
rect 952 62566 1230 62630
rect 1294 62566 1300 62630
rect 21760 62902 21836 62908
rect 21760 62838 21766 62902
rect 21830 62838 21836 62902
rect 21760 62630 21836 62838
rect 21760 62598 21766 62630
rect 952 60998 1300 62566
rect 21765 62566 21766 62598
rect 21830 62598 21836 62630
rect 22576 62902 22652 62908
rect 22576 62838 22582 62902
rect 22646 62838 22652 62902
rect 22576 62630 22652 62838
rect 22576 62598 22582 62630
rect 21830 62566 21831 62598
rect 21765 62565 21831 62566
rect 22581 62566 22582 62598
rect 22646 62598 22652 62630
rect 22984 62902 23060 62908
rect 22984 62838 22990 62902
rect 23054 62838 23060 62902
rect 23397 62902 23463 62903
rect 23397 62870 23398 62902
rect 22984 62630 23060 62838
rect 22984 62598 22990 62630
rect 22646 62566 22647 62598
rect 22581 62565 22647 62566
rect 22989 62566 22990 62598
rect 23054 62598 23060 62630
rect 23392 62838 23398 62870
rect 23462 62870 23463 62902
rect 115197 62902 115263 62903
rect 115197 62870 115198 62902
rect 23462 62838 23468 62870
rect 23392 62630 23468 62838
rect 115192 62838 115198 62870
rect 115262 62870 115263 62902
rect 115605 62902 115671 62903
rect 115605 62870 115606 62902
rect 115262 62838 115268 62870
rect 23054 62566 23055 62598
rect 22989 62565 23055 62566
rect 23392 62566 23398 62630
rect 23462 62566 23468 62630
rect 23392 62560 23468 62566
rect 110160 62630 110236 62636
rect 110160 62566 110166 62630
rect 110230 62566 110236 62630
rect 21760 62494 21836 62500
rect 21760 62430 21766 62494
rect 21830 62430 21836 62494
rect 21760 62222 21836 62430
rect 21760 62190 21766 62222
rect 21765 62158 21766 62190
rect 21830 62190 21836 62222
rect 22168 62494 22244 62500
rect 22168 62430 22174 62494
rect 22238 62430 22244 62494
rect 22989 62494 23055 62495
rect 22989 62462 22990 62494
rect 22168 62222 22244 62430
rect 22168 62190 22174 62222
rect 21830 62158 21831 62190
rect 21765 62157 21831 62158
rect 22173 62158 22174 62190
rect 22238 62190 22244 62222
rect 22984 62430 22990 62462
rect 23054 62462 23055 62494
rect 23533 62494 23599 62495
rect 23533 62462 23534 62494
rect 23054 62430 23060 62462
rect 22984 62222 23060 62430
rect 22238 62158 22239 62190
rect 22173 62157 22239 62158
rect 22984 62158 22990 62222
rect 23054 62158 23060 62222
rect 22984 62152 23060 62158
rect 23528 62430 23534 62462
rect 23598 62462 23599 62494
rect 23598 62430 23604 62462
rect 23528 62222 23604 62430
rect 110160 62358 110236 62566
rect 115192 62630 115268 62838
rect 115192 62566 115198 62630
rect 115262 62566 115268 62630
rect 115192 62560 115268 62566
rect 115600 62838 115606 62870
rect 115670 62870 115671 62902
rect 116149 62902 116215 62903
rect 116149 62870 116150 62902
rect 115670 62838 115676 62870
rect 115600 62630 115676 62838
rect 115600 62566 115606 62630
rect 115670 62566 115676 62630
rect 115600 62560 115676 62566
rect 116144 62838 116150 62870
rect 116214 62870 116215 62902
rect 116285 62902 116351 62903
rect 116285 62870 116286 62902
rect 116214 62838 116220 62870
rect 116144 62630 116220 62838
rect 116144 62566 116150 62630
rect 116214 62566 116220 62630
rect 116144 62560 116220 62566
rect 116280 62838 116286 62870
rect 116350 62870 116351 62902
rect 116965 62902 117031 62903
rect 116965 62870 116966 62902
rect 116350 62838 116356 62870
rect 116280 62630 116356 62838
rect 116280 62566 116286 62630
rect 116350 62566 116356 62630
rect 116280 62560 116356 62566
rect 116960 62838 116966 62870
rect 117030 62870 117031 62902
rect 117030 62838 117036 62870
rect 116960 62630 117036 62838
rect 116960 62566 116966 62630
rect 117030 62566 117036 62630
rect 116960 62560 117036 62566
rect 137496 62630 137844 64198
rect 137496 62566 137502 62630
rect 137566 62566 137844 62630
rect 115333 62494 115399 62495
rect 115333 62462 115334 62494
rect 110160 62326 110166 62358
rect 110165 62294 110166 62326
rect 110230 62326 110236 62358
rect 115328 62430 115334 62462
rect 115398 62462 115399 62494
rect 115736 62494 115812 62500
rect 115398 62430 115404 62462
rect 110230 62294 110231 62326
rect 110165 62293 110231 62294
rect 23528 62158 23534 62222
rect 23598 62158 23604 62222
rect 23528 62152 23604 62158
rect 115328 62222 115404 62430
rect 115328 62158 115334 62222
rect 115398 62158 115404 62222
rect 115736 62430 115742 62494
rect 115806 62430 115812 62494
rect 116421 62494 116487 62495
rect 116421 62462 116422 62494
rect 115736 62222 115812 62430
rect 115736 62190 115742 62222
rect 115328 62152 115404 62158
rect 115741 62158 115742 62190
rect 115806 62190 115812 62222
rect 116416 62430 116422 62462
rect 116486 62462 116487 62494
rect 116824 62494 116900 62500
rect 116486 62430 116492 62462
rect 116416 62222 116492 62430
rect 115806 62158 115807 62190
rect 115741 62157 115807 62158
rect 116416 62158 116422 62222
rect 116486 62158 116492 62222
rect 116824 62430 116830 62494
rect 116894 62430 116900 62494
rect 116824 62222 116900 62430
rect 116824 62190 116830 62222
rect 116416 62152 116492 62158
rect 116829 62158 116830 62190
rect 116894 62190 116900 62222
rect 116894 62158 116895 62190
rect 116829 62157 116895 62158
rect 21901 62086 21967 62087
rect 21901 62054 21902 62086
rect 21896 62022 21902 62054
rect 21966 62054 21967 62086
rect 22445 62086 22511 62087
rect 22445 62054 22446 62086
rect 21966 62022 21972 62054
rect 21896 61814 21972 62022
rect 21896 61750 21902 61814
rect 21966 61750 21972 61814
rect 21896 61744 21972 61750
rect 22440 62022 22446 62054
rect 22510 62054 22511 62086
rect 22989 62086 23055 62087
rect 22989 62054 22990 62086
rect 22510 62022 22516 62054
rect 22440 61814 22516 62022
rect 22440 61750 22446 61814
rect 22510 61750 22516 61814
rect 22440 61744 22516 61750
rect 22984 62022 22990 62054
rect 23054 62054 23055 62086
rect 23397 62086 23463 62087
rect 23397 62054 23398 62086
rect 23054 62022 23060 62054
rect 22984 61814 23060 62022
rect 22984 61750 22990 61814
rect 23054 61750 23060 61814
rect 22984 61744 23060 61750
rect 23392 62022 23398 62054
rect 23462 62054 23463 62086
rect 115197 62086 115263 62087
rect 115197 62054 115198 62086
rect 23462 62022 23468 62054
rect 23392 61814 23468 62022
rect 23392 61750 23398 61814
rect 23462 61750 23468 61814
rect 23392 61744 23468 61750
rect 115192 62022 115198 62054
rect 115262 62054 115263 62086
rect 115605 62086 115671 62087
rect 115605 62054 115606 62086
rect 115262 62022 115268 62054
rect 115192 61814 115268 62022
rect 115192 61750 115198 61814
rect 115262 61750 115268 61814
rect 115192 61744 115268 61750
rect 115600 62022 115606 62054
rect 115670 62054 115671 62086
rect 116552 62086 116628 62092
rect 115670 62022 115676 62054
rect 115600 61814 115676 62022
rect 115600 61750 115606 61814
rect 115670 61750 115676 61814
rect 116552 62022 116558 62086
rect 116622 62022 116628 62086
rect 116965 62086 117031 62087
rect 116965 62054 116966 62086
rect 116552 61814 116628 62022
rect 116552 61782 116558 61814
rect 115600 61744 115676 61750
rect 116557 61750 116558 61782
rect 116622 61782 116628 61814
rect 116960 62022 116966 62054
rect 117030 62054 117031 62086
rect 117030 62022 117036 62054
rect 116960 61814 117036 62022
rect 116622 61750 116623 61782
rect 116557 61749 116623 61750
rect 116960 61750 116966 61814
rect 117030 61750 117036 61814
rect 116960 61744 117036 61750
rect 21901 61678 21967 61679
rect 21901 61646 21902 61678
rect 21896 61614 21902 61646
rect 21966 61646 21967 61678
rect 22309 61678 22375 61679
rect 22309 61646 22310 61678
rect 21966 61614 21972 61646
rect 21896 61406 21972 61614
rect 21896 61342 21902 61406
rect 21966 61342 21972 61406
rect 21896 61336 21972 61342
rect 22304 61614 22310 61646
rect 22374 61646 22375 61678
rect 22445 61678 22511 61679
rect 22445 61646 22446 61678
rect 22374 61614 22380 61646
rect 22304 61406 22380 61614
rect 22304 61342 22310 61406
rect 22374 61342 22380 61406
rect 22304 61336 22380 61342
rect 22440 61614 22446 61646
rect 22510 61646 22511 61678
rect 22984 61678 23060 61684
rect 22510 61614 22516 61646
rect 22440 61406 22516 61614
rect 22440 61342 22446 61406
rect 22510 61342 22516 61406
rect 22984 61614 22990 61678
rect 23054 61614 23060 61678
rect 22984 61406 23060 61614
rect 22984 61374 22990 61406
rect 22440 61336 22516 61342
rect 22989 61342 22990 61374
rect 23054 61374 23060 61406
rect 23528 61678 23604 61684
rect 23528 61614 23534 61678
rect 23598 61614 23604 61678
rect 23528 61406 23604 61614
rect 23528 61374 23534 61406
rect 23054 61342 23055 61374
rect 22989 61341 23055 61342
rect 23533 61342 23534 61374
rect 23598 61374 23604 61406
rect 115328 61678 115404 61684
rect 115328 61614 115334 61678
rect 115398 61614 115404 61678
rect 115328 61406 115404 61614
rect 115328 61374 115334 61406
rect 23598 61342 23599 61374
rect 23533 61341 23599 61342
rect 115333 61342 115334 61374
rect 115398 61374 115404 61406
rect 115736 61678 115812 61684
rect 115736 61614 115742 61678
rect 115806 61614 115812 61678
rect 116149 61678 116215 61679
rect 116149 61646 116150 61678
rect 115736 61406 115812 61614
rect 115736 61374 115742 61406
rect 115398 61342 115399 61374
rect 115333 61341 115399 61342
rect 115741 61342 115742 61374
rect 115806 61374 115812 61406
rect 116144 61614 116150 61646
rect 116214 61646 116215 61678
rect 116824 61678 116900 61684
rect 116214 61614 116220 61646
rect 116144 61406 116220 61614
rect 115806 61342 115807 61374
rect 115741 61341 115807 61342
rect 116144 61342 116150 61406
rect 116214 61342 116220 61406
rect 116824 61614 116830 61678
rect 116894 61614 116900 61678
rect 116824 61406 116900 61614
rect 116824 61374 116830 61406
rect 116144 61336 116220 61342
rect 116829 61342 116830 61374
rect 116894 61374 116900 61406
rect 116894 61342 116895 61374
rect 116829 61341 116895 61342
rect 22712 61270 22788 61276
rect 22712 61206 22718 61270
rect 22782 61206 22788 61270
rect 952 60934 1230 60998
rect 1294 60934 1300 60998
rect 22445 60998 22511 60999
rect 22445 60966 22446 60998
rect 952 59230 1300 60934
rect 22440 60934 22446 60966
rect 22510 60966 22511 60998
rect 22712 60998 22788 61206
rect 22712 60966 22718 60998
rect 22510 60934 22516 60966
rect 22440 60726 22516 60934
rect 22717 60934 22718 60966
rect 22782 60966 22788 60998
rect 22984 61270 23060 61276
rect 22984 61206 22990 61270
rect 23054 61206 23060 61270
rect 23533 61270 23599 61271
rect 23533 61238 23534 61270
rect 22984 60998 23060 61206
rect 22984 60966 22990 60998
rect 22782 60934 22783 60966
rect 22717 60933 22783 60934
rect 22989 60934 22990 60966
rect 23054 60966 23060 60998
rect 23528 61206 23534 61238
rect 23598 61238 23599 61270
rect 115192 61270 115268 61276
rect 23598 61206 23604 61238
rect 23528 60998 23604 61206
rect 115192 61206 115198 61270
rect 115262 61206 115268 61270
rect 115741 61270 115807 61271
rect 115741 61238 115742 61270
rect 23054 60934 23055 60966
rect 22989 60933 23055 60934
rect 23528 60934 23534 60998
rect 23598 60934 23604 60998
rect 23528 60928 23604 60934
rect 110432 61134 110508 61140
rect 110432 61070 110438 61134
rect 110502 61070 110508 61134
rect 22440 60662 22446 60726
rect 22510 60662 22516 60726
rect 22440 60656 22516 60662
rect 23120 60862 23196 60868
rect 23120 60798 23126 60862
rect 23190 60798 23196 60862
rect 23120 60590 23196 60798
rect 23120 60558 23126 60590
rect 23125 60526 23126 60558
rect 23190 60558 23196 60590
rect 23392 60862 23468 60868
rect 23392 60798 23398 60862
rect 23462 60798 23468 60862
rect 110432 60862 110508 61070
rect 115192 60998 115268 61206
rect 115192 60966 115198 60998
rect 115197 60934 115198 60966
rect 115262 60966 115268 60998
rect 115736 61206 115742 61238
rect 115806 61238 115807 61270
rect 116013 61270 116079 61271
rect 116013 61238 116014 61270
rect 115806 61206 115812 61238
rect 115736 60998 115812 61206
rect 115262 60934 115263 60966
rect 115197 60933 115263 60934
rect 115736 60934 115742 60998
rect 115806 60934 115812 60998
rect 115736 60928 115812 60934
rect 116008 61206 116014 61238
rect 116078 61238 116079 61270
rect 116552 61270 116628 61276
rect 116078 61206 116084 61238
rect 116008 60998 116084 61206
rect 116008 60934 116014 60998
rect 116078 60934 116084 60998
rect 116552 61206 116558 61270
rect 116622 61206 116628 61270
rect 116552 60998 116628 61206
rect 116552 60966 116558 60998
rect 116008 60928 116084 60934
rect 116557 60934 116558 60966
rect 116622 60966 116628 60998
rect 137496 60998 137844 62566
rect 116622 60934 116623 60966
rect 116557 60933 116623 60934
rect 137496 60934 137502 60998
rect 137566 60934 137844 60998
rect 110432 60830 110438 60862
rect 23392 60590 23468 60798
rect 110437 60798 110438 60830
rect 110502 60830 110508 60862
rect 115197 60862 115263 60863
rect 115197 60830 115198 60862
rect 110502 60798 110503 60830
rect 110437 60797 110503 60798
rect 115192 60798 115198 60830
rect 115262 60830 115263 60862
rect 115600 60862 115676 60868
rect 115262 60798 115268 60830
rect 23392 60558 23398 60590
rect 23190 60526 23191 60558
rect 23125 60525 23191 60526
rect 23397 60526 23398 60558
rect 23462 60558 23468 60590
rect 115192 60590 115268 60798
rect 23462 60526 23463 60558
rect 23397 60525 23463 60526
rect 115192 60526 115198 60590
rect 115262 60526 115268 60590
rect 115600 60798 115606 60862
rect 115670 60798 115676 60862
rect 115600 60590 115676 60798
rect 115600 60558 115606 60590
rect 115192 60520 115268 60526
rect 115605 60526 115606 60558
rect 115670 60558 115676 60590
rect 115670 60526 115671 60558
rect 115605 60525 115671 60526
rect 22168 60454 22244 60460
rect 22168 60390 22174 60454
rect 22238 60390 22244 60454
rect 21896 60182 21972 60188
rect 21896 60118 21902 60182
rect 21966 60118 21972 60182
rect 22168 60182 22244 60390
rect 22168 60150 22174 60182
rect 21896 59910 21972 60118
rect 22173 60118 22174 60150
rect 22238 60150 22244 60182
rect 23120 60454 23196 60460
rect 23120 60390 23126 60454
rect 23190 60390 23196 60454
rect 23533 60454 23599 60455
rect 23533 60422 23534 60454
rect 23120 60182 23196 60390
rect 23120 60150 23126 60182
rect 22238 60118 22239 60150
rect 22173 60117 22239 60118
rect 23125 60118 23126 60150
rect 23190 60150 23196 60182
rect 23528 60390 23534 60422
rect 23598 60422 23599 60454
rect 115328 60454 115404 60460
rect 23598 60390 23604 60422
rect 23528 60182 23604 60390
rect 115328 60390 115334 60454
rect 115398 60390 115404 60454
rect 23190 60118 23191 60150
rect 23125 60117 23191 60118
rect 23528 60118 23534 60182
rect 23598 60118 23604 60182
rect 23528 60112 23604 60118
rect 28560 60318 28636 60324
rect 28560 60254 28566 60318
rect 28630 60254 28636 60318
rect 28293 60046 28359 60047
rect 28293 60014 28294 60046
rect 21896 59878 21902 59910
rect 21901 59846 21902 59878
rect 21966 59878 21972 59910
rect 28288 59982 28294 60014
rect 28358 60014 28359 60046
rect 28560 60046 28636 60254
rect 115328 60182 115404 60390
rect 115328 60150 115334 60182
rect 115333 60118 115334 60150
rect 115398 60150 115404 60182
rect 115736 60454 115812 60460
rect 115736 60390 115742 60454
rect 115806 60390 115812 60454
rect 116013 60454 116079 60455
rect 116013 60422 116014 60454
rect 115736 60182 115812 60390
rect 115736 60150 115742 60182
rect 115398 60118 115399 60150
rect 115333 60117 115399 60118
rect 115741 60118 115742 60150
rect 115806 60150 115812 60182
rect 116008 60390 116014 60422
rect 116078 60422 116079 60454
rect 116421 60454 116487 60455
rect 116421 60422 116422 60454
rect 116078 60390 116084 60422
rect 116008 60182 116084 60390
rect 115806 60118 115807 60150
rect 115741 60117 115807 60118
rect 116008 60118 116014 60182
rect 116078 60118 116084 60182
rect 116008 60112 116084 60118
rect 116416 60390 116422 60422
rect 116486 60422 116487 60454
rect 116486 60390 116492 60422
rect 116416 60182 116492 60390
rect 116416 60118 116422 60182
rect 116486 60118 116492 60182
rect 116829 60182 116895 60183
rect 116829 60150 116830 60182
rect 116416 60112 116492 60118
rect 116824 60118 116830 60150
rect 116894 60150 116895 60182
rect 116894 60118 116900 60150
rect 28560 60014 28566 60046
rect 28358 59982 28364 60014
rect 21966 59846 21967 59878
rect 21901 59845 21967 59846
rect 21901 59774 21967 59775
rect 21901 59742 21902 59774
rect 21896 59710 21902 59742
rect 21966 59742 21967 59774
rect 22309 59774 22375 59775
rect 22309 59742 22310 59774
rect 21966 59710 21972 59742
rect 21896 59502 21972 59710
rect 21896 59438 21902 59502
rect 21966 59438 21972 59502
rect 21896 59432 21972 59438
rect 22304 59710 22310 59742
rect 22374 59742 22375 59774
rect 22374 59710 22380 59742
rect 22304 59502 22380 59710
rect 28288 59638 28364 59982
rect 28565 59982 28566 60014
rect 28630 60014 28636 60046
rect 28630 59982 28631 60014
rect 28565 59981 28631 59982
rect 110165 59910 110231 59911
rect 110165 59878 110166 59910
rect 28288 59574 28294 59638
rect 28358 59574 28364 59638
rect 28288 59568 28364 59574
rect 110160 59846 110166 59878
rect 110230 59878 110231 59910
rect 116824 59910 116900 60118
rect 110230 59846 110236 59878
rect 110160 59638 110236 59846
rect 116824 59846 116830 59910
rect 116894 59846 116900 59910
rect 116824 59840 116900 59846
rect 116557 59774 116623 59775
rect 116557 59742 116558 59774
rect 110160 59574 110166 59638
rect 110230 59574 110236 59638
rect 110160 59568 110236 59574
rect 116552 59710 116558 59742
rect 116622 59742 116623 59774
rect 116960 59774 117036 59780
rect 116622 59710 116628 59742
rect 22304 59438 22310 59502
rect 22374 59438 22380 59502
rect 22304 59432 22380 59438
rect 110432 59502 110508 59508
rect 110432 59438 110438 59502
rect 110502 59438 110508 59502
rect 21765 59366 21831 59367
rect 21765 59334 21766 59366
rect 952 59166 1230 59230
rect 1294 59166 1300 59230
rect 952 57462 1300 59166
rect 21760 59302 21766 59334
rect 21830 59334 21831 59366
rect 22989 59366 23055 59367
rect 22989 59334 22990 59366
rect 21830 59302 21836 59334
rect 21760 59094 21836 59302
rect 21760 59030 21766 59094
rect 21830 59030 21836 59094
rect 21760 59024 21836 59030
rect 22984 59302 22990 59334
rect 23054 59334 23055 59366
rect 23533 59366 23599 59367
rect 23533 59334 23534 59366
rect 23054 59302 23060 59334
rect 22984 59094 23060 59302
rect 22984 59030 22990 59094
rect 23054 59030 23060 59094
rect 22984 59024 23060 59030
rect 23528 59302 23534 59334
rect 23598 59334 23599 59366
rect 23598 59302 23604 59334
rect 23528 59094 23604 59302
rect 110432 59230 110508 59438
rect 116552 59502 116628 59710
rect 116552 59438 116558 59502
rect 116622 59438 116628 59502
rect 116960 59710 116966 59774
rect 117030 59710 117036 59774
rect 116960 59502 117036 59710
rect 116960 59470 116966 59502
rect 116552 59432 116628 59438
rect 116965 59438 116966 59470
rect 117030 59470 117036 59502
rect 117030 59438 117031 59470
rect 116965 59437 117031 59438
rect 110432 59198 110438 59230
rect 110437 59166 110438 59198
rect 110502 59198 110508 59230
rect 115328 59366 115404 59372
rect 115328 59302 115334 59366
rect 115398 59302 115404 59366
rect 110502 59166 110503 59198
rect 110437 59165 110503 59166
rect 23528 59030 23534 59094
rect 23598 59030 23604 59094
rect 115328 59094 115404 59302
rect 115328 59062 115334 59094
rect 23528 59024 23604 59030
rect 115333 59030 115334 59062
rect 115398 59062 115404 59094
rect 115736 59366 115812 59372
rect 115736 59302 115742 59366
rect 115806 59302 115812 59366
rect 115736 59094 115812 59302
rect 115736 59062 115742 59094
rect 115398 59030 115399 59062
rect 115333 59029 115399 59030
rect 115741 59030 115742 59062
rect 115806 59062 115812 59094
rect 116824 59366 116900 59372
rect 116824 59302 116830 59366
rect 116894 59302 116900 59366
rect 116824 59094 116900 59302
rect 116824 59062 116830 59094
rect 115806 59030 115807 59062
rect 115741 59029 115807 59030
rect 116829 59030 116830 59062
rect 116894 59062 116900 59094
rect 137496 59094 137844 60934
rect 116894 59030 116895 59062
rect 116829 59029 116895 59030
rect 137496 59030 137502 59094
rect 137566 59030 137844 59094
rect 21896 58958 21972 58964
rect 21896 58894 21902 58958
rect 21966 58894 21972 58958
rect 21896 58686 21972 58894
rect 21896 58654 21902 58686
rect 21901 58622 21902 58654
rect 21966 58654 21972 58686
rect 22304 58958 22380 58964
rect 22304 58894 22310 58958
rect 22374 58894 22380 58958
rect 22304 58686 22380 58894
rect 22304 58654 22310 58686
rect 21966 58622 21967 58654
rect 21901 58621 21967 58622
rect 22309 58622 22310 58654
rect 22374 58654 22380 58686
rect 22984 58958 23060 58964
rect 22984 58894 22990 58958
rect 23054 58894 23060 58958
rect 22984 58686 23060 58894
rect 22984 58654 22990 58686
rect 22374 58622 22375 58654
rect 22309 58621 22375 58622
rect 22989 58622 22990 58654
rect 23054 58654 23060 58686
rect 23392 58958 23468 58964
rect 23392 58894 23398 58958
rect 23462 58894 23468 58958
rect 23392 58686 23468 58894
rect 115192 58958 115268 58964
rect 115192 58894 115198 58958
rect 115262 58894 115268 58958
rect 115741 58958 115807 58959
rect 115741 58926 115742 58958
rect 23392 58654 23398 58686
rect 23054 58622 23055 58654
rect 22989 58621 23055 58622
rect 23397 58622 23398 58654
rect 23462 58654 23468 58686
rect 28565 58686 28631 58687
rect 28565 58654 28566 58686
rect 23462 58622 23463 58654
rect 23397 58621 23463 58622
rect 28560 58622 28566 58654
rect 28630 58654 28631 58686
rect 110432 58686 110508 58692
rect 28630 58622 28636 58654
rect 21901 58550 21967 58551
rect 21901 58518 21902 58550
rect 21896 58486 21902 58518
rect 21966 58518 21967 58550
rect 22168 58550 22244 58556
rect 21966 58486 21972 58518
rect 21896 58278 21972 58486
rect 21896 58214 21902 58278
rect 21966 58214 21972 58278
rect 22168 58486 22174 58550
rect 22238 58486 22244 58550
rect 22717 58550 22783 58551
rect 22717 58518 22718 58550
rect 22168 58278 22244 58486
rect 22168 58246 22174 58278
rect 21896 58208 21972 58214
rect 22173 58214 22174 58246
rect 22238 58246 22244 58278
rect 22712 58486 22718 58518
rect 22782 58518 22783 58550
rect 22989 58550 23055 58551
rect 22989 58518 22990 58550
rect 22782 58486 22788 58518
rect 22712 58278 22788 58486
rect 22238 58214 22239 58246
rect 22173 58213 22239 58214
rect 22712 58214 22718 58278
rect 22782 58214 22788 58278
rect 22712 58208 22788 58214
rect 22984 58486 22990 58518
rect 23054 58518 23055 58550
rect 23397 58550 23463 58551
rect 23397 58518 23398 58550
rect 23054 58486 23060 58518
rect 22984 58278 23060 58486
rect 22984 58214 22990 58278
rect 23054 58214 23060 58278
rect 22984 58208 23060 58214
rect 23392 58486 23398 58518
rect 23462 58518 23463 58550
rect 23462 58486 23468 58518
rect 23392 58278 23468 58486
rect 28560 58414 28636 58622
rect 28560 58350 28566 58414
rect 28630 58350 28636 58414
rect 110432 58622 110438 58686
rect 110502 58622 110508 58686
rect 115192 58686 115268 58894
rect 115192 58654 115198 58686
rect 110432 58414 110508 58622
rect 115197 58622 115198 58654
rect 115262 58654 115268 58686
rect 115736 58894 115742 58926
rect 115806 58926 115807 58958
rect 116149 58958 116215 58959
rect 116149 58926 116150 58958
rect 115806 58894 115812 58926
rect 115736 58686 115812 58894
rect 115262 58622 115263 58654
rect 115197 58621 115263 58622
rect 115736 58622 115742 58686
rect 115806 58622 115812 58686
rect 115736 58616 115812 58622
rect 116144 58894 116150 58926
rect 116214 58926 116215 58958
rect 116552 58958 116628 58964
rect 116214 58894 116220 58926
rect 116144 58686 116220 58894
rect 116144 58622 116150 58686
rect 116214 58622 116220 58686
rect 116552 58894 116558 58958
rect 116622 58894 116628 58958
rect 116829 58958 116895 58959
rect 116829 58926 116830 58958
rect 116552 58686 116628 58894
rect 116552 58654 116558 58686
rect 116144 58616 116220 58622
rect 116557 58622 116558 58654
rect 116622 58654 116628 58686
rect 116824 58894 116830 58926
rect 116894 58926 116895 58958
rect 116894 58894 116900 58926
rect 116824 58686 116900 58894
rect 116622 58622 116623 58654
rect 116557 58621 116623 58622
rect 116824 58622 116830 58686
rect 116894 58622 116900 58686
rect 116824 58616 116900 58622
rect 115197 58550 115263 58551
rect 115197 58518 115198 58550
rect 110432 58382 110438 58414
rect 28560 58344 28636 58350
rect 110437 58350 110438 58382
rect 110502 58382 110508 58414
rect 115192 58486 115198 58518
rect 115262 58518 115263 58550
rect 115736 58550 115812 58556
rect 115262 58486 115268 58518
rect 110502 58350 110503 58382
rect 110437 58349 110503 58350
rect 23392 58214 23398 58278
rect 23462 58214 23468 58278
rect 23392 58208 23468 58214
rect 115192 58278 115268 58486
rect 115192 58214 115198 58278
rect 115262 58214 115268 58278
rect 115736 58486 115742 58550
rect 115806 58486 115812 58550
rect 115736 58278 115812 58486
rect 115736 58246 115742 58278
rect 115192 58208 115268 58214
rect 115741 58214 115742 58246
rect 115806 58246 115812 58278
rect 116008 58550 116084 58556
rect 116008 58486 116014 58550
rect 116078 58486 116084 58550
rect 116008 58278 116084 58486
rect 116008 58246 116014 58278
rect 115806 58214 115807 58246
rect 115741 58213 115807 58214
rect 116013 58214 116014 58246
rect 116078 58246 116084 58278
rect 116824 58550 116900 58556
rect 116824 58486 116830 58550
rect 116894 58486 116900 58550
rect 116824 58278 116900 58486
rect 116824 58246 116830 58278
rect 116078 58214 116079 58246
rect 116013 58213 116079 58214
rect 116829 58214 116830 58246
rect 116894 58246 116900 58278
rect 116894 58214 116895 58246
rect 116829 58213 116895 58214
rect 21765 58142 21831 58143
rect 21765 58110 21766 58142
rect 21760 58078 21766 58110
rect 21830 58110 21831 58142
rect 22440 58142 22516 58148
rect 21830 58078 21836 58110
rect 21760 57870 21836 58078
rect 21760 57806 21766 57870
rect 21830 57806 21836 57870
rect 22440 58078 22446 58142
rect 22510 58078 22516 58142
rect 22989 58142 23055 58143
rect 22989 58110 22990 58142
rect 22440 57870 22516 58078
rect 22440 57838 22446 57870
rect 21760 57800 21836 57806
rect 22445 57806 22446 57838
rect 22510 57838 22516 57870
rect 22984 58078 22990 58110
rect 23054 58110 23055 58142
rect 23528 58142 23604 58148
rect 23054 58078 23060 58110
rect 22984 57870 23060 58078
rect 22510 57806 22511 57838
rect 22445 57805 22511 57806
rect 22984 57806 22990 57870
rect 23054 57806 23060 57870
rect 23528 58078 23534 58142
rect 23598 58078 23604 58142
rect 23528 57870 23604 58078
rect 23528 57838 23534 57870
rect 22984 57800 23060 57806
rect 23533 57806 23534 57838
rect 23598 57838 23604 57870
rect 115192 58142 115268 58148
rect 115192 58078 115198 58142
rect 115262 58078 115268 58142
rect 115192 57870 115268 58078
rect 115192 57838 115198 57870
rect 23598 57806 23599 57838
rect 23533 57805 23599 57806
rect 115197 57806 115198 57838
rect 115262 57838 115268 57870
rect 115736 58142 115812 58148
rect 115736 58078 115742 58142
rect 115806 58078 115812 58142
rect 116829 58142 116895 58143
rect 116829 58110 116830 58142
rect 115736 57870 115812 58078
rect 115736 57838 115742 57870
rect 115262 57806 115263 57838
rect 115197 57805 115263 57806
rect 115741 57806 115742 57838
rect 115806 57838 115812 57870
rect 116824 58078 116830 58110
rect 116894 58110 116895 58142
rect 116894 58078 116900 58110
rect 116824 57870 116900 58078
rect 115806 57806 115807 57838
rect 115741 57805 115807 57806
rect 116824 57806 116830 57870
rect 116894 57806 116900 57870
rect 116824 57800 116900 57806
rect 952 57398 1230 57462
rect 1294 57398 1300 57462
rect 21896 57734 21972 57740
rect 21896 57670 21902 57734
rect 21966 57670 21972 57734
rect 21896 57462 21972 57670
rect 21896 57430 21902 57462
rect 952 55830 1300 57398
rect 21901 57398 21902 57430
rect 21966 57430 21972 57462
rect 22712 57734 22788 57740
rect 22712 57670 22718 57734
rect 22782 57670 22788 57734
rect 22712 57462 22788 57670
rect 22712 57430 22718 57462
rect 21966 57398 21967 57430
rect 21901 57397 21967 57398
rect 22717 57398 22718 57430
rect 22782 57430 22788 57462
rect 23120 57734 23196 57740
rect 23120 57670 23126 57734
rect 23190 57670 23196 57734
rect 23397 57734 23463 57735
rect 23397 57702 23398 57734
rect 23120 57462 23196 57670
rect 23120 57430 23126 57462
rect 22782 57398 22783 57430
rect 22717 57397 22783 57398
rect 23125 57398 23126 57430
rect 23190 57430 23196 57462
rect 23392 57670 23398 57702
rect 23462 57702 23463 57734
rect 115197 57734 115263 57735
rect 115197 57702 115198 57734
rect 23462 57670 23468 57702
rect 23392 57462 23468 57670
rect 23190 57398 23191 57430
rect 23125 57397 23191 57398
rect 23392 57398 23398 57462
rect 23462 57398 23468 57462
rect 23392 57392 23468 57398
rect 115192 57670 115198 57702
rect 115262 57702 115263 57734
rect 115605 57734 115671 57735
rect 115605 57702 115606 57734
rect 115262 57670 115268 57702
rect 115192 57462 115268 57670
rect 115192 57398 115198 57462
rect 115262 57398 115268 57462
rect 115192 57392 115268 57398
rect 115600 57670 115606 57702
rect 115670 57702 115671 57734
rect 116557 57734 116623 57735
rect 116557 57702 116558 57734
rect 115670 57670 115676 57702
rect 115600 57462 115676 57670
rect 115600 57398 115606 57462
rect 115670 57398 115676 57462
rect 115600 57392 115676 57398
rect 116552 57670 116558 57702
rect 116622 57702 116623 57734
rect 116960 57734 117036 57740
rect 116622 57670 116628 57702
rect 116552 57462 116628 57670
rect 116552 57398 116558 57462
rect 116622 57398 116628 57462
rect 116960 57670 116966 57734
rect 117030 57670 117036 57734
rect 116960 57462 117036 57670
rect 116960 57430 116966 57462
rect 116552 57392 116628 57398
rect 116965 57398 116966 57430
rect 117030 57430 117036 57462
rect 137496 57462 137844 59030
rect 117030 57398 117031 57430
rect 116965 57397 117031 57398
rect 137496 57398 137502 57462
rect 137566 57398 137844 57462
rect 23125 57326 23191 57327
rect 23125 57294 23126 57326
rect 23120 57262 23126 57294
rect 23190 57294 23191 57326
rect 23528 57326 23604 57332
rect 23190 57262 23196 57294
rect 23120 57054 23196 57262
rect 23120 56990 23126 57054
rect 23190 56990 23196 57054
rect 23528 57262 23534 57326
rect 23598 57262 23604 57326
rect 23528 57054 23604 57262
rect 23528 57022 23534 57054
rect 23120 56984 23196 56990
rect 23533 56990 23534 57022
rect 23598 57022 23604 57054
rect 115328 57326 115404 57332
rect 115328 57262 115334 57326
rect 115398 57262 115404 57326
rect 115328 57054 115404 57262
rect 115328 57022 115334 57054
rect 23598 56990 23599 57022
rect 23533 56989 23599 56990
rect 115333 56990 115334 57022
rect 115398 57022 115404 57054
rect 115736 57326 115812 57332
rect 115736 57262 115742 57326
rect 115806 57262 115812 57326
rect 116149 57326 116215 57327
rect 116149 57294 116150 57326
rect 115736 57054 115812 57262
rect 115736 57022 115742 57054
rect 115398 56990 115399 57022
rect 115333 56989 115399 56990
rect 115741 56990 115742 57022
rect 115806 57022 115812 57054
rect 116144 57262 116150 57294
rect 116214 57294 116215 57326
rect 116285 57326 116351 57327
rect 116285 57294 116286 57326
rect 116214 57262 116220 57294
rect 116144 57054 116220 57262
rect 115806 56990 115807 57022
rect 115741 56989 115807 56990
rect 116144 56990 116150 57054
rect 116214 56990 116220 57054
rect 116144 56984 116220 56990
rect 116280 57262 116286 57294
rect 116350 57294 116351 57326
rect 116350 57262 116356 57294
rect 116280 57054 116356 57262
rect 116280 56990 116286 57054
rect 116350 56990 116356 57054
rect 116280 56984 116356 56990
rect 22440 56918 22516 56924
rect 22440 56854 22446 56918
rect 22510 56854 22516 56918
rect 22440 56646 22516 56854
rect 22440 56614 22446 56646
rect 22445 56582 22446 56614
rect 22510 56614 22516 56646
rect 22984 56918 23060 56924
rect 22984 56854 22990 56918
rect 23054 56854 23060 56918
rect 23533 56918 23599 56919
rect 23533 56886 23534 56918
rect 22984 56646 23060 56854
rect 22984 56614 22990 56646
rect 22510 56582 22511 56614
rect 22445 56581 22511 56582
rect 22989 56582 22990 56614
rect 23054 56614 23060 56646
rect 23528 56854 23534 56886
rect 23598 56886 23599 56918
rect 115192 56918 115268 56924
rect 23598 56854 23604 56886
rect 23528 56646 23604 56854
rect 23054 56582 23055 56614
rect 22989 56581 23055 56582
rect 23528 56582 23534 56646
rect 23598 56582 23604 56646
rect 115192 56854 115198 56918
rect 115262 56854 115268 56918
rect 115192 56646 115268 56854
rect 115192 56614 115198 56646
rect 23528 56576 23604 56582
rect 115197 56582 115198 56614
rect 115262 56614 115268 56646
rect 115600 56918 115676 56924
rect 115600 56854 115606 56918
rect 115670 56854 115676 56918
rect 115600 56646 115676 56854
rect 115600 56614 115606 56646
rect 115262 56582 115263 56614
rect 115197 56581 115263 56582
rect 115605 56582 115606 56614
rect 115670 56614 115676 56646
rect 115670 56582 115671 56614
rect 115605 56581 115671 56582
rect 22440 56510 22516 56516
rect 22440 56446 22446 56510
rect 22510 56446 22516 56510
rect 21901 56238 21967 56239
rect 21901 56206 21902 56238
rect 21896 56174 21902 56206
rect 21966 56206 21967 56238
rect 22440 56238 22516 56446
rect 22440 56206 22446 56238
rect 21966 56174 21972 56206
rect 21896 55966 21972 56174
rect 22445 56174 22446 56206
rect 22510 56206 22516 56238
rect 22712 56510 22788 56516
rect 22712 56446 22718 56510
rect 22782 56446 22788 56510
rect 22989 56510 23055 56511
rect 22989 56478 22990 56510
rect 22712 56238 22788 56446
rect 22712 56206 22718 56238
rect 22510 56174 22511 56206
rect 22445 56173 22511 56174
rect 22717 56174 22718 56206
rect 22782 56206 22788 56238
rect 22984 56446 22990 56478
rect 23054 56478 23055 56510
rect 23392 56510 23468 56516
rect 23054 56446 23060 56478
rect 22984 56238 23060 56446
rect 22782 56174 22783 56206
rect 22717 56173 22783 56174
rect 22984 56174 22990 56238
rect 23054 56174 23060 56238
rect 23392 56446 23398 56510
rect 23462 56446 23468 56510
rect 23392 56238 23468 56446
rect 115192 56510 115268 56516
rect 115192 56446 115198 56510
rect 115262 56446 115268 56510
rect 115605 56510 115671 56511
rect 115605 56478 115606 56510
rect 110437 56374 110503 56375
rect 110437 56342 110438 56374
rect 23392 56206 23398 56238
rect 22984 56168 23060 56174
rect 23397 56174 23398 56206
rect 23462 56206 23468 56238
rect 110432 56310 110438 56342
rect 110502 56342 110503 56374
rect 110502 56310 110508 56342
rect 23462 56174 23463 56206
rect 23397 56173 23463 56174
rect 110432 56102 110508 56310
rect 115192 56238 115268 56446
rect 115192 56206 115198 56238
rect 115197 56174 115198 56206
rect 115262 56206 115268 56238
rect 115600 56446 115606 56478
rect 115670 56478 115671 56510
rect 116557 56510 116623 56511
rect 116557 56478 116558 56510
rect 115670 56446 115676 56478
rect 115600 56238 115676 56446
rect 115262 56174 115263 56206
rect 115197 56173 115263 56174
rect 115600 56174 115606 56238
rect 115670 56174 115676 56238
rect 115600 56168 115676 56174
rect 116552 56446 116558 56478
rect 116622 56478 116623 56510
rect 116622 56446 116628 56478
rect 116552 56238 116628 56446
rect 116552 56174 116558 56238
rect 116622 56174 116628 56238
rect 116965 56238 117031 56239
rect 116965 56206 116966 56238
rect 116552 56168 116628 56174
rect 116960 56174 116966 56206
rect 117030 56206 117031 56238
rect 117030 56174 117036 56206
rect 110432 56038 110438 56102
rect 110502 56038 110508 56102
rect 110432 56032 110508 56038
rect 21896 55902 21902 55966
rect 21966 55902 21972 55966
rect 28565 55966 28631 55967
rect 28565 55934 28566 55966
rect 21896 55896 21972 55902
rect 28560 55902 28566 55934
rect 28630 55934 28631 55966
rect 110432 55966 110508 55972
rect 28630 55902 28636 55934
rect 952 55766 1230 55830
rect 1294 55766 1300 55830
rect 21765 55830 21831 55831
rect 21765 55798 21766 55830
rect 952 54198 1300 55766
rect 21760 55766 21766 55798
rect 21830 55798 21831 55830
rect 22581 55830 22647 55831
rect 22581 55798 22582 55830
rect 21830 55766 21836 55798
rect 21760 55558 21836 55766
rect 21760 55494 21766 55558
rect 21830 55494 21836 55558
rect 21760 55488 21836 55494
rect 22576 55766 22582 55798
rect 22646 55798 22647 55830
rect 22646 55766 22652 55798
rect 22576 55558 22652 55766
rect 28560 55694 28636 55902
rect 28560 55630 28566 55694
rect 28630 55630 28636 55694
rect 110432 55902 110438 55966
rect 110502 55902 110508 55966
rect 110432 55694 110508 55902
rect 116960 55966 117036 56174
rect 116960 55902 116966 55966
rect 117030 55902 117036 55966
rect 116960 55896 117036 55902
rect 110432 55662 110438 55694
rect 28560 55624 28636 55630
rect 110437 55630 110438 55662
rect 110502 55662 110508 55694
rect 116552 55830 116628 55836
rect 116552 55766 116558 55830
rect 116622 55766 116628 55830
rect 110502 55630 110503 55662
rect 110437 55629 110503 55630
rect 22576 55494 22582 55558
rect 22646 55494 22652 55558
rect 28565 55558 28631 55559
rect 28565 55526 28566 55558
rect 22576 55488 22652 55494
rect 28560 55494 28566 55526
rect 28630 55526 28631 55558
rect 110432 55558 110508 55564
rect 28630 55494 28636 55526
rect 21896 55422 21972 55428
rect 21896 55358 21902 55422
rect 21966 55358 21972 55422
rect 21896 55150 21972 55358
rect 28560 55286 28636 55494
rect 28560 55222 28566 55286
rect 28630 55222 28636 55286
rect 110432 55494 110438 55558
rect 110502 55494 110508 55558
rect 116552 55558 116628 55766
rect 116552 55526 116558 55558
rect 110432 55286 110508 55494
rect 116557 55494 116558 55526
rect 116622 55526 116628 55558
rect 116960 55830 117036 55836
rect 116960 55766 116966 55830
rect 117030 55766 117036 55830
rect 116960 55558 117036 55766
rect 116960 55526 116966 55558
rect 116622 55494 116623 55526
rect 116557 55493 116623 55494
rect 116965 55494 116966 55526
rect 117030 55526 117036 55558
rect 137496 55830 137844 57398
rect 137496 55766 137502 55830
rect 137566 55766 137844 55830
rect 117030 55494 117031 55526
rect 116965 55493 117031 55494
rect 116965 55422 117031 55423
rect 116965 55390 116966 55422
rect 110432 55254 110438 55286
rect 28560 55216 28636 55222
rect 110437 55222 110438 55254
rect 110502 55254 110508 55286
rect 116960 55358 116966 55390
rect 117030 55390 117031 55422
rect 117030 55358 117036 55390
rect 110502 55222 110503 55254
rect 110437 55221 110503 55222
rect 21896 55118 21902 55150
rect 21901 55086 21902 55118
rect 21966 55118 21972 55150
rect 116960 55150 117036 55358
rect 21966 55086 21967 55118
rect 21901 55085 21967 55086
rect 116960 55086 116966 55150
rect 117030 55086 117036 55150
rect 116960 55080 117036 55086
rect 21765 55014 21831 55015
rect 21765 54982 21766 55014
rect 21760 54950 21766 54982
rect 21830 54982 21831 55014
rect 22173 55014 22239 55015
rect 22173 54982 22174 55014
rect 21830 54950 21836 54982
rect 21760 54742 21836 54950
rect 21760 54678 21766 54742
rect 21830 54678 21836 54742
rect 21760 54672 21836 54678
rect 22168 54950 22174 54982
rect 22238 54982 22239 55014
rect 22989 55014 23055 55015
rect 22989 54982 22990 55014
rect 22238 54950 22244 54982
rect 22168 54742 22244 54950
rect 22168 54678 22174 54742
rect 22238 54678 22244 54742
rect 22168 54672 22244 54678
rect 22984 54950 22990 54982
rect 23054 54982 23055 55014
rect 23528 55014 23604 55020
rect 23054 54950 23060 54982
rect 22984 54742 23060 54950
rect 22984 54678 22990 54742
rect 23054 54678 23060 54742
rect 23528 54950 23534 55014
rect 23598 54950 23604 55014
rect 115197 55014 115263 55015
rect 115197 54982 115198 55014
rect 23528 54742 23604 54950
rect 115192 54950 115198 54982
rect 115262 54982 115263 55014
rect 115741 55014 115807 55015
rect 115741 54982 115742 55014
rect 115262 54950 115268 54982
rect 23528 54710 23534 54742
rect 22984 54672 23060 54678
rect 23533 54678 23534 54710
rect 23598 54710 23604 54742
rect 28293 54742 28359 54743
rect 28293 54710 28294 54742
rect 23598 54678 23599 54710
rect 23533 54677 23599 54678
rect 28288 54678 28294 54710
rect 28358 54710 28359 54742
rect 115192 54742 115268 54950
rect 28358 54678 28364 54710
rect 21896 54606 21972 54612
rect 21896 54542 21902 54606
rect 21966 54542 21972 54606
rect 21896 54334 21972 54542
rect 21896 54302 21902 54334
rect 21901 54270 21902 54302
rect 21966 54302 21972 54334
rect 22304 54606 22380 54612
rect 22304 54542 22310 54606
rect 22374 54542 22380 54606
rect 22304 54334 22380 54542
rect 22304 54302 22310 54334
rect 21966 54270 21967 54302
rect 21901 54269 21967 54270
rect 22309 54270 22310 54302
rect 22374 54302 22380 54334
rect 22440 54606 22516 54612
rect 22440 54542 22446 54606
rect 22510 54542 22516 54606
rect 22440 54334 22516 54542
rect 22440 54302 22446 54334
rect 22374 54270 22375 54302
rect 22309 54269 22375 54270
rect 22445 54270 22446 54302
rect 22510 54302 22516 54334
rect 22984 54606 23060 54612
rect 22984 54542 22990 54606
rect 23054 54542 23060 54606
rect 23533 54606 23599 54607
rect 23533 54574 23534 54606
rect 22984 54334 23060 54542
rect 22984 54302 22990 54334
rect 22510 54270 22511 54302
rect 22445 54269 22511 54270
rect 22989 54270 22990 54302
rect 23054 54302 23060 54334
rect 23528 54542 23534 54574
rect 23598 54574 23599 54606
rect 23598 54542 23604 54574
rect 23528 54334 23604 54542
rect 28288 54470 28364 54678
rect 115192 54678 115198 54742
rect 115262 54678 115268 54742
rect 115192 54672 115268 54678
rect 115736 54950 115742 54982
rect 115806 54982 115807 55014
rect 116285 55014 116351 55015
rect 116285 54982 116286 55014
rect 115806 54950 115812 54982
rect 115736 54742 115812 54950
rect 115736 54678 115742 54742
rect 115806 54678 115812 54742
rect 115736 54672 115812 54678
rect 116280 54950 116286 54982
rect 116350 54982 116351 55014
rect 116824 55014 116900 55020
rect 116350 54950 116356 54982
rect 116280 54742 116356 54950
rect 116280 54678 116286 54742
rect 116350 54678 116356 54742
rect 116824 54950 116830 55014
rect 116894 54950 116900 55014
rect 116824 54742 116900 54950
rect 116824 54710 116830 54742
rect 116280 54672 116356 54678
rect 116829 54678 116830 54710
rect 116894 54710 116900 54742
rect 116894 54678 116895 54710
rect 116829 54677 116895 54678
rect 115333 54606 115399 54607
rect 115333 54574 115334 54606
rect 28288 54406 28294 54470
rect 28358 54406 28364 54470
rect 28288 54400 28364 54406
rect 115328 54542 115334 54574
rect 115398 54574 115399 54606
rect 115741 54606 115807 54607
rect 115741 54574 115742 54606
rect 115398 54542 115404 54574
rect 23054 54270 23055 54302
rect 22989 54269 23055 54270
rect 23528 54270 23534 54334
rect 23598 54270 23604 54334
rect 23528 54264 23604 54270
rect 115328 54334 115404 54542
rect 115328 54270 115334 54334
rect 115398 54270 115404 54334
rect 115328 54264 115404 54270
rect 115736 54542 115742 54574
rect 115806 54574 115807 54606
rect 116149 54606 116215 54607
rect 116149 54574 116150 54606
rect 115806 54542 115812 54574
rect 115736 54334 115812 54542
rect 115736 54270 115742 54334
rect 115806 54270 115812 54334
rect 115736 54264 115812 54270
rect 116144 54542 116150 54574
rect 116214 54574 116215 54606
rect 116280 54606 116356 54612
rect 116214 54542 116220 54574
rect 116144 54334 116220 54542
rect 116144 54270 116150 54334
rect 116214 54270 116220 54334
rect 116280 54542 116286 54606
rect 116350 54542 116356 54606
rect 116829 54606 116895 54607
rect 116829 54574 116830 54606
rect 116280 54334 116356 54542
rect 116280 54302 116286 54334
rect 116144 54264 116220 54270
rect 116285 54270 116286 54302
rect 116350 54302 116356 54334
rect 116824 54542 116830 54574
rect 116894 54574 116895 54606
rect 116894 54542 116900 54574
rect 116824 54334 116900 54542
rect 116350 54270 116351 54302
rect 116285 54269 116351 54270
rect 116824 54270 116830 54334
rect 116894 54270 116900 54334
rect 116824 54264 116900 54270
rect 952 54134 1230 54198
rect 1294 54134 1300 54198
rect 21901 54198 21967 54199
rect 21901 54166 21902 54198
rect 952 52566 1300 54134
rect 21896 54134 21902 54166
rect 21966 54166 21967 54198
rect 22168 54198 22244 54204
rect 21966 54134 21972 54166
rect 21896 53926 21972 54134
rect 21896 53862 21902 53926
rect 21966 53862 21972 53926
rect 22168 54134 22174 54198
rect 22238 54134 22244 54198
rect 22168 53926 22244 54134
rect 22168 53894 22174 53926
rect 21896 53856 21972 53862
rect 22173 53862 22174 53894
rect 22238 53894 22244 53926
rect 22984 54198 23060 54204
rect 22984 54134 22990 54198
rect 23054 54134 23060 54198
rect 23397 54198 23463 54199
rect 23397 54166 23398 54198
rect 22984 53926 23060 54134
rect 22984 53894 22990 53926
rect 22238 53862 22239 53894
rect 22173 53861 22239 53862
rect 22989 53862 22990 53894
rect 23054 53894 23060 53926
rect 23392 54134 23398 54166
rect 23462 54166 23463 54198
rect 115328 54198 115404 54204
rect 23462 54134 23468 54166
rect 23392 53926 23468 54134
rect 23054 53862 23055 53894
rect 22989 53861 23055 53862
rect 23392 53862 23398 53926
rect 23462 53862 23468 53926
rect 115328 54134 115334 54198
rect 115398 54134 115404 54198
rect 115605 54198 115671 54199
rect 115605 54166 115606 54198
rect 115328 53926 115404 54134
rect 115328 53894 115334 53926
rect 23392 53856 23468 53862
rect 115333 53862 115334 53894
rect 115398 53894 115404 53926
rect 115600 54134 115606 54166
rect 115670 54166 115671 54198
rect 116008 54198 116084 54204
rect 115670 54134 115676 54166
rect 115600 53926 115676 54134
rect 115398 53862 115399 53894
rect 115333 53861 115399 53862
rect 115600 53862 115606 53926
rect 115670 53862 115676 53926
rect 116008 54134 116014 54198
rect 116078 54134 116084 54198
rect 116008 53926 116084 54134
rect 116008 53894 116014 53926
rect 115600 53856 115676 53862
rect 116013 53862 116014 53894
rect 116078 53894 116084 53926
rect 116416 54198 116492 54204
rect 116416 54134 116422 54198
rect 116486 54134 116492 54198
rect 116416 53926 116492 54134
rect 116416 53894 116422 53926
rect 116078 53862 116079 53894
rect 116013 53861 116079 53862
rect 116421 53862 116422 53894
rect 116486 53894 116492 53926
rect 116824 54198 116900 54204
rect 116824 54134 116830 54198
rect 116894 54134 116900 54198
rect 116824 53926 116900 54134
rect 116824 53894 116830 53926
rect 116486 53862 116487 53894
rect 116421 53861 116487 53862
rect 116829 53862 116830 53894
rect 116894 53894 116900 53926
rect 137496 54198 137844 55766
rect 137496 54134 137502 54198
rect 137566 54134 137844 54198
rect 116894 53862 116895 53894
rect 116829 53861 116895 53862
rect 21765 53790 21831 53791
rect 21765 53758 21766 53790
rect 21760 53726 21766 53758
rect 21830 53758 21831 53790
rect 22173 53790 22239 53791
rect 22173 53758 22174 53790
rect 21830 53726 21836 53758
rect 21760 53518 21836 53726
rect 21760 53454 21766 53518
rect 21830 53454 21836 53518
rect 21760 53448 21836 53454
rect 22168 53726 22174 53758
rect 22238 53758 22239 53790
rect 22581 53790 22647 53791
rect 22581 53758 22582 53790
rect 22238 53726 22244 53758
rect 22168 53518 22244 53726
rect 22168 53454 22174 53518
rect 22238 53454 22244 53518
rect 22168 53448 22244 53454
rect 22576 53726 22582 53758
rect 22646 53758 22647 53790
rect 23120 53790 23196 53796
rect 22646 53726 22652 53758
rect 22576 53518 22652 53726
rect 22576 53454 22582 53518
rect 22646 53454 22652 53518
rect 23120 53726 23126 53790
rect 23190 53726 23196 53790
rect 23120 53518 23196 53726
rect 23120 53486 23126 53518
rect 22576 53448 22652 53454
rect 23125 53454 23126 53486
rect 23190 53486 23196 53518
rect 23528 53790 23604 53796
rect 23528 53726 23534 53790
rect 23598 53726 23604 53790
rect 115333 53790 115399 53791
rect 115333 53758 115334 53790
rect 23528 53518 23604 53726
rect 23528 53486 23534 53518
rect 23190 53454 23191 53486
rect 23125 53453 23191 53454
rect 23533 53454 23534 53486
rect 23598 53486 23604 53518
rect 115328 53726 115334 53758
rect 115398 53758 115399 53790
rect 115736 53790 115812 53796
rect 115398 53726 115404 53758
rect 115328 53518 115404 53726
rect 23598 53454 23599 53486
rect 23533 53453 23599 53454
rect 115328 53454 115334 53518
rect 115398 53454 115404 53518
rect 115736 53726 115742 53790
rect 115806 53726 115812 53790
rect 115736 53518 115812 53726
rect 115736 53486 115742 53518
rect 115328 53448 115404 53454
rect 115741 53454 115742 53486
rect 115806 53486 115812 53518
rect 116280 53790 116356 53796
rect 116280 53726 116286 53790
rect 116350 53726 116356 53790
rect 116829 53790 116895 53791
rect 116829 53758 116830 53790
rect 116280 53518 116356 53726
rect 116280 53486 116286 53518
rect 115806 53454 115807 53486
rect 115741 53453 115807 53454
rect 116285 53454 116286 53486
rect 116350 53486 116356 53518
rect 116824 53726 116830 53758
rect 116894 53758 116895 53790
rect 116894 53726 116900 53758
rect 116824 53518 116900 53726
rect 116350 53454 116351 53486
rect 116285 53453 116351 53454
rect 116824 53454 116830 53518
rect 116894 53454 116900 53518
rect 116824 53448 116900 53454
rect 22717 53382 22783 53383
rect 22717 53350 22718 53382
rect 22712 53318 22718 53350
rect 22782 53350 22783 53382
rect 22989 53382 23055 53383
rect 22989 53350 22990 53382
rect 22782 53318 22788 53350
rect 22712 53110 22788 53318
rect 22712 53046 22718 53110
rect 22782 53046 22788 53110
rect 22712 53040 22788 53046
rect 22984 53318 22990 53350
rect 23054 53350 23055 53382
rect 23397 53382 23463 53383
rect 23397 53350 23398 53382
rect 23054 53318 23060 53350
rect 22984 53110 23060 53318
rect 22984 53046 22990 53110
rect 23054 53046 23060 53110
rect 22984 53040 23060 53046
rect 23392 53318 23398 53350
rect 23462 53350 23463 53382
rect 115192 53382 115268 53388
rect 23462 53318 23468 53350
rect 23392 53110 23468 53318
rect 23392 53046 23398 53110
rect 23462 53046 23468 53110
rect 115192 53318 115198 53382
rect 115262 53318 115268 53382
rect 115605 53382 115671 53383
rect 115605 53350 115606 53382
rect 115192 53110 115268 53318
rect 115192 53078 115198 53110
rect 23392 53040 23468 53046
rect 115197 53046 115198 53078
rect 115262 53078 115268 53110
rect 115600 53318 115606 53350
rect 115670 53350 115671 53382
rect 116557 53382 116623 53383
rect 116557 53350 116558 53382
rect 115670 53318 115676 53350
rect 115600 53110 115676 53318
rect 115262 53046 115263 53078
rect 115197 53045 115263 53046
rect 115600 53046 115606 53110
rect 115670 53046 115676 53110
rect 115600 53040 115676 53046
rect 116552 53318 116558 53350
rect 116622 53350 116623 53382
rect 116622 53318 116628 53350
rect 116552 53110 116628 53318
rect 116552 53046 116558 53110
rect 116622 53046 116628 53110
rect 116552 53040 116628 53046
rect 21760 52974 21836 52980
rect 21760 52910 21766 52974
rect 21830 52910 21836 52974
rect 22445 52974 22511 52975
rect 22445 52942 22446 52974
rect 21760 52702 21836 52910
rect 21760 52670 21766 52702
rect 21765 52638 21766 52670
rect 21830 52670 21836 52702
rect 22440 52910 22446 52942
rect 22510 52942 22511 52974
rect 23120 52974 23196 52980
rect 22510 52910 22516 52942
rect 22440 52702 22516 52910
rect 21830 52638 21831 52670
rect 21765 52637 21831 52638
rect 22440 52638 22446 52702
rect 22510 52638 22516 52702
rect 23120 52910 23126 52974
rect 23190 52910 23196 52974
rect 23120 52702 23196 52910
rect 23120 52670 23126 52702
rect 22440 52632 22516 52638
rect 23125 52638 23126 52670
rect 23190 52670 23196 52702
rect 23528 52974 23604 52980
rect 23528 52910 23534 52974
rect 23598 52910 23604 52974
rect 23528 52702 23604 52910
rect 23528 52670 23534 52702
rect 23190 52638 23191 52670
rect 23125 52637 23191 52638
rect 23533 52638 23534 52670
rect 23598 52670 23604 52702
rect 115328 52974 115404 52980
rect 115328 52910 115334 52974
rect 115398 52910 115404 52974
rect 115328 52702 115404 52910
rect 115328 52670 115334 52702
rect 23598 52638 23599 52670
rect 23533 52637 23599 52638
rect 115333 52638 115334 52670
rect 115398 52670 115404 52702
rect 115736 52974 115812 52980
rect 115736 52910 115742 52974
rect 115806 52910 115812 52974
rect 116149 52974 116215 52975
rect 116149 52942 116150 52974
rect 115736 52702 115812 52910
rect 115736 52670 115742 52702
rect 115398 52638 115399 52670
rect 115333 52637 115399 52638
rect 115741 52638 115742 52670
rect 115806 52670 115812 52702
rect 116144 52910 116150 52942
rect 116214 52942 116215 52974
rect 116285 52974 116351 52975
rect 116285 52942 116286 52974
rect 116214 52910 116220 52942
rect 116144 52702 116220 52910
rect 115806 52638 115807 52670
rect 115741 52637 115807 52638
rect 116144 52638 116150 52702
rect 116214 52638 116220 52702
rect 116144 52632 116220 52638
rect 116280 52910 116286 52942
rect 116350 52942 116351 52974
rect 116416 52974 116492 52980
rect 116350 52910 116356 52942
rect 116280 52702 116356 52910
rect 116280 52638 116286 52702
rect 116350 52638 116356 52702
rect 116416 52910 116422 52974
rect 116486 52910 116492 52974
rect 116416 52702 116492 52910
rect 116416 52670 116422 52702
rect 116280 52632 116356 52638
rect 116421 52638 116422 52670
rect 116486 52670 116492 52702
rect 116824 52974 116900 52980
rect 116824 52910 116830 52974
rect 116894 52910 116900 52974
rect 116824 52702 116900 52910
rect 116824 52670 116830 52702
rect 116486 52638 116487 52670
rect 116421 52637 116487 52638
rect 116829 52638 116830 52670
rect 116894 52670 116900 52702
rect 116894 52638 116895 52670
rect 116829 52637 116895 52638
rect 952 52502 1230 52566
rect 1294 52502 1300 52566
rect 22173 52566 22239 52567
rect 22173 52534 22174 52566
rect 952 50934 1300 52502
rect 22168 52502 22174 52534
rect 22238 52534 22239 52566
rect 22712 52566 22788 52572
rect 22238 52502 22244 52534
rect 21896 52294 21972 52300
rect 21896 52230 21902 52294
rect 21966 52230 21972 52294
rect 21896 52022 21972 52230
rect 22168 52294 22244 52502
rect 22168 52230 22174 52294
rect 22238 52230 22244 52294
rect 22712 52502 22718 52566
rect 22782 52502 22788 52566
rect 22989 52566 23055 52567
rect 22989 52534 22990 52566
rect 22712 52294 22788 52502
rect 22712 52262 22718 52294
rect 22168 52224 22244 52230
rect 22717 52230 22718 52262
rect 22782 52262 22788 52294
rect 22984 52502 22990 52534
rect 23054 52534 23055 52566
rect 23392 52566 23468 52572
rect 23054 52502 23060 52534
rect 22984 52294 23060 52502
rect 22782 52230 22783 52262
rect 22717 52229 22783 52230
rect 22984 52230 22990 52294
rect 23054 52230 23060 52294
rect 23392 52502 23398 52566
rect 23462 52502 23468 52566
rect 115333 52566 115399 52567
rect 115333 52534 115334 52566
rect 23392 52294 23468 52502
rect 115328 52502 115334 52534
rect 115398 52534 115399 52566
rect 115741 52566 115807 52567
rect 115741 52534 115742 52566
rect 115398 52502 115404 52534
rect 110437 52430 110503 52431
rect 110437 52398 110438 52430
rect 23392 52262 23398 52294
rect 22984 52224 23060 52230
rect 23397 52230 23398 52262
rect 23462 52262 23468 52294
rect 110432 52366 110438 52398
rect 110502 52398 110503 52430
rect 110502 52366 110508 52398
rect 23462 52230 23463 52262
rect 23397 52229 23463 52230
rect 22989 52158 23055 52159
rect 22989 52126 22990 52158
rect 21896 51990 21902 52022
rect 21901 51958 21902 51990
rect 21966 51990 21972 52022
rect 22984 52094 22990 52126
rect 23054 52126 23055 52158
rect 23397 52158 23463 52159
rect 23397 52126 23398 52158
rect 23054 52094 23060 52126
rect 21966 51958 21967 51990
rect 21901 51957 21967 51958
rect 22984 51886 23060 52094
rect 22984 51822 22990 51886
rect 23054 51822 23060 51886
rect 22984 51816 23060 51822
rect 23392 52094 23398 52126
rect 23462 52126 23463 52158
rect 110432 52158 110508 52366
rect 115328 52294 115404 52502
rect 115328 52230 115334 52294
rect 115398 52230 115404 52294
rect 115328 52224 115404 52230
rect 115736 52502 115742 52534
rect 115806 52534 115807 52566
rect 116008 52566 116084 52572
rect 115806 52502 115812 52534
rect 115736 52294 115812 52502
rect 115736 52230 115742 52294
rect 115806 52230 115812 52294
rect 116008 52502 116014 52566
rect 116078 52502 116084 52566
rect 116285 52566 116351 52567
rect 116285 52534 116286 52566
rect 116008 52294 116084 52502
rect 116008 52262 116014 52294
rect 115736 52224 115812 52230
rect 116013 52230 116014 52262
rect 116078 52262 116084 52294
rect 116280 52502 116286 52534
rect 116350 52534 116351 52566
rect 137496 52566 137844 54134
rect 116350 52502 116356 52534
rect 116280 52294 116356 52502
rect 137496 52502 137502 52566
rect 137566 52502 137844 52566
rect 116078 52230 116079 52262
rect 116013 52229 116079 52230
rect 116280 52230 116286 52294
rect 116350 52230 116356 52294
rect 116965 52294 117031 52295
rect 116965 52262 116966 52294
rect 116280 52224 116356 52230
rect 116960 52230 116966 52262
rect 117030 52262 117031 52294
rect 117030 52230 117036 52262
rect 23462 52094 23468 52126
rect 23392 51886 23468 52094
rect 110432 52094 110438 52158
rect 110502 52094 110508 52158
rect 110432 52088 110508 52094
rect 115192 52158 115268 52164
rect 115192 52094 115198 52158
rect 115262 52094 115268 52158
rect 115605 52158 115671 52159
rect 115605 52126 115606 52158
rect 23392 51822 23398 51886
rect 23462 51822 23468 51886
rect 28429 51886 28495 51887
rect 28429 51854 28430 51886
rect 23392 51816 23468 51822
rect 28424 51822 28430 51854
rect 28494 51854 28495 51886
rect 115192 51886 115268 52094
rect 115192 51854 115198 51886
rect 28494 51822 28500 51854
rect 22168 51750 22244 51756
rect 22168 51686 22174 51750
rect 22238 51686 22244 51750
rect 21765 51478 21831 51479
rect 21765 51446 21766 51478
rect 21760 51414 21766 51446
rect 21830 51446 21831 51478
rect 22168 51478 22244 51686
rect 28424 51614 28500 51822
rect 115197 51822 115198 51854
rect 115262 51854 115268 51886
rect 115600 52094 115606 52126
rect 115670 52126 115671 52158
rect 115670 52094 115676 52126
rect 115600 51886 115676 52094
rect 116960 52022 117036 52230
rect 116960 51958 116966 52022
rect 117030 51958 117036 52022
rect 116960 51952 117036 51958
rect 115262 51822 115263 51854
rect 115197 51821 115263 51822
rect 115600 51822 115606 51886
rect 115670 51822 115676 51886
rect 115600 51816 115676 51822
rect 116013 51750 116079 51751
rect 116013 51718 116014 51750
rect 116008 51686 116014 51718
rect 116078 51718 116079 51750
rect 116421 51750 116487 51751
rect 116421 51718 116422 51750
rect 116078 51686 116084 51718
rect 28424 51550 28430 51614
rect 28494 51550 28500 51614
rect 28565 51614 28631 51615
rect 28565 51582 28566 51614
rect 28424 51544 28500 51550
rect 28560 51550 28566 51582
rect 28630 51582 28631 51614
rect 28630 51550 28636 51582
rect 22168 51446 22174 51478
rect 21830 51414 21836 51446
rect 21760 51206 21836 51414
rect 22173 51414 22174 51446
rect 22238 51446 22244 51478
rect 22238 51414 22239 51446
rect 22173 51413 22239 51414
rect 28560 51342 28636 51550
rect 116008 51478 116084 51686
rect 116008 51414 116014 51478
rect 116078 51414 116084 51478
rect 116008 51408 116084 51414
rect 116416 51686 116422 51718
rect 116486 51718 116487 51750
rect 116486 51686 116492 51718
rect 116416 51478 116492 51686
rect 116416 51414 116422 51478
rect 116486 51414 116492 51478
rect 116829 51478 116895 51479
rect 116829 51446 116830 51478
rect 116416 51408 116492 51414
rect 116824 51414 116830 51446
rect 116894 51446 116895 51478
rect 116894 51414 116900 51446
rect 28560 51278 28566 51342
rect 28630 51278 28636 51342
rect 28560 51272 28636 51278
rect 21760 51142 21766 51206
rect 21830 51142 21836 51206
rect 21760 51136 21836 51142
rect 116824 51206 116900 51414
rect 116824 51142 116830 51206
rect 116894 51142 116900 51206
rect 116824 51136 116900 51142
rect 952 50870 1230 50934
rect 1294 50870 1300 50934
rect 952 49166 1300 50870
rect 21896 51070 21972 51076
rect 21896 51006 21902 51070
rect 21966 51006 21972 51070
rect 22309 51070 22375 51071
rect 22309 51038 22310 51070
rect 21896 50798 21972 51006
rect 21896 50766 21902 50798
rect 21901 50734 21902 50766
rect 21966 50766 21972 50798
rect 22304 51006 22310 51038
rect 22374 51038 22375 51070
rect 22445 51070 22511 51071
rect 22445 51038 22446 51070
rect 22374 51006 22380 51038
rect 22304 50798 22380 51006
rect 21966 50734 21967 50766
rect 21901 50733 21967 50734
rect 22304 50734 22310 50798
rect 22374 50734 22380 50798
rect 22304 50728 22380 50734
rect 22440 51006 22446 51038
rect 22510 51038 22511 51070
rect 22989 51070 23055 51071
rect 22989 51038 22990 51070
rect 22510 51006 22516 51038
rect 22440 50798 22516 51006
rect 22440 50734 22446 50798
rect 22510 50734 22516 50798
rect 22440 50728 22516 50734
rect 22984 51006 22990 51038
rect 23054 51038 23055 51070
rect 23392 51070 23468 51076
rect 23054 51006 23060 51038
rect 22984 50798 23060 51006
rect 22984 50734 22990 50798
rect 23054 50734 23060 50798
rect 23392 51006 23398 51070
rect 23462 51006 23468 51070
rect 23392 50798 23468 51006
rect 115192 51070 115268 51076
rect 115192 51006 115198 51070
rect 115262 51006 115268 51070
rect 115605 51070 115671 51071
rect 115605 51038 115606 51070
rect 23392 50766 23398 50798
rect 22984 50728 23060 50734
rect 23397 50734 23398 50766
rect 23462 50766 23468 50798
rect 110432 50798 110508 50804
rect 23462 50734 23463 50766
rect 23397 50733 23463 50734
rect 110432 50734 110438 50798
rect 110502 50734 110508 50798
rect 115192 50798 115268 51006
rect 115192 50766 115198 50798
rect 21760 50662 21836 50668
rect 21760 50598 21766 50662
rect 21830 50598 21836 50662
rect 21760 50390 21836 50598
rect 21760 50358 21766 50390
rect 21765 50326 21766 50358
rect 21830 50358 21836 50390
rect 22168 50662 22244 50668
rect 22168 50598 22174 50662
rect 22238 50598 22244 50662
rect 22168 50390 22244 50598
rect 22168 50358 22174 50390
rect 21830 50326 21831 50358
rect 21765 50325 21831 50326
rect 22173 50326 22174 50358
rect 22238 50358 22244 50390
rect 22576 50662 22652 50668
rect 22576 50598 22582 50662
rect 22646 50598 22652 50662
rect 22989 50662 23055 50663
rect 22989 50630 22990 50662
rect 22576 50390 22652 50598
rect 22576 50358 22582 50390
rect 22238 50326 22239 50358
rect 22173 50325 22239 50326
rect 22581 50326 22582 50358
rect 22646 50358 22652 50390
rect 22984 50598 22990 50630
rect 23054 50630 23055 50662
rect 23533 50662 23599 50663
rect 23533 50630 23534 50662
rect 23054 50598 23060 50630
rect 22984 50390 23060 50598
rect 22646 50326 22647 50358
rect 22581 50325 22647 50326
rect 22984 50326 22990 50390
rect 23054 50326 23060 50390
rect 22984 50320 23060 50326
rect 23528 50598 23534 50630
rect 23598 50630 23599 50662
rect 23598 50598 23604 50630
rect 23528 50390 23604 50598
rect 110432 50526 110508 50734
rect 115197 50734 115198 50766
rect 115262 50766 115268 50798
rect 115600 51006 115606 51038
rect 115670 51038 115671 51070
rect 116552 51070 116628 51076
rect 115670 51006 115676 51038
rect 115600 50798 115676 51006
rect 115262 50734 115263 50766
rect 115197 50733 115263 50734
rect 115600 50734 115606 50798
rect 115670 50734 115676 50798
rect 116552 51006 116558 51070
rect 116622 51006 116628 51070
rect 116552 50798 116628 51006
rect 116552 50766 116558 50798
rect 115600 50728 115676 50734
rect 116557 50734 116558 50766
rect 116622 50766 116628 50798
rect 116824 51070 116900 51076
rect 116824 51006 116830 51070
rect 116894 51006 116900 51070
rect 116824 50798 116900 51006
rect 116824 50766 116830 50798
rect 116622 50734 116623 50766
rect 116557 50733 116623 50734
rect 116829 50734 116830 50766
rect 116894 50766 116900 50798
rect 137496 50934 137844 52502
rect 137496 50870 137502 50934
rect 137566 50870 137844 50934
rect 116894 50734 116895 50766
rect 116829 50733 116895 50734
rect 110432 50494 110438 50526
rect 110437 50462 110438 50494
rect 110502 50494 110508 50526
rect 115328 50662 115404 50668
rect 115328 50598 115334 50662
rect 115398 50598 115404 50662
rect 115741 50662 115807 50663
rect 115741 50630 115742 50662
rect 110502 50462 110503 50494
rect 110437 50461 110503 50462
rect 23528 50326 23534 50390
rect 23598 50326 23604 50390
rect 115328 50390 115404 50598
rect 115328 50358 115334 50390
rect 23528 50320 23604 50326
rect 115333 50326 115334 50358
rect 115398 50358 115404 50390
rect 115736 50598 115742 50630
rect 115806 50630 115807 50662
rect 116013 50662 116079 50663
rect 116013 50630 116014 50662
rect 115806 50598 115812 50630
rect 115736 50390 115812 50598
rect 115398 50326 115399 50358
rect 115333 50325 115399 50326
rect 115736 50326 115742 50390
rect 115806 50326 115812 50390
rect 115736 50320 115812 50326
rect 116008 50598 116014 50630
rect 116078 50630 116079 50662
rect 116421 50662 116487 50663
rect 116421 50630 116422 50662
rect 116078 50598 116084 50630
rect 116008 50390 116084 50598
rect 116008 50326 116014 50390
rect 116078 50326 116084 50390
rect 116008 50320 116084 50326
rect 116416 50598 116422 50630
rect 116486 50630 116487 50662
rect 116829 50662 116895 50663
rect 116829 50630 116830 50662
rect 116486 50598 116492 50630
rect 116416 50390 116492 50598
rect 116416 50326 116422 50390
rect 116486 50326 116492 50390
rect 116416 50320 116492 50326
rect 116824 50598 116830 50630
rect 116894 50630 116895 50662
rect 116894 50598 116900 50630
rect 116824 50390 116900 50598
rect 116824 50326 116830 50390
rect 116894 50326 116900 50390
rect 116824 50320 116900 50326
rect 21896 50254 21972 50260
rect 21896 50190 21902 50254
rect 21966 50190 21972 50254
rect 21896 49982 21972 50190
rect 21896 49950 21902 49982
rect 21901 49918 21902 49950
rect 21966 49950 21972 49982
rect 22440 50254 22516 50260
rect 22440 50190 22446 50254
rect 22510 50190 22516 50254
rect 23125 50254 23191 50255
rect 23125 50222 23126 50254
rect 22440 49982 22516 50190
rect 22440 49950 22446 49982
rect 21966 49918 21967 49950
rect 21901 49917 21967 49918
rect 22445 49918 22446 49950
rect 22510 49950 22516 49982
rect 23120 50190 23126 50222
rect 23190 50222 23191 50254
rect 23533 50254 23599 50255
rect 23533 50222 23534 50254
rect 23190 50190 23196 50222
rect 23120 49982 23196 50190
rect 22510 49918 22511 49950
rect 22445 49917 22511 49918
rect 23120 49918 23126 49982
rect 23190 49918 23196 49982
rect 23120 49912 23196 49918
rect 23528 50190 23534 50222
rect 23598 50222 23599 50254
rect 115333 50254 115399 50255
rect 115333 50222 115334 50254
rect 23598 50190 23604 50222
rect 23528 49982 23604 50190
rect 23528 49918 23534 49982
rect 23598 49918 23604 49982
rect 23528 49912 23604 49918
rect 115328 50190 115334 50222
rect 115398 50222 115399 50254
rect 115600 50254 115676 50260
rect 115398 50190 115404 50222
rect 115328 49982 115404 50190
rect 115328 49918 115334 49982
rect 115398 49918 115404 49982
rect 115600 50190 115606 50254
rect 115670 50190 115676 50254
rect 115600 49982 115676 50190
rect 115600 49950 115606 49982
rect 115328 49912 115404 49918
rect 115605 49918 115606 49950
rect 115670 49950 115676 49982
rect 116144 50254 116220 50260
rect 116144 50190 116150 50254
rect 116214 50190 116220 50254
rect 116144 49982 116220 50190
rect 116144 49950 116150 49982
rect 115670 49918 115671 49950
rect 115605 49917 115671 49918
rect 116149 49918 116150 49950
rect 116214 49950 116220 49982
rect 116280 50254 116356 50260
rect 116280 50190 116286 50254
rect 116350 50190 116356 50254
rect 116280 49982 116356 50190
rect 116280 49950 116286 49982
rect 116214 49918 116215 49950
rect 116149 49917 116215 49918
rect 116285 49918 116286 49950
rect 116350 49950 116356 49982
rect 116960 50254 117036 50260
rect 116960 50190 116966 50254
rect 117030 50190 117036 50254
rect 116960 49982 117036 50190
rect 116960 49950 116966 49982
rect 116350 49918 116351 49950
rect 116285 49917 116351 49918
rect 116965 49918 116966 49950
rect 117030 49950 117036 49982
rect 117030 49918 117031 49950
rect 116965 49917 117031 49918
rect 21901 49846 21967 49847
rect 21901 49814 21902 49846
rect 21896 49782 21902 49814
rect 21966 49814 21967 49846
rect 22168 49846 22244 49852
rect 21966 49782 21972 49814
rect 21896 49574 21972 49782
rect 21896 49510 21902 49574
rect 21966 49510 21972 49574
rect 22168 49782 22174 49846
rect 22238 49782 22244 49846
rect 22168 49574 22244 49782
rect 22168 49542 22174 49574
rect 21896 49504 21972 49510
rect 22173 49510 22174 49542
rect 22238 49542 22244 49574
rect 22576 49846 22652 49852
rect 22576 49782 22582 49846
rect 22646 49782 22652 49846
rect 22576 49574 22652 49782
rect 22576 49542 22582 49574
rect 22238 49510 22239 49542
rect 22173 49509 22239 49510
rect 22581 49510 22582 49542
rect 22646 49542 22652 49574
rect 22984 49846 23060 49852
rect 22984 49782 22990 49846
rect 23054 49782 23060 49846
rect 22984 49574 23060 49782
rect 22984 49542 22990 49574
rect 22646 49510 22647 49542
rect 22581 49509 22647 49510
rect 22989 49510 22990 49542
rect 23054 49542 23060 49574
rect 23528 49846 23604 49852
rect 23528 49782 23534 49846
rect 23598 49782 23604 49846
rect 23528 49574 23604 49782
rect 23528 49542 23534 49574
rect 23054 49510 23055 49542
rect 22989 49509 23055 49510
rect 23533 49510 23534 49542
rect 23598 49542 23604 49574
rect 115328 49846 115404 49852
rect 115328 49782 115334 49846
rect 115398 49782 115404 49846
rect 115328 49574 115404 49782
rect 115328 49542 115334 49574
rect 23598 49510 23599 49542
rect 23533 49509 23599 49510
rect 115333 49510 115334 49542
rect 115398 49542 115404 49574
rect 115736 49846 115812 49852
rect 115736 49782 115742 49846
rect 115806 49782 115812 49846
rect 116013 49846 116079 49847
rect 116013 49814 116014 49846
rect 115736 49574 115812 49782
rect 115736 49542 115742 49574
rect 115398 49510 115399 49542
rect 115333 49509 115399 49510
rect 115741 49510 115742 49542
rect 115806 49542 115812 49574
rect 116008 49782 116014 49814
rect 116078 49814 116079 49846
rect 116965 49846 117031 49847
rect 116965 49814 116966 49846
rect 116078 49782 116084 49814
rect 116008 49574 116084 49782
rect 115806 49510 115807 49542
rect 115741 49509 115807 49510
rect 116008 49510 116014 49574
rect 116078 49510 116084 49574
rect 116008 49504 116084 49510
rect 116960 49782 116966 49814
rect 117030 49814 117031 49846
rect 117030 49782 117036 49814
rect 116960 49574 117036 49782
rect 116960 49510 116966 49574
rect 117030 49510 117036 49574
rect 116960 49504 117036 49510
rect 952 49102 1230 49166
rect 1294 49102 1300 49166
rect 21760 49438 21836 49444
rect 21760 49374 21766 49438
rect 21830 49374 21836 49438
rect 21760 49166 21836 49374
rect 21760 49134 21766 49166
rect 952 47398 1300 49102
rect 21765 49102 21766 49134
rect 21830 49134 21836 49166
rect 22576 49438 22652 49444
rect 22576 49374 22582 49438
rect 22646 49374 22652 49438
rect 22989 49438 23055 49439
rect 22989 49406 22990 49438
rect 22576 49166 22652 49374
rect 22576 49134 22582 49166
rect 21830 49102 21831 49134
rect 21765 49101 21831 49102
rect 22581 49102 22582 49134
rect 22646 49134 22652 49166
rect 22984 49374 22990 49406
rect 23054 49406 23055 49438
rect 23528 49438 23604 49444
rect 23054 49374 23060 49406
rect 22984 49166 23060 49374
rect 22646 49102 22647 49134
rect 22581 49101 22647 49102
rect 22984 49102 22990 49166
rect 23054 49102 23060 49166
rect 23528 49374 23534 49438
rect 23598 49374 23604 49438
rect 115333 49438 115399 49439
rect 115333 49406 115334 49438
rect 23528 49166 23604 49374
rect 23528 49134 23534 49166
rect 22984 49096 23060 49102
rect 23533 49102 23534 49134
rect 23598 49134 23604 49166
rect 115328 49374 115334 49406
rect 115398 49406 115399 49438
rect 115741 49438 115807 49439
rect 115741 49406 115742 49438
rect 115398 49374 115404 49406
rect 115328 49166 115404 49374
rect 23598 49102 23599 49134
rect 23533 49101 23599 49102
rect 115328 49102 115334 49166
rect 115398 49102 115404 49166
rect 115328 49096 115404 49102
rect 115736 49374 115742 49406
rect 115806 49406 115807 49438
rect 116421 49438 116487 49439
rect 116421 49406 116422 49438
rect 115806 49374 115812 49406
rect 115736 49166 115812 49374
rect 115736 49102 115742 49166
rect 115806 49102 115812 49166
rect 115736 49096 115812 49102
rect 116416 49374 116422 49406
rect 116486 49406 116487 49438
rect 116824 49438 116900 49444
rect 116486 49374 116492 49406
rect 116416 49166 116492 49374
rect 116416 49102 116422 49166
rect 116486 49102 116492 49166
rect 116824 49374 116830 49438
rect 116894 49374 116900 49438
rect 116824 49166 116900 49374
rect 116824 49134 116830 49166
rect 116416 49096 116492 49102
rect 116829 49102 116830 49134
rect 116894 49134 116900 49166
rect 116894 49102 116895 49134
rect 116829 49101 116895 49102
rect 21896 49030 21972 49036
rect 21896 48966 21902 49030
rect 21966 48966 21972 49030
rect 21896 48758 21972 48966
rect 21896 48726 21902 48758
rect 21901 48694 21902 48726
rect 21966 48726 21972 48758
rect 22712 49030 22788 49036
rect 22712 48966 22718 49030
rect 22782 48966 22788 49030
rect 22712 48758 22788 48966
rect 22712 48726 22718 48758
rect 21966 48694 21967 48726
rect 21901 48693 21967 48694
rect 22717 48694 22718 48726
rect 22782 48726 22788 48758
rect 23120 49030 23196 49036
rect 23120 48966 23126 49030
rect 23190 48966 23196 49030
rect 23397 49030 23463 49031
rect 23397 48998 23398 49030
rect 23120 48758 23196 48966
rect 23120 48726 23126 48758
rect 22782 48694 22783 48726
rect 22717 48693 22783 48694
rect 23125 48694 23126 48726
rect 23190 48726 23196 48758
rect 23392 48966 23398 48998
rect 23462 48998 23463 49030
rect 115197 49030 115263 49031
rect 115197 48998 115198 49030
rect 23462 48966 23468 48998
rect 23392 48758 23468 48966
rect 23190 48694 23191 48726
rect 23125 48693 23191 48694
rect 23392 48694 23398 48758
rect 23462 48694 23468 48758
rect 23392 48688 23468 48694
rect 115192 48966 115198 48998
rect 115262 48998 115263 49030
rect 115600 49030 115676 49036
rect 115262 48966 115268 48998
rect 115192 48758 115268 48966
rect 115192 48694 115198 48758
rect 115262 48694 115268 48758
rect 115600 48966 115606 49030
rect 115670 48966 115676 49030
rect 115600 48758 115676 48966
rect 115600 48726 115606 48758
rect 115192 48688 115268 48694
rect 115605 48694 115606 48726
rect 115670 48726 115676 48758
rect 116552 49030 116628 49036
rect 116552 48966 116558 49030
rect 116622 48966 116628 49030
rect 116965 49030 117031 49031
rect 116965 48998 116966 49030
rect 116552 48758 116628 48966
rect 116552 48726 116558 48758
rect 115670 48694 115671 48726
rect 115605 48693 115671 48694
rect 116557 48694 116558 48726
rect 116622 48726 116628 48758
rect 116960 48966 116966 48998
rect 117030 48998 117031 49030
rect 137496 49030 137844 50870
rect 117030 48966 117036 48998
rect 116960 48758 117036 48966
rect 116622 48694 116623 48726
rect 116557 48693 116623 48694
rect 116960 48694 116966 48758
rect 117030 48694 117036 48758
rect 116960 48688 117036 48694
rect 137496 48966 137502 49030
rect 137566 48966 137844 49030
rect 22309 48622 22375 48623
rect 22309 48590 22310 48622
rect 22304 48558 22310 48590
rect 22374 48590 22375 48622
rect 23125 48622 23191 48623
rect 23125 48590 23126 48622
rect 22374 48558 22380 48590
rect 21765 48350 21831 48351
rect 21765 48318 21766 48350
rect 21760 48286 21766 48318
rect 21830 48318 21831 48350
rect 22304 48350 22380 48558
rect 21830 48286 21836 48318
rect 21760 48078 21836 48286
rect 22304 48286 22310 48350
rect 22374 48286 22380 48350
rect 22304 48280 22380 48286
rect 23120 48558 23126 48590
rect 23190 48590 23191 48622
rect 23397 48622 23463 48623
rect 23397 48590 23398 48622
rect 23190 48558 23196 48590
rect 23120 48350 23196 48558
rect 23120 48286 23126 48350
rect 23190 48286 23196 48350
rect 23120 48280 23196 48286
rect 23392 48558 23398 48590
rect 23462 48590 23463 48622
rect 115328 48622 115404 48628
rect 23462 48558 23468 48590
rect 23392 48350 23468 48558
rect 23392 48286 23398 48350
rect 23462 48286 23468 48350
rect 115328 48558 115334 48622
rect 115398 48558 115404 48622
rect 115328 48350 115404 48558
rect 115328 48318 115334 48350
rect 23392 48280 23468 48286
rect 115333 48286 115334 48318
rect 115398 48318 115404 48350
rect 115736 48622 115812 48628
rect 115736 48558 115742 48622
rect 115806 48558 115812 48622
rect 116149 48622 116215 48623
rect 116149 48590 116150 48622
rect 115736 48350 115812 48558
rect 115736 48318 115742 48350
rect 115398 48286 115399 48318
rect 115333 48285 115399 48286
rect 115741 48286 115742 48318
rect 115806 48318 115812 48350
rect 116144 48558 116150 48590
rect 116214 48590 116215 48622
rect 116280 48622 116356 48628
rect 116214 48558 116220 48590
rect 116144 48350 116220 48558
rect 115806 48286 115807 48318
rect 115741 48285 115807 48286
rect 116144 48286 116150 48350
rect 116214 48286 116220 48350
rect 116280 48558 116286 48622
rect 116350 48558 116356 48622
rect 116280 48350 116356 48558
rect 116280 48318 116286 48350
rect 116144 48280 116220 48286
rect 116285 48286 116286 48318
rect 116350 48318 116356 48350
rect 116829 48350 116895 48351
rect 116829 48318 116830 48350
rect 116350 48286 116351 48318
rect 116285 48285 116351 48286
rect 116824 48286 116830 48318
rect 116894 48318 116895 48350
rect 116894 48286 116900 48318
rect 21760 48014 21766 48078
rect 21830 48014 21836 48078
rect 21760 48008 21836 48014
rect 22984 48214 23060 48220
rect 22984 48150 22990 48214
rect 23054 48150 23060 48214
rect 22984 47942 23060 48150
rect 22984 47910 22990 47942
rect 22989 47878 22990 47910
rect 23054 47910 23060 47942
rect 23392 48214 23468 48220
rect 23392 48150 23398 48214
rect 23462 48150 23468 48214
rect 23392 47942 23468 48150
rect 23392 47910 23398 47942
rect 23054 47878 23055 47910
rect 22989 47877 23055 47878
rect 23397 47878 23398 47910
rect 23462 47910 23468 47942
rect 115192 48214 115268 48220
rect 115192 48150 115198 48214
rect 115262 48150 115268 48214
rect 115741 48214 115807 48215
rect 115741 48182 115742 48214
rect 115192 47942 115268 48150
rect 115192 47910 115198 47942
rect 23462 47878 23463 47910
rect 23397 47877 23463 47878
rect 115197 47878 115198 47910
rect 115262 47910 115268 47942
rect 115736 48150 115742 48182
rect 115806 48182 115807 48214
rect 116149 48214 116215 48215
rect 116149 48182 116150 48214
rect 115806 48150 115812 48182
rect 115736 47942 115812 48150
rect 116144 48150 116150 48182
rect 116214 48182 116215 48214
rect 116214 48150 116220 48182
rect 116144 48084 116220 48150
rect 116144 48078 116356 48084
rect 116144 48014 116286 48078
rect 116350 48014 116356 48078
rect 116144 48008 116356 48014
rect 116824 48078 116900 48286
rect 116824 48014 116830 48078
rect 116894 48014 116900 48078
rect 116824 48008 116900 48014
rect 115262 47878 115263 47910
rect 115197 47877 115263 47878
rect 115736 47878 115742 47942
rect 115806 47878 115812 47942
rect 115736 47872 115812 47878
rect 22712 47806 22788 47812
rect 22712 47742 22718 47806
rect 22782 47742 22788 47806
rect 116557 47806 116623 47807
rect 116557 47774 116558 47806
rect 952 47334 1230 47398
rect 1294 47334 1300 47398
rect 952 45630 1300 47334
rect 21760 47534 21836 47540
rect 21760 47470 21766 47534
rect 21830 47470 21836 47534
rect 22712 47534 22788 47742
rect 116552 47742 116558 47774
rect 116622 47774 116623 47806
rect 116622 47742 116628 47774
rect 22712 47502 22718 47534
rect 21760 47262 21836 47470
rect 22717 47470 22718 47502
rect 22782 47502 22788 47534
rect 110160 47670 110236 47676
rect 110160 47606 110166 47670
rect 110230 47606 110236 47670
rect 22782 47470 22783 47502
rect 22717 47469 22783 47470
rect 110160 47398 110236 47606
rect 116552 47534 116628 47742
rect 116552 47470 116558 47534
rect 116622 47470 116628 47534
rect 116965 47534 117031 47535
rect 116965 47502 116966 47534
rect 116552 47464 116628 47470
rect 116960 47470 116966 47502
rect 117030 47502 117031 47534
rect 137496 47534 137844 48966
rect 117030 47470 117036 47502
rect 110160 47366 110166 47398
rect 110165 47334 110166 47366
rect 110230 47366 110236 47398
rect 110230 47334 110231 47366
rect 110165 47333 110231 47334
rect 21760 47230 21766 47262
rect 21765 47198 21766 47230
rect 21830 47230 21836 47262
rect 28288 47262 28364 47268
rect 21830 47198 21831 47230
rect 21765 47197 21831 47198
rect 28288 47198 28294 47262
rect 28358 47198 28364 47262
rect 110301 47262 110367 47263
rect 110301 47230 110302 47262
rect 21765 47126 21831 47127
rect 21765 47094 21766 47126
rect 21760 47062 21766 47094
rect 21830 47094 21831 47126
rect 22445 47126 22511 47127
rect 22445 47094 22446 47126
rect 21830 47062 21836 47094
rect 21760 46854 21836 47062
rect 21760 46790 21766 46854
rect 21830 46790 21836 46854
rect 21760 46784 21836 46790
rect 22440 47062 22446 47094
rect 22510 47094 22511 47126
rect 22510 47062 22516 47094
rect 22440 46854 22516 47062
rect 28288 46990 28364 47198
rect 28288 46958 28294 46990
rect 28293 46926 28294 46958
rect 28358 46958 28364 46990
rect 110296 47198 110302 47230
rect 110366 47230 110367 47262
rect 116960 47262 117036 47470
rect 110366 47198 110372 47230
rect 110296 46990 110372 47198
rect 116960 47198 116966 47262
rect 117030 47198 117036 47262
rect 116960 47192 117036 47198
rect 137496 47470 137502 47534
rect 137566 47470 137844 47534
rect 116149 47126 116215 47127
rect 116149 47094 116150 47126
rect 28358 46926 28359 46958
rect 28293 46925 28359 46926
rect 110296 46926 110302 46990
rect 110366 46926 110372 46990
rect 110296 46920 110372 46926
rect 116144 47062 116150 47094
rect 116214 47094 116215 47126
rect 116285 47126 116351 47127
rect 116285 47094 116286 47126
rect 116214 47062 116220 47094
rect 22440 46790 22446 46854
rect 22510 46790 22516 46854
rect 22440 46784 22516 46790
rect 110432 46854 110508 46860
rect 110432 46790 110438 46854
rect 110502 46790 110508 46854
rect 21901 46718 21967 46719
rect 21901 46686 21902 46718
rect 21896 46654 21902 46686
rect 21966 46686 21967 46718
rect 22989 46718 23055 46719
rect 22989 46686 22990 46718
rect 21966 46654 21972 46686
rect 21896 46446 21972 46654
rect 21896 46382 21902 46446
rect 21966 46382 21972 46446
rect 21896 46376 21972 46382
rect 22984 46654 22990 46686
rect 23054 46686 23055 46718
rect 23392 46718 23468 46724
rect 23054 46654 23060 46686
rect 22984 46446 23060 46654
rect 22984 46382 22990 46446
rect 23054 46382 23060 46446
rect 23392 46654 23398 46718
rect 23462 46654 23468 46718
rect 23392 46446 23468 46654
rect 110432 46582 110508 46790
rect 116144 46854 116220 47062
rect 116144 46790 116150 46854
rect 116214 46790 116220 46854
rect 116144 46784 116220 46790
rect 116280 47062 116286 47094
rect 116350 47094 116351 47126
rect 116829 47126 116895 47127
rect 116829 47094 116830 47126
rect 116350 47062 116356 47094
rect 116280 46854 116356 47062
rect 116280 46790 116286 46854
rect 116350 46790 116356 46854
rect 116280 46784 116356 46790
rect 116824 47062 116830 47094
rect 116894 47094 116895 47126
rect 116894 47062 116900 47094
rect 116824 46854 116900 47062
rect 116824 46790 116830 46854
rect 116894 46790 116900 46854
rect 116824 46784 116900 46790
rect 115197 46718 115263 46719
rect 115197 46686 115198 46718
rect 110432 46550 110438 46582
rect 110437 46518 110438 46550
rect 110502 46550 110508 46582
rect 115192 46654 115198 46686
rect 115262 46686 115263 46718
rect 115605 46718 115671 46719
rect 115605 46686 115606 46718
rect 115262 46654 115268 46686
rect 110502 46518 110503 46550
rect 110437 46517 110503 46518
rect 23392 46414 23398 46446
rect 22984 46376 23060 46382
rect 23397 46382 23398 46414
rect 23462 46414 23468 46446
rect 28288 46446 28364 46452
rect 23462 46382 23463 46414
rect 23397 46381 23463 46382
rect 28288 46382 28294 46446
rect 28358 46382 28364 46446
rect 21760 46310 21836 46316
rect 21760 46246 21766 46310
rect 21830 46246 21836 46310
rect 22173 46310 22239 46311
rect 22173 46278 22174 46310
rect 21760 46038 21836 46246
rect 21760 46006 21766 46038
rect 21765 45974 21766 46006
rect 21830 46006 21836 46038
rect 22168 46246 22174 46278
rect 22238 46278 22239 46310
rect 23120 46310 23196 46316
rect 22238 46246 22244 46278
rect 22168 46038 22244 46246
rect 21830 45974 21831 46006
rect 21765 45973 21831 45974
rect 22168 45974 22174 46038
rect 22238 45974 22244 46038
rect 23120 46246 23126 46310
rect 23190 46246 23196 46310
rect 23533 46310 23599 46311
rect 23533 46278 23534 46310
rect 23120 46038 23196 46246
rect 23120 46006 23126 46038
rect 22168 45968 22244 45974
rect 23125 45974 23126 46006
rect 23190 46006 23196 46038
rect 23528 46246 23534 46278
rect 23598 46278 23599 46310
rect 23598 46246 23604 46278
rect 23528 46038 23604 46246
rect 23190 45974 23191 46006
rect 23125 45973 23191 45974
rect 23528 45974 23534 46038
rect 23598 45974 23604 46038
rect 28288 46038 28364 46382
rect 115192 46446 115268 46654
rect 115192 46382 115198 46446
rect 115262 46382 115268 46446
rect 115192 46376 115268 46382
rect 115600 46654 115606 46686
rect 115670 46686 115671 46718
rect 116824 46718 116900 46724
rect 115670 46654 115676 46686
rect 115600 46446 115676 46654
rect 115600 46382 115606 46446
rect 115670 46382 115676 46446
rect 116824 46654 116830 46718
rect 116894 46654 116900 46718
rect 116824 46446 116900 46654
rect 116824 46414 116830 46446
rect 115600 46376 115676 46382
rect 116829 46382 116830 46414
rect 116894 46414 116900 46446
rect 116894 46382 116895 46414
rect 116829 46381 116895 46382
rect 28288 46006 28294 46038
rect 23528 45968 23604 45974
rect 28293 45974 28294 46006
rect 28358 46006 28364 46038
rect 115328 46310 115404 46316
rect 115328 46246 115334 46310
rect 115398 46246 115404 46310
rect 115741 46310 115807 46311
rect 115741 46278 115742 46310
rect 115328 46038 115404 46246
rect 115328 46006 115334 46038
rect 28358 45974 28359 46006
rect 28293 45973 28359 45974
rect 115333 45974 115334 46006
rect 115398 46006 115404 46038
rect 115736 46246 115742 46278
rect 115806 46278 115807 46310
rect 116013 46310 116079 46311
rect 116013 46278 116014 46310
rect 115806 46246 115812 46278
rect 115736 46038 115812 46246
rect 115398 45974 115399 46006
rect 115333 45973 115399 45974
rect 115736 45974 115742 46038
rect 115806 45974 115812 46038
rect 115736 45968 115812 45974
rect 116008 46246 116014 46278
rect 116078 46278 116079 46310
rect 116824 46310 116900 46316
rect 116078 46246 116084 46278
rect 116008 46038 116084 46246
rect 116008 45974 116014 46038
rect 116078 45974 116084 46038
rect 116824 46246 116830 46310
rect 116894 46246 116900 46310
rect 116824 46038 116900 46246
rect 116824 46006 116830 46038
rect 116008 45968 116084 45974
rect 116829 45974 116830 46006
rect 116894 46006 116900 46038
rect 116894 45974 116895 46006
rect 116829 45973 116895 45974
rect 952 45566 1230 45630
rect 1294 45566 1300 45630
rect 21896 45902 21972 45908
rect 21896 45838 21902 45902
rect 21966 45838 21972 45902
rect 21896 45630 21972 45838
rect 21896 45598 21902 45630
rect 952 44134 1300 45566
rect 21901 45566 21902 45598
rect 21966 45598 21972 45630
rect 22304 45902 22380 45908
rect 22304 45838 22310 45902
rect 22374 45838 22380 45902
rect 23125 45902 23191 45903
rect 23125 45870 23126 45902
rect 22304 45630 22380 45838
rect 22304 45598 22310 45630
rect 21966 45566 21967 45598
rect 21901 45565 21967 45566
rect 22309 45566 22310 45598
rect 22374 45598 22380 45630
rect 23120 45838 23126 45870
rect 23190 45870 23191 45902
rect 23392 45902 23468 45908
rect 23190 45838 23196 45870
rect 23120 45630 23196 45838
rect 22374 45566 22375 45598
rect 22309 45565 22375 45566
rect 23120 45566 23126 45630
rect 23190 45566 23196 45630
rect 23392 45838 23398 45902
rect 23462 45838 23468 45902
rect 23392 45630 23468 45838
rect 23392 45598 23398 45630
rect 23120 45560 23196 45566
rect 23397 45566 23398 45598
rect 23462 45598 23468 45630
rect 115192 45902 115268 45908
rect 115192 45838 115198 45902
rect 115262 45838 115268 45902
rect 115192 45630 115268 45838
rect 115192 45598 115198 45630
rect 23462 45566 23463 45598
rect 23397 45565 23463 45566
rect 115197 45566 115198 45598
rect 115262 45598 115268 45630
rect 115600 45902 115676 45908
rect 115600 45838 115606 45902
rect 115670 45838 115676 45902
rect 116421 45902 116487 45903
rect 116421 45870 116422 45902
rect 115600 45630 115676 45838
rect 115600 45598 115606 45630
rect 115262 45566 115263 45598
rect 115197 45565 115263 45566
rect 115605 45566 115606 45598
rect 115670 45598 115676 45630
rect 116416 45838 116422 45870
rect 116486 45870 116487 45902
rect 116960 45902 117036 45908
rect 116486 45838 116492 45870
rect 116416 45630 116492 45838
rect 115670 45566 115671 45598
rect 115605 45565 115671 45566
rect 116416 45566 116422 45630
rect 116486 45566 116492 45630
rect 116960 45838 116966 45902
rect 117030 45838 117036 45902
rect 116960 45630 117036 45838
rect 116960 45598 116966 45630
rect 116416 45560 116492 45566
rect 116965 45566 116966 45598
rect 117030 45598 117036 45630
rect 137496 45630 137844 47470
rect 117030 45566 117031 45598
rect 116965 45565 117031 45566
rect 137496 45566 137502 45630
rect 137566 45566 137844 45630
rect 21901 45494 21967 45495
rect 21901 45462 21902 45494
rect 21896 45430 21902 45462
rect 21966 45462 21967 45494
rect 22576 45494 22652 45500
rect 21966 45430 21972 45462
rect 21896 45222 21972 45430
rect 21896 45158 21902 45222
rect 21966 45158 21972 45222
rect 22576 45430 22582 45494
rect 22646 45430 22652 45494
rect 22989 45494 23055 45495
rect 22989 45462 22990 45494
rect 22576 45222 22652 45430
rect 22576 45190 22582 45222
rect 21896 45152 21972 45158
rect 22581 45158 22582 45190
rect 22646 45190 22652 45222
rect 22984 45430 22990 45462
rect 23054 45462 23055 45494
rect 23397 45494 23463 45495
rect 23397 45462 23398 45494
rect 23054 45430 23060 45462
rect 22984 45222 23060 45430
rect 22646 45158 22647 45190
rect 22581 45157 22647 45158
rect 22984 45158 22990 45222
rect 23054 45158 23060 45222
rect 22984 45152 23060 45158
rect 23392 45430 23398 45462
rect 23462 45462 23463 45494
rect 115328 45494 115404 45500
rect 23462 45430 23468 45462
rect 23392 45222 23468 45430
rect 23392 45158 23398 45222
rect 23462 45158 23468 45222
rect 115328 45430 115334 45494
rect 115398 45430 115404 45494
rect 115328 45222 115404 45430
rect 115328 45190 115334 45222
rect 23392 45152 23468 45158
rect 115333 45158 115334 45190
rect 115398 45190 115404 45222
rect 115736 45494 115812 45500
rect 115736 45430 115742 45494
rect 115806 45430 115812 45494
rect 116149 45494 116215 45495
rect 116149 45462 116150 45494
rect 115736 45222 115812 45430
rect 115736 45190 115742 45222
rect 115398 45158 115399 45190
rect 115333 45157 115399 45158
rect 115741 45158 115742 45190
rect 115806 45190 115812 45222
rect 116144 45430 116150 45462
rect 116214 45462 116215 45494
rect 116285 45494 116351 45495
rect 116285 45462 116286 45494
rect 116214 45430 116220 45462
rect 116144 45222 116220 45430
rect 115806 45158 115807 45190
rect 115741 45157 115807 45158
rect 116144 45158 116150 45222
rect 116214 45158 116220 45222
rect 116144 45152 116220 45158
rect 116280 45430 116286 45462
rect 116350 45462 116351 45494
rect 116965 45494 117031 45495
rect 116965 45462 116966 45494
rect 116350 45430 116356 45462
rect 116280 45222 116356 45430
rect 116280 45158 116286 45222
rect 116350 45158 116356 45222
rect 116280 45152 116356 45158
rect 116960 45430 116966 45462
rect 117030 45462 117031 45494
rect 117030 45430 117036 45462
rect 116960 45222 117036 45430
rect 116960 45158 116966 45222
rect 117030 45158 117036 45222
rect 116960 45152 117036 45158
rect 21760 45086 21836 45092
rect 21760 45022 21766 45086
rect 21830 45022 21836 45086
rect 21760 44814 21836 45022
rect 21760 44782 21766 44814
rect 21765 44750 21766 44782
rect 21830 44782 21836 44814
rect 22168 45086 22244 45092
rect 22168 45022 22174 45086
rect 22238 45022 22244 45086
rect 22581 45086 22647 45087
rect 22581 45054 22582 45086
rect 22168 44814 22244 45022
rect 22168 44782 22174 44814
rect 21830 44750 21831 44782
rect 21765 44749 21831 44750
rect 22173 44750 22174 44782
rect 22238 44782 22244 44814
rect 22576 45022 22582 45054
rect 22646 45054 22647 45086
rect 22989 45086 23055 45087
rect 22989 45054 22990 45086
rect 22646 45022 22652 45054
rect 22576 44814 22652 45022
rect 22238 44750 22239 44782
rect 22173 44749 22239 44750
rect 22576 44750 22582 44814
rect 22646 44750 22652 44814
rect 22576 44744 22652 44750
rect 22984 45022 22990 45054
rect 23054 45054 23055 45086
rect 23528 45086 23604 45092
rect 23054 45022 23060 45054
rect 22984 44814 23060 45022
rect 22984 44750 22990 44814
rect 23054 44750 23060 44814
rect 23528 45022 23534 45086
rect 23598 45022 23604 45086
rect 115333 45086 115399 45087
rect 115333 45054 115334 45086
rect 23528 44814 23604 45022
rect 23528 44782 23534 44814
rect 22984 44744 23060 44750
rect 23533 44750 23534 44782
rect 23598 44782 23604 44814
rect 115328 45022 115334 45054
rect 115398 45054 115399 45086
rect 115741 45086 115807 45087
rect 115741 45054 115742 45086
rect 115398 45022 115404 45054
rect 115328 44814 115404 45022
rect 23598 44750 23599 44782
rect 23533 44749 23599 44750
rect 115328 44750 115334 44814
rect 115398 44750 115404 44814
rect 115328 44744 115404 44750
rect 115736 45022 115742 45054
rect 115806 45054 115807 45086
rect 116421 45086 116487 45087
rect 116421 45054 116422 45086
rect 115806 45022 115812 45054
rect 115736 44814 115812 45022
rect 115736 44750 115742 44814
rect 115806 44750 115812 44814
rect 115736 44744 115812 44750
rect 116416 45022 116422 45054
rect 116486 45054 116487 45086
rect 116824 45086 116900 45092
rect 116486 45022 116492 45054
rect 116416 44814 116492 45022
rect 116416 44750 116422 44814
rect 116486 44750 116492 44814
rect 116824 45022 116830 45086
rect 116894 45022 116900 45086
rect 116824 44814 116900 45022
rect 116824 44782 116830 44814
rect 116416 44744 116492 44750
rect 116829 44750 116830 44782
rect 116894 44782 116900 44814
rect 116894 44750 116895 44782
rect 116829 44749 116895 44750
rect 22309 44678 22375 44679
rect 22309 44646 22310 44678
rect 22304 44614 22310 44646
rect 22374 44646 22375 44678
rect 22717 44678 22783 44679
rect 22717 44646 22718 44678
rect 22374 44614 22380 44646
rect 22304 44406 22380 44614
rect 22304 44342 22310 44406
rect 22374 44342 22380 44406
rect 22304 44336 22380 44342
rect 22712 44614 22718 44646
rect 22782 44646 22783 44678
rect 23120 44678 23196 44684
rect 22782 44614 22788 44646
rect 22712 44406 22788 44614
rect 22712 44342 22718 44406
rect 22782 44342 22788 44406
rect 23120 44614 23126 44678
rect 23190 44614 23196 44678
rect 23120 44406 23196 44614
rect 23120 44374 23126 44406
rect 22712 44336 22788 44342
rect 23125 44342 23126 44374
rect 23190 44374 23196 44406
rect 23392 44678 23468 44684
rect 23392 44614 23398 44678
rect 23462 44614 23468 44678
rect 23392 44406 23468 44614
rect 115192 44678 115268 44684
rect 115192 44614 115198 44678
rect 115262 44614 115268 44678
rect 110165 44542 110231 44543
rect 110165 44510 110166 44542
rect 23392 44374 23398 44406
rect 23190 44342 23191 44374
rect 23125 44341 23191 44342
rect 23397 44342 23398 44374
rect 23462 44374 23468 44406
rect 110160 44478 110166 44510
rect 110230 44510 110231 44542
rect 110230 44478 110236 44510
rect 23462 44342 23463 44374
rect 23397 44341 23463 44342
rect 952 44070 1230 44134
rect 1294 44070 1300 44134
rect 952 42502 1300 44070
rect 22984 44270 23060 44276
rect 22984 44206 22990 44270
rect 23054 44206 23060 44270
rect 23397 44270 23463 44271
rect 23397 44238 23398 44270
rect 22984 43998 23060 44206
rect 22984 43966 22990 43998
rect 22989 43934 22990 43966
rect 23054 43966 23060 43998
rect 23392 44206 23398 44238
rect 23462 44238 23463 44270
rect 110160 44270 110236 44478
rect 115192 44406 115268 44614
rect 115192 44374 115198 44406
rect 115197 44342 115198 44374
rect 115262 44374 115268 44406
rect 115600 44678 115676 44684
rect 115600 44614 115606 44678
rect 115670 44614 115676 44678
rect 115600 44406 115676 44614
rect 116552 44678 116628 44684
rect 116552 44614 116558 44678
rect 116622 44614 116628 44678
rect 115600 44374 115606 44406
rect 115262 44342 115263 44374
rect 115197 44341 115263 44342
rect 115605 44342 115606 44374
rect 115670 44374 115676 44406
rect 116285 44406 116351 44407
rect 116285 44374 116286 44406
rect 115670 44342 115671 44374
rect 115605 44341 115671 44342
rect 116280 44342 116286 44374
rect 116350 44374 116351 44406
rect 116552 44406 116628 44614
rect 116552 44374 116558 44406
rect 116350 44342 116356 44374
rect 23462 44206 23468 44238
rect 23392 43998 23468 44206
rect 110160 44206 110166 44270
rect 110230 44206 110236 44270
rect 115197 44270 115263 44271
rect 115197 44238 115198 44270
rect 110160 44200 110236 44206
rect 115192 44206 115198 44238
rect 115262 44238 115263 44270
rect 115605 44270 115671 44271
rect 115605 44238 115606 44270
rect 115262 44206 115268 44238
rect 23054 43934 23055 43966
rect 22989 43933 23055 43934
rect 23392 43934 23398 43998
rect 23462 43934 23468 43998
rect 23392 43928 23468 43934
rect 115192 43998 115268 44206
rect 115192 43934 115198 43998
rect 115262 43934 115268 43998
rect 115192 43928 115268 43934
rect 115600 44206 115606 44238
rect 115670 44238 115671 44270
rect 115670 44206 115676 44238
rect 115600 43998 115676 44206
rect 116280 44134 116356 44342
rect 116557 44342 116558 44374
rect 116622 44374 116628 44406
rect 116622 44342 116623 44374
rect 116557 44341 116623 44342
rect 116280 44070 116286 44134
rect 116350 44070 116356 44134
rect 116280 44064 116356 44070
rect 137496 44134 137844 45566
rect 137496 44070 137502 44134
rect 137566 44070 137844 44134
rect 115600 43934 115606 43998
rect 115670 43934 115676 43998
rect 115600 43928 115676 43934
rect 22173 43862 22239 43863
rect 22173 43830 22174 43862
rect 22168 43798 22174 43830
rect 22238 43830 22239 43862
rect 22581 43862 22647 43863
rect 22581 43830 22582 43862
rect 22238 43798 22244 43830
rect 21901 43590 21967 43591
rect 21901 43558 21902 43590
rect 21896 43526 21902 43558
rect 21966 43558 21967 43590
rect 22168 43590 22244 43798
rect 22576 43798 22582 43830
rect 22646 43830 22647 43862
rect 22984 43862 23060 43868
rect 22646 43798 22652 43830
rect 21966 43526 21972 43558
rect 21896 43318 21972 43526
rect 22168 43526 22174 43590
rect 22238 43526 22244 43590
rect 22445 43590 22511 43591
rect 22445 43558 22446 43590
rect 22168 43520 22244 43526
rect 22440 43526 22446 43558
rect 22510 43558 22511 43590
rect 22576 43590 22652 43798
rect 22510 43526 22516 43558
rect 21896 43254 21902 43318
rect 21966 43254 21972 43318
rect 21896 43248 21972 43254
rect 22440 43324 22516 43526
rect 22576 43526 22582 43590
rect 22646 43526 22652 43590
rect 22984 43798 22990 43862
rect 23054 43798 23060 43862
rect 22984 43590 23060 43798
rect 22984 43558 22990 43590
rect 22576 43520 22652 43526
rect 22989 43526 22990 43558
rect 23054 43558 23060 43590
rect 23392 43862 23468 43868
rect 23392 43798 23398 43862
rect 23462 43798 23468 43862
rect 23392 43590 23468 43798
rect 115192 43862 115268 43868
rect 115192 43798 115198 43862
rect 115262 43798 115268 43862
rect 23392 43558 23398 43590
rect 23054 43526 23055 43558
rect 22989 43525 23055 43526
rect 23397 43526 23398 43558
rect 23462 43558 23468 43590
rect 110432 43726 110508 43732
rect 110432 43662 110438 43726
rect 110502 43662 110508 43726
rect 23462 43526 23463 43558
rect 23397 43525 23463 43526
rect 110432 43454 110508 43662
rect 115192 43590 115268 43798
rect 115192 43558 115198 43590
rect 115197 43526 115198 43558
rect 115262 43558 115268 43590
rect 115600 43862 115676 43868
rect 115600 43798 115606 43862
rect 115670 43798 115676 43862
rect 115600 43590 115676 43798
rect 115600 43558 115606 43590
rect 115262 43526 115263 43558
rect 115197 43525 115263 43526
rect 115605 43526 115606 43558
rect 115670 43558 115676 43590
rect 116008 43862 116084 43868
rect 116008 43798 116014 43862
rect 116078 43798 116084 43862
rect 116008 43590 116084 43798
rect 116008 43558 116014 43590
rect 115670 43526 115671 43558
rect 115605 43525 115671 43526
rect 116013 43526 116014 43558
rect 116078 43558 116084 43590
rect 116552 43862 116628 43868
rect 116552 43798 116558 43862
rect 116622 43798 116628 43862
rect 116552 43590 116628 43798
rect 116552 43558 116558 43590
rect 116078 43526 116079 43558
rect 116013 43525 116079 43526
rect 116557 43526 116558 43558
rect 116622 43558 116628 43590
rect 116960 43590 117036 43596
rect 116622 43526 116623 43558
rect 116557 43525 116623 43526
rect 116960 43526 116966 43590
rect 117030 43526 117036 43590
rect 110432 43422 110438 43454
rect 110437 43390 110438 43422
rect 110502 43422 110508 43454
rect 110502 43390 110503 43422
rect 110437 43389 110503 43390
rect 22440 43318 22652 43324
rect 22440 43254 22582 43318
rect 22646 43254 22652 43318
rect 28293 43318 28359 43319
rect 28293 43286 28294 43318
rect 22440 43248 22652 43254
rect 28288 43254 28294 43286
rect 28358 43286 28359 43318
rect 110160 43318 110236 43324
rect 28358 43254 28364 43286
rect 21760 43182 21836 43188
rect 21760 43118 21766 43182
rect 21830 43118 21836 43182
rect 22445 43182 22511 43183
rect 22445 43150 22446 43182
rect 21760 42910 21836 43118
rect 21760 42878 21766 42910
rect 21765 42846 21766 42878
rect 21830 42878 21836 42910
rect 22440 43118 22446 43150
rect 22510 43150 22511 43182
rect 22510 43118 22516 43150
rect 22440 42910 22516 43118
rect 28288 43046 28364 43254
rect 28288 42982 28294 43046
rect 28358 42982 28364 43046
rect 110160 43254 110166 43318
rect 110230 43254 110236 43318
rect 116960 43318 117036 43526
rect 116960 43286 116966 43318
rect 110160 43046 110236 43254
rect 116965 43254 116966 43286
rect 117030 43286 117036 43318
rect 117030 43254 117031 43286
rect 116965 43253 117031 43254
rect 116965 43182 117031 43183
rect 116965 43150 116966 43182
rect 110160 43014 110166 43046
rect 28288 42976 28364 42982
rect 110165 42982 110166 43014
rect 110230 43014 110236 43046
rect 116960 43118 116966 43150
rect 117030 43150 117031 43182
rect 117030 43118 117036 43150
rect 110230 42982 110231 43014
rect 110165 42981 110231 42982
rect 21830 42846 21831 42878
rect 21765 42845 21831 42846
rect 22440 42846 22446 42910
rect 22510 42846 22516 42910
rect 22440 42840 22516 42846
rect 28288 42910 28364 42916
rect 28288 42846 28294 42910
rect 28358 42846 28364 42910
rect 21765 42774 21831 42775
rect 21765 42742 21766 42774
rect 952 42438 1230 42502
rect 1294 42438 1300 42502
rect 952 40734 1300 42438
rect 21760 42710 21766 42742
rect 21830 42742 21831 42774
rect 23125 42774 23191 42775
rect 23125 42742 23126 42774
rect 21830 42710 21836 42742
rect 21760 42502 21836 42710
rect 21760 42438 21766 42502
rect 21830 42438 21836 42502
rect 21760 42432 21836 42438
rect 23120 42710 23126 42742
rect 23190 42742 23191 42774
rect 23392 42774 23468 42780
rect 23190 42710 23196 42742
rect 23120 42502 23196 42710
rect 23120 42438 23126 42502
rect 23190 42438 23196 42502
rect 23392 42710 23398 42774
rect 23462 42710 23468 42774
rect 23392 42502 23468 42710
rect 28288 42638 28364 42846
rect 116960 42910 117036 43118
rect 116960 42846 116966 42910
rect 117030 42846 117036 42910
rect 116960 42840 117036 42846
rect 115333 42774 115399 42775
rect 115333 42742 115334 42774
rect 28288 42606 28294 42638
rect 28293 42574 28294 42606
rect 28358 42606 28364 42638
rect 115328 42710 115334 42742
rect 115398 42742 115399 42774
rect 115600 42774 115676 42780
rect 115398 42710 115404 42742
rect 28358 42574 28359 42606
rect 28293 42573 28359 42574
rect 23392 42470 23398 42502
rect 23120 42432 23196 42438
rect 23397 42438 23398 42470
rect 23462 42470 23468 42502
rect 115328 42502 115404 42710
rect 23462 42438 23463 42470
rect 23397 42437 23463 42438
rect 115328 42438 115334 42502
rect 115398 42438 115404 42502
rect 115600 42710 115606 42774
rect 115670 42710 115676 42774
rect 115600 42502 115676 42710
rect 115600 42470 115606 42502
rect 115328 42432 115404 42438
rect 115605 42438 115606 42470
rect 115670 42470 115676 42502
rect 116960 42774 117036 42780
rect 116960 42710 116966 42774
rect 117030 42710 117036 42774
rect 116960 42502 117036 42710
rect 116960 42470 116966 42502
rect 115670 42438 115671 42470
rect 115605 42437 115671 42438
rect 116965 42438 116966 42470
rect 117030 42470 117036 42502
rect 137496 42502 137844 44070
rect 117030 42438 117031 42470
rect 116965 42437 117031 42438
rect 137496 42438 137502 42502
rect 137566 42438 137844 42502
rect 21896 42366 21972 42372
rect 21896 42302 21902 42366
rect 21966 42302 21972 42366
rect 21896 42094 21972 42302
rect 21896 42062 21902 42094
rect 21901 42030 21902 42062
rect 21966 42062 21972 42094
rect 23120 42366 23196 42372
rect 23120 42302 23126 42366
rect 23190 42302 23196 42366
rect 23120 42094 23196 42302
rect 23120 42062 23126 42094
rect 21966 42030 21967 42062
rect 21901 42029 21967 42030
rect 23125 42030 23126 42062
rect 23190 42062 23196 42094
rect 23392 42366 23468 42372
rect 23392 42302 23398 42366
rect 23462 42302 23468 42366
rect 23392 42094 23468 42302
rect 115192 42366 115268 42372
rect 115192 42302 115198 42366
rect 115262 42302 115268 42366
rect 115605 42366 115671 42367
rect 115605 42334 115606 42366
rect 23392 42062 23398 42094
rect 23190 42030 23191 42062
rect 23125 42029 23191 42030
rect 23397 42030 23398 42062
rect 23462 42062 23468 42094
rect 110432 42094 110508 42100
rect 23462 42030 23463 42062
rect 23397 42029 23463 42030
rect 110432 42030 110438 42094
rect 110502 42030 110508 42094
rect 115192 42094 115268 42302
rect 115192 42062 115198 42094
rect 21760 41958 21836 41964
rect 21760 41894 21766 41958
rect 21830 41894 21836 41958
rect 21760 41686 21836 41894
rect 21760 41654 21766 41686
rect 21765 41622 21766 41654
rect 21830 41654 21836 41686
rect 22168 41958 22244 41964
rect 22168 41894 22174 41958
rect 22238 41894 22244 41958
rect 22445 41958 22511 41959
rect 22445 41926 22446 41958
rect 22168 41686 22244 41894
rect 22168 41654 22174 41686
rect 21830 41622 21831 41654
rect 21765 41621 21831 41622
rect 22173 41622 22174 41654
rect 22238 41654 22244 41686
rect 22440 41894 22446 41926
rect 22510 41926 22511 41958
rect 23120 41958 23196 41964
rect 22510 41894 22516 41926
rect 22440 41686 22516 41894
rect 22238 41622 22239 41654
rect 22173 41621 22239 41622
rect 22440 41622 22446 41686
rect 22510 41622 22516 41686
rect 23120 41894 23126 41958
rect 23190 41894 23196 41958
rect 23533 41958 23599 41959
rect 23533 41926 23534 41958
rect 23120 41686 23196 41894
rect 23120 41654 23126 41686
rect 22440 41616 22516 41622
rect 23125 41622 23126 41654
rect 23190 41654 23196 41686
rect 23528 41894 23534 41926
rect 23598 41926 23599 41958
rect 23598 41894 23604 41926
rect 23528 41686 23604 41894
rect 110432 41822 110508 42030
rect 115197 42030 115198 42062
rect 115262 42062 115268 42094
rect 115600 42302 115606 42334
rect 115670 42334 115671 42366
rect 116144 42366 116220 42372
rect 115670 42302 115676 42334
rect 115600 42094 115676 42302
rect 115262 42030 115263 42062
rect 115197 42029 115263 42030
rect 115600 42030 115606 42094
rect 115670 42030 115676 42094
rect 116144 42302 116150 42366
rect 116214 42302 116220 42366
rect 116965 42366 117031 42367
rect 116965 42334 116966 42366
rect 116144 42094 116220 42302
rect 116144 42062 116150 42094
rect 115600 42024 115676 42030
rect 116149 42030 116150 42062
rect 116214 42062 116220 42094
rect 116960 42302 116966 42334
rect 117030 42334 117031 42366
rect 117030 42302 117036 42334
rect 116960 42094 117036 42302
rect 116214 42030 116215 42062
rect 116149 42029 116215 42030
rect 116960 42030 116966 42094
rect 117030 42030 117036 42094
rect 116960 42024 117036 42030
rect 110432 41790 110438 41822
rect 110437 41758 110438 41790
rect 110502 41790 110508 41822
rect 115328 41958 115404 41964
rect 115328 41894 115334 41958
rect 115398 41894 115404 41958
rect 115741 41958 115807 41959
rect 115741 41926 115742 41958
rect 110502 41758 110503 41790
rect 110437 41757 110503 41758
rect 23190 41622 23191 41654
rect 23125 41621 23191 41622
rect 23528 41622 23534 41686
rect 23598 41622 23604 41686
rect 115328 41686 115404 41894
rect 115328 41654 115334 41686
rect 23528 41616 23604 41622
rect 115333 41622 115334 41654
rect 115398 41654 115404 41686
rect 115736 41894 115742 41926
rect 115806 41926 115807 41958
rect 116013 41958 116079 41959
rect 116013 41926 116014 41958
rect 115806 41894 115812 41926
rect 115736 41686 115812 41894
rect 115398 41622 115399 41654
rect 115333 41621 115399 41622
rect 115736 41622 115742 41686
rect 115806 41622 115812 41686
rect 115736 41616 115812 41622
rect 116008 41894 116014 41926
rect 116078 41926 116079 41958
rect 116421 41958 116487 41959
rect 116421 41926 116422 41958
rect 116078 41894 116084 41926
rect 116008 41686 116084 41894
rect 116008 41622 116014 41686
rect 116078 41622 116084 41686
rect 116008 41616 116084 41622
rect 116416 41894 116422 41926
rect 116486 41926 116487 41958
rect 116824 41958 116900 41964
rect 116486 41894 116492 41926
rect 116416 41686 116492 41894
rect 116416 41622 116422 41686
rect 116486 41622 116492 41686
rect 116824 41894 116830 41958
rect 116894 41894 116900 41958
rect 116824 41686 116900 41894
rect 116824 41654 116830 41686
rect 116416 41616 116492 41622
rect 116829 41622 116830 41654
rect 116894 41654 116900 41686
rect 116894 41622 116895 41654
rect 116829 41621 116895 41622
rect 21765 41550 21831 41551
rect 21765 41518 21766 41550
rect 21760 41486 21766 41518
rect 21830 41518 21831 41550
rect 23125 41550 23191 41551
rect 23125 41518 23126 41550
rect 21830 41486 21836 41518
rect 21760 41278 21836 41486
rect 21760 41214 21766 41278
rect 21830 41214 21836 41278
rect 21760 41208 21836 41214
rect 23120 41486 23126 41518
rect 23190 41518 23191 41550
rect 23392 41550 23468 41556
rect 23190 41486 23196 41518
rect 23120 41278 23196 41486
rect 23120 41214 23126 41278
rect 23190 41214 23196 41278
rect 23392 41486 23398 41550
rect 23462 41486 23468 41550
rect 23392 41278 23468 41486
rect 23392 41246 23398 41278
rect 23120 41208 23196 41214
rect 23397 41214 23398 41246
rect 23462 41246 23468 41278
rect 115192 41550 115268 41556
rect 115192 41486 115198 41550
rect 115262 41486 115268 41550
rect 115192 41278 115268 41486
rect 115192 41246 115198 41278
rect 23462 41214 23463 41246
rect 23397 41213 23463 41214
rect 115197 41214 115198 41246
rect 115262 41246 115268 41278
rect 115600 41550 115676 41556
rect 115600 41486 115606 41550
rect 115670 41486 115676 41550
rect 115600 41278 115676 41486
rect 115600 41246 115606 41278
rect 115262 41214 115263 41246
rect 115197 41213 115263 41214
rect 115605 41214 115606 41246
rect 115670 41246 115676 41278
rect 116008 41550 116084 41556
rect 116008 41486 116014 41550
rect 116078 41486 116084 41550
rect 116008 41278 116084 41486
rect 116008 41246 116014 41278
rect 115670 41214 115671 41246
rect 115605 41213 115671 41214
rect 116013 41214 116014 41246
rect 116078 41246 116084 41278
rect 116280 41550 116356 41556
rect 116280 41486 116286 41550
rect 116350 41486 116356 41550
rect 116280 41278 116356 41486
rect 116280 41246 116286 41278
rect 116078 41214 116079 41246
rect 116013 41213 116079 41214
rect 116285 41214 116286 41246
rect 116350 41246 116356 41278
rect 116552 41550 116628 41556
rect 116552 41486 116558 41550
rect 116622 41486 116628 41550
rect 116552 41278 116628 41486
rect 116552 41246 116558 41278
rect 116350 41214 116351 41246
rect 116285 41213 116351 41214
rect 116557 41214 116558 41246
rect 116622 41246 116628 41278
rect 116960 41550 117036 41556
rect 116960 41486 116966 41550
rect 117030 41486 117036 41550
rect 116960 41278 117036 41486
rect 116960 41246 116966 41278
rect 116622 41214 116623 41246
rect 116557 41213 116623 41214
rect 116965 41214 116966 41246
rect 117030 41246 117036 41278
rect 117030 41214 117031 41246
rect 116965 41213 117031 41214
rect 21760 41142 21836 41148
rect 21760 41078 21766 41142
rect 21830 41078 21836 41142
rect 21760 40870 21836 41078
rect 21760 40838 21766 40870
rect 21765 40806 21766 40838
rect 21830 40838 21836 40870
rect 22168 41142 22244 41148
rect 22168 41078 22174 41142
rect 22238 41078 22244 41142
rect 22717 41142 22783 41143
rect 22717 41110 22718 41142
rect 22168 40870 22244 41078
rect 22168 40838 22174 40870
rect 21830 40806 21831 40838
rect 21765 40805 21831 40806
rect 22173 40806 22174 40838
rect 22238 40838 22244 40870
rect 22712 41078 22718 41110
rect 22782 41110 22783 41142
rect 22984 41142 23060 41148
rect 22782 41078 22788 41110
rect 22712 40870 22788 41078
rect 22238 40806 22239 40838
rect 22173 40805 22239 40806
rect 22712 40806 22718 40870
rect 22782 40806 22788 40870
rect 22984 41078 22990 41142
rect 23054 41078 23060 41142
rect 22984 40870 23060 41078
rect 22984 40838 22990 40870
rect 22712 40800 22788 40806
rect 22989 40806 22990 40838
rect 23054 40838 23060 40870
rect 23528 41142 23604 41148
rect 23528 41078 23534 41142
rect 23598 41078 23604 41142
rect 115197 41142 115263 41143
rect 115197 41110 115198 41142
rect 23528 40870 23604 41078
rect 23528 40838 23534 40870
rect 23054 40806 23055 40838
rect 22989 40805 23055 40806
rect 23533 40806 23534 40838
rect 23598 40838 23604 40870
rect 115192 41078 115198 41110
rect 115262 41110 115263 41142
rect 115736 41142 115812 41148
rect 115262 41078 115268 41110
rect 115192 40870 115268 41078
rect 23598 40806 23599 40838
rect 23533 40805 23599 40806
rect 115192 40806 115198 40870
rect 115262 40806 115268 40870
rect 115736 41078 115742 41142
rect 115806 41078 115812 41142
rect 115736 40870 115812 41078
rect 115736 40838 115742 40870
rect 115192 40800 115268 40806
rect 115741 40806 115742 40838
rect 115806 40838 115812 40870
rect 116008 41142 116084 41148
rect 116008 41078 116014 41142
rect 116078 41078 116084 41142
rect 116965 41142 117031 41143
rect 116965 41110 116966 41142
rect 116008 40870 116084 41078
rect 116008 40838 116014 40870
rect 115806 40806 115807 40838
rect 115741 40805 115807 40806
rect 116013 40806 116014 40838
rect 116078 40838 116084 40870
rect 116960 41078 116966 41110
rect 117030 41110 117031 41142
rect 117030 41078 117036 41110
rect 116960 40870 117036 41078
rect 116078 40806 116079 40838
rect 116013 40805 116079 40806
rect 116960 40806 116966 40870
rect 117030 40806 117036 40870
rect 116960 40800 117036 40806
rect 952 40670 1230 40734
rect 1294 40670 1300 40734
rect 952 39102 1300 40670
rect 22576 40734 22652 40740
rect 22576 40670 22582 40734
rect 22646 40670 22652 40734
rect 14688 40598 14764 40604
rect 14688 40534 14694 40598
rect 14758 40534 14764 40598
rect 14557 39238 14623 39239
rect 14557 39206 14558 39238
rect 952 39038 1230 39102
rect 1294 39038 1300 39102
rect 952 37470 1300 39038
rect 952 37406 1230 37470
rect 1294 37406 1300 37470
rect 952 35838 1300 37406
rect 14552 39174 14558 39206
rect 14622 39206 14623 39238
rect 14622 39174 14628 39206
rect 14552 36518 14628 39174
rect 14688 37878 14764 40534
rect 22576 40462 22652 40670
rect 22576 40430 22582 40462
rect 22581 40398 22582 40430
rect 22646 40430 22652 40462
rect 23120 40734 23196 40740
rect 23120 40670 23126 40734
rect 23190 40670 23196 40734
rect 23533 40734 23599 40735
rect 23533 40702 23534 40734
rect 23120 40462 23196 40670
rect 23120 40430 23126 40462
rect 22646 40398 22647 40430
rect 22581 40397 22647 40398
rect 23125 40398 23126 40430
rect 23190 40430 23196 40462
rect 23528 40670 23534 40702
rect 23598 40702 23599 40734
rect 115192 40734 115268 40740
rect 23598 40670 23604 40702
rect 23528 40462 23604 40670
rect 115192 40670 115198 40734
rect 115262 40670 115268 40734
rect 115741 40734 115807 40735
rect 115741 40702 115742 40734
rect 110165 40598 110231 40599
rect 110165 40566 110166 40598
rect 23190 40398 23191 40430
rect 23125 40397 23191 40398
rect 23528 40398 23534 40462
rect 23598 40398 23604 40462
rect 23528 40392 23604 40398
rect 110160 40534 110166 40566
rect 110230 40566 110231 40598
rect 110230 40534 110236 40566
rect 22989 40326 23055 40327
rect 22989 40294 22990 40326
rect 22984 40262 22990 40294
rect 23054 40294 23055 40326
rect 23392 40326 23468 40332
rect 23054 40262 23060 40294
rect 22984 40054 23060 40262
rect 22984 39990 22990 40054
rect 23054 39990 23060 40054
rect 23392 40262 23398 40326
rect 23462 40262 23468 40326
rect 23392 40054 23468 40262
rect 110160 40326 110236 40534
rect 115192 40462 115268 40670
rect 115192 40430 115198 40462
rect 115197 40398 115198 40430
rect 115262 40430 115268 40462
rect 115736 40670 115742 40702
rect 115806 40702 115807 40734
rect 116013 40734 116079 40735
rect 116013 40702 116014 40734
rect 115806 40670 115812 40702
rect 115736 40462 115812 40670
rect 115262 40398 115263 40430
rect 115197 40397 115263 40398
rect 115736 40398 115742 40462
rect 115806 40398 115812 40462
rect 115736 40392 115812 40398
rect 116008 40670 116014 40702
rect 116078 40702 116079 40734
rect 137496 40734 137844 42438
rect 116078 40670 116084 40702
rect 116008 40462 116084 40670
rect 116008 40398 116014 40462
rect 116078 40398 116084 40462
rect 116008 40392 116084 40398
rect 137496 40670 137502 40734
rect 137566 40670 137844 40734
rect 110160 40262 110166 40326
rect 110230 40262 110236 40326
rect 115197 40326 115263 40327
rect 115197 40294 115198 40326
rect 110160 40256 110236 40262
rect 115192 40262 115198 40294
rect 115262 40294 115263 40326
rect 115600 40326 115676 40332
rect 115262 40262 115268 40294
rect 23392 40022 23398 40054
rect 22984 39984 23060 39990
rect 23397 39990 23398 40022
rect 23462 40022 23468 40054
rect 115192 40054 115268 40262
rect 23462 39990 23463 40022
rect 23397 39989 23463 39990
rect 115192 39990 115198 40054
rect 115262 39990 115268 40054
rect 115600 40262 115606 40326
rect 115670 40262 115676 40326
rect 115600 40054 115676 40262
rect 115600 40022 115606 40054
rect 115192 39984 115268 39990
rect 115605 39990 115606 40022
rect 115670 40022 115676 40054
rect 115670 39990 115671 40022
rect 115605 39989 115671 39990
rect 22576 39918 22652 39924
rect 22576 39854 22582 39918
rect 22646 39854 22652 39918
rect 21765 39646 21831 39647
rect 21765 39614 21766 39646
rect 21760 39582 21766 39614
rect 21830 39614 21831 39646
rect 22576 39646 22652 39854
rect 22576 39614 22582 39646
rect 21830 39582 21836 39614
rect 21760 39374 21836 39582
rect 22581 39582 22582 39614
rect 22646 39614 22652 39646
rect 23120 39918 23196 39924
rect 23120 39854 23126 39918
rect 23190 39854 23196 39918
rect 23120 39646 23196 39854
rect 23120 39614 23126 39646
rect 22646 39582 22647 39614
rect 22581 39581 22647 39582
rect 23125 39582 23126 39614
rect 23190 39614 23196 39646
rect 23528 39918 23604 39924
rect 23528 39854 23534 39918
rect 23598 39854 23604 39918
rect 115197 39918 115263 39919
rect 115197 39886 115198 39918
rect 23528 39646 23604 39854
rect 115192 39854 115198 39886
rect 115262 39886 115263 39918
rect 115605 39918 115671 39919
rect 115605 39886 115606 39918
rect 115262 39854 115268 39886
rect 23528 39614 23534 39646
rect 23190 39582 23191 39614
rect 23125 39581 23191 39582
rect 23533 39582 23534 39614
rect 23598 39614 23604 39646
rect 28424 39782 28500 39788
rect 28424 39718 28430 39782
rect 28494 39718 28500 39782
rect 23598 39582 23599 39614
rect 23533 39581 23599 39582
rect 28424 39510 28500 39718
rect 115192 39646 115268 39854
rect 115192 39582 115198 39646
rect 115262 39582 115268 39646
rect 115192 39576 115268 39582
rect 115600 39854 115606 39886
rect 115670 39886 115671 39918
rect 116416 39918 116492 39924
rect 115670 39854 115676 39886
rect 115600 39646 115676 39854
rect 115600 39582 115606 39646
rect 115670 39582 115676 39646
rect 116416 39854 116422 39918
rect 116486 39854 116492 39918
rect 116416 39646 116492 39854
rect 116416 39614 116422 39646
rect 115600 39576 115676 39582
rect 116421 39582 116422 39614
rect 116486 39614 116492 39646
rect 116824 39646 116900 39652
rect 116486 39582 116487 39614
rect 116421 39581 116487 39582
rect 116824 39582 116830 39646
rect 116894 39582 116900 39646
rect 28424 39478 28430 39510
rect 28429 39446 28430 39478
rect 28494 39478 28500 39510
rect 28494 39446 28495 39478
rect 28429 39445 28495 39446
rect 21760 39310 21766 39374
rect 21830 39310 21836 39374
rect 21760 39304 21836 39310
rect 28288 39374 28364 39380
rect 28288 39310 28294 39374
rect 28358 39310 28364 39374
rect 110437 39374 110503 39375
rect 110437 39342 110438 39374
rect 21901 39238 21967 39239
rect 21901 39206 21902 39238
rect 21896 39174 21902 39206
rect 21966 39206 21967 39238
rect 22309 39238 22375 39239
rect 22309 39206 22310 39238
rect 21966 39174 21972 39206
rect 21896 38966 21972 39174
rect 21896 38902 21902 38966
rect 21966 38902 21972 38966
rect 21896 38896 21972 38902
rect 22304 39174 22310 39206
rect 22374 39206 22375 39238
rect 22445 39238 22511 39239
rect 22445 39206 22446 39238
rect 22374 39174 22380 39206
rect 22304 38966 22380 39174
rect 22304 38902 22310 38966
rect 22374 38902 22380 38966
rect 22304 38896 22380 38902
rect 22440 39174 22446 39206
rect 22510 39206 22511 39238
rect 22510 39174 22516 39206
rect 22440 38966 22516 39174
rect 28288 39102 28364 39310
rect 28288 39070 28294 39102
rect 28293 39038 28294 39070
rect 28358 39070 28364 39102
rect 110432 39310 110438 39342
rect 110502 39342 110503 39374
rect 116824 39374 116900 39582
rect 116824 39342 116830 39374
rect 110502 39310 110508 39342
rect 110432 39102 110508 39310
rect 116829 39310 116830 39342
rect 116894 39342 116900 39374
rect 116894 39310 116895 39342
rect 116829 39309 116895 39310
rect 116557 39238 116623 39239
rect 116557 39206 116558 39238
rect 28358 39038 28359 39070
rect 28293 39037 28359 39038
rect 110432 39038 110438 39102
rect 110502 39038 110508 39102
rect 110432 39032 110508 39038
rect 116552 39174 116558 39206
rect 116622 39206 116623 39238
rect 116960 39238 117036 39244
rect 116622 39174 116628 39206
rect 22440 38902 22446 38966
rect 22510 38902 22516 38966
rect 28293 38966 28359 38967
rect 28293 38934 28294 38966
rect 22440 38896 22516 38902
rect 28288 38902 28294 38934
rect 28358 38934 28359 38966
rect 116552 38966 116628 39174
rect 28358 38902 28364 38934
rect 21901 38830 21967 38831
rect 21901 38798 21902 38830
rect 21896 38766 21902 38798
rect 21966 38798 21967 38830
rect 21966 38766 21972 38798
rect 21896 38558 21972 38766
rect 28288 38694 28364 38902
rect 116552 38902 116558 38966
rect 116622 38902 116628 38966
rect 116960 39174 116966 39238
rect 117030 39174 117036 39238
rect 116960 38966 117036 39174
rect 116960 38934 116966 38966
rect 116552 38896 116628 38902
rect 116965 38902 116966 38934
rect 117030 38934 117036 38966
rect 137496 38966 137844 40670
rect 117030 38902 117031 38934
rect 116965 38901 117031 38902
rect 137496 38902 137502 38966
rect 137566 38902 137844 38966
rect 116965 38830 117031 38831
rect 116965 38798 116966 38830
rect 116960 38766 116966 38798
rect 117030 38798 117031 38830
rect 117030 38766 117036 38798
rect 28288 38630 28294 38694
rect 28358 38630 28364 38694
rect 110165 38694 110231 38695
rect 110165 38662 110166 38694
rect 28288 38624 28364 38630
rect 110160 38630 110166 38662
rect 110230 38662 110231 38694
rect 110230 38630 110236 38662
rect 21896 38494 21902 38558
rect 21966 38494 21972 38558
rect 21896 38488 21972 38494
rect 21896 38422 21972 38428
rect 21896 38358 21902 38422
rect 21966 38358 21972 38422
rect 22173 38422 22239 38423
rect 22173 38390 22174 38422
rect 21896 38150 21972 38358
rect 21896 38118 21902 38150
rect 21901 38086 21902 38118
rect 21966 38118 21972 38150
rect 22168 38358 22174 38390
rect 22238 38390 22239 38422
rect 22712 38422 22788 38428
rect 22238 38358 22244 38390
rect 22168 38150 22244 38358
rect 21966 38086 21967 38118
rect 21901 38085 21967 38086
rect 22168 38086 22174 38150
rect 22238 38086 22244 38150
rect 22712 38358 22718 38422
rect 22782 38358 22788 38422
rect 22712 38150 22788 38358
rect 22712 38118 22718 38150
rect 22168 38080 22244 38086
rect 22717 38086 22718 38118
rect 22782 38118 22788 38150
rect 22984 38422 23060 38428
rect 22984 38358 22990 38422
rect 23054 38358 23060 38422
rect 22984 38150 23060 38358
rect 22984 38118 22990 38150
rect 22782 38086 22783 38118
rect 22717 38085 22783 38086
rect 22989 38086 22990 38118
rect 23054 38118 23060 38150
rect 23392 38422 23468 38428
rect 23392 38358 23398 38422
rect 23462 38358 23468 38422
rect 23392 38150 23468 38358
rect 110160 38422 110236 38630
rect 116960 38558 117036 38766
rect 116960 38494 116966 38558
rect 117030 38494 117036 38558
rect 116960 38488 117036 38494
rect 110160 38358 110166 38422
rect 110230 38358 110236 38422
rect 115333 38422 115399 38423
rect 115333 38390 115334 38422
rect 110160 38352 110236 38358
rect 115328 38358 115334 38390
rect 115398 38390 115399 38422
rect 115741 38422 115807 38423
rect 115741 38390 115742 38422
rect 115398 38358 115404 38390
rect 23392 38118 23398 38150
rect 23054 38086 23055 38118
rect 22989 38085 23055 38086
rect 23397 38086 23398 38118
rect 23462 38118 23468 38150
rect 115328 38150 115404 38358
rect 23462 38086 23463 38118
rect 23397 38085 23463 38086
rect 115328 38086 115334 38150
rect 115398 38086 115404 38150
rect 115328 38080 115404 38086
rect 115736 38358 115742 38390
rect 115806 38390 115807 38422
rect 116013 38422 116079 38423
rect 116013 38390 116014 38422
rect 115806 38358 115812 38390
rect 115736 38150 115812 38358
rect 115736 38086 115742 38150
rect 115806 38086 115812 38150
rect 115736 38080 115812 38086
rect 116008 38358 116014 38390
rect 116078 38390 116079 38422
rect 116829 38422 116895 38423
rect 116829 38390 116830 38422
rect 116078 38358 116084 38390
rect 116008 38150 116084 38358
rect 116008 38086 116014 38150
rect 116078 38086 116084 38150
rect 116008 38080 116084 38086
rect 116824 38358 116830 38390
rect 116894 38390 116895 38422
rect 116894 38358 116900 38390
rect 116824 38150 116900 38358
rect 116824 38086 116830 38150
rect 116894 38086 116900 38150
rect 116824 38080 116900 38086
rect 21901 38014 21967 38015
rect 21901 37982 21902 38014
rect 14688 37846 14694 37878
rect 14693 37814 14694 37846
rect 14758 37846 14764 37878
rect 21896 37950 21902 37982
rect 21966 37982 21967 38014
rect 22989 38014 23055 38015
rect 22989 37982 22990 38014
rect 21966 37950 21972 37982
rect 14758 37814 14759 37846
rect 14693 37813 14759 37814
rect 14829 37742 14895 37743
rect 14829 37710 14830 37742
rect 14552 36454 14558 36518
rect 14622 36454 14628 36518
rect 14552 36448 14628 36454
rect 14824 37678 14830 37710
rect 14894 37710 14895 37742
rect 21896 37742 21972 37950
rect 14894 37678 14900 37710
rect 952 35774 1230 35838
rect 1294 35774 1300 35838
rect 952 34070 1300 35774
rect 14688 36382 14764 36388
rect 14688 36318 14694 36382
rect 14758 36318 14764 36382
rect 14557 34886 14623 34887
rect 14557 34854 14558 34886
rect 952 34006 1230 34070
rect 1294 34006 1300 34070
rect 952 32438 1300 34006
rect 952 32374 1230 32438
rect 1294 32374 1300 32438
rect 952 30670 1300 32374
rect 14552 34822 14558 34854
rect 14622 34854 14623 34886
rect 14622 34822 14628 34854
rect 14552 32302 14628 34822
rect 14688 33662 14764 36318
rect 14824 35158 14900 37678
rect 21896 37678 21902 37742
rect 21966 37678 21972 37742
rect 21896 37672 21972 37678
rect 22984 37950 22990 37982
rect 23054 37982 23055 38014
rect 23397 38014 23463 38015
rect 23397 37982 23398 38014
rect 23054 37950 23060 37982
rect 22984 37742 23060 37950
rect 22984 37678 22990 37742
rect 23054 37678 23060 37742
rect 22984 37672 23060 37678
rect 23392 37950 23398 37982
rect 23462 37982 23463 38014
rect 115192 38014 115268 38020
rect 23462 37950 23468 37982
rect 23392 37742 23468 37950
rect 23392 37678 23398 37742
rect 23462 37678 23468 37742
rect 115192 37950 115198 38014
rect 115262 37950 115268 38014
rect 115192 37742 115268 37950
rect 115192 37710 115198 37742
rect 23392 37672 23468 37678
rect 115197 37678 115198 37710
rect 115262 37710 115268 37742
rect 115600 38014 115676 38020
rect 115600 37950 115606 38014
rect 115670 37950 115676 38014
rect 116013 38014 116079 38015
rect 116013 37982 116014 38014
rect 115600 37742 115676 37950
rect 115600 37710 115606 37742
rect 115262 37678 115263 37710
rect 115197 37677 115263 37678
rect 115605 37678 115606 37710
rect 115670 37710 115676 37742
rect 116008 37950 116014 37982
rect 116078 37982 116079 38014
rect 116965 38014 117031 38015
rect 116965 37982 116966 38014
rect 116078 37950 116084 37982
rect 116008 37742 116084 37950
rect 115670 37678 115671 37710
rect 115605 37677 115671 37678
rect 116008 37678 116014 37742
rect 116078 37678 116084 37742
rect 116008 37672 116084 37678
rect 116960 37950 116966 37982
rect 117030 37982 117031 38014
rect 117030 37950 117036 37982
rect 116960 37742 117036 37950
rect 116960 37678 116966 37742
rect 117030 37678 117036 37742
rect 116960 37672 117036 37678
rect 21760 37606 21836 37612
rect 21760 37542 21766 37606
rect 21830 37542 21836 37606
rect 21760 37334 21836 37542
rect 21760 37302 21766 37334
rect 21765 37270 21766 37302
rect 21830 37302 21836 37334
rect 22168 37606 22244 37612
rect 22168 37542 22174 37606
rect 22238 37542 22244 37606
rect 22445 37606 22511 37607
rect 22445 37574 22446 37606
rect 22168 37334 22244 37542
rect 22168 37302 22174 37334
rect 21830 37270 21831 37302
rect 21765 37269 21831 37270
rect 22173 37270 22174 37302
rect 22238 37302 22244 37334
rect 22440 37542 22446 37574
rect 22510 37574 22511 37606
rect 23120 37606 23196 37612
rect 22510 37542 22516 37574
rect 22440 37334 22516 37542
rect 22238 37270 22239 37302
rect 22173 37269 22239 37270
rect 22440 37270 22446 37334
rect 22510 37270 22516 37334
rect 23120 37542 23126 37606
rect 23190 37542 23196 37606
rect 23533 37606 23599 37607
rect 23533 37574 23534 37606
rect 23120 37334 23196 37542
rect 23120 37302 23126 37334
rect 22440 37264 22516 37270
rect 23125 37270 23126 37302
rect 23190 37302 23196 37334
rect 23528 37542 23534 37574
rect 23598 37574 23599 37606
rect 115328 37606 115404 37612
rect 23598 37542 23604 37574
rect 23528 37334 23604 37542
rect 23190 37270 23191 37302
rect 23125 37269 23191 37270
rect 23528 37270 23534 37334
rect 23598 37270 23604 37334
rect 115328 37542 115334 37606
rect 115398 37542 115404 37606
rect 115328 37334 115404 37542
rect 115328 37302 115334 37334
rect 23528 37264 23604 37270
rect 115333 37270 115334 37302
rect 115398 37302 115404 37334
rect 115736 37606 115812 37612
rect 115736 37542 115742 37606
rect 115806 37542 115812 37606
rect 115736 37334 115812 37542
rect 115736 37302 115742 37334
rect 115398 37270 115399 37302
rect 115333 37269 115399 37270
rect 115741 37270 115742 37302
rect 115806 37302 115812 37334
rect 116144 37606 116220 37612
rect 116144 37542 116150 37606
rect 116214 37542 116220 37606
rect 116144 37334 116220 37542
rect 116144 37302 116150 37334
rect 115806 37270 115807 37302
rect 115741 37269 115807 37270
rect 116149 37270 116150 37302
rect 116214 37302 116220 37334
rect 116280 37606 116356 37612
rect 116280 37542 116286 37606
rect 116350 37542 116356 37606
rect 116280 37334 116356 37542
rect 116280 37302 116286 37334
rect 116214 37270 116215 37302
rect 116149 37269 116215 37270
rect 116285 37270 116286 37302
rect 116350 37302 116356 37334
rect 116824 37606 116900 37612
rect 116824 37542 116830 37606
rect 116894 37542 116900 37606
rect 116824 37334 116900 37542
rect 116824 37302 116830 37334
rect 116350 37270 116351 37302
rect 116285 37269 116351 37270
rect 116829 37270 116830 37302
rect 116894 37302 116900 37334
rect 137496 37334 137844 38902
rect 116894 37270 116895 37302
rect 116829 37269 116895 37270
rect 137496 37270 137502 37334
rect 137566 37270 137844 37334
rect 21896 37198 21972 37204
rect 21896 37134 21902 37198
rect 21966 37134 21972 37198
rect 21896 36926 21972 37134
rect 21896 36894 21902 36926
rect 21901 36862 21902 36894
rect 21966 36894 21972 36926
rect 22984 37198 23060 37204
rect 22984 37134 22990 37198
rect 23054 37134 23060 37198
rect 22984 36926 23060 37134
rect 22984 36894 22990 36926
rect 21966 36862 21967 36894
rect 21901 36861 21967 36862
rect 22989 36862 22990 36894
rect 23054 36894 23060 36926
rect 23392 37198 23468 37204
rect 23392 37134 23398 37198
rect 23462 37134 23468 37198
rect 115333 37198 115399 37199
rect 115333 37166 115334 37198
rect 23392 36926 23468 37134
rect 23392 36894 23398 36926
rect 23054 36862 23055 36894
rect 22989 36861 23055 36862
rect 23397 36862 23398 36894
rect 23462 36894 23468 36926
rect 115328 37134 115334 37166
rect 115398 37166 115399 37198
rect 115600 37198 115676 37204
rect 115398 37134 115404 37166
rect 115328 36926 115404 37134
rect 23462 36862 23463 36894
rect 23397 36861 23463 36862
rect 115328 36862 115334 36926
rect 115398 36862 115404 36926
rect 115600 37134 115606 37198
rect 115670 37134 115676 37198
rect 116149 37198 116215 37199
rect 116149 37166 116150 37198
rect 115600 36926 115676 37134
rect 115600 36894 115606 36926
rect 115328 36856 115404 36862
rect 115605 36862 115606 36894
rect 115670 36894 115676 36926
rect 116144 37134 116150 37166
rect 116214 37166 116215 37198
rect 116285 37198 116351 37199
rect 116285 37166 116286 37198
rect 116214 37134 116220 37166
rect 116144 36926 116220 37134
rect 115670 36862 115671 36894
rect 115605 36861 115671 36862
rect 116144 36862 116150 36926
rect 116214 36862 116220 36926
rect 116144 36856 116220 36862
rect 116280 37134 116286 37166
rect 116350 37166 116351 37198
rect 116552 37198 116628 37204
rect 116350 37134 116356 37166
rect 116280 36926 116356 37134
rect 116280 36862 116286 36926
rect 116350 36862 116356 36926
rect 116552 37134 116558 37198
rect 116622 37134 116628 37198
rect 116829 37198 116895 37199
rect 116829 37166 116830 37198
rect 116552 36926 116628 37134
rect 116552 36894 116558 36926
rect 116280 36856 116356 36862
rect 116557 36862 116558 36894
rect 116622 36894 116628 36926
rect 116824 37134 116830 37166
rect 116894 37166 116895 37198
rect 116894 37134 116900 37166
rect 116824 36926 116900 37134
rect 116622 36862 116623 36894
rect 116557 36861 116623 36862
rect 116824 36862 116830 36926
rect 116894 36862 116900 36926
rect 116824 36856 116900 36862
rect 22168 36790 22244 36796
rect 22168 36726 22174 36790
rect 22238 36726 22244 36790
rect 22717 36790 22783 36791
rect 22717 36758 22718 36790
rect 22168 36518 22244 36726
rect 22168 36486 22174 36518
rect 22173 36454 22174 36486
rect 22238 36486 22244 36518
rect 22712 36726 22718 36758
rect 22782 36758 22783 36790
rect 22989 36790 23055 36791
rect 22989 36758 22990 36790
rect 22782 36726 22788 36758
rect 22712 36518 22788 36726
rect 22238 36454 22239 36486
rect 22173 36453 22239 36454
rect 22712 36454 22718 36518
rect 22782 36454 22788 36518
rect 22712 36448 22788 36454
rect 22984 36726 22990 36758
rect 23054 36758 23055 36790
rect 23397 36790 23463 36791
rect 23397 36758 23398 36790
rect 23054 36726 23060 36758
rect 22984 36518 23060 36726
rect 22984 36454 22990 36518
rect 23054 36454 23060 36518
rect 22984 36448 23060 36454
rect 23392 36726 23398 36758
rect 23462 36758 23463 36790
rect 115197 36790 115263 36791
rect 115197 36758 115198 36790
rect 23462 36726 23468 36758
rect 23392 36518 23468 36726
rect 23392 36454 23398 36518
rect 23462 36454 23468 36518
rect 23392 36448 23468 36454
rect 115192 36726 115198 36758
rect 115262 36758 115263 36790
rect 115605 36790 115671 36791
rect 115605 36758 115606 36790
rect 115262 36726 115268 36758
rect 115192 36518 115268 36726
rect 115192 36454 115198 36518
rect 115262 36454 115268 36518
rect 115192 36448 115268 36454
rect 115600 36726 115606 36758
rect 115670 36758 115671 36790
rect 116013 36790 116079 36791
rect 116013 36758 116014 36790
rect 115670 36726 115676 36758
rect 115600 36518 115676 36726
rect 115600 36454 115606 36518
rect 115670 36454 115676 36518
rect 115600 36448 115676 36454
rect 116008 36726 116014 36758
rect 116078 36758 116079 36790
rect 116285 36790 116351 36791
rect 116285 36758 116286 36790
rect 116078 36726 116084 36758
rect 116008 36518 116084 36726
rect 116008 36454 116014 36518
rect 116078 36454 116084 36518
rect 116008 36448 116084 36454
rect 116280 36726 116286 36758
rect 116350 36758 116351 36790
rect 116350 36726 116356 36758
rect 116280 36518 116356 36726
rect 116280 36454 116286 36518
rect 116350 36454 116356 36518
rect 116280 36448 116356 36454
rect 21901 36382 21967 36383
rect 21901 36350 21902 36382
rect 21896 36318 21902 36350
rect 21966 36350 21967 36382
rect 22173 36382 22239 36383
rect 22173 36350 22174 36382
rect 21966 36318 21972 36350
rect 21896 36110 21972 36318
rect 21896 36046 21902 36110
rect 21966 36046 21972 36110
rect 21896 36040 21972 36046
rect 22168 36318 22174 36350
rect 22238 36350 22239 36382
rect 22581 36382 22647 36383
rect 22581 36350 22582 36382
rect 22238 36318 22244 36350
rect 22168 36110 22244 36318
rect 22168 36046 22174 36110
rect 22238 36046 22244 36110
rect 22168 36040 22244 36046
rect 22576 36318 22582 36350
rect 22646 36350 22647 36382
rect 22989 36382 23055 36383
rect 22989 36350 22990 36382
rect 22646 36318 22652 36350
rect 22576 36110 22652 36318
rect 22576 36046 22582 36110
rect 22646 36046 22652 36110
rect 22576 36040 22652 36046
rect 22984 36318 22990 36350
rect 23054 36350 23055 36382
rect 23528 36382 23604 36388
rect 23054 36318 23060 36350
rect 22984 36110 23060 36318
rect 22984 36046 22990 36110
rect 23054 36046 23060 36110
rect 23528 36318 23534 36382
rect 23598 36318 23604 36382
rect 23528 36110 23604 36318
rect 23528 36078 23534 36110
rect 22984 36040 23060 36046
rect 23533 36046 23534 36078
rect 23598 36078 23604 36110
rect 115328 36382 115404 36388
rect 115328 36318 115334 36382
rect 115398 36318 115404 36382
rect 115741 36382 115807 36383
rect 115741 36350 115742 36382
rect 115328 36110 115404 36318
rect 115328 36078 115334 36110
rect 23598 36046 23599 36078
rect 23533 36045 23599 36046
rect 115333 36046 115334 36078
rect 115398 36078 115404 36110
rect 115736 36318 115742 36350
rect 115806 36350 115807 36382
rect 116280 36382 116356 36388
rect 115806 36318 115812 36350
rect 115736 36110 115812 36318
rect 115398 36046 115399 36078
rect 115333 36045 115399 36046
rect 115736 36046 115742 36110
rect 115806 36046 115812 36110
rect 116280 36318 116286 36382
rect 116350 36318 116356 36382
rect 116280 36110 116356 36318
rect 116280 36078 116286 36110
rect 115736 36040 115812 36046
rect 116285 36046 116286 36078
rect 116350 36078 116356 36110
rect 116960 36382 117036 36388
rect 116960 36318 116966 36382
rect 117030 36318 117036 36382
rect 116960 36110 117036 36318
rect 116960 36078 116966 36110
rect 116350 36046 116351 36078
rect 116285 36045 116351 36046
rect 116965 36046 116966 36078
rect 117030 36078 117036 36110
rect 117030 36046 117031 36078
rect 116965 36045 117031 36046
rect 22712 35974 22788 35980
rect 22712 35910 22718 35974
rect 22782 35910 22788 35974
rect 21901 35702 21967 35703
rect 21901 35670 21902 35702
rect 21896 35638 21902 35670
rect 21966 35670 21967 35702
rect 22712 35702 22788 35910
rect 22712 35670 22718 35702
rect 21966 35638 21972 35670
rect 21896 35430 21972 35638
rect 22717 35638 22718 35670
rect 22782 35670 22788 35702
rect 23120 35974 23196 35980
rect 23120 35910 23126 35974
rect 23190 35910 23196 35974
rect 23120 35702 23196 35910
rect 23120 35670 23126 35702
rect 22782 35638 22783 35670
rect 22717 35637 22783 35638
rect 23125 35638 23126 35670
rect 23190 35670 23196 35702
rect 23392 35974 23468 35980
rect 23392 35910 23398 35974
rect 23462 35910 23468 35974
rect 115333 35974 115399 35975
rect 115333 35942 115334 35974
rect 23392 35702 23468 35910
rect 115328 35910 115334 35942
rect 115398 35942 115399 35974
rect 115600 35974 115676 35980
rect 115398 35910 115404 35942
rect 23392 35670 23398 35702
rect 23190 35638 23191 35670
rect 23125 35637 23191 35638
rect 23397 35638 23398 35670
rect 23462 35670 23468 35702
rect 28560 35838 28636 35844
rect 28560 35774 28566 35838
rect 28630 35774 28636 35838
rect 23462 35638 23463 35670
rect 23397 35637 23463 35638
rect 28560 35566 28636 35774
rect 28560 35534 28566 35566
rect 28565 35502 28566 35534
rect 28630 35534 28636 35566
rect 110296 35838 110372 35844
rect 110296 35774 110302 35838
rect 110366 35774 110372 35838
rect 110296 35566 110372 35774
rect 115328 35702 115404 35910
rect 115328 35638 115334 35702
rect 115398 35638 115404 35702
rect 115600 35910 115606 35974
rect 115670 35910 115676 35974
rect 116557 35974 116623 35975
rect 116557 35942 116558 35974
rect 115600 35702 115676 35910
rect 116552 35910 116558 35942
rect 116622 35942 116623 35974
rect 116622 35910 116628 35942
rect 115600 35670 115606 35702
rect 115328 35632 115404 35638
rect 115605 35638 115606 35670
rect 115670 35670 115676 35702
rect 116285 35702 116351 35703
rect 116285 35670 116286 35702
rect 115670 35638 115671 35670
rect 115605 35637 115671 35638
rect 116280 35638 116286 35670
rect 116350 35670 116351 35702
rect 116552 35702 116628 35910
rect 116350 35638 116356 35670
rect 110296 35534 110302 35566
rect 28630 35502 28631 35534
rect 28565 35501 28631 35502
rect 110301 35502 110302 35534
rect 110366 35534 110372 35566
rect 110366 35502 110367 35534
rect 110301 35501 110367 35502
rect 21896 35366 21902 35430
rect 21966 35366 21972 35430
rect 21896 35360 21972 35366
rect 116280 35430 116356 35638
rect 116552 35638 116558 35702
rect 116622 35638 116628 35702
rect 116965 35702 117031 35703
rect 116965 35670 116966 35702
rect 116552 35632 116628 35638
rect 116960 35638 116966 35670
rect 117030 35670 117031 35702
rect 137496 35702 137844 37270
rect 117030 35638 117036 35670
rect 116280 35366 116286 35430
rect 116350 35366 116356 35430
rect 116280 35360 116356 35366
rect 116960 35430 117036 35638
rect 116960 35366 116966 35430
rect 117030 35366 117036 35430
rect 116960 35360 117036 35366
rect 137496 35638 137502 35702
rect 137566 35638 137844 35702
rect 14824 35094 14830 35158
rect 14894 35094 14900 35158
rect 14824 35088 14900 35094
rect 21760 35294 21836 35300
rect 21760 35230 21766 35294
rect 21830 35230 21836 35294
rect 22581 35294 22647 35295
rect 22581 35262 22582 35294
rect 21760 35022 21836 35230
rect 21760 34990 21766 35022
rect 21765 34958 21766 34990
rect 21830 34990 21836 35022
rect 22576 35230 22582 35262
rect 22646 35262 22647 35294
rect 116552 35294 116628 35300
rect 22646 35230 22652 35262
rect 21830 34958 21831 34990
rect 21765 34957 21831 34958
rect 21896 34886 21972 34892
rect 21896 34822 21902 34886
rect 21966 34822 21972 34886
rect 21896 34614 21972 34822
rect 22576 34886 22652 35230
rect 116552 35230 116558 35294
rect 116622 35230 116628 35294
rect 110437 35022 110503 35023
rect 110437 34990 110438 35022
rect 22576 34822 22582 34886
rect 22646 34822 22652 34886
rect 22576 34816 22652 34822
rect 110432 34958 110438 34990
rect 110502 34990 110503 35022
rect 110502 34958 110508 34990
rect 110165 34750 110231 34751
rect 110165 34718 110166 34750
rect 21896 34582 21902 34614
rect 21901 34550 21902 34582
rect 21966 34582 21972 34614
rect 110160 34686 110166 34718
rect 110230 34718 110231 34750
rect 110432 34750 110508 34958
rect 116552 34886 116628 35230
rect 116824 35294 116900 35300
rect 116824 35230 116830 35294
rect 116894 35230 116900 35294
rect 116824 35022 116900 35230
rect 116824 34990 116830 35022
rect 116829 34958 116830 34990
rect 116894 34990 116900 35022
rect 116894 34958 116895 34990
rect 116829 34957 116895 34958
rect 116552 34854 116558 34886
rect 116557 34822 116558 34854
rect 116622 34854 116628 34886
rect 116960 34886 117036 34892
rect 116622 34822 116623 34854
rect 116557 34821 116623 34822
rect 116960 34822 116966 34886
rect 117030 34822 117036 34886
rect 110230 34686 110236 34718
rect 21966 34550 21967 34582
rect 21901 34549 21967 34550
rect 21901 34478 21967 34479
rect 21901 34446 21902 34478
rect 21896 34414 21902 34446
rect 21966 34446 21967 34478
rect 22445 34478 22511 34479
rect 22445 34446 22446 34478
rect 21966 34414 21972 34446
rect 21896 34206 21972 34414
rect 21896 34142 21902 34206
rect 21966 34142 21972 34206
rect 21896 34136 21972 34142
rect 22440 34414 22446 34446
rect 22510 34446 22511 34478
rect 23125 34478 23191 34479
rect 23125 34446 23126 34478
rect 22510 34414 22516 34446
rect 22440 34206 22516 34414
rect 22440 34142 22446 34206
rect 22510 34142 22516 34206
rect 22440 34136 22516 34142
rect 23120 34414 23126 34446
rect 23190 34446 23191 34478
rect 23397 34478 23463 34479
rect 23397 34446 23398 34478
rect 23190 34414 23196 34446
rect 23120 34206 23196 34414
rect 23120 34142 23126 34206
rect 23190 34142 23196 34206
rect 23120 34136 23196 34142
rect 23392 34414 23398 34446
rect 23462 34446 23463 34478
rect 110160 34478 110236 34686
rect 110432 34686 110438 34750
rect 110502 34686 110508 34750
rect 110432 34680 110508 34686
rect 116960 34614 117036 34822
rect 116960 34582 116966 34614
rect 116965 34550 116966 34582
rect 117030 34582 117036 34614
rect 117030 34550 117031 34582
rect 116965 34549 117031 34550
rect 23462 34414 23468 34446
rect 23392 34206 23468 34414
rect 110160 34414 110166 34478
rect 110230 34414 110236 34478
rect 110160 34408 110236 34414
rect 115328 34478 115404 34484
rect 115328 34414 115334 34478
rect 115398 34414 115404 34478
rect 115605 34478 115671 34479
rect 115605 34446 115606 34478
rect 23392 34142 23398 34206
rect 23462 34142 23468 34206
rect 23392 34136 23468 34142
rect 28288 34206 28364 34212
rect 28288 34142 28294 34206
rect 28358 34142 28364 34206
rect 115328 34206 115404 34414
rect 115328 34174 115334 34206
rect 21765 34070 21831 34071
rect 21765 34038 21766 34070
rect 21760 34006 21766 34038
rect 21830 34038 21831 34070
rect 22173 34070 22239 34071
rect 22173 34038 22174 34070
rect 21830 34006 21836 34038
rect 21760 33798 21836 34006
rect 21760 33734 21766 33798
rect 21830 33734 21836 33798
rect 21760 33728 21836 33734
rect 22168 34006 22174 34038
rect 22238 34038 22239 34070
rect 22712 34070 22788 34076
rect 22238 34006 22244 34038
rect 22168 33798 22244 34006
rect 22168 33734 22174 33798
rect 22238 33734 22244 33798
rect 22712 34006 22718 34070
rect 22782 34006 22788 34070
rect 22712 33798 22788 34006
rect 22712 33766 22718 33798
rect 22168 33728 22244 33734
rect 22717 33734 22718 33766
rect 22782 33766 22788 33798
rect 22984 34070 23060 34076
rect 22984 34006 22990 34070
rect 23054 34006 23060 34070
rect 23533 34070 23599 34071
rect 23533 34038 23534 34070
rect 22984 33798 23060 34006
rect 22984 33766 22990 33798
rect 22782 33734 22783 33766
rect 22717 33733 22783 33734
rect 22989 33734 22990 33766
rect 23054 33766 23060 33798
rect 23528 34006 23534 34038
rect 23598 34038 23599 34070
rect 23598 34006 23604 34038
rect 23528 33798 23604 34006
rect 28288 33934 28364 34142
rect 115333 34142 115334 34174
rect 115398 34174 115404 34206
rect 115600 34414 115606 34446
rect 115670 34446 115671 34478
rect 116008 34478 116084 34484
rect 115670 34414 115676 34446
rect 115600 34206 115676 34414
rect 115398 34142 115399 34174
rect 115333 34141 115399 34142
rect 115600 34142 115606 34206
rect 115670 34142 115676 34206
rect 116008 34414 116014 34478
rect 116078 34414 116084 34478
rect 116965 34478 117031 34479
rect 116965 34446 116966 34478
rect 116008 34206 116084 34414
rect 116008 34174 116014 34206
rect 115600 34136 115676 34142
rect 116013 34142 116014 34174
rect 116078 34174 116084 34206
rect 116960 34414 116966 34446
rect 117030 34446 117031 34478
rect 117030 34414 117036 34446
rect 116960 34206 117036 34414
rect 116078 34142 116079 34174
rect 116013 34141 116079 34142
rect 116960 34142 116966 34206
rect 117030 34142 117036 34206
rect 116960 34136 117036 34142
rect 115333 34070 115399 34071
rect 115333 34038 115334 34070
rect 28288 33902 28294 33934
rect 28293 33870 28294 33902
rect 28358 33902 28364 33934
rect 115328 34006 115334 34038
rect 115398 34038 115399 34070
rect 115600 34070 115676 34076
rect 115398 34006 115404 34038
rect 28358 33870 28359 33902
rect 28293 33869 28359 33870
rect 23054 33734 23055 33766
rect 22989 33733 23055 33734
rect 23528 33734 23534 33798
rect 23598 33734 23604 33798
rect 23528 33728 23604 33734
rect 115328 33798 115404 34006
rect 115328 33734 115334 33798
rect 115398 33734 115404 33798
rect 115600 34006 115606 34070
rect 115670 34006 115676 34070
rect 115600 33798 115676 34006
rect 115600 33766 115606 33798
rect 115328 33728 115404 33734
rect 115605 33734 115606 33766
rect 115670 33766 115676 33798
rect 116280 34070 116356 34076
rect 116280 34006 116286 34070
rect 116350 34006 116356 34070
rect 116280 33798 116356 34006
rect 116280 33766 116286 33798
rect 115670 33734 115671 33766
rect 115605 33733 115671 33734
rect 116285 33734 116286 33766
rect 116350 33766 116356 33798
rect 116552 34070 116628 34076
rect 116552 34006 116558 34070
rect 116622 34006 116628 34070
rect 116829 34070 116895 34071
rect 116829 34038 116830 34070
rect 116552 33798 116628 34006
rect 116552 33766 116558 33798
rect 116350 33734 116351 33766
rect 116285 33733 116351 33734
rect 116557 33734 116558 33766
rect 116622 33766 116628 33798
rect 116824 34006 116830 34038
rect 116894 34038 116895 34070
rect 137496 34070 137844 35638
rect 116894 34006 116900 34038
rect 116824 33798 116900 34006
rect 116622 33734 116623 33766
rect 116557 33733 116623 33734
rect 116824 33734 116830 33798
rect 116894 33734 116900 33798
rect 116824 33728 116900 33734
rect 137496 34006 137502 34070
rect 137566 34006 137844 34070
rect 14688 33630 14694 33662
rect 14693 33598 14694 33630
rect 14758 33630 14764 33662
rect 21896 33662 21972 33668
rect 14758 33598 14759 33630
rect 14693 33597 14759 33598
rect 21896 33598 21902 33662
rect 21966 33598 21972 33662
rect 14693 33526 14759 33527
rect 14693 33494 14694 33526
rect 14552 32238 14558 32302
rect 14622 32238 14628 32302
rect 14552 32232 14628 32238
rect 14688 33462 14694 33494
rect 14758 33494 14759 33526
rect 14758 33462 14764 33494
rect 14557 32166 14623 32167
rect 14557 32134 14558 32166
rect 952 30606 1230 30670
rect 1294 30606 1300 30670
rect 952 28902 1300 30606
rect 14552 32102 14558 32134
rect 14622 32134 14623 32166
rect 14622 32102 14628 32134
rect 14552 29446 14628 32102
rect 14688 30806 14764 33462
rect 21896 33390 21972 33598
rect 21896 33358 21902 33390
rect 21901 33326 21902 33358
rect 21966 33358 21972 33390
rect 23120 33662 23196 33668
rect 23120 33598 23126 33662
rect 23190 33598 23196 33662
rect 23120 33390 23196 33598
rect 23120 33358 23126 33390
rect 21966 33326 21967 33358
rect 21901 33325 21967 33326
rect 23125 33326 23126 33358
rect 23190 33358 23196 33390
rect 23392 33662 23468 33668
rect 23392 33598 23398 33662
rect 23462 33598 23468 33662
rect 23392 33390 23468 33598
rect 23392 33358 23398 33390
rect 23190 33326 23191 33358
rect 23125 33325 23191 33326
rect 23397 33326 23398 33358
rect 23462 33358 23468 33390
rect 115192 33662 115268 33668
rect 115192 33598 115198 33662
rect 115262 33598 115268 33662
rect 115192 33390 115268 33598
rect 115192 33358 115198 33390
rect 23462 33326 23463 33358
rect 23397 33325 23463 33326
rect 115197 33326 115198 33358
rect 115262 33358 115268 33390
rect 115600 33662 115676 33668
rect 115600 33598 115606 33662
rect 115670 33598 115676 33662
rect 115600 33390 115676 33598
rect 115600 33358 115606 33390
rect 115262 33326 115263 33358
rect 115197 33325 115263 33326
rect 115605 33326 115606 33358
rect 115670 33358 115676 33390
rect 116144 33662 116220 33668
rect 116144 33598 116150 33662
rect 116214 33598 116220 33662
rect 116144 33390 116220 33598
rect 116144 33358 116150 33390
rect 115670 33326 115671 33358
rect 115605 33325 115671 33326
rect 116149 33326 116150 33358
rect 116214 33358 116220 33390
rect 116960 33662 117036 33668
rect 116960 33598 116966 33662
rect 117030 33598 117036 33662
rect 116960 33390 117036 33598
rect 116960 33358 116966 33390
rect 116214 33326 116215 33358
rect 116149 33325 116215 33326
rect 116965 33326 116966 33358
rect 117030 33358 117036 33390
rect 117030 33326 117031 33358
rect 116965 33325 117031 33326
rect 21765 33254 21831 33255
rect 21765 33222 21766 33254
rect 21760 33190 21766 33222
rect 21830 33222 21831 33254
rect 22173 33254 22239 33255
rect 22173 33222 22174 33254
rect 21830 33190 21836 33222
rect 21760 32982 21836 33190
rect 21760 32918 21766 32982
rect 21830 32918 21836 32982
rect 21760 32912 21836 32918
rect 22168 33190 22174 33222
rect 22238 33222 22239 33254
rect 22576 33254 22652 33260
rect 22238 33190 22244 33222
rect 22168 32982 22244 33190
rect 22168 32918 22174 32982
rect 22238 32918 22244 32982
rect 22576 33190 22582 33254
rect 22646 33190 22652 33254
rect 22989 33254 23055 33255
rect 22989 33222 22990 33254
rect 22576 32982 22652 33190
rect 22576 32950 22582 32982
rect 22168 32912 22244 32918
rect 22581 32918 22582 32950
rect 22646 32950 22652 32982
rect 22984 33190 22990 33222
rect 23054 33222 23055 33254
rect 23528 33254 23604 33260
rect 23054 33190 23060 33222
rect 22984 32982 23060 33190
rect 22646 32918 22647 32950
rect 22581 32917 22647 32918
rect 22984 32918 22990 32982
rect 23054 32918 23060 32982
rect 23528 33190 23534 33254
rect 23598 33190 23604 33254
rect 23528 32982 23604 33190
rect 23528 32950 23534 32982
rect 22984 32912 23060 32918
rect 23533 32918 23534 32950
rect 23598 32950 23604 32982
rect 115328 33254 115404 33260
rect 115328 33190 115334 33254
rect 115398 33190 115404 33254
rect 115741 33254 115807 33255
rect 115741 33222 115742 33254
rect 115328 32982 115404 33190
rect 115328 32950 115334 32982
rect 23598 32918 23599 32950
rect 23533 32917 23599 32918
rect 115333 32918 115334 32950
rect 115398 32950 115404 32982
rect 115736 33190 115742 33222
rect 115806 33222 115807 33254
rect 116144 33254 116220 33260
rect 115806 33190 115812 33222
rect 115736 32982 115812 33190
rect 115398 32918 115399 32950
rect 115333 32917 115399 32918
rect 115736 32918 115742 32982
rect 115806 32918 115812 32982
rect 116144 33190 116150 33254
rect 116214 33190 116220 33254
rect 116421 33254 116487 33255
rect 116421 33222 116422 33254
rect 116144 32982 116220 33190
rect 116144 32950 116150 32982
rect 115736 32912 115812 32918
rect 116149 32918 116150 32950
rect 116214 32950 116220 32982
rect 116416 33190 116422 33222
rect 116486 33222 116487 33254
rect 116829 33254 116895 33255
rect 116829 33222 116830 33254
rect 116486 33190 116492 33222
rect 116416 32982 116492 33190
rect 116214 32918 116215 32950
rect 116149 32917 116215 32918
rect 116416 32918 116422 32982
rect 116486 32918 116492 32982
rect 116416 32912 116492 32918
rect 116824 33190 116830 33222
rect 116894 33222 116895 33254
rect 116894 33190 116900 33222
rect 116824 32982 116900 33190
rect 116824 32918 116830 32982
rect 116894 32918 116900 32982
rect 116824 32912 116900 32918
rect 21896 32846 21972 32852
rect 21896 32782 21902 32846
rect 21966 32782 21972 32846
rect 21896 32574 21972 32782
rect 21896 32542 21902 32574
rect 21901 32510 21902 32542
rect 21966 32542 21972 32574
rect 22304 32846 22380 32852
rect 22304 32782 22310 32846
rect 22374 32782 22380 32846
rect 22304 32574 22380 32782
rect 22304 32542 22310 32574
rect 21966 32510 21967 32542
rect 21901 32509 21967 32510
rect 22309 32510 22310 32542
rect 22374 32542 22380 32574
rect 22440 32846 22516 32852
rect 22440 32782 22446 32846
rect 22510 32782 22516 32846
rect 22440 32574 22516 32782
rect 22440 32542 22446 32574
rect 22374 32510 22375 32542
rect 22309 32509 22375 32510
rect 22445 32510 22446 32542
rect 22510 32542 22516 32574
rect 22984 32846 23060 32852
rect 22984 32782 22990 32846
rect 23054 32782 23060 32846
rect 23533 32846 23599 32847
rect 23533 32814 23534 32846
rect 22984 32574 23060 32782
rect 22984 32542 22990 32574
rect 22510 32510 22511 32542
rect 22445 32509 22511 32510
rect 22989 32510 22990 32542
rect 23054 32542 23060 32574
rect 23528 32782 23534 32814
rect 23598 32814 23599 32846
rect 115333 32846 115399 32847
rect 115333 32814 115334 32846
rect 23598 32782 23604 32814
rect 23528 32574 23604 32782
rect 23054 32510 23055 32542
rect 22989 32509 23055 32510
rect 23528 32510 23534 32574
rect 23598 32510 23604 32574
rect 23528 32504 23604 32510
rect 115328 32782 115334 32814
rect 115398 32814 115399 32846
rect 115600 32846 115676 32852
rect 115398 32782 115404 32814
rect 115328 32574 115404 32782
rect 115328 32510 115334 32574
rect 115398 32510 115404 32574
rect 115600 32782 115606 32846
rect 115670 32782 115676 32846
rect 115600 32574 115676 32782
rect 115600 32542 115606 32574
rect 115328 32504 115404 32510
rect 115605 32510 115606 32542
rect 115670 32542 115676 32574
rect 116008 32846 116084 32852
rect 116008 32782 116014 32846
rect 116078 32782 116084 32846
rect 116285 32846 116351 32847
rect 116285 32814 116286 32846
rect 116008 32574 116084 32782
rect 116008 32542 116014 32574
rect 115670 32510 115671 32542
rect 115605 32509 115671 32510
rect 116013 32510 116014 32542
rect 116078 32542 116084 32574
rect 116280 32782 116286 32814
rect 116350 32814 116351 32846
rect 116829 32846 116895 32847
rect 116829 32814 116830 32846
rect 116350 32782 116356 32814
rect 116280 32574 116356 32782
rect 116078 32510 116079 32542
rect 116013 32509 116079 32510
rect 116280 32510 116286 32574
rect 116350 32510 116356 32574
rect 116280 32504 116356 32510
rect 116824 32782 116830 32814
rect 116894 32814 116895 32846
rect 116894 32782 116900 32814
rect 116824 32574 116900 32782
rect 116824 32510 116830 32574
rect 116894 32510 116900 32574
rect 116824 32504 116900 32510
rect 21901 32438 21967 32439
rect 21901 32406 21902 32438
rect 21896 32374 21902 32406
rect 21966 32406 21967 32438
rect 22989 32438 23055 32439
rect 22989 32406 22990 32438
rect 21966 32374 21972 32406
rect 21896 32166 21972 32374
rect 21896 32102 21902 32166
rect 21966 32102 21972 32166
rect 21896 32096 21972 32102
rect 22984 32374 22990 32406
rect 23054 32406 23055 32438
rect 23397 32438 23463 32439
rect 23397 32406 23398 32438
rect 23054 32374 23060 32406
rect 22984 32166 23060 32374
rect 22984 32102 22990 32166
rect 23054 32102 23060 32166
rect 22984 32096 23060 32102
rect 23392 32374 23398 32406
rect 23462 32406 23463 32438
rect 115197 32438 115263 32439
rect 115197 32406 115198 32438
rect 23462 32374 23468 32406
rect 23392 32166 23468 32374
rect 23392 32102 23398 32166
rect 23462 32102 23468 32166
rect 23392 32096 23468 32102
rect 115192 32374 115198 32406
rect 115262 32406 115263 32438
rect 115605 32438 115671 32439
rect 115605 32406 115606 32438
rect 115262 32374 115268 32406
rect 115192 32166 115268 32374
rect 115192 32102 115198 32166
rect 115262 32102 115268 32166
rect 115192 32096 115268 32102
rect 115600 32374 115606 32406
rect 115670 32406 115671 32438
rect 116008 32438 116084 32444
rect 115670 32374 115676 32406
rect 115600 32166 115676 32374
rect 115600 32102 115606 32166
rect 115670 32102 115676 32166
rect 116008 32374 116014 32438
rect 116078 32374 116084 32438
rect 116285 32438 116351 32439
rect 116285 32406 116286 32438
rect 116008 32166 116084 32374
rect 116008 32134 116014 32166
rect 115600 32096 115676 32102
rect 116013 32102 116014 32134
rect 116078 32134 116084 32166
rect 116280 32374 116286 32406
rect 116350 32406 116351 32438
rect 116965 32438 117031 32439
rect 116965 32406 116966 32438
rect 116350 32374 116356 32406
rect 116280 32166 116356 32374
rect 116078 32102 116079 32134
rect 116013 32101 116079 32102
rect 116280 32102 116286 32166
rect 116350 32102 116356 32166
rect 116280 32096 116356 32102
rect 116960 32374 116966 32406
rect 117030 32406 117031 32438
rect 137496 32438 137844 34006
rect 117030 32374 117036 32406
rect 116960 32166 117036 32374
rect 116960 32102 116966 32166
rect 117030 32102 117036 32166
rect 116960 32096 117036 32102
rect 137496 32374 137502 32438
rect 137566 32374 137844 32438
rect 22581 32030 22647 32031
rect 22581 31998 22582 32030
rect 22576 31966 22582 31998
rect 22646 31998 22647 32030
rect 23120 32030 23196 32036
rect 22646 31966 22652 31998
rect 21765 31758 21831 31759
rect 21765 31726 21766 31758
rect 21760 31694 21766 31726
rect 21830 31726 21831 31758
rect 22576 31758 22652 31966
rect 21830 31694 21836 31726
rect 21760 31486 21836 31694
rect 22576 31694 22582 31758
rect 22646 31694 22652 31758
rect 23120 31966 23126 32030
rect 23190 31966 23196 32030
rect 23120 31758 23196 31966
rect 23120 31726 23126 31758
rect 22576 31688 22652 31694
rect 23125 31694 23126 31726
rect 23190 31726 23196 31758
rect 23528 32030 23604 32036
rect 23528 31966 23534 32030
rect 23598 31966 23604 32030
rect 23528 31758 23604 31966
rect 115328 32030 115404 32036
rect 115328 31966 115334 32030
rect 115398 31966 115404 32030
rect 110165 31894 110231 31895
rect 110165 31862 110166 31894
rect 23528 31726 23534 31758
rect 23190 31694 23191 31726
rect 23125 31693 23191 31694
rect 23533 31694 23534 31726
rect 23598 31726 23604 31758
rect 110160 31830 110166 31862
rect 110230 31862 110231 31894
rect 110230 31830 110236 31862
rect 23598 31694 23599 31726
rect 23533 31693 23599 31694
rect 22989 31622 23055 31623
rect 22989 31590 22990 31622
rect 21760 31422 21766 31486
rect 21830 31422 21836 31486
rect 21760 31416 21836 31422
rect 22984 31558 22990 31590
rect 23054 31590 23055 31622
rect 23397 31622 23463 31623
rect 23397 31590 23398 31622
rect 23054 31558 23060 31590
rect 22984 31350 23060 31558
rect 22984 31286 22990 31350
rect 23054 31286 23060 31350
rect 22984 31280 23060 31286
rect 23392 31558 23398 31590
rect 23462 31590 23463 31622
rect 110160 31622 110236 31830
rect 115328 31758 115404 31966
rect 115328 31726 115334 31758
rect 115333 31694 115334 31726
rect 115398 31726 115404 31758
rect 115736 32030 115812 32036
rect 115736 31966 115742 32030
rect 115806 31966 115812 32030
rect 115736 31758 115812 31966
rect 115736 31726 115742 31758
rect 115398 31694 115399 31726
rect 115333 31693 115399 31694
rect 115741 31694 115742 31726
rect 115806 31726 115812 31758
rect 116144 31824 116492 31900
rect 116144 31758 116220 31824
rect 116144 31726 116150 31758
rect 115806 31694 115807 31726
rect 115741 31693 115807 31694
rect 116149 31694 116150 31726
rect 116214 31726 116220 31758
rect 116285 31758 116351 31759
rect 116285 31726 116286 31758
rect 116214 31694 116215 31726
rect 116149 31693 116215 31694
rect 116280 31694 116286 31726
rect 116350 31726 116351 31758
rect 116416 31758 116492 31824
rect 116350 31694 116356 31726
rect 23462 31558 23468 31590
rect 23392 31350 23468 31558
rect 110160 31558 110166 31622
rect 110230 31558 110236 31622
rect 110160 31552 110236 31558
rect 115192 31622 115268 31628
rect 115192 31558 115198 31622
rect 115262 31558 115268 31622
rect 115605 31622 115671 31623
rect 115605 31590 115606 31622
rect 23392 31286 23398 31350
rect 23462 31286 23468 31350
rect 115192 31350 115268 31558
rect 115192 31318 115198 31350
rect 23392 31280 23468 31286
rect 115197 31286 115198 31318
rect 115262 31318 115268 31350
rect 115600 31558 115606 31590
rect 115670 31590 115671 31622
rect 115670 31558 115676 31590
rect 115600 31350 115676 31558
rect 116280 31492 116356 31694
rect 116416 31694 116422 31758
rect 116486 31694 116492 31758
rect 116829 31758 116895 31759
rect 116829 31726 116830 31758
rect 116416 31688 116492 31694
rect 116824 31694 116830 31726
rect 116894 31726 116895 31758
rect 116894 31694 116900 31726
rect 116280 31486 116492 31492
rect 116280 31422 116422 31486
rect 116486 31422 116492 31486
rect 116280 31416 116492 31422
rect 116824 31486 116900 31694
rect 116824 31422 116830 31486
rect 116894 31422 116900 31486
rect 116824 31416 116900 31422
rect 115262 31286 115263 31318
rect 115197 31285 115263 31286
rect 115600 31286 115606 31350
rect 115670 31286 115676 31350
rect 115600 31280 115676 31286
rect 22576 31214 22652 31220
rect 22576 31150 22582 31214
rect 22646 31150 22652 31214
rect 14688 30742 14694 30806
rect 14758 30742 14764 30806
rect 14688 30736 14764 30742
rect 21760 30942 21836 30948
rect 21760 30878 21766 30942
rect 21830 30878 21836 30942
rect 22576 30942 22652 31150
rect 116008 31214 116084 31220
rect 116008 31150 116014 31214
rect 116078 31150 116084 31214
rect 28293 31078 28359 31079
rect 28293 31046 28294 31078
rect 22576 30910 22582 30942
rect 18501 30670 18567 30671
rect 18501 30638 18502 30670
rect 14552 29382 14558 29446
rect 14622 29382 14628 29446
rect 14552 29376 14628 29382
rect 18496 30606 18502 30638
rect 18566 30638 18567 30670
rect 21760 30670 21836 30878
rect 22581 30878 22582 30910
rect 22646 30910 22652 30942
rect 28288 31014 28294 31046
rect 28358 31046 28359 31078
rect 28358 31014 28364 31046
rect 22646 30878 22647 30910
rect 22581 30877 22647 30878
rect 28288 30806 28364 31014
rect 116008 30942 116084 31150
rect 116008 30910 116014 30942
rect 116013 30878 116014 30910
rect 116078 30910 116084 30942
rect 116829 30942 116895 30943
rect 116829 30910 116830 30942
rect 116078 30878 116079 30910
rect 116013 30877 116079 30878
rect 116824 30878 116830 30910
rect 116894 30910 116895 30942
rect 116894 30878 116900 30910
rect 28288 30742 28294 30806
rect 28358 30742 28364 30806
rect 28288 30736 28364 30742
rect 21760 30638 21766 30670
rect 18566 30606 18572 30638
rect 16597 29310 16663 29311
rect 16597 29278 16598 29310
rect 952 28838 1230 28902
rect 1294 28838 1300 28902
rect 952 27406 1300 28838
rect 952 27342 1230 27406
rect 1294 27342 1300 27406
rect 952 25638 1300 27342
rect 16592 29246 16598 29278
rect 16662 29278 16663 29310
rect 16662 29246 16668 29278
rect 16592 26726 16668 29246
rect 18496 29038 18572 30606
rect 21765 30606 21766 30638
rect 21830 30638 21836 30670
rect 28288 30670 28364 30676
rect 21830 30606 21831 30638
rect 21765 30605 21831 30606
rect 28288 30606 28294 30670
rect 28358 30606 28364 30670
rect 110437 30670 110503 30671
rect 110437 30638 110438 30670
rect 21901 30534 21967 30535
rect 21901 30502 21902 30534
rect 21896 30470 21902 30502
rect 21966 30502 21967 30534
rect 22440 30534 22516 30540
rect 21966 30470 21972 30502
rect 21896 30262 21972 30470
rect 21896 30198 21902 30262
rect 21966 30198 21972 30262
rect 22440 30470 22446 30534
rect 22510 30470 22516 30534
rect 22440 30262 22516 30470
rect 22440 30230 22446 30262
rect 21896 30192 21972 30198
rect 22445 30198 22446 30230
rect 22510 30230 22516 30262
rect 22712 30534 22788 30540
rect 22712 30470 22718 30534
rect 22782 30470 22788 30534
rect 22712 30262 22788 30470
rect 28288 30398 28364 30606
rect 28288 30366 28294 30398
rect 28293 30334 28294 30366
rect 28358 30366 28364 30398
rect 110432 30606 110438 30638
rect 110502 30638 110503 30670
rect 116824 30670 116900 30878
rect 110502 30606 110508 30638
rect 110432 30398 110508 30606
rect 116824 30606 116830 30670
rect 116894 30606 116900 30670
rect 116824 30600 116900 30606
rect 116285 30534 116351 30535
rect 116285 30502 116286 30534
rect 28358 30334 28359 30366
rect 28293 30333 28359 30334
rect 110432 30334 110438 30398
rect 110502 30334 110508 30398
rect 110432 30328 110508 30334
rect 116280 30470 116286 30502
rect 116350 30502 116351 30534
rect 116960 30534 117036 30540
rect 116350 30470 116356 30502
rect 22712 30230 22718 30262
rect 22510 30198 22511 30230
rect 22445 30197 22511 30198
rect 22717 30198 22718 30230
rect 22782 30230 22788 30262
rect 28288 30262 28364 30268
rect 22782 30198 22783 30230
rect 22717 30197 22783 30198
rect 28288 30198 28294 30262
rect 28358 30198 28364 30262
rect 21760 30126 21836 30132
rect 21760 30062 21766 30126
rect 21830 30062 21836 30126
rect 23125 30126 23191 30127
rect 23125 30094 23126 30126
rect 21760 29854 21836 30062
rect 21760 29822 21766 29854
rect 21765 29790 21766 29822
rect 21830 29822 21836 29854
rect 23120 30062 23126 30094
rect 23190 30094 23191 30126
rect 23397 30126 23463 30127
rect 23397 30094 23398 30126
rect 23190 30062 23196 30094
rect 23120 29854 23196 30062
rect 21830 29790 21831 29822
rect 21765 29789 21831 29790
rect 23120 29790 23126 29854
rect 23190 29790 23196 29854
rect 23120 29784 23196 29790
rect 23392 30062 23398 30094
rect 23462 30094 23463 30126
rect 23462 30062 23468 30094
rect 23392 29854 23468 30062
rect 28288 29990 28364 30198
rect 28288 29958 28294 29990
rect 28293 29926 28294 29958
rect 28358 29958 28364 29990
rect 110160 30262 110236 30268
rect 110160 30198 110166 30262
rect 110230 30198 110236 30262
rect 110160 29990 110236 30198
rect 116280 30262 116356 30470
rect 116280 30198 116286 30262
rect 116350 30198 116356 30262
rect 116960 30470 116966 30534
rect 117030 30470 117036 30534
rect 116960 30262 117036 30470
rect 116960 30230 116966 30262
rect 116280 30192 116356 30198
rect 116965 30198 116966 30230
rect 117030 30230 117036 30262
rect 137496 30534 137844 32374
rect 137496 30470 137502 30534
rect 137566 30470 137844 30534
rect 117030 30198 117031 30230
rect 116965 30197 117031 30198
rect 110160 29958 110166 29990
rect 28358 29926 28359 29958
rect 28293 29925 28359 29926
rect 110165 29926 110166 29958
rect 110230 29958 110236 29990
rect 115328 30126 115404 30132
rect 115328 30062 115334 30126
rect 115398 30062 115404 30126
rect 110230 29926 110231 29958
rect 110165 29925 110231 29926
rect 23392 29790 23398 29854
rect 23462 29790 23468 29854
rect 115328 29854 115404 30062
rect 115328 29822 115334 29854
rect 23392 29784 23468 29790
rect 115333 29790 115334 29822
rect 115398 29822 115404 29854
rect 115736 30126 115812 30132
rect 115736 30062 115742 30126
rect 115806 30062 115812 30126
rect 116965 30126 117031 30127
rect 116965 30094 116966 30126
rect 115736 29854 115812 30062
rect 115736 29822 115742 29854
rect 115398 29790 115399 29822
rect 115333 29789 115399 29790
rect 115741 29790 115742 29822
rect 115806 29822 115812 29854
rect 116960 30062 116966 30094
rect 117030 30094 117031 30126
rect 117030 30062 117036 30094
rect 116960 29854 117036 30062
rect 115806 29790 115807 29822
rect 115741 29789 115807 29790
rect 116960 29790 116966 29854
rect 117030 29790 117036 29854
rect 116960 29784 117036 29790
rect 21765 29718 21831 29719
rect 21765 29686 21766 29718
rect 21760 29654 21766 29686
rect 21830 29686 21831 29718
rect 22581 29718 22647 29719
rect 22581 29686 22582 29718
rect 21830 29654 21836 29686
rect 21760 29446 21836 29654
rect 21760 29382 21766 29446
rect 21830 29382 21836 29446
rect 21760 29376 21836 29382
rect 22576 29654 22582 29686
rect 22646 29686 22647 29718
rect 22984 29718 23060 29724
rect 22646 29654 22652 29686
rect 22576 29446 22652 29654
rect 22576 29382 22582 29446
rect 22646 29382 22652 29446
rect 22984 29654 22990 29718
rect 23054 29654 23060 29718
rect 22984 29446 23060 29654
rect 22984 29414 22990 29446
rect 22576 29376 22652 29382
rect 22989 29382 22990 29414
rect 23054 29414 23060 29446
rect 23392 29718 23468 29724
rect 23392 29654 23398 29718
rect 23462 29654 23468 29718
rect 23392 29446 23468 29654
rect 23392 29414 23398 29446
rect 23054 29382 23055 29414
rect 22989 29381 23055 29382
rect 23397 29382 23398 29414
rect 23462 29414 23468 29446
rect 115192 29718 115268 29724
rect 115192 29654 115198 29718
rect 115262 29654 115268 29718
rect 115192 29446 115268 29654
rect 115192 29414 115198 29446
rect 23462 29382 23463 29414
rect 23397 29381 23463 29382
rect 115197 29382 115198 29414
rect 115262 29414 115268 29446
rect 115600 29718 115676 29724
rect 115600 29654 115606 29718
rect 115670 29654 115676 29718
rect 116013 29718 116079 29719
rect 116013 29686 116014 29718
rect 115600 29446 115676 29654
rect 115600 29414 115606 29446
rect 115262 29382 115263 29414
rect 115197 29381 115263 29382
rect 115605 29382 115606 29414
rect 115670 29414 115676 29446
rect 116008 29654 116014 29686
rect 116078 29686 116079 29718
rect 116960 29718 117036 29724
rect 116078 29654 116084 29686
rect 116008 29446 116084 29654
rect 115670 29382 115671 29414
rect 115605 29381 115671 29382
rect 116008 29382 116014 29446
rect 116078 29382 116084 29446
rect 116960 29654 116966 29718
rect 117030 29654 117036 29718
rect 116960 29446 117036 29654
rect 116960 29414 116966 29446
rect 116008 29376 116084 29382
rect 116965 29382 116966 29414
rect 117030 29414 117036 29446
rect 117030 29382 117031 29414
rect 116965 29381 117031 29382
rect 18496 28974 18502 29038
rect 18566 28974 18572 29038
rect 21896 29310 21972 29316
rect 21896 29246 21902 29310
rect 21966 29246 21972 29310
rect 21896 29038 21972 29246
rect 21896 29006 21902 29038
rect 18496 28968 18572 28974
rect 21901 28974 21902 29006
rect 21966 29006 21972 29038
rect 22712 29310 22788 29316
rect 22712 29246 22718 29310
rect 22782 29246 22788 29310
rect 22989 29310 23055 29311
rect 22989 29278 22990 29310
rect 22712 29038 22788 29246
rect 22712 29006 22718 29038
rect 21966 28974 21967 29006
rect 21901 28973 21967 28974
rect 22717 28974 22718 29006
rect 22782 29006 22788 29038
rect 22984 29246 22990 29278
rect 23054 29278 23055 29310
rect 23392 29310 23468 29316
rect 23054 29246 23060 29278
rect 22984 29038 23060 29246
rect 22782 28974 22783 29006
rect 22717 28973 22783 28974
rect 22984 28974 22990 29038
rect 23054 28974 23060 29038
rect 23392 29246 23398 29310
rect 23462 29246 23468 29310
rect 115197 29310 115263 29311
rect 115197 29278 115198 29310
rect 23392 29038 23468 29246
rect 23392 29006 23398 29038
rect 22984 28968 23060 28974
rect 23397 28974 23398 29006
rect 23462 29006 23468 29038
rect 115192 29246 115198 29278
rect 115262 29278 115263 29310
rect 115605 29310 115671 29311
rect 115605 29278 115606 29310
rect 115262 29246 115268 29278
rect 115192 29038 115268 29246
rect 23462 28974 23463 29006
rect 23397 28973 23463 28974
rect 115192 28974 115198 29038
rect 115262 28974 115268 29038
rect 115192 28968 115268 28974
rect 115600 29246 115606 29278
rect 115670 29278 115671 29310
rect 116144 29310 116220 29316
rect 115670 29246 115676 29278
rect 115600 29038 115676 29246
rect 115600 28974 115606 29038
rect 115670 28974 115676 29038
rect 116144 29246 116150 29310
rect 116214 29246 116220 29310
rect 116144 29038 116220 29246
rect 116144 29006 116150 29038
rect 115600 28968 115676 28974
rect 116149 28974 116150 29006
rect 116214 29006 116220 29038
rect 116960 29310 117036 29316
rect 116960 29246 116966 29310
rect 117030 29246 117036 29310
rect 116960 29038 117036 29246
rect 116960 29006 116966 29038
rect 116214 28974 116215 29006
rect 116149 28973 116215 28974
rect 116965 28974 116966 29006
rect 117030 29006 117036 29038
rect 137496 29038 137844 30470
rect 117030 28974 117031 29006
rect 116965 28973 117031 28974
rect 137496 28974 137502 29038
rect 137566 28974 137844 29038
rect 18093 28902 18159 28903
rect 18093 28870 18094 28902
rect 18088 28838 18094 28870
rect 18158 28870 18159 28902
rect 18909 28902 18975 28903
rect 18909 28870 18910 28902
rect 18158 28838 18164 28870
rect 18088 28222 18164 28838
rect 18088 28158 18094 28222
rect 18158 28158 18164 28222
rect 18088 28152 18164 28158
rect 18904 28838 18910 28870
rect 18974 28870 18975 28902
rect 19448 28902 19524 28908
rect 18974 28838 18980 28870
rect 18904 28222 18980 28838
rect 18904 28158 18910 28222
rect 18974 28158 18980 28222
rect 19448 28838 19454 28902
rect 19518 28838 19524 28902
rect 21765 28902 21831 28903
rect 21765 28870 21766 28902
rect 19448 28222 19524 28838
rect 21760 28838 21766 28870
rect 21830 28870 21831 28902
rect 22168 28902 22244 28908
rect 21830 28838 21836 28870
rect 21760 28630 21836 28838
rect 21760 28566 21766 28630
rect 21830 28566 21836 28630
rect 22168 28838 22174 28902
rect 22238 28838 22244 28902
rect 22445 28902 22511 28903
rect 22445 28870 22446 28902
rect 22168 28630 22244 28838
rect 22168 28598 22174 28630
rect 21760 28560 21836 28566
rect 22173 28566 22174 28598
rect 22238 28598 22244 28630
rect 22440 28838 22446 28870
rect 22510 28870 22511 28902
rect 22989 28902 23055 28903
rect 22989 28870 22990 28902
rect 22510 28838 22516 28870
rect 22440 28630 22516 28838
rect 22238 28566 22239 28598
rect 22173 28565 22239 28566
rect 22440 28566 22446 28630
rect 22510 28566 22516 28630
rect 22440 28560 22516 28566
rect 22984 28838 22990 28870
rect 23054 28870 23055 28902
rect 23533 28902 23599 28903
rect 23533 28870 23534 28902
rect 23054 28838 23060 28870
rect 22984 28630 23060 28838
rect 22984 28566 22990 28630
rect 23054 28566 23060 28630
rect 22984 28560 23060 28566
rect 23528 28838 23534 28870
rect 23598 28870 23599 28902
rect 115328 28902 115404 28908
rect 23598 28838 23604 28870
rect 23528 28630 23604 28838
rect 23528 28566 23534 28630
rect 23598 28566 23604 28630
rect 115328 28838 115334 28902
rect 115398 28838 115404 28902
rect 115328 28630 115404 28838
rect 115328 28598 115334 28630
rect 23528 28560 23604 28566
rect 115333 28566 115334 28598
rect 115398 28598 115404 28630
rect 115736 28902 115812 28908
rect 115736 28838 115742 28902
rect 115806 28838 115812 28902
rect 116013 28902 116079 28903
rect 116013 28870 116014 28902
rect 115736 28630 115812 28838
rect 115736 28598 115742 28630
rect 115398 28566 115399 28598
rect 115333 28565 115399 28566
rect 115741 28566 115742 28598
rect 115806 28598 115812 28630
rect 116008 28838 116014 28870
rect 116078 28870 116079 28902
rect 116829 28902 116895 28903
rect 116829 28870 116830 28902
rect 116078 28838 116084 28870
rect 116008 28630 116084 28838
rect 115806 28566 115807 28598
rect 115741 28565 115807 28566
rect 116008 28566 116014 28630
rect 116078 28566 116084 28630
rect 116008 28560 116084 28566
rect 116824 28838 116830 28870
rect 116894 28870 116895 28902
rect 119005 28902 119071 28903
rect 119005 28870 119006 28902
rect 116894 28838 116900 28870
rect 116824 28630 116900 28838
rect 116824 28566 116830 28630
rect 116894 28566 116900 28630
rect 116824 28560 116900 28566
rect 119000 28838 119006 28870
rect 119070 28870 119071 28902
rect 119272 28902 119348 28908
rect 119070 28838 119076 28870
rect 21765 28494 21831 28495
rect 21765 28462 21766 28494
rect 19448 28190 19454 28222
rect 18904 28152 18980 28158
rect 19453 28158 19454 28190
rect 19518 28190 19524 28222
rect 21760 28430 21766 28462
rect 21830 28462 21831 28494
rect 22984 28494 23060 28500
rect 21830 28430 21836 28462
rect 21760 28222 21836 28430
rect 19518 28158 19519 28190
rect 19453 28157 19519 28158
rect 21760 28158 21766 28222
rect 21830 28158 21836 28222
rect 22984 28430 22990 28494
rect 23054 28430 23060 28494
rect 22984 28222 23060 28430
rect 22984 28190 22990 28222
rect 21760 28152 21836 28158
rect 22989 28158 22990 28190
rect 23054 28190 23060 28222
rect 23392 28494 23468 28500
rect 23392 28430 23398 28494
rect 23462 28430 23468 28494
rect 115333 28494 115399 28495
rect 115333 28462 115334 28494
rect 23392 28222 23468 28430
rect 23392 28190 23398 28222
rect 23054 28158 23055 28190
rect 22989 28157 23055 28158
rect 23397 28158 23398 28190
rect 23462 28190 23468 28222
rect 115328 28430 115334 28462
rect 115398 28462 115399 28494
rect 115741 28494 115807 28495
rect 115741 28462 115742 28494
rect 115398 28430 115404 28462
rect 115328 28222 115404 28430
rect 23462 28158 23463 28190
rect 23397 28157 23463 28158
rect 115328 28158 115334 28222
rect 115398 28158 115404 28222
rect 115328 28152 115404 28158
rect 115736 28430 115742 28462
rect 115806 28462 115807 28494
rect 116960 28494 117036 28500
rect 115806 28430 115812 28462
rect 115736 28222 115812 28430
rect 115736 28158 115742 28222
rect 115806 28158 115812 28222
rect 116960 28430 116966 28494
rect 117030 28430 117036 28494
rect 116960 28222 117036 28430
rect 116960 28190 116966 28222
rect 115736 28152 115812 28158
rect 116965 28158 116966 28190
rect 117030 28190 117036 28222
rect 119000 28222 119076 28838
rect 117030 28158 117031 28190
rect 116965 28157 117031 28158
rect 119000 28158 119006 28222
rect 119070 28158 119076 28222
rect 119272 28838 119278 28902
rect 119342 28838 119348 28902
rect 119272 28222 119348 28838
rect 119272 28190 119278 28222
rect 119000 28152 119076 28158
rect 119277 28158 119278 28190
rect 119342 28190 119348 28222
rect 119952 28902 120028 28908
rect 119952 28838 119958 28902
rect 120022 28838 120028 28902
rect 120501 28902 120567 28903
rect 120501 28870 120502 28902
rect 119952 28222 120028 28838
rect 119952 28190 119958 28222
rect 119342 28158 119343 28190
rect 119277 28157 119343 28158
rect 119957 28158 119958 28190
rect 120022 28190 120028 28222
rect 120496 28838 120502 28870
rect 120566 28870 120567 28902
rect 120566 28838 120572 28870
rect 120496 28222 120572 28838
rect 120022 28158 120023 28190
rect 119957 28157 120023 28158
rect 120496 28158 120502 28222
rect 120566 28158 120572 28222
rect 120496 28152 120572 28158
rect 18088 28086 18164 28092
rect 18088 28022 18094 28086
rect 18158 28022 18164 28086
rect 18088 27542 18164 28022
rect 18088 27510 18094 27542
rect 18093 27478 18094 27510
rect 18158 27510 18164 27542
rect 19040 28086 19116 28092
rect 19040 28022 19046 28086
rect 19110 28022 19116 28086
rect 19453 28086 19519 28087
rect 19453 28054 19454 28086
rect 19040 27542 19116 28022
rect 19448 28022 19454 28054
rect 19518 28054 19519 28086
rect 19725 28086 19791 28087
rect 19725 28054 19726 28086
rect 19518 28022 19524 28054
rect 19317 27678 19383 27679
rect 19317 27646 19318 27678
rect 19040 27510 19046 27542
rect 18158 27478 18159 27510
rect 18093 27477 18159 27478
rect 19045 27478 19046 27510
rect 19110 27510 19116 27542
rect 19312 27614 19318 27646
rect 19382 27646 19383 27678
rect 19382 27614 19388 27646
rect 19110 27478 19111 27510
rect 19045 27477 19111 27478
rect 19312 27406 19388 27614
rect 19312 27342 19318 27406
rect 19382 27342 19388 27406
rect 19312 27336 19388 27342
rect 19448 27406 19524 28022
rect 19448 27342 19454 27406
rect 19518 27342 19524 27406
rect 19448 27336 19524 27342
rect 19720 28022 19726 28054
rect 19790 28054 19791 28086
rect 22309 28086 22375 28087
rect 22309 28054 22310 28086
rect 19790 28022 19796 28054
rect 19720 27406 19796 28022
rect 22304 28022 22310 28054
rect 22374 28054 22375 28086
rect 22717 28086 22783 28087
rect 22717 28054 22718 28086
rect 22374 28022 22380 28054
rect 22304 27814 22380 28022
rect 22304 27750 22310 27814
rect 22374 27750 22380 27814
rect 22304 27744 22380 27750
rect 22712 28022 22718 28054
rect 22782 28054 22783 28086
rect 22989 28086 23055 28087
rect 22989 28054 22990 28086
rect 22782 28022 22788 28054
rect 22712 27814 22788 28022
rect 22712 27750 22718 27814
rect 22782 27750 22788 27814
rect 22712 27744 22788 27750
rect 22984 28022 22990 28054
rect 23054 28054 23055 28086
rect 23397 28086 23463 28087
rect 23397 28054 23398 28086
rect 23054 28022 23060 28054
rect 22984 27814 23060 28022
rect 22984 27750 22990 27814
rect 23054 27750 23060 27814
rect 22984 27744 23060 27750
rect 23392 28022 23398 28054
rect 23462 28054 23463 28086
rect 115328 28086 115404 28092
rect 23462 28022 23468 28054
rect 23392 27814 23468 28022
rect 115328 28022 115334 28086
rect 115398 28022 115404 28086
rect 23392 27750 23398 27814
rect 23462 27750 23468 27814
rect 23392 27744 23468 27750
rect 28288 27950 28364 27956
rect 28288 27886 28294 27950
rect 28358 27886 28364 27950
rect 19720 27342 19726 27406
rect 19790 27342 19796 27406
rect 23120 27678 23196 27684
rect 23120 27614 23126 27678
rect 23190 27614 23196 27678
rect 23120 27406 23196 27614
rect 23120 27374 23126 27406
rect 19720 27336 19796 27342
rect 23125 27342 23126 27374
rect 23190 27374 23196 27406
rect 23528 27678 23604 27684
rect 23528 27614 23534 27678
rect 23598 27614 23604 27678
rect 28288 27678 28364 27886
rect 115328 27814 115404 28022
rect 115328 27782 115334 27814
rect 115333 27750 115334 27782
rect 115398 27782 115404 27814
rect 115736 28086 115812 28092
rect 115736 28022 115742 28086
rect 115806 28022 115812 28086
rect 115736 27814 115812 28022
rect 115736 27782 115742 27814
rect 115398 27750 115399 27782
rect 115333 27749 115399 27750
rect 115741 27750 115742 27782
rect 115806 27782 115812 27814
rect 116008 28086 116084 28092
rect 116008 28022 116014 28086
rect 116078 28022 116084 28086
rect 116008 27814 116084 28022
rect 116008 27782 116014 27814
rect 115806 27750 115807 27782
rect 115741 27749 115807 27750
rect 116013 27750 116014 27782
rect 116078 27782 116084 27814
rect 119000 28086 119076 28092
rect 119000 28022 119006 28086
rect 119070 28022 119076 28086
rect 116078 27750 116079 27782
rect 116013 27749 116079 27750
rect 28288 27646 28294 27678
rect 23528 27406 23604 27614
rect 28293 27614 28294 27646
rect 28358 27646 28364 27678
rect 115328 27678 115404 27684
rect 28358 27614 28359 27646
rect 28293 27613 28359 27614
rect 115328 27614 115334 27678
rect 115398 27614 115404 27678
rect 115741 27678 115807 27679
rect 115741 27646 115742 27678
rect 23528 27374 23534 27406
rect 23190 27342 23191 27374
rect 23125 27341 23191 27342
rect 23533 27342 23534 27374
rect 23598 27374 23604 27406
rect 28424 27406 28500 27412
rect 23598 27342 23599 27374
rect 23533 27341 23599 27342
rect 28424 27342 28430 27406
rect 28494 27342 28500 27406
rect 16592 26662 16598 26726
rect 16662 26662 16668 26726
rect 18088 27270 18164 27276
rect 18088 27206 18094 27270
rect 18158 27206 18164 27270
rect 18088 26726 18164 27206
rect 18088 26694 18094 26726
rect 16592 26656 16668 26662
rect 18093 26662 18094 26694
rect 18158 26694 18164 26726
rect 18496 27270 18572 27276
rect 18496 27206 18502 27270
rect 18566 27206 18572 27270
rect 18158 26662 18159 26694
rect 18093 26661 18159 26662
rect 18496 26454 18572 27206
rect 19312 27270 19388 27276
rect 19312 27206 19318 27270
rect 19382 27206 19388 27270
rect 18909 27134 18975 27135
rect 18909 27102 18910 27134
rect 18904 27070 18910 27102
rect 18974 27102 18975 27134
rect 18974 27070 18980 27102
rect 18904 26726 18980 27070
rect 18904 26662 18910 26726
rect 18974 26662 18980 26726
rect 19312 26726 19388 27206
rect 19312 26694 19318 26726
rect 18904 26656 18980 26662
rect 19317 26662 19318 26694
rect 19382 26694 19388 26726
rect 19856 27270 19932 27276
rect 19856 27206 19862 27270
rect 19926 27206 19932 27270
rect 19856 26726 19932 27206
rect 22304 27270 22380 27276
rect 22304 27206 22310 27270
rect 22374 27206 22380 27270
rect 21901 26998 21967 26999
rect 21901 26966 21902 26998
rect 19856 26694 19862 26726
rect 19382 26662 19383 26694
rect 19317 26661 19383 26662
rect 19861 26662 19862 26694
rect 19926 26694 19932 26726
rect 21896 26934 21902 26966
rect 21966 26966 21967 26998
rect 22304 26998 22380 27206
rect 28424 27134 28500 27342
rect 110160 27406 110236 27412
rect 110160 27342 110166 27406
rect 110230 27342 110236 27406
rect 115328 27406 115404 27614
rect 115328 27374 115334 27406
rect 28424 27102 28430 27134
rect 28429 27070 28430 27102
rect 28494 27102 28500 27134
rect 28565 27134 28631 27135
rect 28565 27102 28566 27134
rect 28494 27070 28495 27102
rect 28429 27069 28495 27070
rect 28560 27070 28566 27102
rect 28630 27102 28631 27134
rect 110160 27134 110236 27342
rect 115333 27342 115334 27374
rect 115398 27374 115404 27406
rect 115736 27614 115742 27646
rect 115806 27646 115807 27678
rect 115806 27614 115812 27646
rect 115736 27406 115812 27614
rect 115398 27342 115399 27374
rect 115333 27341 115399 27342
rect 115736 27342 115742 27406
rect 115806 27342 115812 27406
rect 119000 27406 119076 28022
rect 119000 27374 119006 27406
rect 115736 27336 115812 27342
rect 119005 27342 119006 27374
rect 119070 27374 119076 27406
rect 119408 28086 119484 28092
rect 119408 28022 119414 28086
rect 119478 28022 119484 28086
rect 119957 28086 120023 28087
rect 119957 28054 119958 28086
rect 119408 27406 119484 28022
rect 119952 28022 119958 28054
rect 120022 28054 120023 28086
rect 120637 28086 120703 28087
rect 120637 28054 120638 28086
rect 120022 28022 120028 28054
rect 119952 27542 120028 28022
rect 119952 27478 119958 27542
rect 120022 27478 120028 27542
rect 119952 27472 120028 27478
rect 120632 28022 120638 28054
rect 120702 28054 120703 28086
rect 120702 28022 120708 28054
rect 120632 27542 120708 28022
rect 120632 27478 120638 27542
rect 120702 27478 120708 27542
rect 120632 27472 120708 27478
rect 119408 27374 119414 27406
rect 119070 27342 119071 27374
rect 119005 27341 119071 27342
rect 119413 27342 119414 27374
rect 119478 27374 119484 27406
rect 119478 27342 119479 27374
rect 119413 27341 119479 27342
rect 116552 27270 116628 27276
rect 116552 27206 116558 27270
rect 116622 27206 116628 27270
rect 119277 27270 119343 27271
rect 119277 27238 119278 27270
rect 110160 27102 110166 27134
rect 28630 27070 28636 27102
rect 22304 26966 22310 26998
rect 21966 26934 21972 26966
rect 21896 26726 21972 26934
rect 22309 26934 22310 26966
rect 22374 26966 22380 26998
rect 22374 26934 22375 26966
rect 22309 26933 22375 26934
rect 28560 26862 28636 27070
rect 110165 27070 110166 27102
rect 110230 27102 110236 27134
rect 110296 27134 110372 27140
rect 110230 27070 110231 27102
rect 110165 27069 110231 27070
rect 110296 27070 110302 27134
rect 110366 27070 110372 27134
rect 28560 26798 28566 26862
rect 28630 26798 28636 26862
rect 110296 26862 110372 27070
rect 116552 26998 116628 27206
rect 119272 27206 119278 27238
rect 119342 27238 119343 27270
rect 120088 27270 120164 27276
rect 119342 27206 119348 27238
rect 116552 26966 116558 26998
rect 116557 26934 116558 26966
rect 116622 26966 116628 26998
rect 116824 26998 116900 27004
rect 116622 26934 116623 26966
rect 116557 26933 116623 26934
rect 116824 26934 116830 26998
rect 116894 26934 116900 26998
rect 110296 26830 110302 26862
rect 28560 26792 28636 26798
rect 110301 26798 110302 26830
rect 110366 26830 110372 26862
rect 110366 26798 110367 26830
rect 110301 26797 110367 26798
rect 19926 26662 19927 26694
rect 19861 26661 19927 26662
rect 21896 26662 21902 26726
rect 21966 26662 21972 26726
rect 28293 26726 28359 26727
rect 28293 26694 28294 26726
rect 21896 26656 21972 26662
rect 28288 26662 28294 26694
rect 28358 26694 28359 26726
rect 110301 26726 110367 26727
rect 110301 26694 110302 26726
rect 28358 26662 28364 26694
rect 21760 26590 21836 26596
rect 21760 26526 21766 26590
rect 21830 26526 21836 26590
rect 18496 26422 18502 26454
rect 18501 26390 18502 26422
rect 18566 26422 18572 26454
rect 19453 26454 19519 26455
rect 19453 26422 19454 26454
rect 18566 26390 18567 26422
rect 18501 26389 18567 26390
rect 19448 26390 19454 26422
rect 19518 26422 19519 26454
rect 19725 26454 19791 26455
rect 19725 26422 19726 26454
rect 19518 26390 19524 26422
rect 952 25574 1230 25638
rect 1294 25574 1300 25638
rect 952 24006 1300 25574
rect 3808 25910 3884 25916
rect 3808 25846 3814 25910
rect 3878 25846 3884 25910
rect 2540 25365 2606 25366
rect 2540 25301 2541 25365
rect 2605 25301 2606 25365
rect 2540 25300 2606 25301
rect 952 23942 1230 24006
rect 1294 23942 1300 24006
rect 2312 24550 2388 24556
rect 2312 24486 2318 24550
rect 2382 24486 2388 24550
rect 2312 24006 2388 24486
rect 2312 23974 2318 24006
rect 952 22374 1300 23942
rect 2317 23942 2318 23974
rect 2382 23974 2388 24006
rect 2382 23942 2383 23974
rect 2317 23941 2383 23942
rect 952 22310 1230 22374
rect 1294 22310 1300 22374
rect 952 20470 1300 22310
rect 952 20406 1230 20470
rect 1294 20406 1300 20470
rect 952 18974 1300 20406
rect 952 18910 1230 18974
rect 1294 18910 1300 18974
rect 952 17070 1300 18910
rect 2543 17959 2603 25300
rect 3808 23326 3884 25846
rect 19448 25094 19524 26390
rect 19720 26390 19726 26422
rect 19790 26422 19791 26454
rect 19790 26390 19796 26422
rect 19448 25030 19454 25094
rect 19518 25030 19524 25094
rect 19584 25366 19660 25372
rect 19584 25302 19590 25366
rect 19654 25302 19660 25366
rect 19584 25094 19660 25302
rect 19584 25062 19590 25094
rect 19448 25024 19524 25030
rect 19589 25030 19590 25062
rect 19654 25062 19660 25094
rect 19720 25094 19796 26390
rect 21760 26318 21836 26526
rect 21760 26286 21766 26318
rect 21765 26254 21766 26286
rect 21830 26286 21836 26318
rect 22712 26590 22788 26596
rect 22712 26526 22718 26590
rect 22782 26526 22788 26590
rect 22712 26318 22788 26526
rect 28288 26454 28364 26662
rect 28288 26390 28294 26454
rect 28358 26390 28364 26454
rect 28288 26384 28364 26390
rect 110296 26662 110302 26694
rect 110366 26694 110367 26726
rect 116824 26726 116900 26934
rect 116824 26694 116830 26726
rect 110366 26662 110372 26694
rect 110296 26454 110372 26662
rect 116829 26662 116830 26694
rect 116894 26694 116900 26726
rect 119272 26726 119348 27206
rect 116894 26662 116895 26694
rect 116829 26661 116895 26662
rect 119272 26662 119278 26726
rect 119342 26662 119348 26726
rect 120088 27206 120094 27270
rect 120158 27206 120164 27270
rect 120088 26726 120164 27206
rect 120088 26694 120094 26726
rect 119272 26656 119348 26662
rect 120093 26662 120094 26694
rect 120158 26694 120164 26726
rect 120496 27270 120572 27276
rect 120496 27206 120502 27270
rect 120566 27206 120572 27270
rect 120496 26726 120572 27206
rect 120496 26694 120502 26726
rect 120158 26662 120159 26694
rect 120093 26661 120159 26662
rect 120501 26662 120502 26694
rect 120566 26694 120572 26726
rect 137496 27270 137844 28974
rect 137496 27206 137502 27270
rect 137566 27206 137844 27270
rect 120566 26662 120567 26694
rect 120501 26661 120567 26662
rect 116013 26590 116079 26591
rect 116013 26558 116014 26590
rect 110296 26390 110302 26454
rect 110366 26390 110372 26454
rect 110296 26384 110372 26390
rect 116008 26526 116014 26558
rect 116078 26558 116079 26590
rect 116829 26590 116895 26591
rect 116829 26558 116830 26590
rect 116078 26526 116084 26558
rect 22712 26286 22718 26318
rect 21830 26254 21831 26286
rect 21765 26253 21831 26254
rect 22717 26254 22718 26286
rect 22782 26286 22788 26318
rect 110432 26318 110508 26324
rect 22782 26254 22783 26286
rect 22717 26253 22783 26254
rect 110432 26254 110438 26318
rect 110502 26254 110508 26318
rect 21896 26182 21972 26188
rect 21896 26118 21902 26182
rect 21966 26118 21972 26182
rect 22989 26182 23055 26183
rect 22989 26150 22990 26182
rect 21896 25910 21972 26118
rect 22984 26118 22990 26150
rect 23054 26150 23055 26182
rect 23392 26182 23468 26188
rect 23054 26118 23060 26150
rect 22445 26046 22511 26047
rect 22445 26014 22446 26046
rect 21896 25878 21902 25910
rect 21901 25846 21902 25878
rect 21966 25878 21972 25910
rect 22440 25982 22446 26014
rect 22510 26014 22511 26046
rect 22510 25982 22516 26014
rect 22440 25916 22516 25982
rect 22440 25910 22652 25916
rect 21966 25846 21967 25878
rect 21901 25845 21967 25846
rect 22440 25846 22582 25910
rect 22646 25846 22652 25910
rect 22440 25840 22652 25846
rect 22984 25910 23060 26118
rect 22984 25846 22990 25910
rect 23054 25846 23060 25910
rect 23392 26118 23398 26182
rect 23462 26118 23468 26182
rect 23392 25910 23468 26118
rect 110432 26046 110508 26254
rect 116008 26318 116084 26526
rect 116008 26254 116014 26318
rect 116078 26254 116084 26318
rect 116008 26248 116084 26254
rect 116824 26526 116830 26558
rect 116894 26558 116895 26590
rect 119816 26590 119892 26596
rect 116894 26526 116900 26558
rect 116824 26318 116900 26526
rect 119816 26526 119822 26590
rect 119886 26526 119892 26590
rect 116824 26254 116830 26318
rect 116894 26254 116900 26318
rect 116824 26248 116900 26254
rect 119408 26454 119484 26460
rect 119408 26390 119414 26454
rect 119478 26390 119484 26454
rect 115197 26182 115263 26183
rect 115197 26150 115198 26182
rect 110432 26014 110438 26046
rect 110437 25982 110438 26014
rect 110502 26014 110508 26046
rect 115192 26118 115198 26150
rect 115262 26150 115263 26182
rect 115600 26182 115676 26188
rect 115262 26118 115268 26150
rect 110502 25982 110503 26014
rect 110437 25981 110503 25982
rect 23392 25878 23398 25910
rect 22984 25840 23060 25846
rect 23397 25846 23398 25878
rect 23462 25878 23468 25910
rect 28565 25910 28631 25911
rect 28565 25878 28566 25910
rect 23462 25846 23463 25878
rect 23397 25845 23463 25846
rect 28560 25846 28566 25878
rect 28630 25878 28631 25910
rect 115192 25910 115268 26118
rect 28630 25846 28636 25878
rect 21901 25774 21967 25775
rect 21901 25742 21902 25774
rect 21896 25710 21902 25742
rect 21966 25742 21967 25774
rect 22445 25774 22511 25775
rect 22445 25742 22446 25774
rect 21966 25710 21972 25742
rect 21896 25502 21972 25710
rect 21896 25438 21902 25502
rect 21966 25438 21972 25502
rect 21896 25432 21972 25438
rect 22440 25710 22446 25742
rect 22510 25742 22511 25774
rect 23120 25774 23196 25780
rect 22510 25710 22516 25742
rect 22440 25502 22516 25710
rect 22440 25438 22446 25502
rect 22510 25438 22516 25502
rect 23120 25710 23126 25774
rect 23190 25710 23196 25774
rect 23120 25502 23196 25710
rect 23120 25470 23126 25502
rect 22440 25432 22516 25438
rect 23125 25438 23126 25470
rect 23190 25470 23196 25502
rect 23528 25774 23604 25780
rect 23528 25710 23534 25774
rect 23598 25710 23604 25774
rect 23528 25502 23604 25710
rect 23528 25470 23534 25502
rect 23190 25438 23191 25470
rect 23125 25437 23191 25438
rect 23533 25438 23534 25470
rect 23598 25470 23604 25502
rect 28560 25502 28636 25846
rect 115192 25846 115198 25910
rect 115262 25846 115268 25910
rect 115600 26118 115606 26182
rect 115670 26118 115676 26182
rect 116965 26182 117031 26183
rect 116965 26150 116966 26182
rect 115600 25910 115676 26118
rect 115600 25878 115606 25910
rect 115192 25840 115268 25846
rect 115605 25846 115606 25878
rect 115670 25878 115676 25910
rect 116960 26118 116966 26150
rect 117030 26150 117031 26182
rect 117030 26118 117036 26150
rect 116960 25910 117036 26118
rect 115670 25846 115671 25878
rect 115605 25845 115671 25846
rect 116960 25846 116966 25910
rect 117030 25846 117036 25910
rect 116960 25840 117036 25846
rect 23598 25438 23599 25470
rect 23533 25437 23599 25438
rect 28560 25438 28566 25502
rect 28630 25438 28636 25502
rect 115328 25774 115404 25780
rect 115328 25710 115334 25774
rect 115398 25710 115404 25774
rect 115328 25502 115404 25710
rect 115328 25470 115334 25502
rect 28560 25432 28636 25438
rect 115333 25438 115334 25470
rect 115398 25470 115404 25502
rect 115736 25774 115812 25780
rect 115736 25710 115742 25774
rect 115806 25710 115812 25774
rect 115736 25502 115812 25710
rect 115736 25470 115742 25502
rect 115398 25438 115399 25470
rect 115333 25437 115399 25438
rect 115741 25438 115742 25470
rect 115806 25470 115812 25502
rect 116280 25774 116356 25780
rect 116280 25710 116286 25774
rect 116350 25710 116356 25774
rect 116280 25502 116356 25710
rect 116280 25470 116286 25502
rect 115806 25438 115807 25470
rect 115741 25437 115807 25438
rect 116285 25438 116286 25470
rect 116350 25470 116356 25502
rect 116416 25774 116492 25780
rect 116416 25710 116422 25774
rect 116486 25710 116492 25774
rect 116965 25774 117031 25775
rect 116965 25742 116966 25774
rect 116416 25502 116492 25710
rect 116416 25470 116422 25502
rect 116350 25438 116351 25470
rect 116285 25437 116351 25438
rect 116421 25438 116422 25470
rect 116486 25470 116492 25502
rect 116960 25710 116966 25742
rect 117030 25742 117031 25774
rect 119277 25774 119343 25775
rect 119277 25742 119278 25774
rect 117030 25710 117036 25742
rect 116960 25502 117036 25710
rect 116486 25438 116487 25470
rect 116421 25437 116487 25438
rect 116960 25438 116966 25502
rect 117030 25438 117036 25502
rect 116960 25432 117036 25438
rect 119272 25710 119278 25742
rect 119342 25742 119343 25774
rect 119342 25710 119348 25742
rect 21765 25366 21831 25367
rect 21765 25334 21766 25366
rect 19654 25030 19655 25062
rect 19589 25029 19655 25030
rect 19720 25030 19726 25094
rect 19790 25030 19796 25094
rect 19720 25024 19796 25030
rect 21760 25302 21766 25334
rect 21830 25334 21831 25366
rect 22173 25366 22239 25367
rect 22173 25334 22174 25366
rect 21830 25302 21836 25334
rect 21760 25094 21836 25302
rect 21760 25030 21766 25094
rect 21830 25030 21836 25094
rect 21760 25024 21836 25030
rect 22168 25302 22174 25334
rect 22238 25334 22239 25366
rect 22712 25366 22788 25372
rect 22238 25302 22244 25334
rect 22168 25094 22244 25302
rect 22168 25030 22174 25094
rect 22238 25030 22244 25094
rect 22712 25302 22718 25366
rect 22782 25302 22788 25366
rect 22989 25366 23055 25367
rect 22989 25334 22990 25366
rect 22712 25094 22788 25302
rect 22712 25062 22718 25094
rect 22168 25024 22244 25030
rect 22717 25030 22718 25062
rect 22782 25062 22788 25094
rect 22984 25302 22990 25334
rect 23054 25334 23055 25366
rect 23533 25366 23599 25367
rect 23533 25334 23534 25366
rect 23054 25302 23060 25334
rect 22984 25094 23060 25302
rect 22782 25030 22783 25062
rect 22717 25029 22783 25030
rect 22984 25030 22990 25094
rect 23054 25030 23060 25094
rect 22984 25024 23060 25030
rect 23528 25302 23534 25334
rect 23598 25334 23599 25366
rect 115192 25366 115268 25372
rect 23598 25302 23604 25334
rect 23528 25094 23604 25302
rect 23528 25030 23534 25094
rect 23598 25030 23604 25094
rect 115192 25302 115198 25366
rect 115262 25302 115268 25366
rect 115741 25366 115807 25367
rect 115741 25334 115742 25366
rect 115192 25094 115268 25302
rect 115192 25062 115198 25094
rect 23528 25024 23604 25030
rect 115197 25030 115198 25062
rect 115262 25062 115268 25094
rect 115736 25302 115742 25334
rect 115806 25334 115807 25366
rect 116552 25366 116628 25372
rect 115806 25302 115812 25334
rect 115736 25094 115812 25302
rect 115262 25030 115263 25062
rect 115197 25029 115263 25030
rect 115736 25030 115742 25094
rect 115806 25030 115812 25094
rect 116552 25302 116558 25366
rect 116622 25302 116628 25366
rect 116552 25094 116628 25302
rect 116552 25062 116558 25094
rect 115736 25024 115812 25030
rect 116557 25030 116558 25062
rect 116622 25062 116628 25094
rect 116960 25366 117036 25372
rect 116960 25302 116966 25366
rect 117030 25302 117036 25366
rect 116960 25094 117036 25302
rect 116960 25062 116966 25094
rect 116622 25030 116623 25062
rect 116557 25029 116623 25030
rect 116965 25030 116966 25062
rect 117030 25062 117036 25094
rect 119272 25094 119348 25710
rect 117030 25030 117031 25062
rect 116965 25029 117031 25030
rect 119272 25030 119278 25094
rect 119342 25030 119348 25094
rect 119408 25094 119484 26390
rect 119408 25062 119414 25094
rect 119272 25024 119348 25030
rect 119413 25030 119414 25062
rect 119478 25062 119484 25094
rect 119816 25094 119892 26526
rect 119816 25062 119822 25094
rect 119478 25030 119479 25062
rect 119413 25029 119479 25030
rect 119821 25030 119822 25062
rect 119886 25062 119892 25094
rect 137496 25638 137844 27206
rect 137496 25574 137502 25638
rect 137566 25574 137844 25638
rect 119886 25030 119887 25062
rect 119821 25029 119887 25030
rect 18224 24958 18300 24964
rect 18224 24894 18230 24958
rect 18294 24894 18300 24958
rect 18224 24278 18300 24894
rect 18224 24246 18230 24278
rect 18229 24214 18230 24246
rect 18294 24246 18300 24278
rect 18904 24958 18980 24964
rect 18904 24894 18910 24958
rect 18974 24894 18980 24958
rect 18904 24278 18980 24894
rect 18904 24246 18910 24278
rect 18294 24214 18295 24246
rect 18229 24213 18295 24214
rect 18909 24214 18910 24246
rect 18974 24246 18980 24278
rect 19312 24958 19388 24964
rect 19312 24894 19318 24958
rect 19382 24894 19388 24958
rect 19312 24278 19388 24894
rect 21896 24958 21972 24964
rect 21896 24894 21902 24958
rect 21966 24894 21972 24958
rect 21896 24686 21972 24894
rect 21896 24654 21902 24686
rect 21901 24622 21902 24654
rect 21966 24654 21972 24686
rect 22168 24958 22244 24964
rect 22168 24894 22174 24958
rect 22238 24894 22244 24958
rect 22168 24686 22244 24894
rect 22168 24654 22174 24686
rect 21966 24622 21967 24654
rect 21901 24621 21967 24622
rect 22173 24622 22174 24654
rect 22238 24654 22244 24686
rect 23120 24958 23196 24964
rect 23120 24894 23126 24958
rect 23190 24894 23196 24958
rect 23397 24958 23463 24959
rect 23397 24926 23398 24958
rect 23120 24686 23196 24894
rect 23120 24654 23126 24686
rect 22238 24622 22239 24654
rect 22173 24621 22239 24622
rect 23125 24622 23126 24654
rect 23190 24654 23196 24686
rect 23392 24894 23398 24926
rect 23462 24926 23463 24958
rect 115197 24958 115263 24959
rect 115197 24926 115198 24958
rect 23462 24894 23468 24926
rect 23392 24686 23468 24894
rect 23190 24622 23191 24654
rect 23125 24621 23191 24622
rect 23392 24622 23398 24686
rect 23462 24622 23468 24686
rect 23392 24616 23468 24622
rect 115192 24894 115198 24926
rect 115262 24926 115263 24958
rect 115600 24958 115676 24964
rect 115262 24894 115268 24926
rect 115192 24686 115268 24894
rect 115192 24622 115198 24686
rect 115262 24622 115268 24686
rect 115600 24894 115606 24958
rect 115670 24894 115676 24958
rect 115600 24686 115676 24894
rect 115600 24654 115606 24686
rect 115192 24616 115268 24622
rect 115605 24622 115606 24654
rect 115670 24654 115676 24686
rect 116144 24958 116220 24964
rect 116144 24894 116150 24958
rect 116214 24894 116220 24958
rect 116965 24958 117031 24959
rect 116965 24926 116966 24958
rect 116144 24686 116220 24894
rect 116144 24654 116150 24686
rect 115670 24622 115671 24654
rect 115605 24621 115671 24622
rect 116149 24622 116150 24654
rect 116214 24654 116220 24686
rect 116960 24894 116966 24926
rect 117030 24926 117031 24958
rect 119000 24958 119076 24964
rect 117030 24894 117036 24926
rect 116960 24686 117036 24894
rect 116214 24622 116215 24654
rect 116149 24621 116215 24622
rect 116960 24622 116966 24686
rect 117030 24622 117036 24686
rect 116960 24616 117036 24622
rect 119000 24894 119006 24958
rect 119070 24894 119076 24958
rect 19312 24246 19318 24278
rect 18974 24214 18975 24246
rect 18909 24213 18975 24214
rect 19317 24214 19318 24246
rect 19382 24246 19388 24278
rect 21760 24550 21836 24556
rect 21760 24486 21766 24550
rect 21830 24486 21836 24550
rect 22309 24550 22375 24551
rect 22309 24518 22310 24550
rect 21760 24278 21836 24486
rect 21760 24246 21766 24278
rect 19382 24214 19383 24246
rect 19317 24213 19383 24214
rect 21765 24214 21766 24246
rect 21830 24246 21836 24278
rect 22304 24486 22310 24518
rect 22374 24518 22375 24550
rect 23120 24550 23196 24556
rect 22374 24486 22380 24518
rect 22304 24278 22380 24486
rect 21830 24214 21831 24246
rect 21765 24213 21831 24214
rect 22304 24214 22310 24278
rect 22374 24214 22380 24278
rect 23120 24486 23126 24550
rect 23190 24486 23196 24550
rect 23533 24550 23599 24551
rect 23533 24518 23534 24550
rect 23120 24278 23196 24486
rect 23120 24246 23126 24278
rect 22304 24208 22380 24214
rect 23125 24214 23126 24246
rect 23190 24246 23196 24278
rect 23528 24486 23534 24518
rect 23598 24518 23599 24550
rect 115197 24550 115263 24551
rect 115197 24518 115198 24550
rect 23598 24486 23604 24518
rect 23528 24278 23604 24486
rect 23190 24214 23191 24246
rect 23125 24213 23191 24214
rect 23528 24214 23534 24278
rect 23598 24214 23604 24278
rect 23528 24208 23604 24214
rect 115192 24486 115198 24518
rect 115262 24518 115263 24550
rect 115741 24550 115807 24551
rect 115741 24518 115742 24550
rect 115262 24486 115268 24518
rect 115192 24278 115268 24486
rect 115192 24214 115198 24278
rect 115262 24214 115268 24278
rect 115192 24208 115268 24214
rect 115736 24486 115742 24518
rect 115806 24518 115807 24550
rect 116013 24550 116079 24551
rect 116013 24518 116014 24550
rect 115806 24486 115812 24518
rect 115736 24278 115812 24486
rect 115736 24214 115742 24278
rect 115806 24214 115812 24278
rect 115736 24208 115812 24214
rect 116008 24486 116014 24518
rect 116078 24518 116079 24550
rect 116824 24550 116900 24556
rect 116078 24486 116084 24518
rect 116008 24278 116084 24486
rect 116008 24214 116014 24278
rect 116078 24214 116084 24278
rect 116824 24486 116830 24550
rect 116894 24486 116900 24550
rect 116824 24278 116900 24486
rect 116824 24246 116830 24278
rect 116008 24208 116084 24214
rect 116829 24214 116830 24246
rect 116894 24246 116900 24278
rect 119000 24278 119076 24894
rect 119000 24246 119006 24278
rect 116894 24214 116895 24246
rect 116829 24213 116895 24214
rect 119005 24214 119006 24246
rect 119070 24246 119076 24278
rect 119408 24958 119484 24964
rect 119408 24894 119414 24958
rect 119478 24894 119484 24958
rect 119408 24278 119484 24894
rect 119408 24246 119414 24278
rect 119070 24214 119071 24246
rect 119005 24213 119071 24214
rect 119413 24214 119414 24246
rect 119478 24246 119484 24278
rect 120088 24958 120164 24964
rect 120088 24894 120094 24958
rect 120158 24894 120164 24958
rect 120637 24958 120703 24959
rect 120637 24926 120638 24958
rect 120088 24278 120164 24894
rect 120088 24246 120094 24278
rect 119478 24214 119479 24246
rect 119413 24213 119479 24214
rect 120093 24214 120094 24246
rect 120158 24246 120164 24278
rect 120632 24894 120638 24926
rect 120702 24926 120703 24958
rect 120702 24894 120708 24926
rect 120632 24278 120708 24894
rect 120158 24214 120159 24246
rect 120093 24213 120159 24214
rect 120632 24214 120638 24278
rect 120702 24214 120708 24278
rect 120632 24208 120708 24214
rect 18224 24142 18300 24148
rect 18224 24078 18230 24142
rect 18294 24078 18300 24142
rect 18501 24142 18567 24143
rect 18501 24110 18502 24142
rect 18224 23598 18300 24078
rect 18224 23566 18230 23598
rect 18229 23534 18230 23566
rect 18294 23566 18300 23598
rect 18496 24078 18502 24110
rect 18566 24110 18567 24142
rect 19317 24142 19383 24143
rect 19317 24110 19318 24142
rect 18566 24078 18572 24110
rect 18496 23598 18572 24078
rect 18294 23534 18295 23566
rect 18229 23533 18295 23534
rect 18496 23534 18502 23598
rect 18566 23534 18572 23598
rect 18496 23528 18572 23534
rect 19312 24078 19318 24110
rect 19382 24110 19383 24142
rect 19861 24142 19927 24143
rect 19861 24110 19862 24142
rect 19382 24078 19388 24110
rect 19312 23462 19388 24078
rect 19312 23398 19318 23462
rect 19382 23398 19388 23462
rect 19312 23392 19388 23398
rect 19856 24078 19862 24110
rect 19926 24110 19927 24142
rect 22304 24142 22380 24148
rect 19926 24078 19932 24110
rect 19856 23462 19932 24078
rect 22304 24078 22310 24142
rect 22374 24078 22380 24142
rect 22581 24142 22647 24143
rect 22581 24110 22582 24142
rect 22304 23870 22380 24078
rect 22304 23838 22310 23870
rect 22309 23806 22310 23838
rect 22374 23838 22380 23870
rect 22576 24078 22582 24110
rect 22646 24110 22647 24142
rect 22984 24142 23060 24148
rect 22646 24078 22652 24110
rect 22576 23870 22652 24078
rect 22374 23806 22375 23838
rect 22309 23805 22375 23806
rect 22576 23806 22582 23870
rect 22646 23806 22652 23870
rect 22984 24078 22990 24142
rect 23054 24078 23060 24142
rect 22984 23870 23060 24078
rect 22984 23838 22990 23870
rect 22576 23800 22652 23806
rect 22989 23806 22990 23838
rect 23054 23838 23060 23870
rect 23392 24142 23468 24148
rect 23392 24078 23398 24142
rect 23462 24078 23468 24142
rect 115333 24142 115399 24143
rect 115333 24110 115334 24142
rect 23392 23870 23468 24078
rect 115328 24078 115334 24110
rect 115398 24110 115399 24142
rect 115741 24142 115807 24143
rect 115741 24110 115742 24142
rect 115398 24078 115404 24110
rect 23392 23838 23398 23870
rect 23054 23806 23055 23838
rect 22989 23805 23055 23806
rect 23397 23806 23398 23838
rect 23462 23838 23468 23870
rect 28424 24006 28500 24012
rect 28424 23942 28430 24006
rect 28494 23942 28500 24006
rect 110437 24006 110503 24007
rect 110437 23974 110438 24006
rect 23462 23806 23463 23838
rect 23397 23805 23463 23806
rect 22989 23734 23055 23735
rect 22989 23702 22990 23734
rect 19856 23398 19862 23462
rect 19926 23398 19932 23462
rect 19856 23392 19932 23398
rect 22984 23670 22990 23702
rect 23054 23702 23055 23734
rect 23397 23734 23463 23735
rect 23397 23702 23398 23734
rect 23054 23670 23060 23702
rect 22984 23462 23060 23670
rect 22984 23398 22990 23462
rect 23054 23398 23060 23462
rect 22984 23392 23060 23398
rect 23392 23670 23398 23702
rect 23462 23702 23463 23734
rect 28424 23734 28500 23942
rect 28424 23702 28430 23734
rect 23462 23670 23468 23702
rect 23392 23462 23468 23670
rect 28429 23670 28430 23702
rect 28494 23702 28500 23734
rect 110432 23942 110438 23974
rect 110502 23974 110503 24006
rect 110502 23942 110508 23974
rect 110432 23734 110508 23942
rect 115328 23870 115404 24078
rect 115328 23806 115334 23870
rect 115398 23806 115404 23870
rect 115328 23800 115404 23806
rect 115736 24078 115742 24110
rect 115806 24110 115807 24142
rect 116149 24142 116215 24143
rect 116149 24110 116150 24142
rect 115806 24078 115812 24110
rect 115736 23870 115812 24078
rect 115736 23806 115742 23870
rect 115806 23806 115812 23870
rect 115736 23800 115812 23806
rect 116144 24078 116150 24110
rect 116214 24110 116215 24142
rect 116552 24142 116628 24148
rect 116214 24078 116220 24110
rect 116144 23870 116220 24078
rect 116144 23806 116150 23870
rect 116214 23806 116220 23870
rect 116552 24078 116558 24142
rect 116622 24078 116628 24142
rect 116552 23870 116628 24078
rect 116552 23838 116558 23870
rect 116144 23800 116220 23806
rect 116557 23806 116558 23838
rect 116622 23838 116628 23870
rect 119000 24142 119076 24148
rect 119000 24078 119006 24142
rect 119070 24078 119076 24142
rect 116622 23806 116623 23838
rect 116557 23805 116623 23806
rect 28494 23670 28495 23702
rect 28429 23669 28495 23670
rect 110432 23670 110438 23734
rect 110502 23670 110508 23734
rect 110432 23664 110508 23670
rect 115328 23734 115404 23740
rect 115328 23670 115334 23734
rect 115398 23670 115404 23734
rect 23392 23398 23398 23462
rect 23462 23398 23468 23462
rect 115328 23462 115404 23670
rect 115328 23430 115334 23462
rect 23392 23392 23468 23398
rect 115333 23398 115334 23430
rect 115398 23430 115404 23462
rect 115736 23734 115812 23740
rect 115736 23670 115742 23734
rect 115806 23670 115812 23734
rect 115736 23462 115812 23670
rect 115736 23430 115742 23462
rect 115398 23398 115399 23430
rect 115333 23397 115399 23398
rect 115741 23398 115742 23430
rect 115806 23430 115812 23462
rect 119000 23462 119076 24078
rect 119000 23430 119006 23462
rect 115806 23398 115807 23430
rect 115741 23397 115807 23398
rect 119005 23398 119006 23430
rect 119070 23430 119076 23462
rect 119272 24142 119348 24148
rect 119272 24078 119278 24142
rect 119342 24078 119348 24142
rect 119685 24142 119751 24143
rect 119685 24110 119686 24142
rect 119272 23462 119348 24078
rect 119680 24078 119686 24110
rect 119750 24110 119751 24142
rect 120637 24142 120703 24143
rect 120637 24110 120638 24142
rect 119750 24078 119756 24110
rect 119680 23598 119756 24078
rect 120632 24078 120638 24110
rect 120702 24110 120703 24142
rect 120702 24078 120708 24110
rect 120501 24006 120567 24007
rect 120501 23974 120502 24006
rect 119680 23534 119686 23598
rect 119750 23534 119756 23598
rect 119680 23528 119756 23534
rect 120496 23942 120502 23974
rect 120566 23974 120567 24006
rect 120566 23942 120572 23974
rect 120496 23598 120572 23942
rect 120496 23534 120502 23598
rect 120566 23534 120572 23598
rect 120496 23528 120572 23534
rect 120632 23598 120708 24078
rect 120632 23534 120638 23598
rect 120702 23534 120708 23598
rect 120632 23528 120708 23534
rect 137496 24006 137844 25574
rect 137496 23942 137502 24006
rect 137566 23942 137844 24006
rect 119272 23430 119278 23462
rect 119070 23398 119071 23430
rect 119005 23397 119071 23398
rect 119277 23398 119278 23430
rect 119342 23430 119348 23462
rect 119342 23398 119343 23430
rect 119277 23397 119343 23398
rect 3808 23294 3814 23326
rect 3813 23262 3814 23294
rect 3878 23294 3884 23326
rect 18229 23326 18295 23327
rect 18229 23294 18230 23326
rect 3878 23262 3879 23294
rect 3813 23261 3879 23262
rect 18224 23262 18230 23294
rect 18294 23294 18295 23326
rect 18632 23326 18708 23332
rect 18294 23262 18300 23294
rect 18224 22782 18300 23262
rect 18632 23262 18638 23326
rect 18702 23262 18708 23326
rect 19317 23326 19383 23327
rect 19317 23294 19318 23326
rect 18224 22718 18230 22782
rect 18294 22718 18300 22782
rect 18360 23190 18436 23196
rect 18360 23126 18366 23190
rect 18430 23126 18436 23190
rect 18360 22782 18436 23126
rect 18360 22750 18366 22782
rect 18224 22712 18300 22718
rect 18365 22718 18366 22750
rect 18430 22750 18436 22782
rect 18632 22782 18708 23262
rect 18632 22750 18638 22782
rect 18430 22718 18431 22750
rect 18365 22717 18431 22718
rect 18637 22718 18638 22750
rect 18702 22750 18708 22782
rect 19312 23262 19318 23294
rect 19382 23294 19383 23326
rect 19725 23326 19791 23327
rect 19725 23294 19726 23326
rect 19382 23262 19388 23294
rect 19312 22782 19388 23262
rect 18702 22718 18703 22750
rect 18637 22717 18703 22718
rect 19312 22718 19318 22782
rect 19382 22718 19388 22782
rect 19312 22712 19388 22718
rect 19720 23262 19726 23294
rect 19790 23294 19791 23326
rect 22173 23326 22239 23327
rect 22173 23294 22174 23326
rect 19790 23262 19796 23294
rect 19720 22782 19796 23262
rect 22168 23262 22174 23294
rect 22238 23294 22239 23326
rect 22576 23326 22652 23332
rect 22238 23262 22244 23294
rect 21765 23054 21831 23055
rect 21765 23022 21766 23054
rect 19720 22718 19726 22782
rect 19790 22718 19796 22782
rect 19720 22712 19796 22718
rect 21760 22990 21766 23022
rect 21830 23022 21831 23054
rect 22168 23054 22244 23262
rect 21830 22990 21836 23022
rect 21760 22782 21836 22990
rect 22168 22990 22174 23054
rect 22238 22990 22244 23054
rect 22576 23262 22582 23326
rect 22646 23262 22652 23326
rect 22576 23054 22652 23262
rect 22576 23022 22582 23054
rect 22168 22984 22244 22990
rect 22581 22990 22582 23022
rect 22646 23022 22652 23054
rect 23120 23326 23196 23332
rect 23120 23262 23126 23326
rect 23190 23262 23196 23326
rect 23120 23054 23196 23262
rect 23120 23022 23126 23054
rect 22646 22990 22647 23022
rect 22581 22989 22647 22990
rect 23125 22990 23126 23022
rect 23190 23022 23196 23054
rect 23528 23326 23604 23332
rect 23528 23262 23534 23326
rect 23598 23262 23604 23326
rect 23528 23054 23604 23262
rect 115328 23326 115404 23332
rect 115328 23262 115334 23326
rect 115398 23262 115404 23326
rect 23528 23022 23534 23054
rect 23190 22990 23191 23022
rect 23125 22989 23191 22990
rect 23533 22990 23534 23022
rect 23598 23022 23604 23054
rect 110432 23190 110508 23196
rect 110432 23126 110438 23190
rect 110502 23126 110508 23190
rect 23598 22990 23599 23022
rect 23533 22989 23599 22990
rect 110432 22918 110508 23126
rect 115328 23054 115404 23262
rect 115328 23022 115334 23054
rect 115333 22990 115334 23022
rect 115398 23022 115404 23054
rect 115736 23326 115812 23332
rect 115736 23262 115742 23326
rect 115806 23262 115812 23326
rect 115736 23054 115812 23262
rect 115736 23022 115742 23054
rect 115398 22990 115399 23022
rect 115333 22989 115399 22990
rect 115741 22990 115742 23022
rect 115806 23022 115812 23054
rect 116280 23326 116356 23332
rect 116280 23262 116286 23326
rect 116350 23262 116356 23326
rect 119005 23326 119071 23327
rect 119005 23294 119006 23326
rect 116280 23054 116356 23262
rect 119000 23262 119006 23294
rect 119070 23294 119071 23326
rect 119277 23326 119343 23327
rect 119277 23294 119278 23326
rect 119070 23262 119076 23294
rect 116280 23022 116286 23054
rect 115806 22990 115807 23022
rect 115741 22989 115807 22990
rect 116285 22990 116286 23022
rect 116350 23022 116356 23054
rect 116829 23054 116895 23055
rect 116829 23022 116830 23054
rect 116350 22990 116351 23022
rect 116285 22989 116351 22990
rect 116824 22990 116830 23022
rect 116894 23022 116895 23054
rect 116894 22990 116900 23022
rect 110432 22886 110438 22918
rect 110437 22854 110438 22886
rect 110502 22886 110508 22918
rect 110502 22854 110503 22886
rect 110437 22853 110503 22854
rect 21760 22718 21766 22782
rect 21830 22718 21836 22782
rect 21760 22712 21836 22718
rect 28560 22782 28636 22788
rect 28560 22718 28566 22782
rect 28630 22718 28636 22782
rect 110165 22782 110231 22783
rect 110165 22750 110166 22782
rect 21760 22646 21836 22652
rect 21760 22582 21766 22646
rect 21830 22582 21836 22646
rect 22445 22646 22511 22647
rect 22445 22614 22446 22646
rect 18632 22510 18708 22516
rect 18632 22446 18638 22510
rect 18702 22446 18708 22510
rect 19861 22510 19927 22511
rect 19861 22478 19862 22510
rect 3133 22238 3199 22239
rect 3133 22206 3134 22238
rect 3128 22174 3134 22206
rect 3198 22206 3199 22238
rect 3198 22174 3204 22206
rect 3128 21830 3204 22174
rect 3128 21766 3134 21830
rect 3198 21766 3204 21830
rect 3128 21760 3204 21766
rect 18632 21150 18708 22446
rect 18632 21118 18638 21150
rect 18637 21086 18638 21118
rect 18702 21118 18708 21150
rect 19856 22446 19862 22478
rect 19926 22478 19927 22510
rect 19926 22446 19932 22478
rect 19856 21150 19932 22446
rect 21760 22374 21836 22582
rect 21760 22342 21766 22374
rect 21765 22310 21766 22342
rect 21830 22342 21836 22374
rect 22440 22582 22446 22614
rect 22510 22614 22511 22646
rect 22510 22582 22516 22614
rect 22440 22374 22516 22582
rect 21830 22310 21831 22342
rect 21765 22309 21831 22310
rect 22440 22310 22446 22374
rect 22510 22310 22516 22374
rect 28293 22374 28359 22375
rect 28293 22342 28294 22374
rect 22440 22304 22516 22310
rect 28288 22310 28294 22342
rect 28358 22342 28359 22374
rect 28560 22374 28636 22718
rect 110160 22718 110166 22750
rect 110230 22750 110231 22782
rect 116824 22782 116900 22990
rect 110230 22718 110236 22750
rect 110160 22510 110236 22718
rect 116824 22718 116830 22782
rect 116894 22718 116900 22782
rect 116824 22712 116900 22718
rect 119000 22782 119076 23262
rect 119000 22718 119006 22782
rect 119070 22718 119076 22782
rect 119000 22712 119076 22718
rect 119272 23262 119278 23294
rect 119342 23294 119343 23326
rect 119685 23326 119751 23327
rect 119685 23294 119686 23326
rect 119342 23262 119348 23294
rect 119272 22782 119348 23262
rect 119272 22718 119278 22782
rect 119342 22718 119348 22782
rect 119272 22712 119348 22718
rect 119680 23262 119686 23294
rect 119750 23294 119751 23326
rect 120632 23326 120708 23332
rect 119750 23262 119756 23294
rect 119680 22782 119756 23262
rect 119680 22718 119686 22782
rect 119750 22718 119756 22782
rect 120632 23262 120638 23326
rect 120702 23262 120708 23326
rect 120632 22782 120708 23262
rect 120632 22750 120638 22782
rect 119680 22712 119756 22718
rect 120637 22718 120638 22750
rect 120702 22750 120708 22782
rect 120702 22718 120703 22750
rect 120637 22717 120703 22718
rect 116285 22646 116351 22647
rect 116285 22614 116286 22646
rect 110160 22446 110166 22510
rect 110230 22446 110236 22510
rect 110160 22440 110236 22446
rect 116280 22582 116286 22614
rect 116350 22614 116351 22646
rect 116824 22646 116900 22652
rect 116350 22582 116356 22614
rect 28560 22342 28566 22374
rect 28358 22310 28364 22342
rect 21765 22238 21831 22239
rect 21765 22206 21766 22238
rect 21760 22174 21766 22206
rect 21830 22206 21831 22238
rect 21830 22174 21836 22206
rect 21760 21966 21836 22174
rect 28288 22102 28364 22310
rect 28565 22310 28566 22342
rect 28630 22342 28636 22374
rect 116280 22374 116356 22582
rect 28630 22310 28631 22342
rect 28565 22309 28631 22310
rect 116280 22310 116286 22374
rect 116350 22310 116356 22374
rect 116824 22582 116830 22646
rect 116894 22582 116900 22646
rect 116824 22374 116900 22582
rect 120496 22646 120572 22652
rect 120496 22582 120502 22646
rect 120566 22582 120572 22646
rect 119005 22510 119071 22511
rect 119005 22478 119006 22510
rect 116824 22342 116830 22374
rect 116280 22304 116356 22310
rect 116829 22310 116830 22342
rect 116894 22342 116900 22374
rect 119000 22446 119006 22478
rect 119070 22478 119071 22510
rect 119070 22446 119076 22478
rect 116894 22310 116895 22342
rect 116829 22309 116895 22310
rect 116829 22238 116895 22239
rect 116829 22206 116830 22238
rect 116824 22174 116830 22206
rect 116894 22206 116895 22238
rect 116894 22174 116900 22206
rect 28288 22038 28294 22102
rect 28358 22038 28364 22102
rect 28288 22032 28364 22038
rect 28424 22102 28500 22108
rect 28424 22038 28430 22102
rect 28494 22038 28500 22102
rect 21760 21902 21766 21966
rect 21830 21902 21836 21966
rect 21760 21896 21836 21902
rect 21896 21830 21972 21836
rect 21896 21766 21902 21830
rect 21966 21766 21972 21830
rect 21896 21558 21972 21766
rect 21896 21526 21902 21558
rect 21901 21494 21902 21526
rect 21966 21526 21972 21558
rect 22304 21830 22380 21836
rect 22304 21766 22310 21830
rect 22374 21766 22380 21830
rect 22304 21558 22380 21766
rect 22304 21526 22310 21558
rect 21966 21494 21967 21526
rect 21901 21493 21967 21494
rect 22309 21494 22310 21526
rect 22374 21526 22380 21558
rect 23120 21830 23196 21836
rect 23120 21766 23126 21830
rect 23190 21766 23196 21830
rect 23120 21558 23196 21766
rect 23120 21526 23126 21558
rect 22374 21494 22375 21526
rect 22309 21493 22375 21494
rect 23125 21494 23126 21526
rect 23190 21526 23196 21558
rect 23392 21830 23468 21836
rect 23392 21766 23398 21830
rect 23462 21766 23468 21830
rect 28424 21830 28500 22038
rect 116824 21966 116900 22174
rect 116824 21902 116830 21966
rect 116894 21902 116900 21966
rect 116824 21896 116900 21902
rect 28424 21798 28430 21830
rect 23392 21558 23468 21766
rect 28429 21766 28430 21798
rect 28494 21798 28500 21830
rect 115197 21830 115263 21831
rect 115197 21798 115198 21830
rect 28494 21766 28495 21798
rect 28429 21765 28495 21766
rect 115192 21766 115198 21798
rect 115262 21798 115263 21830
rect 115600 21830 115676 21836
rect 115262 21766 115268 21798
rect 23392 21526 23398 21558
rect 23190 21494 23191 21526
rect 23125 21493 23191 21494
rect 23397 21494 23398 21526
rect 23462 21526 23468 21558
rect 115192 21558 115268 21766
rect 23462 21494 23463 21526
rect 23397 21493 23463 21494
rect 115192 21494 115198 21558
rect 115262 21494 115268 21558
rect 115600 21766 115606 21830
rect 115670 21766 115676 21830
rect 115600 21558 115676 21766
rect 115600 21526 115606 21558
rect 115192 21488 115268 21494
rect 115605 21494 115606 21526
rect 115670 21526 115676 21558
rect 116552 21830 116628 21836
rect 116552 21766 116558 21830
rect 116622 21766 116628 21830
rect 116552 21558 116628 21766
rect 116552 21526 116558 21558
rect 115670 21494 115671 21526
rect 115605 21493 115671 21494
rect 116557 21494 116558 21526
rect 116622 21526 116628 21558
rect 116960 21830 117036 21836
rect 116960 21766 116966 21830
rect 117030 21766 117036 21830
rect 116960 21558 117036 21766
rect 116960 21526 116966 21558
rect 116622 21494 116623 21526
rect 116557 21493 116623 21494
rect 116965 21494 116966 21526
rect 117030 21526 117036 21558
rect 117030 21494 117031 21526
rect 116965 21493 117031 21494
rect 21901 21422 21967 21423
rect 21901 21390 21902 21422
rect 18702 21086 18703 21118
rect 18637 21085 18703 21086
rect 19856 21086 19862 21150
rect 19926 21086 19932 21150
rect 19856 21080 19932 21086
rect 21896 21358 21902 21390
rect 21966 21390 21967 21422
rect 22309 21422 22375 21423
rect 22309 21390 22310 21422
rect 21966 21358 21972 21390
rect 21896 21150 21972 21358
rect 21896 21086 21902 21150
rect 21966 21086 21972 21150
rect 21896 21080 21972 21086
rect 22304 21358 22310 21390
rect 22374 21390 22375 21422
rect 22445 21422 22511 21423
rect 22445 21390 22446 21422
rect 22374 21358 22380 21390
rect 22304 21150 22380 21358
rect 22304 21086 22310 21150
rect 22374 21086 22380 21150
rect 22304 21080 22380 21086
rect 22440 21358 22446 21390
rect 22510 21390 22511 21422
rect 22984 21422 23060 21428
rect 22510 21358 22516 21390
rect 22440 21150 22516 21358
rect 22440 21086 22446 21150
rect 22510 21086 22516 21150
rect 22984 21358 22990 21422
rect 23054 21358 23060 21422
rect 23397 21422 23463 21423
rect 23397 21390 23398 21422
rect 22984 21150 23060 21358
rect 22984 21118 22990 21150
rect 22440 21080 22516 21086
rect 22989 21086 22990 21118
rect 23054 21118 23060 21150
rect 23392 21358 23398 21390
rect 23462 21390 23463 21422
rect 115328 21422 115404 21428
rect 23462 21358 23468 21390
rect 23392 21150 23468 21358
rect 23054 21086 23055 21118
rect 22989 21085 23055 21086
rect 23392 21086 23398 21150
rect 23462 21086 23468 21150
rect 115328 21358 115334 21422
rect 115398 21358 115404 21422
rect 115605 21422 115671 21423
rect 115605 21390 115606 21422
rect 115328 21150 115404 21358
rect 115328 21118 115334 21150
rect 23392 21080 23468 21086
rect 115333 21086 115334 21118
rect 115398 21118 115404 21150
rect 115600 21358 115606 21390
rect 115670 21390 115671 21422
rect 116008 21422 116084 21428
rect 115670 21358 115676 21390
rect 115600 21150 115676 21358
rect 115398 21086 115399 21118
rect 115333 21085 115399 21086
rect 115600 21086 115606 21150
rect 115670 21086 115676 21150
rect 116008 21358 116014 21422
rect 116078 21358 116084 21422
rect 116965 21422 117031 21423
rect 116965 21390 116966 21422
rect 116008 21150 116084 21358
rect 116008 21118 116014 21150
rect 115600 21080 115676 21086
rect 116013 21086 116014 21118
rect 116078 21118 116084 21150
rect 116960 21358 116966 21390
rect 117030 21390 117031 21422
rect 117030 21358 117036 21390
rect 116960 21150 117036 21358
rect 116078 21086 116079 21118
rect 116013 21085 116079 21086
rect 116960 21086 116966 21150
rect 117030 21086 117036 21150
rect 116960 21080 117036 21086
rect 119000 21150 119076 22446
rect 119000 21086 119006 21150
rect 119070 21086 119076 21150
rect 120496 21150 120572 22582
rect 120496 21118 120502 21150
rect 119000 21080 119076 21086
rect 120501 21086 120502 21118
rect 120566 21118 120572 21150
rect 137496 22374 137844 23942
rect 137496 22310 137502 22374
rect 137566 22310 137844 22374
rect 120566 21086 120567 21118
rect 120501 21085 120567 21086
rect 18909 21014 18975 21015
rect 18909 20982 18910 21014
rect 18904 20950 18910 20982
rect 18974 20982 18975 21014
rect 19317 21014 19383 21015
rect 19317 20982 19318 21014
rect 18974 20950 18980 20982
rect 3808 20334 4020 20340
rect 3808 20270 3950 20334
rect 4014 20270 4020 20334
rect 3808 20264 4020 20270
rect 18904 20334 18980 20950
rect 18904 20270 18910 20334
rect 18974 20270 18980 20334
rect 18904 20264 18980 20270
rect 19312 20950 19318 20982
rect 19382 20982 19383 21014
rect 19856 21014 19932 21020
rect 19382 20950 19388 20982
rect 19312 20334 19388 20950
rect 19312 20270 19318 20334
rect 19382 20270 19388 20334
rect 19856 20950 19862 21014
rect 19926 20950 19932 21014
rect 21765 21014 21831 21015
rect 21765 20982 21766 21014
rect 19856 20334 19932 20950
rect 21760 20950 21766 20982
rect 21830 20982 21831 21014
rect 22712 21014 22788 21020
rect 21830 20950 21836 20982
rect 21760 20742 21836 20950
rect 21760 20678 21766 20742
rect 21830 20678 21836 20742
rect 22712 20950 22718 21014
rect 22782 20950 22788 21014
rect 22989 21014 23055 21015
rect 22989 20982 22990 21014
rect 22712 20742 22788 20950
rect 22712 20710 22718 20742
rect 21760 20672 21836 20678
rect 22717 20678 22718 20710
rect 22782 20710 22788 20742
rect 22984 20950 22990 20982
rect 23054 20982 23055 21014
rect 23533 21014 23599 21015
rect 23533 20982 23534 21014
rect 23054 20950 23060 20982
rect 22984 20742 23060 20950
rect 22782 20678 22783 20710
rect 22717 20677 22783 20678
rect 22984 20678 22990 20742
rect 23054 20678 23060 20742
rect 22984 20672 23060 20678
rect 23528 20950 23534 20982
rect 23598 20982 23599 21014
rect 115192 21014 115268 21020
rect 23598 20950 23604 20982
rect 23528 20742 23604 20950
rect 23528 20678 23534 20742
rect 23598 20678 23604 20742
rect 115192 20950 115198 21014
rect 115262 20950 115268 21014
rect 115192 20742 115268 20950
rect 115192 20710 115198 20742
rect 23528 20672 23604 20678
rect 115197 20678 115198 20710
rect 115262 20710 115268 20742
rect 115600 21014 115676 21020
rect 115600 20950 115606 21014
rect 115670 20950 115676 21014
rect 115600 20742 115676 20950
rect 115600 20710 115606 20742
rect 115262 20678 115263 20710
rect 115197 20677 115263 20678
rect 115605 20678 115606 20710
rect 115670 20710 115676 20742
rect 116008 21014 116084 21020
rect 116008 20950 116014 21014
rect 116078 20950 116084 21014
rect 116829 21014 116895 21015
rect 116829 20982 116830 21014
rect 116008 20742 116084 20950
rect 116008 20710 116014 20742
rect 115670 20678 115671 20710
rect 115605 20677 115671 20678
rect 116013 20678 116014 20710
rect 116078 20710 116084 20742
rect 116824 20950 116830 20982
rect 116894 20982 116895 21014
rect 118864 21014 118940 21020
rect 116894 20950 116900 20982
rect 116824 20742 116900 20950
rect 116078 20678 116079 20710
rect 116013 20677 116079 20678
rect 116824 20678 116830 20742
rect 116894 20678 116900 20742
rect 116824 20672 116900 20678
rect 118864 20950 118870 21014
rect 118934 20950 118940 21014
rect 119413 21014 119479 21015
rect 119413 20982 119414 21014
rect 21901 20606 21967 20607
rect 21901 20574 21902 20606
rect 19856 20302 19862 20334
rect 19312 20264 19388 20270
rect 19861 20270 19862 20302
rect 19926 20302 19932 20334
rect 21896 20542 21902 20574
rect 21966 20574 21967 20606
rect 22309 20606 22375 20607
rect 22309 20574 22310 20606
rect 21966 20542 21972 20574
rect 21896 20334 21972 20542
rect 19926 20270 19927 20302
rect 19861 20269 19927 20270
rect 21896 20270 21902 20334
rect 21966 20270 21972 20334
rect 21896 20264 21972 20270
rect 22304 20542 22310 20574
rect 22374 20574 22375 20606
rect 22712 20606 22788 20612
rect 22374 20542 22380 20574
rect 22304 20334 22380 20542
rect 22304 20270 22310 20334
rect 22374 20270 22380 20334
rect 22712 20542 22718 20606
rect 22782 20542 22788 20606
rect 22989 20606 23055 20607
rect 22989 20574 22990 20606
rect 22712 20334 22788 20542
rect 22712 20302 22718 20334
rect 22304 20264 22380 20270
rect 22717 20270 22718 20302
rect 22782 20302 22788 20334
rect 22984 20542 22990 20574
rect 23054 20574 23055 20606
rect 23392 20606 23468 20612
rect 23054 20542 23060 20574
rect 22984 20334 23060 20542
rect 22782 20270 22783 20302
rect 22717 20269 22783 20270
rect 22984 20270 22990 20334
rect 23054 20270 23060 20334
rect 23392 20542 23398 20606
rect 23462 20542 23468 20606
rect 23392 20334 23468 20542
rect 23392 20302 23398 20334
rect 22984 20264 23060 20270
rect 23397 20270 23398 20302
rect 23462 20302 23468 20334
rect 115192 20606 115268 20612
rect 115192 20542 115198 20606
rect 115262 20542 115268 20606
rect 115192 20334 115268 20542
rect 115192 20302 115198 20334
rect 23462 20270 23463 20302
rect 23397 20269 23463 20270
rect 115197 20270 115198 20302
rect 115262 20302 115268 20334
rect 115600 20606 115676 20612
rect 115600 20542 115606 20606
rect 115670 20542 115676 20606
rect 116013 20606 116079 20607
rect 116013 20574 116014 20606
rect 115600 20334 115676 20542
rect 115600 20302 115606 20334
rect 115262 20270 115263 20302
rect 115197 20269 115263 20270
rect 115605 20270 115606 20302
rect 115670 20302 115676 20334
rect 116008 20542 116014 20574
rect 116078 20574 116079 20606
rect 116960 20606 117036 20612
rect 116078 20542 116084 20574
rect 116008 20334 116084 20542
rect 115670 20270 115671 20302
rect 115605 20269 115671 20270
rect 116008 20270 116014 20334
rect 116078 20270 116084 20334
rect 116960 20542 116966 20606
rect 117030 20542 117036 20606
rect 116960 20334 117036 20542
rect 116960 20302 116966 20334
rect 116008 20264 116084 20270
rect 116965 20270 116966 20302
rect 117030 20302 117036 20334
rect 118864 20334 118940 20950
rect 118864 20302 118870 20334
rect 117030 20270 117031 20302
rect 116965 20269 117031 20270
rect 118869 20270 118870 20302
rect 118934 20302 118940 20334
rect 119408 20950 119414 20982
rect 119478 20982 119479 21014
rect 119816 21014 119892 21020
rect 119478 20950 119484 20982
rect 119408 20334 119484 20950
rect 118934 20270 118935 20302
rect 118869 20269 118935 20270
rect 119408 20270 119414 20334
rect 119478 20270 119484 20334
rect 119816 20950 119822 21014
rect 119886 20950 119892 21014
rect 119816 20334 119892 20950
rect 119816 20302 119822 20334
rect 119408 20264 119484 20270
rect 119821 20270 119822 20302
rect 119886 20302 119892 20334
rect 137496 20470 137844 22310
rect 137496 20406 137502 20470
rect 137566 20406 137844 20470
rect 119886 20270 119887 20302
rect 119821 20269 119887 20270
rect 2540 17958 2606 17959
rect 2540 17894 2541 17958
rect 2605 17894 2606 17958
rect 2540 17893 2606 17894
rect 3808 17614 3884 20264
rect 17136 20198 17212 20204
rect 17136 20134 17142 20198
rect 17206 20134 17212 20198
rect 17136 19110 17212 20134
rect 17136 19078 17142 19110
rect 17141 19046 17142 19078
rect 17206 19078 17212 19110
rect 17544 20198 17620 20204
rect 17544 20134 17550 20198
rect 17614 20134 17620 20198
rect 17206 19046 17207 19078
rect 17141 19045 17207 19046
rect 3808 17582 3814 17614
rect 3813 17550 3814 17582
rect 3878 17582 3884 17614
rect 15232 18838 15308 18844
rect 15232 18774 15238 18838
rect 15302 18774 15308 18838
rect 3878 17550 3879 17582
rect 3813 17549 3879 17550
rect 952 17006 1230 17070
rect 1294 17006 1300 17070
rect 952 15574 1300 17006
rect 15096 17478 15172 17484
rect 15096 17414 15102 17478
rect 15166 17414 15172 17478
rect 952 15510 1230 15574
rect 1294 15510 1300 15574
rect 3128 16118 3204 16124
rect 3128 16054 3134 16118
rect 3198 16054 3204 16118
rect 3128 15574 3204 16054
rect 3128 15542 3134 15574
rect 952 13942 1300 15510
rect 3133 15510 3134 15542
rect 3198 15542 3204 15574
rect 3198 15510 3199 15542
rect 3133 15509 3199 15510
rect 15096 14758 15172 17414
rect 15232 16254 15308 18774
rect 17544 17614 17620 20134
rect 17544 17582 17550 17614
rect 17549 17550 17550 17582
rect 17614 17582 17620 17614
rect 21760 20198 21836 20204
rect 21760 20134 21766 20198
rect 21830 20134 21836 20198
rect 23533 20198 23599 20199
rect 23533 20166 23534 20198
rect 17614 17550 17615 17582
rect 17549 17549 17615 17550
rect 21760 17342 21836 20134
rect 23528 20134 23534 20166
rect 23598 20166 23599 20198
rect 24213 20198 24279 20199
rect 24213 20166 24214 20198
rect 23598 20134 23604 20166
rect 23528 19790 23604 20134
rect 23528 19726 23534 19790
rect 23598 19726 23604 19790
rect 23528 19720 23604 19726
rect 24208 20134 24214 20166
rect 24278 20166 24279 20198
rect 121317 20198 121383 20199
rect 121317 20166 121318 20198
rect 24278 20134 24284 20166
rect 24208 19790 24284 20134
rect 121312 20134 121318 20166
rect 121382 20166 121383 20198
rect 124173 20198 124239 20199
rect 124173 20166 124174 20198
rect 121382 20134 121388 20166
rect 24208 19726 24214 19790
rect 24278 19726 24284 19790
rect 24208 19720 24284 19726
rect 28288 20062 28364 20068
rect 28288 19998 28294 20062
rect 28358 19998 28364 20062
rect 21760 17310 21766 17342
rect 21765 17278 21766 17310
rect 21830 17310 21836 17342
rect 23392 19654 23468 19660
rect 23392 19590 23398 19654
rect 23462 19590 23468 19654
rect 27885 19654 27951 19655
rect 27885 19622 27886 19654
rect 21830 17278 21831 17310
rect 21765 17277 21831 17278
rect 15232 16222 15238 16254
rect 15237 16190 15238 16222
rect 15302 16222 15308 16254
rect 21080 17206 21156 17212
rect 21080 17142 21086 17206
rect 21150 17142 21156 17206
rect 15302 16190 15303 16222
rect 15237 16189 15303 16190
rect 15096 14726 15102 14758
rect 15101 14694 15102 14726
rect 15166 14726 15172 14758
rect 15232 16118 15308 16124
rect 15232 16054 15238 16118
rect 15302 16054 15308 16118
rect 15166 14694 15167 14726
rect 15101 14693 15167 14694
rect 952 13878 1230 13942
rect 1294 13878 1300 13942
rect 952 12174 1300 13878
rect 15096 14622 15172 14628
rect 15096 14558 15102 14622
rect 15166 14558 15172 14622
rect 3133 13806 3199 13807
rect 3133 13774 3134 13806
rect 3128 13742 3134 13774
rect 3198 13774 3199 13806
rect 3198 13742 3204 13774
rect 3128 13398 3204 13742
rect 3128 13334 3134 13398
rect 3198 13334 3204 13398
rect 3128 13328 3204 13334
rect 952 12110 1230 12174
rect 1294 12110 1300 12174
rect 952 10406 1300 12110
rect 15096 12038 15172 14558
rect 15232 13398 15308 16054
rect 21080 14622 21156 17142
rect 21080 14590 21086 14622
rect 21085 14558 21086 14590
rect 21150 14590 21156 14622
rect 22304 15846 22380 15852
rect 22304 15782 22310 15846
rect 22374 15782 22380 15846
rect 23392 15846 23468 19590
rect 27880 19590 27886 19622
rect 27950 19622 27951 19654
rect 28288 19654 28364 19998
rect 28288 19622 28294 19654
rect 27950 19590 27956 19622
rect 27880 19382 27956 19590
rect 28293 19590 28294 19622
rect 28358 19622 28364 19654
rect 110160 19790 110236 19796
rect 110160 19726 110166 19790
rect 110230 19726 110236 19790
rect 28358 19590 28359 19622
rect 28293 19589 28359 19590
rect 27880 19318 27886 19382
rect 27950 19318 27956 19382
rect 27880 19312 27956 19318
rect 60520 19382 60596 19388
rect 60520 19318 60526 19382
rect 60590 19318 60596 19382
rect 29109 19246 29175 19247
rect 29109 19214 29110 19246
rect 29104 19182 29110 19214
rect 29174 19214 29175 19246
rect 30469 19246 30535 19247
rect 30469 19214 30470 19246
rect 29174 19182 29180 19214
rect 29104 18838 29180 19182
rect 29104 18774 29110 18838
rect 29174 18774 29180 18838
rect 29104 18768 29180 18774
rect 30464 19182 30470 19214
rect 30534 19214 30535 19246
rect 32232 19246 32308 19252
rect 30534 19182 30540 19214
rect 30464 18838 30540 19182
rect 30464 18774 30470 18838
rect 30534 18774 30540 18838
rect 32232 19182 32238 19246
rect 32302 19182 32308 19246
rect 32232 18838 32308 19182
rect 32232 18806 32238 18838
rect 30464 18768 30540 18774
rect 32237 18774 32238 18806
rect 32302 18806 32308 18838
rect 32776 19246 32852 19252
rect 32776 19182 32782 19246
rect 32846 19182 32852 19246
rect 32917 19246 32983 19247
rect 32917 19214 32918 19246
rect 32776 18838 32852 19182
rect 32776 18806 32782 18838
rect 32302 18774 32303 18806
rect 32237 18773 32303 18774
rect 32781 18774 32782 18806
rect 32846 18806 32852 18838
rect 32912 19182 32918 19214
rect 32982 19214 32983 19246
rect 34141 19246 34207 19247
rect 34141 19214 34142 19246
rect 32982 19182 32988 19214
rect 32912 18838 32988 19182
rect 32846 18774 32847 18806
rect 32781 18773 32847 18774
rect 32912 18774 32918 18838
rect 32982 18774 32988 18838
rect 32912 18768 32988 18774
rect 34136 19182 34142 19214
rect 34206 19214 34207 19246
rect 34680 19246 34756 19252
rect 34206 19182 34212 19214
rect 34136 18838 34212 19182
rect 34136 18774 34142 18838
rect 34206 18774 34212 18838
rect 34680 19182 34686 19246
rect 34750 19182 34756 19246
rect 35501 19246 35567 19247
rect 35501 19214 35502 19246
rect 34680 18838 34756 19182
rect 34680 18806 34686 18838
rect 34136 18768 34212 18774
rect 34685 18774 34686 18806
rect 34750 18806 34756 18838
rect 35496 19182 35502 19214
rect 35566 19214 35567 19246
rect 35904 19246 35980 19252
rect 35566 19182 35572 19214
rect 35496 18838 35572 19182
rect 35904 19182 35910 19246
rect 35974 19182 35980 19246
rect 36725 19246 36791 19247
rect 36725 19214 36726 19246
rect 35904 18974 35980 19182
rect 35904 18942 35910 18974
rect 35909 18910 35910 18942
rect 35974 18942 35980 18974
rect 36720 19182 36726 19214
rect 36790 19214 36791 19246
rect 38488 19246 38564 19252
rect 36790 19182 36796 19214
rect 35974 18910 35975 18942
rect 35909 18909 35975 18910
rect 34750 18774 34751 18806
rect 34685 18773 34751 18774
rect 35496 18774 35502 18838
rect 35566 18774 35572 18838
rect 35496 18768 35572 18774
rect 36720 18838 36796 19182
rect 36720 18774 36726 18838
rect 36790 18774 36796 18838
rect 38488 19182 38494 19246
rect 38558 19182 38564 19246
rect 39173 19246 39239 19247
rect 39173 19214 39174 19246
rect 38488 18838 38564 19182
rect 38488 18806 38494 18838
rect 36720 18768 36796 18774
rect 38493 18774 38494 18806
rect 38558 18806 38564 18838
rect 39168 19182 39174 19214
rect 39238 19214 39239 19246
rect 39576 19246 39652 19252
rect 39238 19182 39244 19214
rect 39168 18838 39244 19182
rect 38558 18774 38559 18806
rect 38493 18773 38559 18774
rect 39168 18774 39174 18838
rect 39238 18774 39244 18838
rect 39576 19182 39582 19246
rect 39646 19182 39652 19246
rect 39576 18838 39652 19182
rect 39576 18806 39582 18838
rect 39168 18768 39244 18774
rect 39581 18774 39582 18806
rect 39646 18806 39652 18838
rect 40936 19246 41012 19252
rect 40936 19182 40942 19246
rect 41006 19182 41012 19246
rect 41621 19246 41687 19247
rect 41621 19214 41622 19246
rect 40936 18838 41012 19182
rect 40936 18806 40942 18838
rect 39646 18774 39647 18806
rect 39581 18773 39647 18774
rect 40941 18774 40942 18806
rect 41006 18806 41012 18838
rect 41616 19182 41622 19214
rect 41686 19214 41687 19246
rect 42845 19246 42911 19247
rect 42845 19214 42846 19246
rect 41686 19182 41692 19214
rect 41616 18838 41692 19182
rect 41006 18774 41007 18806
rect 40941 18773 41007 18774
rect 41616 18774 41622 18838
rect 41686 18774 41692 18838
rect 41616 18768 41692 18774
rect 42840 19182 42846 19214
rect 42910 19214 42911 19246
rect 43384 19246 43460 19252
rect 42910 19182 42916 19214
rect 42840 18838 42916 19182
rect 42840 18774 42846 18838
rect 42910 18774 42916 18838
rect 43384 19182 43390 19246
rect 43454 19182 43460 19246
rect 44069 19246 44135 19247
rect 44069 19214 44070 19246
rect 43384 18838 43460 19182
rect 43384 18806 43390 18838
rect 42840 18768 42916 18774
rect 43389 18774 43390 18806
rect 43454 18806 43460 18838
rect 44064 19182 44070 19214
rect 44134 19214 44135 19246
rect 45701 19246 45767 19247
rect 45701 19214 45702 19246
rect 44134 19182 44140 19214
rect 44064 18838 44140 19182
rect 43454 18774 43455 18806
rect 43389 18773 43455 18774
rect 44064 18774 44070 18838
rect 44134 18774 44140 18838
rect 44064 18768 44140 18774
rect 45696 19182 45702 19214
rect 45766 19214 45767 19246
rect 46653 19246 46719 19247
rect 46653 19214 46654 19246
rect 45766 19182 45772 19214
rect 45696 18838 45772 19182
rect 45696 18774 45702 18838
rect 45766 18774 45772 18838
rect 45696 18768 45772 18774
rect 46648 19182 46654 19214
rect 46718 19214 46719 19246
rect 47192 19246 47268 19252
rect 46718 19182 46724 19214
rect 46648 18838 46724 19182
rect 46648 18774 46654 18838
rect 46718 18774 46724 18838
rect 47192 19182 47198 19246
rect 47262 19182 47268 19246
rect 47877 19246 47943 19247
rect 47877 19214 47878 19246
rect 47192 18838 47268 19182
rect 47192 18806 47198 18838
rect 46648 18768 46724 18774
rect 47197 18774 47198 18806
rect 47262 18806 47268 18838
rect 47872 19182 47878 19214
rect 47942 19214 47943 19246
rect 48416 19246 48492 19252
rect 47942 19182 47948 19214
rect 47872 18838 47948 19182
rect 47262 18774 47263 18806
rect 47197 18773 47263 18774
rect 47872 18774 47878 18838
rect 47942 18774 47948 18838
rect 48416 19182 48422 19246
rect 48486 19182 48492 19246
rect 49101 19246 49167 19247
rect 49101 19214 49102 19246
rect 48416 18838 48492 19182
rect 48416 18806 48422 18838
rect 47872 18768 47948 18774
rect 48421 18774 48422 18806
rect 48486 18806 48492 18838
rect 49096 19182 49102 19214
rect 49166 19214 49167 19246
rect 49640 19246 49716 19252
rect 49166 19182 49172 19214
rect 49096 18838 49172 19182
rect 48486 18774 48487 18806
rect 48421 18773 48487 18774
rect 49096 18774 49102 18838
rect 49166 18774 49172 18838
rect 49640 19182 49646 19246
rect 49710 19182 49716 19246
rect 50461 19246 50527 19247
rect 50461 19214 50462 19246
rect 49640 18838 49716 19182
rect 49640 18806 49646 18838
rect 49096 18768 49172 18774
rect 49645 18774 49646 18806
rect 49710 18806 49716 18838
rect 50456 19182 50462 19214
rect 50526 19214 50527 19246
rect 52088 19246 52164 19252
rect 50526 19182 50532 19214
rect 50456 18838 50532 19182
rect 49710 18774 49711 18806
rect 49645 18773 49711 18774
rect 50456 18774 50462 18838
rect 50526 18774 50532 18838
rect 52088 19182 52094 19246
rect 52158 19182 52164 19246
rect 52909 19246 52975 19247
rect 52909 19214 52910 19246
rect 52088 18838 52164 19182
rect 52088 18806 52094 18838
rect 50456 18768 50532 18774
rect 52093 18774 52094 18806
rect 52158 18806 52164 18838
rect 52904 19182 52910 19214
rect 52974 19214 52975 19246
rect 54133 19246 54199 19247
rect 54133 19214 54134 19246
rect 52974 19182 52980 19214
rect 52904 18838 52980 19182
rect 52158 18774 52159 18806
rect 52093 18773 52159 18774
rect 52904 18774 52910 18838
rect 52974 18774 52980 18838
rect 52904 18768 52980 18774
rect 54128 19182 54134 19214
rect 54198 19214 54199 19246
rect 54672 19246 54748 19252
rect 54198 19182 54204 19214
rect 54128 18838 54204 19182
rect 54128 18774 54134 18838
rect 54198 18774 54204 18838
rect 54672 19182 54678 19246
rect 54742 19182 54748 19246
rect 55357 19246 55423 19247
rect 55357 19214 55358 19246
rect 54672 18838 54748 19182
rect 54672 18806 54678 18838
rect 54128 18768 54204 18774
rect 54677 18774 54678 18806
rect 54742 18806 54748 18838
rect 55352 19182 55358 19214
rect 55422 19214 55423 19246
rect 55896 19246 55972 19252
rect 55422 19182 55428 19214
rect 55352 18838 55428 19182
rect 54742 18774 54743 18806
rect 54677 18773 54743 18774
rect 55352 18774 55358 18838
rect 55422 18774 55428 18838
rect 55896 19182 55902 19246
rect 55966 19182 55972 19246
rect 56717 19246 56783 19247
rect 56717 19214 56718 19246
rect 55896 18838 55972 19182
rect 55896 18806 55902 18838
rect 55352 18768 55428 18774
rect 55901 18774 55902 18806
rect 55966 18806 55972 18838
rect 56712 19182 56718 19214
rect 56782 19214 56783 19246
rect 57120 19246 57196 19252
rect 56782 19182 56788 19214
rect 56712 18838 56788 19182
rect 55966 18774 55967 18806
rect 55901 18773 55967 18774
rect 56712 18774 56718 18838
rect 56782 18774 56788 18838
rect 57120 19182 57126 19246
rect 57190 19182 57196 19246
rect 57669 19246 57735 19247
rect 57669 19214 57670 19246
rect 57120 18838 57196 19182
rect 57120 18806 57126 18838
rect 56712 18768 56788 18774
rect 57125 18774 57126 18806
rect 57190 18806 57196 18838
rect 57664 19182 57670 19214
rect 57734 19214 57735 19246
rect 58344 19246 58420 19252
rect 57734 19182 57740 19214
rect 57664 18838 57740 19182
rect 57190 18774 57191 18806
rect 57125 18773 57191 18774
rect 57664 18774 57670 18838
rect 57734 18774 57740 18838
rect 58344 19182 58350 19246
rect 58414 19182 58420 19246
rect 59165 19246 59231 19247
rect 59165 19214 59166 19246
rect 58344 18838 58420 19182
rect 58344 18806 58350 18838
rect 57664 18768 57740 18774
rect 58349 18774 58350 18806
rect 58414 18806 58420 18838
rect 59160 19182 59166 19214
rect 59230 19214 59231 19246
rect 59704 19246 59780 19252
rect 59230 19182 59236 19214
rect 59160 18838 59236 19182
rect 58414 18774 58415 18806
rect 58349 18773 58415 18774
rect 59160 18774 59166 18838
rect 59230 18774 59236 18838
rect 59704 19182 59710 19246
rect 59774 19182 59780 19246
rect 59704 18838 59780 19182
rect 59704 18806 59710 18838
rect 59160 18768 59236 18774
rect 59709 18774 59710 18806
rect 59774 18806 59780 18838
rect 60520 18838 60596 19318
rect 94248 19382 94324 19388
rect 94248 19318 94254 19382
rect 94318 19318 94324 19382
rect 61613 19246 61679 19247
rect 61613 19214 61614 19246
rect 60520 18806 60526 18838
rect 59774 18774 59775 18806
rect 59709 18773 59775 18774
rect 60525 18774 60526 18806
rect 60590 18806 60596 18838
rect 61608 19182 61614 19214
rect 61678 19214 61679 19246
rect 62152 19246 62228 19252
rect 61678 19182 61684 19214
rect 61608 18838 61684 19182
rect 60590 18774 60591 18806
rect 60525 18773 60591 18774
rect 61608 18774 61614 18838
rect 61678 18774 61684 18838
rect 62152 19182 62158 19246
rect 62222 19182 62228 19246
rect 62837 19246 62903 19247
rect 62837 19214 62838 19246
rect 62152 18838 62228 19182
rect 62152 18806 62158 18838
rect 61608 18768 61684 18774
rect 62157 18774 62158 18806
rect 62222 18806 62228 18838
rect 62832 19182 62838 19214
rect 62902 19214 62903 19246
rect 63376 19246 63452 19252
rect 62902 19182 62908 19214
rect 62832 18838 62908 19182
rect 62222 18774 62223 18806
rect 62157 18773 62223 18774
rect 62832 18774 62838 18838
rect 62902 18774 62908 18838
rect 63376 19182 63382 19246
rect 63446 19182 63452 19246
rect 64197 19246 64263 19247
rect 64197 19214 64198 19246
rect 63376 18838 63452 19182
rect 63376 18806 63382 18838
rect 62832 18768 62908 18774
rect 63381 18774 63382 18806
rect 63446 18806 63452 18838
rect 64192 19182 64198 19214
rect 64262 19214 64263 19246
rect 64600 19246 64676 19252
rect 64262 19182 64268 19214
rect 64192 18838 64268 19182
rect 63446 18774 63447 18806
rect 63381 18773 63447 18774
rect 64192 18774 64198 18838
rect 64262 18774 64268 18838
rect 64600 19182 64606 19246
rect 64670 19182 64676 19246
rect 64600 18838 64676 19182
rect 64600 18806 64606 18838
rect 64192 18768 64268 18774
rect 64605 18774 64606 18806
rect 64670 18806 64676 18838
rect 65824 19246 65900 19252
rect 65824 19182 65830 19246
rect 65894 19182 65900 19246
rect 65824 18838 65900 19182
rect 65824 18806 65830 18838
rect 64670 18774 64671 18806
rect 64605 18773 64671 18774
rect 65829 18774 65830 18806
rect 65894 18806 65900 18838
rect 67184 19246 67260 19252
rect 67184 19182 67190 19246
rect 67254 19182 67260 19246
rect 67869 19246 67935 19247
rect 67869 19214 67870 19246
rect 67184 18838 67260 19182
rect 67184 18806 67190 18838
rect 65894 18774 65895 18806
rect 65829 18773 65895 18774
rect 67189 18774 67190 18806
rect 67254 18806 67260 18838
rect 67864 19182 67870 19214
rect 67934 19214 67935 19246
rect 68408 19246 68484 19252
rect 67934 19182 67940 19214
rect 67864 18838 67940 19182
rect 67254 18774 67255 18806
rect 67189 18773 67255 18774
rect 67864 18774 67870 18838
rect 67934 18774 67940 18838
rect 68408 19182 68414 19246
rect 68478 19182 68484 19246
rect 69093 19246 69159 19247
rect 69093 19214 69094 19246
rect 68408 18838 68484 19182
rect 68408 18806 68414 18838
rect 67864 18768 67940 18774
rect 68413 18774 68414 18806
rect 68478 18806 68484 18838
rect 69088 19182 69094 19214
rect 69158 19214 69159 19246
rect 70317 19246 70383 19247
rect 70317 19214 70318 19246
rect 69158 19182 69164 19214
rect 69088 18838 69164 19182
rect 68478 18774 68479 18806
rect 68413 18773 68479 18774
rect 69088 18774 69094 18838
rect 69158 18774 69164 18838
rect 69088 18768 69164 18774
rect 70312 19182 70318 19214
rect 70382 19214 70383 19246
rect 70856 19246 70932 19252
rect 70382 19182 70388 19214
rect 70312 18838 70388 19182
rect 70312 18774 70318 18838
rect 70382 18774 70388 18838
rect 70856 19182 70862 19246
rect 70926 19182 70932 19246
rect 71541 19246 71607 19247
rect 71541 19214 71542 19246
rect 70856 18838 70932 19182
rect 70856 18806 70862 18838
rect 70312 18768 70388 18774
rect 70861 18774 70862 18806
rect 70926 18806 70932 18838
rect 71536 19182 71542 19214
rect 71606 19214 71607 19246
rect 73304 19246 73380 19252
rect 71606 19182 71612 19214
rect 71536 18838 71612 19182
rect 70926 18774 70927 18806
rect 70861 18773 70927 18774
rect 71536 18774 71542 18838
rect 71606 18774 71612 18838
rect 73304 19182 73310 19246
rect 73374 19182 73380 19246
rect 73304 18838 73380 19182
rect 73304 18806 73310 18838
rect 71536 18768 71612 18774
rect 73309 18774 73310 18806
rect 73374 18806 73380 18838
rect 74664 19246 74740 19252
rect 74664 19182 74670 19246
rect 74734 19182 74740 19246
rect 74664 18838 74740 19182
rect 74664 18806 74670 18838
rect 73374 18774 73375 18806
rect 73309 18773 73375 18774
rect 74669 18774 74670 18806
rect 74734 18806 74740 18838
rect 75208 19246 75284 19252
rect 75208 19182 75214 19246
rect 75278 19182 75284 19246
rect 75349 19246 75415 19247
rect 75349 19214 75350 19246
rect 75208 18838 75284 19182
rect 75208 18806 75214 18838
rect 74734 18774 74735 18806
rect 74669 18773 74735 18774
rect 75213 18774 75214 18806
rect 75278 18806 75284 18838
rect 75344 19182 75350 19214
rect 75414 19214 75415 19246
rect 75888 19246 75964 19252
rect 75414 19182 75420 19214
rect 75344 18838 75420 19182
rect 75278 18774 75279 18806
rect 75213 18773 75279 18774
rect 75344 18774 75350 18838
rect 75414 18774 75420 18838
rect 75888 19182 75894 19246
rect 75958 19182 75964 19246
rect 76573 19246 76639 19247
rect 76573 19214 76574 19246
rect 75888 18838 75964 19182
rect 75888 18806 75894 18838
rect 75344 18768 75420 18774
rect 75893 18774 75894 18806
rect 75958 18806 75964 18838
rect 76568 19182 76574 19214
rect 76638 19214 76639 19246
rect 77112 19246 77188 19252
rect 76638 19182 76644 19214
rect 76568 18838 76644 19182
rect 75958 18774 75959 18806
rect 75893 18773 75959 18774
rect 76568 18774 76574 18838
rect 76638 18774 76644 18838
rect 77112 19182 77118 19246
rect 77182 19182 77188 19246
rect 77933 19246 77999 19247
rect 77933 19214 77934 19246
rect 77112 18838 77188 19182
rect 77112 18806 77118 18838
rect 76568 18768 76644 18774
rect 77117 18774 77118 18806
rect 77182 18806 77188 18838
rect 77928 19182 77934 19214
rect 77998 19214 77999 19246
rect 78336 19246 78412 19252
rect 77998 19182 78004 19214
rect 77928 18838 78004 19182
rect 78336 19182 78342 19246
rect 78406 19182 78412 19246
rect 79157 19246 79223 19247
rect 79157 19214 79158 19246
rect 78336 18974 78412 19182
rect 78336 18942 78342 18974
rect 78341 18910 78342 18942
rect 78406 18942 78412 18974
rect 79152 19182 79158 19214
rect 79222 19214 79223 19246
rect 80512 19246 80588 19252
rect 79222 19182 79228 19214
rect 78406 18910 78407 18942
rect 78341 18909 78407 18910
rect 77182 18774 77183 18806
rect 77117 18773 77183 18774
rect 77928 18774 77934 18838
rect 77998 18774 78004 18838
rect 77928 18768 78004 18774
rect 79152 18838 79228 19182
rect 79152 18774 79158 18838
rect 79222 18774 79228 18838
rect 80512 19182 80518 19246
rect 80582 19182 80588 19246
rect 80512 18838 80588 19182
rect 80512 18806 80518 18838
rect 79152 18768 79228 18774
rect 80517 18774 80518 18806
rect 80582 18806 80588 18838
rect 81464 19246 81540 19252
rect 81464 19182 81470 19246
rect 81534 19182 81540 19246
rect 81605 19246 81671 19247
rect 81605 19214 81606 19246
rect 81464 18838 81540 19182
rect 81464 18806 81470 18838
rect 80582 18774 80583 18806
rect 80517 18773 80583 18774
rect 81469 18774 81470 18806
rect 81534 18806 81540 18838
rect 81600 19182 81606 19214
rect 81670 19214 81671 19246
rect 82008 19246 82084 19252
rect 81670 19182 81676 19214
rect 81600 18838 81676 19182
rect 81534 18774 81535 18806
rect 81469 18773 81535 18774
rect 81600 18774 81606 18838
rect 81670 18774 81676 18838
rect 82008 19182 82014 19246
rect 82078 19182 82084 19246
rect 82829 19246 82895 19247
rect 82829 19214 82830 19246
rect 82008 18838 82084 19182
rect 82008 18806 82014 18838
rect 81600 18768 81676 18774
rect 82013 18774 82014 18806
rect 82078 18806 82084 18838
rect 82824 19182 82830 19214
rect 82894 19214 82895 19246
rect 83368 19246 83444 19252
rect 82894 19182 82900 19214
rect 82824 18838 82900 19182
rect 82078 18774 82079 18806
rect 82013 18773 82079 18774
rect 82824 18774 82830 18838
rect 82894 18774 82900 18838
rect 83368 19182 83374 19246
rect 83438 19182 83444 19246
rect 84053 19246 84119 19247
rect 84053 19214 84054 19246
rect 83368 18838 83444 19182
rect 83368 18806 83374 18838
rect 82824 18768 82900 18774
rect 83373 18774 83374 18806
rect 83438 18806 83444 18838
rect 84048 19182 84054 19214
rect 84118 19214 84119 19246
rect 84592 19246 84668 19252
rect 84118 19182 84124 19214
rect 84048 18838 84124 19182
rect 83438 18774 83439 18806
rect 83373 18773 83439 18774
rect 84048 18774 84054 18838
rect 84118 18774 84124 18838
rect 84592 19182 84598 19246
rect 84662 19182 84668 19246
rect 85277 19246 85343 19247
rect 85277 19214 85278 19246
rect 84592 18838 84668 19182
rect 84592 18806 84598 18838
rect 84048 18768 84124 18774
rect 84597 18774 84598 18806
rect 84662 18806 84668 18838
rect 85272 19182 85278 19214
rect 85342 19214 85343 19246
rect 85816 19246 85892 19252
rect 85342 19182 85348 19214
rect 85272 18838 85348 19182
rect 84662 18774 84663 18806
rect 84597 18773 84663 18774
rect 85272 18774 85278 18838
rect 85342 18774 85348 18838
rect 85816 19182 85822 19246
rect 85886 19182 85892 19246
rect 86501 19246 86567 19247
rect 86501 19214 86502 19246
rect 85816 18838 85892 19182
rect 85816 18806 85822 18838
rect 85272 18768 85348 18774
rect 85821 18774 85822 18806
rect 85886 18806 85892 18838
rect 86496 19182 86502 19214
rect 86566 19214 86567 19246
rect 86768 19246 86844 19252
rect 86566 19182 86572 19214
rect 86496 18838 86572 19182
rect 85886 18774 85887 18806
rect 85821 18773 85887 18774
rect 86496 18774 86502 18838
rect 86566 18774 86572 18838
rect 86768 19182 86774 19246
rect 86838 19182 86844 19246
rect 88133 19246 88199 19247
rect 88133 19214 88134 19246
rect 86768 18838 86844 19182
rect 86768 18806 86774 18838
rect 86496 18768 86572 18774
rect 86773 18774 86774 18806
rect 86838 18806 86844 18838
rect 88128 19182 88134 19214
rect 88198 19214 88199 19246
rect 89624 19246 89700 19252
rect 88198 19182 88204 19214
rect 88128 18838 88204 19182
rect 86838 18774 86839 18806
rect 86773 18773 86839 18774
rect 88128 18774 88134 18838
rect 88198 18774 88204 18838
rect 89624 19182 89630 19246
rect 89694 19182 89700 19246
rect 90309 19246 90375 19247
rect 90309 19214 90310 19246
rect 89624 18838 89700 19182
rect 89624 18806 89630 18838
rect 88128 18768 88204 18774
rect 89629 18774 89630 18806
rect 89694 18806 89700 18838
rect 90304 19182 90310 19214
rect 90374 19214 90375 19246
rect 90848 19246 90924 19252
rect 90374 19182 90380 19214
rect 90304 18838 90380 19182
rect 89694 18774 89695 18806
rect 89629 18773 89695 18774
rect 90304 18774 90310 18838
rect 90374 18774 90380 18838
rect 90848 19182 90854 19246
rect 90918 19182 90924 19246
rect 90848 18838 90924 19182
rect 90848 18806 90854 18838
rect 90304 18768 90380 18774
rect 90853 18774 90854 18806
rect 90918 18806 90924 18838
rect 92072 19246 92148 19252
rect 92072 19182 92078 19246
rect 92142 19182 92148 19246
rect 92757 19246 92823 19247
rect 92757 19214 92758 19246
rect 92072 18838 92148 19182
rect 92072 18806 92078 18838
rect 90918 18774 90919 18806
rect 90853 18773 90919 18774
rect 92077 18774 92078 18806
rect 92142 18806 92148 18838
rect 92752 19182 92758 19214
rect 92822 19214 92823 19246
rect 92822 19182 92828 19214
rect 92752 18838 92828 19182
rect 92142 18774 92143 18806
rect 92077 18773 92143 18774
rect 92752 18774 92758 18838
rect 92822 18774 92828 18838
rect 94248 18838 94324 19318
rect 102952 19382 103028 19388
rect 102952 19318 102958 19382
rect 103022 19318 103028 19382
rect 94389 19246 94455 19247
rect 94389 19214 94390 19246
rect 94248 18806 94254 18838
rect 92752 18768 92828 18774
rect 94253 18774 94254 18806
rect 94318 18806 94324 18838
rect 94384 19182 94390 19214
rect 94454 19214 94455 19246
rect 95341 19246 95407 19247
rect 95341 19214 95342 19246
rect 94454 19182 94460 19214
rect 94384 18838 94460 19182
rect 94318 18774 94319 18806
rect 94253 18773 94319 18774
rect 94384 18774 94390 18838
rect 94454 18774 94460 18838
rect 94384 18768 94460 18774
rect 95336 19182 95342 19214
rect 95406 19214 95407 19246
rect 95744 19246 95820 19252
rect 95406 19182 95412 19214
rect 95336 18838 95412 19182
rect 95336 18774 95342 18838
rect 95406 18774 95412 18838
rect 95744 19182 95750 19246
rect 95814 19182 95820 19246
rect 96565 19246 96631 19247
rect 96565 19214 96566 19246
rect 95744 18838 95820 19182
rect 95744 18806 95750 18838
rect 95336 18768 95412 18774
rect 95749 18774 95750 18806
rect 95814 18806 95820 18838
rect 96560 19182 96566 19214
rect 96630 19214 96631 19246
rect 98328 19246 98404 19252
rect 96630 19182 96636 19214
rect 96560 18838 96636 19182
rect 95814 18774 95815 18806
rect 95749 18773 95815 18774
rect 96560 18774 96566 18838
rect 96630 18774 96636 18838
rect 98328 19182 98334 19246
rect 98398 19182 98404 19246
rect 99149 19246 99215 19247
rect 99149 19214 99150 19246
rect 98328 18838 98404 19182
rect 98328 18806 98334 18838
rect 96560 18768 96636 18774
rect 98333 18774 98334 18806
rect 98398 18806 98404 18838
rect 99144 19182 99150 19214
rect 99214 19214 99215 19246
rect 99552 19246 99628 19252
rect 99214 19182 99220 19214
rect 99144 18838 99220 19182
rect 98398 18774 98399 18806
rect 98333 18773 98399 18774
rect 99144 18774 99150 18838
rect 99214 18774 99220 18838
rect 99552 19182 99558 19246
rect 99622 19182 99628 19246
rect 100373 19246 100439 19247
rect 100373 19214 100374 19246
rect 99552 18838 99628 19182
rect 99552 18806 99558 18838
rect 99144 18768 99220 18774
rect 99557 18774 99558 18806
rect 99622 18806 99628 18838
rect 100368 19182 100374 19214
rect 100438 19214 100439 19246
rect 101597 19246 101663 19247
rect 101597 19214 101598 19246
rect 100438 19182 100444 19214
rect 100368 18838 100444 19182
rect 99622 18774 99623 18806
rect 99557 18773 99623 18774
rect 100368 18774 100374 18838
rect 100438 18774 100444 18838
rect 100368 18768 100444 18774
rect 101592 19182 101598 19214
rect 101662 19214 101663 19246
rect 102000 19246 102076 19252
rect 101662 19182 101668 19214
rect 101592 18838 101668 19182
rect 101592 18774 101598 18838
rect 101662 18774 101668 18838
rect 102000 19182 102006 19246
rect 102070 19182 102076 19246
rect 102000 18838 102076 19182
rect 102000 18806 102006 18838
rect 101592 18768 101668 18774
rect 102005 18774 102006 18806
rect 102070 18806 102076 18838
rect 102952 18838 103028 19318
rect 104045 19246 104111 19247
rect 104045 19214 104046 19246
rect 102952 18806 102958 18838
rect 102070 18774 102071 18806
rect 102005 18773 102071 18774
rect 102957 18774 102958 18806
rect 103022 18806 103028 18838
rect 104040 19182 104046 19214
rect 104110 19214 104111 19246
rect 104584 19246 104660 19252
rect 104110 19182 104116 19214
rect 104040 18838 104116 19182
rect 103022 18774 103023 18806
rect 102957 18773 103023 18774
rect 104040 18774 104046 18838
rect 104110 18774 104116 18838
rect 104584 19182 104590 19246
rect 104654 19182 104660 19246
rect 105269 19246 105335 19247
rect 105269 19214 105270 19246
rect 104584 18838 104660 19182
rect 104584 18806 104590 18838
rect 104040 18768 104116 18774
rect 104589 18774 104590 18806
rect 104654 18806 104660 18838
rect 105264 19182 105270 19214
rect 105334 19214 105335 19246
rect 105808 19246 105884 19252
rect 105334 19182 105340 19214
rect 105264 18838 105340 19182
rect 104654 18774 104655 18806
rect 104589 18773 104655 18774
rect 105264 18774 105270 18838
rect 105334 18774 105340 18838
rect 105808 19182 105814 19246
rect 105878 19182 105884 19246
rect 106629 19246 106695 19247
rect 106629 19214 106630 19246
rect 105808 18838 105884 19182
rect 105808 18806 105814 18838
rect 105264 18768 105340 18774
rect 105813 18774 105814 18806
rect 105878 18806 105884 18838
rect 106624 19182 106630 19214
rect 106694 19214 106695 19246
rect 107032 19246 107108 19252
rect 106694 19182 106700 19214
rect 106624 18838 106700 19182
rect 105878 18774 105879 18806
rect 105813 18773 105879 18774
rect 106624 18774 106630 18838
rect 106694 18774 106700 18838
rect 107032 19182 107038 19246
rect 107102 19182 107108 19246
rect 107032 18838 107108 19182
rect 107032 18806 107038 18838
rect 106624 18768 106700 18774
rect 107037 18774 107038 18806
rect 107102 18806 107108 18838
rect 108256 19246 108332 19252
rect 108256 19182 108262 19246
rect 108326 19182 108332 19246
rect 109077 19246 109143 19247
rect 109077 19214 109078 19246
rect 108256 18838 108332 19182
rect 108256 18806 108262 18838
rect 107102 18774 107103 18806
rect 107037 18773 107103 18774
rect 108261 18774 108262 18806
rect 108326 18806 108332 18838
rect 109072 19182 109078 19214
rect 109142 19214 109143 19246
rect 109142 19182 109148 19214
rect 109072 18838 109148 19182
rect 108326 18774 108327 18806
rect 108261 18773 108327 18774
rect 109072 18774 109078 18838
rect 109142 18774 109148 18838
rect 109072 18768 109148 18774
rect 77117 18702 77183 18703
rect 77117 18670 77118 18702
rect 77112 18638 77118 18670
rect 77182 18670 77183 18702
rect 77182 18638 77188 18670
rect 23392 15814 23398 15846
rect 21150 14558 21151 14590
rect 21085 14557 21151 14558
rect 22173 14350 22239 14351
rect 22173 14318 22174 14350
rect 15232 13366 15238 13398
rect 15237 13334 15238 13366
rect 15302 13366 15308 13398
rect 22168 14286 22174 14318
rect 22238 14318 22239 14350
rect 22238 14286 22244 14318
rect 15302 13334 15303 13366
rect 15237 13333 15303 13334
rect 15096 12006 15102 12038
rect 15101 11974 15102 12006
rect 15166 12006 15172 12038
rect 15232 13262 15308 13268
rect 15232 13198 15238 13262
rect 15302 13198 15308 13262
rect 15166 11974 15167 12006
rect 15101 11973 15167 11974
rect 952 10342 1230 10406
rect 1294 10342 1300 10406
rect 952 8910 1300 10342
rect 15096 11766 15172 11772
rect 15096 11702 15102 11766
rect 15166 11702 15172 11766
rect 15096 9182 15172 11702
rect 15232 10542 15308 13198
rect 22168 11766 22244 14286
rect 22304 13126 22380 15782
rect 23397 15782 23398 15814
rect 23462 15814 23468 15846
rect 29920 17070 29996 17076
rect 29920 17006 29926 17070
rect 29990 17006 29996 17070
rect 23462 15782 23463 15814
rect 23397 15781 23463 15782
rect 29920 15166 29996 17006
rect 32640 17070 32716 17076
rect 32640 17006 32646 17070
rect 32710 17006 32716 17070
rect 29920 15134 29926 15166
rect 29925 15102 29926 15134
rect 29990 15134 29996 15166
rect 30056 15166 30132 15172
rect 29990 15102 29991 15134
rect 29925 15101 29991 15102
rect 30056 15102 30062 15166
rect 30126 15102 30132 15166
rect 29925 14350 29991 14351
rect 29925 14318 29926 14350
rect 29920 14286 29926 14318
rect 29990 14318 29991 14350
rect 29990 14286 29996 14318
rect 29920 13670 29996 14286
rect 29920 13606 29926 13670
rect 29990 13606 29996 13670
rect 29920 13600 29996 13606
rect 29920 13534 29996 13540
rect 29920 13470 29926 13534
rect 29990 13470 29996 13534
rect 22304 13094 22310 13126
rect 22309 13062 22310 13094
rect 22374 13094 22380 13126
rect 28973 13126 29039 13127
rect 28973 13094 28974 13126
rect 22374 13062 22375 13094
rect 22309 13061 22375 13062
rect 28968 13062 28974 13094
rect 29038 13094 29039 13126
rect 29038 13062 29044 13094
rect 22168 11702 22174 11766
rect 22238 11702 22244 11766
rect 22168 11696 22244 11702
rect 15232 10510 15238 10542
rect 15237 10478 15238 10510
rect 15302 10510 15308 10542
rect 15302 10478 15303 10510
rect 15237 10477 15303 10478
rect 15237 10406 15303 10407
rect 15237 10374 15238 10406
rect 15096 9150 15102 9182
rect 15101 9118 15102 9150
rect 15166 9150 15172 9182
rect 15232 10342 15238 10374
rect 15302 10374 15303 10406
rect 15302 10342 15308 10374
rect 15166 9118 15167 9150
rect 15101 9117 15167 9118
rect 952 8846 1230 8910
rect 1294 8846 1300 8910
rect 952 7006 1300 8846
rect 15232 7686 15308 10342
rect 16869 9046 16935 9047
rect 16869 9014 16870 9046
rect 15232 7622 15238 7686
rect 15302 7622 15308 7686
rect 15232 7616 15308 7622
rect 16864 8982 16870 9014
rect 16934 9014 16935 9046
rect 16934 8982 16940 9014
rect 952 6942 1230 7006
rect 1294 6942 1300 7006
rect 952 5510 1300 6942
rect 952 5446 1230 5510
rect 1294 5446 1300 5510
rect 952 3878 1300 5446
rect 952 3814 1230 3878
rect 1294 3814 1300 3878
rect 952 1294 1300 3814
rect 16864 3878 16940 8982
rect 16864 3814 16870 3878
rect 16934 3814 16940 3878
rect 16864 3808 16940 3814
rect 16597 2926 16663 2927
rect 16597 2894 16598 2926
rect 16592 2862 16598 2894
rect 16662 2894 16663 2926
rect 17685 2926 17751 2927
rect 17685 2894 17686 2926
rect 16662 2862 16668 2894
rect 2045 1702 2111 1703
rect 2045 1670 2046 1702
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 1300 1294
rect 952 1158 1300 1230
rect 2040 1638 2046 1670
rect 2110 1670 2111 1702
rect 3813 1702 3879 1703
rect 3813 1670 3814 1702
rect 2110 1638 2116 1670
rect 2040 1294 2116 1638
rect 2040 1230 2046 1294
rect 2110 1230 2116 1294
rect 2040 1224 2116 1230
rect 3808 1638 3814 1670
rect 3878 1670 3879 1702
rect 5445 1702 5511 1703
rect 5445 1670 5446 1702
rect 3878 1638 3884 1670
rect 3808 1294 3884 1638
rect 3808 1230 3814 1294
rect 3878 1230 3884 1294
rect 3808 1224 3884 1230
rect 5440 1638 5446 1670
rect 5510 1670 5511 1702
rect 7213 1702 7279 1703
rect 7213 1670 7214 1702
rect 5510 1638 5516 1670
rect 5440 1294 5516 1638
rect 5440 1230 5446 1294
rect 5510 1230 5516 1294
rect 5440 1224 5516 1230
rect 7208 1638 7214 1670
rect 7278 1670 7279 1702
rect 8709 1702 8775 1703
rect 8709 1670 8710 1702
rect 7278 1638 7284 1670
rect 7208 1294 7284 1638
rect 7208 1230 7214 1294
rect 7278 1230 7284 1294
rect 7208 1224 7284 1230
rect 8704 1638 8710 1670
rect 8774 1670 8775 1702
rect 10477 1702 10543 1703
rect 10477 1670 10478 1702
rect 8774 1638 8780 1670
rect 8704 1294 8780 1638
rect 8704 1230 8710 1294
rect 8774 1230 8780 1294
rect 8704 1224 8780 1230
rect 10472 1638 10478 1670
rect 10542 1670 10543 1702
rect 12109 1702 12175 1703
rect 12109 1670 12110 1702
rect 10542 1638 10548 1670
rect 10472 1294 10548 1638
rect 10472 1230 10478 1294
rect 10542 1230 10548 1294
rect 10472 1224 10548 1230
rect 12104 1638 12110 1670
rect 12174 1670 12175 1702
rect 13877 1702 13943 1703
rect 13877 1670 13878 1702
rect 12174 1638 12180 1670
rect 12104 1294 12180 1638
rect 12104 1230 12110 1294
rect 12174 1230 12180 1294
rect 12104 1224 12180 1230
rect 13872 1638 13878 1670
rect 13942 1670 13943 1702
rect 15645 1702 15711 1703
rect 15645 1670 15646 1702
rect 13942 1638 13948 1670
rect 13872 1294 13948 1638
rect 13872 1230 13878 1294
rect 13942 1230 13948 1294
rect 13872 1224 13948 1230
rect 15640 1638 15646 1670
rect 15710 1670 15711 1702
rect 15710 1638 15716 1670
rect 15640 1294 15716 1638
rect 15640 1230 15646 1294
rect 15710 1230 15716 1294
rect 15640 1224 15716 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 1300 1158
rect 952 1022 1300 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 1300 1022
rect 952 952 1300 958
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 620 614
rect 272 478 620 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 620 478
rect 272 342 620 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 620 342
rect 272 272 620 278
rect 16592 0 16668 2862
rect 17680 2862 17686 2894
rect 17750 2894 17751 2926
rect 18773 2926 18839 2927
rect 18773 2894 18774 2926
rect 17750 2862 17756 2894
rect 17141 1702 17207 1703
rect 17141 1670 17142 1702
rect 17136 1638 17142 1670
rect 17206 1670 17207 1702
rect 17206 1638 17212 1670
rect 17136 1294 17212 1638
rect 17136 1230 17142 1294
rect 17206 1230 17212 1294
rect 17136 1224 17212 1230
rect 17680 0 17756 2862
rect 18768 2862 18774 2894
rect 18838 2894 18839 2926
rect 20133 2926 20199 2927
rect 20133 2894 20134 2926
rect 18838 2862 18844 2894
rect 18768 0 18844 2862
rect 20128 2862 20134 2894
rect 20198 2894 20199 2926
rect 21085 2926 21151 2927
rect 21085 2894 21086 2926
rect 20198 2862 20204 2894
rect 19317 2382 19383 2383
rect 19317 2350 19318 2382
rect 19312 2318 19318 2350
rect 19382 2350 19383 2382
rect 19382 2318 19388 2350
rect 19045 1702 19111 1703
rect 19045 1670 19046 1702
rect 19040 1638 19046 1670
rect 19110 1670 19111 1702
rect 19110 1638 19116 1670
rect 19040 1294 19116 1638
rect 19040 1230 19046 1294
rect 19110 1230 19116 1294
rect 19040 1224 19116 1230
rect 19312 614 19388 2318
rect 19312 550 19318 614
rect 19382 550 19388 614
rect 19312 544 19388 550
rect 20128 0 20204 2862
rect 21080 2862 21086 2894
rect 21150 2894 21151 2926
rect 22309 2926 22375 2927
rect 22309 2894 22310 2926
rect 21150 2862 21156 2894
rect 20541 1702 20607 1703
rect 20541 1670 20542 1702
rect 20536 1638 20542 1670
rect 20606 1670 20607 1702
rect 20606 1638 20612 1670
rect 20536 1294 20612 1638
rect 20536 1230 20542 1294
rect 20606 1230 20612 1294
rect 20536 1224 20612 1230
rect 21080 0 21156 2862
rect 22304 2862 22310 2894
rect 22374 2894 22375 2926
rect 23669 2926 23735 2927
rect 23669 2894 23670 2926
rect 22374 2862 22380 2894
rect 22173 1702 22239 1703
rect 22173 1670 22174 1702
rect 22168 1638 22174 1670
rect 22238 1670 22239 1702
rect 22238 1638 22244 1670
rect 22168 1294 22244 1638
rect 22168 1230 22174 1294
rect 22238 1230 22244 1294
rect 22168 1224 22244 1230
rect 22304 0 22380 2862
rect 23664 2862 23670 2894
rect 23734 2894 23735 2926
rect 24757 2926 24823 2927
rect 24757 2894 24758 2926
rect 23734 2862 23740 2894
rect 23664 0 23740 2862
rect 24752 2862 24758 2894
rect 24822 2894 24823 2926
rect 25981 2926 26047 2927
rect 25981 2894 25982 2926
rect 24822 2862 24828 2894
rect 23941 1702 24007 1703
rect 23941 1670 23942 1702
rect 23936 1638 23942 1670
rect 24006 1670 24007 1702
rect 24006 1638 24012 1670
rect 23936 1294 24012 1638
rect 23936 1230 23942 1294
rect 24006 1230 24012 1294
rect 23936 1224 24012 1230
rect 24752 0 24828 2862
rect 25976 2862 25982 2894
rect 26046 2894 26047 2926
rect 27069 2926 27135 2927
rect 27069 2894 27070 2926
rect 26046 2862 26052 2894
rect 25709 1702 25775 1703
rect 25709 1670 25710 1702
rect 25704 1638 25710 1670
rect 25774 1670 25775 1702
rect 25774 1638 25780 1670
rect 25704 1294 25780 1638
rect 25704 1230 25710 1294
rect 25774 1230 25780 1294
rect 25704 1224 25780 1230
rect 25976 0 26052 2862
rect 27064 2862 27070 2894
rect 27134 2894 27135 2926
rect 28157 2926 28223 2927
rect 28157 2894 28158 2926
rect 27134 2862 27140 2894
rect 27064 0 27140 2862
rect 28152 2862 28158 2894
rect 28222 2894 28223 2926
rect 28222 2862 28228 2894
rect 27205 1702 27271 1703
rect 27205 1670 27206 1702
rect 27200 1638 27206 1670
rect 27270 1670 27271 1702
rect 27270 1638 27276 1670
rect 27200 1294 27276 1638
rect 27200 1230 27206 1294
rect 27270 1230 27276 1294
rect 27200 1224 27276 1230
rect 28152 0 28228 2862
rect 28837 1702 28903 1703
rect 28837 1670 28838 1702
rect 28832 1638 28838 1670
rect 28902 1670 28903 1702
rect 28902 1638 28908 1670
rect 28832 1294 28908 1638
rect 28832 1230 28838 1294
rect 28902 1230 28908 1294
rect 28832 1224 28908 1230
rect 28968 0 29044 13062
rect 29789 12310 29855 12311
rect 29789 12278 29790 12310
rect 29784 12246 29790 12278
rect 29854 12278 29855 12310
rect 29854 12246 29860 12278
rect 29653 11902 29719 11903
rect 29653 11870 29654 11902
rect 29648 11838 29654 11870
rect 29718 11870 29719 11902
rect 29718 11838 29724 11870
rect 29240 11358 29316 11364
rect 29240 11294 29246 11358
rect 29310 11294 29316 11358
rect 29240 9590 29316 11294
rect 29512 11086 29588 11092
rect 29512 11022 29518 11086
rect 29582 11022 29588 11086
rect 29512 10678 29588 11022
rect 29648 11086 29724 11838
rect 29784 11766 29860 12246
rect 29920 12038 29996 13470
rect 30056 13262 30132 15102
rect 32504 15166 32580 15172
rect 32504 15102 32510 15166
rect 32574 15102 32580 15166
rect 32640 15166 32716 17006
rect 35088 17070 35164 17076
rect 35088 17006 35094 17070
rect 35158 17006 35164 17070
rect 32640 15134 32646 15166
rect 32373 14350 32439 14351
rect 32373 14318 32374 14350
rect 32368 14286 32374 14318
rect 32438 14318 32439 14350
rect 32438 14286 32444 14318
rect 32368 13670 32444 14286
rect 32368 13606 32374 13670
rect 32438 13606 32444 13670
rect 32368 13600 32444 13606
rect 30056 13230 30062 13262
rect 30061 13198 30062 13230
rect 30126 13230 30132 13262
rect 32368 13534 32444 13540
rect 32368 13470 32374 13534
rect 32438 13470 32444 13534
rect 30126 13198 30127 13230
rect 30061 13197 30127 13198
rect 30056 13126 30132 13132
rect 30056 13062 30062 13126
rect 30126 13062 30132 13126
rect 31965 13126 32031 13127
rect 31965 13094 31966 13126
rect 30056 12582 30132 13062
rect 30056 12550 30062 12582
rect 30061 12518 30062 12550
rect 30126 12550 30132 12582
rect 31960 13062 31966 13094
rect 32030 13094 32031 13126
rect 32030 13062 32036 13094
rect 30126 12518 30127 12550
rect 30061 12517 30127 12518
rect 29920 12006 29926 12038
rect 29925 11974 29926 12006
rect 29990 12006 29996 12038
rect 29990 11974 29991 12006
rect 29925 11973 29991 11974
rect 29784 11702 29790 11766
rect 29854 11702 29860 11766
rect 29784 11696 29860 11702
rect 29648 11022 29654 11086
rect 29718 11022 29724 11086
rect 29648 11016 29724 11022
rect 29512 10646 29518 10678
rect 29517 10614 29518 10646
rect 29582 10646 29588 10678
rect 29582 10614 29583 10646
rect 29517 10613 29583 10614
rect 29240 9558 29246 9590
rect 29245 9526 29246 9558
rect 29310 9558 29316 9590
rect 29310 9526 29311 9558
rect 29245 9525 29311 9526
rect 29245 2926 29311 2927
rect 29245 2894 29246 2926
rect 29240 2862 29246 2894
rect 29310 2894 29311 2926
rect 30605 2926 30671 2927
rect 30605 2894 30606 2926
rect 29310 2862 29316 2894
rect 29240 0 29316 2862
rect 30600 2862 30606 2894
rect 30670 2894 30671 2926
rect 31829 2926 31895 2927
rect 31829 2894 31830 2926
rect 30670 2862 30676 2894
rect 30469 1702 30535 1703
rect 30469 1670 30470 1702
rect 30464 1638 30470 1670
rect 30534 1670 30535 1702
rect 30534 1638 30540 1670
rect 30464 1294 30540 1638
rect 30464 1230 30470 1294
rect 30534 1230 30540 1294
rect 30464 1224 30540 1230
rect 30600 0 30676 2862
rect 31824 2862 31830 2894
rect 31894 2894 31895 2926
rect 31894 2862 31900 2894
rect 31824 0 31900 2862
rect 31960 0 32036 13062
rect 32237 12310 32303 12311
rect 32237 12278 32238 12310
rect 32232 12246 32238 12278
rect 32302 12278 32303 12310
rect 32302 12246 32308 12278
rect 32101 11902 32167 11903
rect 32101 11870 32102 11902
rect 32096 11838 32102 11870
rect 32166 11870 32167 11902
rect 32166 11838 32172 11870
rect 32096 11086 32172 11838
rect 32232 11766 32308 12246
rect 32368 12038 32444 13470
rect 32504 13262 32580 15102
rect 32645 15102 32646 15134
rect 32710 15134 32716 15166
rect 34952 15166 35028 15172
rect 32710 15102 32711 15134
rect 32645 15101 32711 15102
rect 34952 15102 34958 15166
rect 35022 15102 35028 15166
rect 35088 15166 35164 17006
rect 35088 15134 35094 15166
rect 34821 14350 34887 14351
rect 34821 14318 34822 14350
rect 34816 14286 34822 14318
rect 34886 14318 34887 14350
rect 34886 14286 34892 14318
rect 32504 13230 32510 13262
rect 32509 13198 32510 13230
rect 32574 13230 32580 13262
rect 34680 13670 34756 13676
rect 34680 13606 34686 13670
rect 34750 13606 34756 13670
rect 32574 13198 32575 13230
rect 32509 13197 32575 13198
rect 32504 13126 32580 13132
rect 32504 13062 32510 13126
rect 32574 13062 32580 13126
rect 34413 13126 34479 13127
rect 34413 13094 34414 13126
rect 32504 12582 32580 13062
rect 32504 12550 32510 12582
rect 32509 12518 32510 12550
rect 32574 12550 32580 12582
rect 34408 13062 34414 13094
rect 34478 13094 34479 13126
rect 34478 13062 34484 13094
rect 32574 12518 32575 12550
rect 32509 12517 32575 12518
rect 32368 12006 32374 12038
rect 32373 11974 32374 12006
rect 32438 12006 32444 12038
rect 32438 11974 32439 12006
rect 32373 11973 32439 11974
rect 32232 11702 32238 11766
rect 32302 11702 32308 11766
rect 32232 11696 32308 11702
rect 32096 11022 32102 11086
rect 32166 11022 32172 11086
rect 32096 11016 32172 11022
rect 32917 2926 32983 2927
rect 32917 2894 32918 2926
rect 32912 2862 32918 2894
rect 32982 2894 32983 2926
rect 34005 2926 34071 2927
rect 34005 2894 34006 2926
rect 32982 2862 32988 2894
rect 32237 1702 32303 1703
rect 32237 1670 32238 1702
rect 32232 1638 32238 1670
rect 32302 1670 32303 1702
rect 32302 1638 32308 1670
rect 32232 1294 32308 1638
rect 32232 1230 32238 1294
rect 32302 1230 32308 1294
rect 32232 1224 32308 1230
rect 32912 0 32988 2862
rect 34000 2862 34006 2894
rect 34070 2894 34071 2926
rect 34070 2862 34076 2894
rect 34000 0 34076 2862
rect 34277 1702 34343 1703
rect 34277 1670 34278 1702
rect 34272 1638 34278 1670
rect 34342 1670 34343 1702
rect 34342 1638 34348 1670
rect 34272 1294 34348 1638
rect 34272 1230 34278 1294
rect 34342 1230 34348 1294
rect 34272 1224 34348 1230
rect 34408 0 34484 13062
rect 34680 12038 34756 13606
rect 34816 13670 34892 14286
rect 34816 13606 34822 13670
rect 34886 13606 34892 13670
rect 34816 13600 34892 13606
rect 34816 13126 34892 13132
rect 34816 13062 34822 13126
rect 34886 13062 34892 13126
rect 34952 13126 35028 15102
rect 35093 15102 35094 15134
rect 35158 15134 35164 15166
rect 37400 17070 37476 17076
rect 37400 17006 37406 17070
rect 37470 17006 37476 17070
rect 37400 15166 37476 17006
rect 40120 17070 40196 17076
rect 40120 17006 40126 17070
rect 40190 17006 40196 17070
rect 37400 15134 37406 15166
rect 35158 15102 35159 15134
rect 35093 15101 35159 15102
rect 37405 15102 37406 15134
rect 37470 15134 37476 15166
rect 37536 15166 37612 15172
rect 37470 15102 37471 15134
rect 37405 15101 37471 15102
rect 37536 15102 37542 15166
rect 37606 15102 37612 15166
rect 37405 14350 37471 14351
rect 37405 14318 37406 14350
rect 37400 14286 37406 14318
rect 37470 14318 37471 14350
rect 37470 14286 37476 14318
rect 37400 13670 37476 14286
rect 37400 13606 37406 13670
rect 37470 13606 37476 13670
rect 37400 13600 37476 13606
rect 37264 13534 37340 13540
rect 37264 13470 37270 13534
rect 37334 13470 37340 13534
rect 34952 13094 34958 13126
rect 34816 12582 34892 13062
rect 34957 13062 34958 13094
rect 35022 13094 35028 13126
rect 36997 13126 37063 13127
rect 36997 13094 36998 13126
rect 35022 13062 35023 13094
rect 34957 13061 35023 13062
rect 36992 13062 36998 13094
rect 37062 13094 37063 13126
rect 37062 13062 37068 13094
rect 34816 12550 34822 12582
rect 34821 12518 34822 12550
rect 34886 12550 34892 12582
rect 34886 12518 34887 12550
rect 34821 12517 34887 12518
rect 34821 12310 34887 12311
rect 34821 12278 34822 12310
rect 34680 12006 34686 12038
rect 34685 11974 34686 12006
rect 34750 12006 34756 12038
rect 34816 12246 34822 12278
rect 34886 12278 34887 12310
rect 34886 12246 34892 12278
rect 34750 11974 34751 12006
rect 34685 11973 34751 11974
rect 34685 11902 34751 11903
rect 34685 11870 34686 11902
rect 34680 11838 34686 11870
rect 34750 11870 34751 11902
rect 34750 11838 34756 11870
rect 34680 11086 34756 11838
rect 34816 11766 34892 12246
rect 34816 11702 34822 11766
rect 34886 11702 34892 11766
rect 34816 11696 34892 11702
rect 34680 11022 34686 11086
rect 34750 11022 34756 11086
rect 34680 11016 34756 11022
rect 36725 3742 36791 3743
rect 36725 3710 36726 3742
rect 36720 3678 36726 3710
rect 36790 3710 36791 3742
rect 36790 3678 36796 3710
rect 35093 2926 35159 2927
rect 35093 2894 35094 2926
rect 35088 2862 35094 2894
rect 35158 2894 35159 2926
rect 36453 2926 36519 2927
rect 36453 2894 36454 2926
rect 35158 2862 35164 2894
rect 35088 0 35164 2862
rect 36448 2862 36454 2894
rect 36518 2894 36519 2926
rect 36518 2862 36524 2894
rect 35637 1702 35703 1703
rect 35637 1670 35638 1702
rect 35632 1638 35638 1670
rect 35702 1670 35703 1702
rect 35702 1638 35708 1670
rect 35632 1294 35708 1638
rect 35632 1230 35638 1294
rect 35702 1230 35708 1294
rect 35632 1224 35708 1230
rect 36448 0 36524 2862
rect 36720 1838 36796 3678
rect 36720 1774 36726 1838
rect 36790 1774 36796 1838
rect 36720 1768 36796 1774
rect 36992 0 37068 13062
rect 37264 12038 37340 13470
rect 37536 13262 37612 15102
rect 39984 15166 40060 15172
rect 39984 15102 39990 15166
rect 40054 15102 40060 15166
rect 40120 15166 40196 17006
rect 40120 15134 40126 15166
rect 39853 14350 39919 14351
rect 39853 14318 39854 14350
rect 39848 14286 39854 14318
rect 39918 14318 39919 14350
rect 39918 14286 39924 14318
rect 39848 13670 39924 14286
rect 39848 13606 39854 13670
rect 39918 13606 39924 13670
rect 39848 13600 39924 13606
rect 37536 13230 37542 13262
rect 37541 13198 37542 13230
rect 37606 13230 37612 13262
rect 39712 13534 39788 13540
rect 39712 13470 39718 13534
rect 39782 13470 39788 13534
rect 37606 13198 37607 13230
rect 37541 13197 37607 13198
rect 37400 13126 37476 13132
rect 37400 13062 37406 13126
rect 37470 13062 37476 13126
rect 39445 13126 39511 13127
rect 39445 13094 39446 13126
rect 37400 12582 37476 13062
rect 37400 12550 37406 12582
rect 37405 12518 37406 12550
rect 37470 12550 37476 12582
rect 39440 13062 39446 13094
rect 39510 13094 39511 13126
rect 39510 13062 39516 13094
rect 37470 12518 37471 12550
rect 37405 12517 37471 12518
rect 37405 12310 37471 12311
rect 37405 12278 37406 12310
rect 37264 12006 37270 12038
rect 37269 11974 37270 12006
rect 37334 12006 37340 12038
rect 37400 12246 37406 12278
rect 37470 12278 37471 12310
rect 37470 12246 37476 12278
rect 37334 11974 37335 12006
rect 37269 11973 37335 11974
rect 37269 11902 37335 11903
rect 37269 11870 37270 11902
rect 37264 11838 37270 11870
rect 37334 11870 37335 11902
rect 37334 11838 37340 11870
rect 37264 11086 37340 11838
rect 37400 11766 37476 12246
rect 37400 11702 37406 11766
rect 37470 11702 37476 11766
rect 37400 11696 37476 11702
rect 37264 11022 37270 11086
rect 37334 11022 37340 11086
rect 37264 11016 37340 11022
rect 37541 2926 37607 2927
rect 37541 2894 37542 2926
rect 37536 2862 37542 2894
rect 37606 2894 37607 2926
rect 38629 2926 38695 2927
rect 38629 2894 38630 2926
rect 37606 2862 37612 2894
rect 37269 1702 37335 1703
rect 37269 1670 37270 1702
rect 37264 1638 37270 1670
rect 37334 1670 37335 1702
rect 37334 1638 37340 1670
rect 37264 1294 37340 1638
rect 37264 1230 37270 1294
rect 37334 1230 37340 1294
rect 37264 1224 37340 1230
rect 37536 0 37612 2862
rect 38624 2862 38630 2894
rect 38694 2894 38695 2926
rect 38694 2862 38700 2894
rect 38624 0 38700 2862
rect 39037 1702 39103 1703
rect 39037 1670 39038 1702
rect 39032 1638 39038 1670
rect 39102 1670 39103 1702
rect 39102 1638 39108 1670
rect 39032 1294 39108 1638
rect 39032 1230 39038 1294
rect 39102 1230 39108 1294
rect 39032 1224 39108 1230
rect 39440 0 39516 13062
rect 39712 12038 39788 13470
rect 39984 13262 40060 15102
rect 40125 15102 40126 15134
rect 40190 15134 40196 15166
rect 42432 17070 42508 17076
rect 42432 17006 42438 17070
rect 42502 17006 42508 17070
rect 42432 15166 42508 17006
rect 44880 17070 44956 17076
rect 44880 17006 44886 17070
rect 44950 17006 44956 17070
rect 42432 15134 42438 15166
rect 40190 15102 40191 15134
rect 40125 15101 40191 15102
rect 42437 15102 42438 15134
rect 42502 15134 42508 15166
rect 42568 15166 42644 15172
rect 42502 15102 42503 15134
rect 42437 15101 42503 15102
rect 42568 15102 42574 15166
rect 42638 15102 42644 15166
rect 44880 15166 44956 17006
rect 47600 17070 47676 17076
rect 47600 17006 47606 17070
rect 47670 17006 47676 17070
rect 44880 15134 44886 15166
rect 42165 14350 42231 14351
rect 42165 14318 42166 14350
rect 42160 14286 42166 14318
rect 42230 14318 42231 14350
rect 42230 14286 42236 14318
rect 42160 13670 42236 14286
rect 42160 13606 42166 13670
rect 42230 13606 42236 13670
rect 42160 13600 42236 13606
rect 39984 13230 39990 13262
rect 39989 13198 39990 13230
rect 40054 13230 40060 13262
rect 42432 13534 42508 13540
rect 42432 13470 42438 13534
rect 42502 13470 42508 13534
rect 40054 13198 40055 13230
rect 39989 13197 40055 13198
rect 39848 13126 39924 13132
rect 39848 13062 39854 13126
rect 39918 13062 39924 13126
rect 41757 13126 41823 13127
rect 41757 13094 41758 13126
rect 39848 12582 39924 13062
rect 39848 12550 39854 12582
rect 39853 12518 39854 12550
rect 39918 12550 39924 12582
rect 41752 13062 41758 13094
rect 41822 13094 41823 13126
rect 42296 13126 42372 13132
rect 41822 13062 41828 13094
rect 39918 12518 39919 12550
rect 39853 12517 39919 12518
rect 39853 12310 39919 12311
rect 39853 12278 39854 12310
rect 39712 12006 39718 12038
rect 39717 11974 39718 12006
rect 39782 12006 39788 12038
rect 39848 12246 39854 12278
rect 39918 12278 39919 12310
rect 39918 12246 39924 12278
rect 39782 11974 39783 12006
rect 39717 11973 39783 11974
rect 39717 11902 39783 11903
rect 39717 11870 39718 11902
rect 39712 11838 39718 11870
rect 39782 11870 39783 11902
rect 39782 11838 39788 11870
rect 39712 11086 39788 11838
rect 39848 11766 39924 12246
rect 39848 11702 39854 11766
rect 39918 11702 39924 11766
rect 39848 11696 39924 11702
rect 39712 11022 39718 11086
rect 39782 11022 39788 11086
rect 39712 11016 39788 11022
rect 39989 2926 40055 2927
rect 39989 2894 39990 2926
rect 39984 2862 39990 2894
rect 40054 2894 40055 2926
rect 41213 2926 41279 2927
rect 41213 2894 41214 2926
rect 40054 2862 40060 2894
rect 39984 0 40060 2862
rect 41208 2862 41214 2894
rect 41278 2894 41279 2926
rect 41278 2862 41284 2894
rect 40669 1702 40735 1703
rect 40669 1670 40670 1702
rect 40664 1638 40670 1670
rect 40734 1670 40735 1702
rect 40734 1638 40740 1670
rect 40664 1294 40740 1638
rect 40664 1230 40670 1294
rect 40734 1230 40740 1294
rect 40664 1224 40740 1230
rect 41208 0 41284 2862
rect 41752 0 41828 13062
rect 42296 13062 42302 13126
rect 42366 13062 42372 13126
rect 42296 12582 42372 13062
rect 42296 12550 42302 12582
rect 42301 12518 42302 12550
rect 42366 12550 42372 12582
rect 42366 12518 42367 12550
rect 42301 12517 42367 12518
rect 42165 12310 42231 12311
rect 42165 12278 42166 12310
rect 42160 12246 42166 12278
rect 42230 12278 42231 12310
rect 42230 12246 42236 12278
rect 42160 11766 42236 12246
rect 42432 12038 42508 13470
rect 42568 13262 42644 15102
rect 44885 15102 44886 15134
rect 44950 15134 44956 15166
rect 45016 15166 45092 15172
rect 44950 15102 44951 15134
rect 44885 15101 44951 15102
rect 45016 15102 45022 15166
rect 45086 15102 45092 15166
rect 44885 14350 44951 14351
rect 44885 14318 44886 14350
rect 44880 14286 44886 14318
rect 44950 14318 44951 14350
rect 44950 14286 44956 14318
rect 44880 13670 44956 14286
rect 44880 13606 44886 13670
rect 44950 13606 44956 13670
rect 44880 13600 44956 13606
rect 42568 13230 42574 13262
rect 42573 13198 42574 13230
rect 42638 13230 42644 13262
rect 44880 13534 44956 13540
rect 44880 13470 44886 13534
rect 44950 13470 44956 13534
rect 42638 13198 42639 13230
rect 42573 13197 42639 13198
rect 44205 13126 44271 13127
rect 44205 13094 44206 13126
rect 42432 12006 42438 12038
rect 42437 11974 42438 12006
rect 42502 12006 42508 12038
rect 44200 13062 44206 13094
rect 44270 13094 44271 13126
rect 44270 13062 44276 13094
rect 42502 11974 42503 12006
rect 42437 11973 42503 11974
rect 42301 11902 42367 11903
rect 42301 11870 42302 11902
rect 42160 11702 42166 11766
rect 42230 11702 42236 11766
rect 42160 11696 42236 11702
rect 42296 11838 42302 11870
rect 42366 11870 42367 11902
rect 42366 11838 42372 11870
rect 42296 11086 42372 11838
rect 42296 11022 42302 11086
rect 42366 11022 42372 11086
rect 42296 11016 42372 11022
rect 42301 2926 42367 2927
rect 42301 2894 42302 2926
rect 42296 2862 42302 2894
rect 42366 2894 42367 2926
rect 43389 2926 43455 2927
rect 43389 2894 43390 2926
rect 42366 2862 42372 2894
rect 42296 0 42372 2862
rect 43384 2862 43390 2894
rect 43454 2894 43455 2926
rect 43454 2862 43460 2894
rect 42437 1702 42503 1703
rect 42437 1670 42438 1702
rect 42432 1638 42438 1670
rect 42502 1670 42503 1702
rect 42502 1638 42508 1670
rect 42432 1294 42508 1638
rect 42432 1230 42438 1294
rect 42502 1230 42508 1294
rect 42432 1224 42508 1230
rect 43384 0 43460 2862
rect 44069 1702 44135 1703
rect 44069 1670 44070 1702
rect 44064 1638 44070 1670
rect 44134 1670 44135 1702
rect 44134 1638 44140 1670
rect 44064 1294 44140 1638
rect 44064 1230 44070 1294
rect 44134 1230 44140 1294
rect 44064 1224 44140 1230
rect 44200 0 44276 13062
rect 44613 12310 44679 12311
rect 44613 12278 44614 12310
rect 44608 12246 44614 12278
rect 44678 12278 44679 12310
rect 44678 12246 44684 12278
rect 44608 11766 44684 12246
rect 44880 12038 44956 13470
rect 45016 13262 45092 15102
rect 47464 15166 47540 15172
rect 47464 15102 47470 15166
rect 47534 15102 47540 15166
rect 47600 15166 47676 17006
rect 47600 15134 47606 15166
rect 47197 14350 47263 14351
rect 47197 14318 47198 14350
rect 47192 14286 47198 14318
rect 47262 14318 47263 14350
rect 47262 14286 47268 14318
rect 47192 13670 47268 14286
rect 47192 13606 47198 13670
rect 47262 13606 47268 13670
rect 47192 13600 47268 13606
rect 45016 13230 45022 13262
rect 45021 13198 45022 13230
rect 45086 13230 45092 13262
rect 47328 13534 47404 13540
rect 47328 13470 47334 13534
rect 47398 13470 47404 13534
rect 45086 13198 45087 13230
rect 45021 13197 45087 13198
rect 45016 13126 45092 13132
rect 45016 13062 45022 13126
rect 45086 13062 45092 13126
rect 46517 13126 46583 13127
rect 46517 13094 46518 13126
rect 45016 12582 45092 13062
rect 45016 12550 45022 12582
rect 45021 12518 45022 12550
rect 45086 12550 45092 12582
rect 46512 13062 46518 13094
rect 46582 13094 46583 13126
rect 46582 13062 46588 13094
rect 45086 12518 45087 12550
rect 45021 12517 45087 12518
rect 44880 12006 44886 12038
rect 44885 11974 44886 12006
rect 44950 12006 44956 12038
rect 44950 11974 44951 12006
rect 44885 11973 44951 11974
rect 44749 11902 44815 11903
rect 44749 11870 44750 11902
rect 44608 11702 44614 11766
rect 44678 11702 44684 11766
rect 44608 11696 44684 11702
rect 44744 11838 44750 11870
rect 44814 11870 44815 11902
rect 44814 11838 44820 11870
rect 44744 11086 44820 11838
rect 44744 11022 44750 11086
rect 44814 11022 44820 11086
rect 44744 11016 44820 11022
rect 44477 2926 44543 2927
rect 44477 2894 44478 2926
rect 44472 2862 44478 2894
rect 44542 2894 44543 2926
rect 45837 2926 45903 2927
rect 45837 2894 45838 2926
rect 44542 2862 44548 2894
rect 44472 0 44548 2862
rect 45832 2862 45838 2894
rect 45902 2894 45903 2926
rect 45902 2862 45908 2894
rect 45701 1702 45767 1703
rect 45701 1670 45702 1702
rect 45696 1638 45702 1670
rect 45766 1670 45767 1702
rect 45766 1638 45772 1670
rect 45696 1294 45772 1638
rect 45696 1230 45702 1294
rect 45766 1230 45772 1294
rect 45696 1224 45772 1230
rect 45832 0 45908 2862
rect 46512 0 46588 13062
rect 47197 12310 47263 12311
rect 47197 12278 47198 12310
rect 47192 12246 47198 12278
rect 47262 12278 47263 12310
rect 47262 12246 47268 12278
rect 47061 11902 47127 11903
rect 47061 11870 47062 11902
rect 47056 11838 47062 11870
rect 47126 11870 47127 11902
rect 47126 11838 47132 11870
rect 47056 11086 47132 11838
rect 47192 11766 47268 12246
rect 47328 12038 47404 13470
rect 47464 13262 47540 15102
rect 47605 15102 47606 15134
rect 47670 15134 47676 15166
rect 49912 17070 49988 17076
rect 49912 17006 49918 17070
rect 49982 17006 49988 17070
rect 49912 15166 49988 17006
rect 52496 17070 52572 17076
rect 52496 17006 52502 17070
rect 52566 17006 52572 17070
rect 49912 15134 49918 15166
rect 47670 15102 47671 15134
rect 47605 15101 47671 15102
rect 49917 15102 49918 15134
rect 49982 15134 49988 15166
rect 50184 15166 50260 15172
rect 49982 15102 49983 15134
rect 49917 15101 49983 15102
rect 50184 15102 50190 15166
rect 50254 15102 50260 15166
rect 49781 14350 49847 14351
rect 49781 14318 49782 14350
rect 49776 14286 49782 14318
rect 49846 14318 49847 14350
rect 49846 14286 49852 14318
rect 47464 13230 47470 13262
rect 47469 13198 47470 13230
rect 47534 13230 47540 13262
rect 49640 13670 49716 13676
rect 49640 13606 49646 13670
rect 49710 13606 49716 13670
rect 47534 13198 47535 13230
rect 47469 13197 47535 13198
rect 47464 13126 47540 13132
rect 47464 13062 47470 13126
rect 47534 13062 47540 13126
rect 47464 12582 47540 13062
rect 47464 12550 47470 12582
rect 47469 12518 47470 12550
rect 47534 12550 47540 12582
rect 47534 12518 47535 12550
rect 47469 12517 47535 12518
rect 49509 12310 49575 12311
rect 49509 12278 49510 12310
rect 47328 12006 47334 12038
rect 47333 11974 47334 12006
rect 47398 12006 47404 12038
rect 49504 12246 49510 12278
rect 49574 12278 49575 12310
rect 49574 12246 49580 12278
rect 47398 11974 47399 12006
rect 47333 11973 47399 11974
rect 47192 11702 47198 11766
rect 47262 11702 47268 11766
rect 47192 11696 47268 11702
rect 49504 11766 49580 12246
rect 49640 12038 49716 13606
rect 49776 13670 49852 14286
rect 49776 13606 49782 13670
rect 49846 13606 49852 13670
rect 49776 13600 49852 13606
rect 49917 13398 49983 13399
rect 49917 13366 49918 13398
rect 49912 13334 49918 13366
rect 49982 13366 49983 13398
rect 49982 13334 49988 13366
rect 49776 13126 49852 13132
rect 49776 13062 49782 13126
rect 49846 13062 49852 13126
rect 49776 12582 49852 13062
rect 49776 12550 49782 12582
rect 49781 12518 49782 12550
rect 49846 12550 49852 12582
rect 49846 12518 49847 12550
rect 49781 12517 49847 12518
rect 49640 12006 49646 12038
rect 49645 11974 49646 12006
rect 49710 12006 49716 12038
rect 49710 11974 49711 12006
rect 49645 11973 49711 11974
rect 49781 11902 49847 11903
rect 49781 11870 49782 11902
rect 49504 11702 49510 11766
rect 49574 11702 49580 11766
rect 49504 11696 49580 11702
rect 49776 11838 49782 11870
rect 49846 11870 49847 11902
rect 49846 11838 49852 11870
rect 47056 11022 47062 11086
rect 47126 11022 47132 11086
rect 47056 11016 47132 11022
rect 49776 11086 49852 11838
rect 49776 11022 49782 11086
rect 49846 11022 49852 11086
rect 49776 11016 49852 11022
rect 46925 2926 46991 2927
rect 46925 2894 46926 2926
rect 46920 2862 46926 2894
rect 46990 2894 46991 2926
rect 48149 2926 48215 2927
rect 48149 2894 48150 2926
rect 46990 2862 46996 2894
rect 46920 0 46996 2862
rect 48144 2862 48150 2894
rect 48214 2894 48215 2926
rect 49237 2926 49303 2927
rect 49237 2894 49238 2926
rect 48214 2862 48220 2894
rect 47469 1702 47535 1703
rect 47469 1670 47470 1702
rect 47464 1638 47470 1670
rect 47534 1670 47535 1702
rect 47534 1638 47540 1670
rect 47464 1294 47540 1638
rect 47464 1230 47470 1294
rect 47534 1230 47540 1294
rect 47464 1224 47540 1230
rect 48144 0 48220 2862
rect 49232 2862 49238 2894
rect 49302 2894 49303 2926
rect 49302 2862 49308 2894
rect 48965 1702 49031 1703
rect 48965 1670 48966 1702
rect 48960 1638 48966 1670
rect 49030 1670 49031 1702
rect 49030 1638 49036 1670
rect 48960 1294 49036 1638
rect 48960 1230 48966 1294
rect 49030 1230 49036 1294
rect 48960 1224 49036 1230
rect 49232 0 49308 2862
rect 49912 0 49988 13334
rect 50184 13126 50260 15102
rect 52360 15166 52436 15172
rect 52360 15102 52366 15166
rect 52430 15102 52436 15166
rect 52496 15166 52572 17006
rect 55080 17070 55156 17076
rect 55080 17006 55086 17070
rect 55150 17006 55156 17070
rect 52496 15134 52502 15166
rect 52229 14350 52295 14351
rect 52229 14318 52230 14350
rect 52224 14286 52230 14318
rect 52294 14318 52295 14350
rect 52294 14286 52300 14318
rect 52224 13670 52300 14286
rect 52224 13606 52230 13670
rect 52294 13606 52300 13670
rect 52224 13600 52300 13606
rect 52224 13534 52300 13540
rect 52224 13470 52230 13534
rect 52294 13470 52300 13534
rect 50184 13094 50190 13126
rect 50189 13062 50190 13094
rect 50254 13094 50260 13126
rect 51957 13126 52023 13127
rect 51957 13094 51958 13126
rect 50254 13062 50255 13094
rect 50189 13061 50255 13062
rect 51952 13062 51958 13094
rect 52022 13094 52023 13126
rect 52022 13062 52028 13094
rect 50325 2926 50391 2927
rect 50325 2894 50326 2926
rect 50320 2862 50326 2894
rect 50390 2894 50391 2926
rect 51685 2926 51751 2927
rect 51685 2894 51686 2926
rect 50390 2862 50396 2894
rect 50320 0 50396 2862
rect 51680 2862 51686 2894
rect 51750 2894 51751 2926
rect 51750 2862 51756 2894
rect 50733 1702 50799 1703
rect 50733 1670 50734 1702
rect 50728 1638 50734 1670
rect 50798 1670 50799 1702
rect 50798 1638 50804 1670
rect 50728 1294 50804 1638
rect 50728 1230 50734 1294
rect 50798 1230 50804 1294
rect 50728 1224 50804 1230
rect 51680 0 51756 2862
rect 51952 0 52028 13062
rect 52224 12038 52300 13470
rect 52360 13262 52436 15102
rect 52501 15102 52502 15134
rect 52566 15134 52572 15166
rect 54944 15166 55020 15172
rect 52566 15102 52567 15134
rect 52501 15101 52567 15102
rect 54944 15102 54950 15166
rect 55014 15102 55020 15166
rect 55080 15166 55156 17006
rect 55080 15134 55086 15166
rect 54813 14350 54879 14351
rect 54813 14318 54814 14350
rect 54808 14286 54814 14318
rect 54878 14318 54879 14350
rect 54878 14286 54884 14318
rect 54808 13670 54884 14286
rect 54808 13606 54814 13670
rect 54878 13606 54884 13670
rect 54808 13600 54884 13606
rect 52360 13230 52366 13262
rect 52365 13198 52366 13230
rect 52430 13230 52436 13262
rect 54808 13534 54884 13540
rect 54808 13470 54814 13534
rect 54878 13470 54884 13534
rect 52430 13198 52431 13230
rect 52365 13197 52431 13198
rect 52360 13126 52436 13132
rect 52360 13062 52366 13126
rect 52430 13062 52436 13126
rect 54541 13126 54607 13127
rect 54541 13094 54542 13126
rect 52360 12582 52436 13062
rect 52360 12550 52366 12582
rect 52365 12518 52366 12550
rect 52430 12550 52436 12582
rect 54536 13062 54542 13094
rect 54606 13094 54607 13126
rect 54606 13062 54612 13094
rect 52430 12518 52431 12550
rect 52365 12517 52431 12518
rect 52365 12310 52431 12311
rect 52365 12278 52366 12310
rect 52224 12006 52230 12038
rect 52229 11974 52230 12006
rect 52294 12006 52300 12038
rect 52360 12246 52366 12278
rect 52430 12278 52431 12310
rect 54400 12310 54476 12316
rect 52430 12246 52436 12278
rect 52294 11974 52295 12006
rect 52229 11973 52295 11974
rect 52229 11902 52295 11903
rect 52229 11870 52230 11902
rect 52224 11838 52230 11870
rect 52294 11870 52295 11902
rect 52294 11838 52300 11870
rect 52224 11086 52300 11838
rect 52360 11766 52436 12246
rect 52360 11702 52366 11766
rect 52430 11702 52436 11766
rect 52360 11696 52436 11702
rect 54400 12246 54406 12310
rect 54470 12246 54476 12310
rect 54400 11494 54476 12246
rect 54400 11462 54406 11494
rect 54405 11430 54406 11462
rect 54470 11462 54476 11494
rect 54470 11430 54471 11462
rect 54405 11429 54471 11430
rect 52224 11022 52230 11086
rect 52294 11022 52300 11086
rect 52224 11016 52300 11022
rect 52773 2926 52839 2927
rect 52773 2894 52774 2926
rect 52768 2862 52774 2894
rect 52838 2894 52839 2926
rect 53861 2926 53927 2927
rect 53861 2894 53862 2926
rect 52838 2862 52844 2894
rect 52501 1702 52567 1703
rect 52501 1670 52502 1702
rect 52496 1638 52502 1670
rect 52566 1670 52567 1702
rect 52566 1638 52572 1670
rect 52496 1294 52572 1638
rect 52496 1230 52502 1294
rect 52566 1230 52572 1294
rect 52496 1224 52572 1230
rect 52768 0 52844 2862
rect 53856 2862 53862 2894
rect 53926 2894 53927 2926
rect 53926 2862 53932 2894
rect 53856 0 53932 2862
rect 54133 1702 54199 1703
rect 54133 1670 54134 1702
rect 54128 1638 54134 1670
rect 54198 1670 54199 1702
rect 54198 1638 54204 1670
rect 54128 1294 54204 1638
rect 54128 1230 54134 1294
rect 54198 1230 54204 1294
rect 54128 1224 54204 1230
rect 54536 0 54612 13062
rect 54808 12038 54884 13470
rect 54944 13262 55020 15102
rect 55085 15102 55086 15134
rect 55150 15134 55156 15166
rect 57392 17070 57468 17076
rect 57392 17006 57398 17070
rect 57462 17006 57468 17070
rect 57392 15166 57468 17006
rect 59840 17070 60052 17076
rect 59840 17006 59982 17070
rect 60046 17006 60052 17070
rect 59840 17000 60052 17006
rect 62560 17070 62636 17076
rect 62560 17006 62566 17070
rect 62630 17006 62636 17070
rect 57392 15134 57398 15166
rect 55150 15102 55151 15134
rect 55085 15101 55151 15102
rect 57397 15102 57398 15134
rect 57462 15134 57468 15166
rect 57528 15166 57604 15172
rect 57462 15102 57463 15134
rect 57397 15101 57463 15102
rect 57528 15102 57534 15166
rect 57598 15102 57604 15166
rect 59840 15166 59916 17000
rect 59840 15134 59846 15166
rect 57397 14350 57463 14351
rect 57397 14318 57398 14350
rect 57392 14286 57398 14318
rect 57462 14318 57463 14350
rect 57462 14286 57468 14318
rect 57392 13670 57468 14286
rect 57392 13606 57398 13670
rect 57462 13606 57468 13670
rect 57392 13600 57468 13606
rect 54944 13230 54950 13262
rect 54949 13198 54950 13230
rect 55014 13230 55020 13262
rect 57392 13534 57468 13540
rect 57392 13470 57398 13534
rect 57462 13470 57468 13534
rect 55014 13198 55015 13230
rect 54949 13197 55015 13198
rect 54944 13126 55020 13132
rect 54944 13062 54950 13126
rect 55014 13062 55020 13126
rect 56989 13126 57055 13127
rect 56989 13094 56990 13126
rect 54944 12582 55020 13062
rect 54944 12550 54950 12582
rect 54949 12518 54950 12550
rect 55014 12550 55020 12582
rect 56984 13062 56990 13094
rect 57054 13094 57055 13126
rect 57256 13126 57332 13132
rect 57054 13062 57060 13094
rect 55014 12518 55015 12550
rect 54949 12517 55015 12518
rect 54808 12006 54814 12038
rect 54813 11974 54814 12006
rect 54878 12006 54884 12038
rect 54878 11974 54879 12006
rect 54813 11973 54879 11974
rect 54813 11902 54879 11903
rect 54813 11870 54814 11902
rect 54808 11838 54814 11870
rect 54878 11870 54879 11902
rect 54878 11838 54884 11870
rect 54808 11086 54884 11838
rect 54808 11022 54814 11086
rect 54878 11022 54884 11086
rect 54808 11016 54884 11022
rect 54949 2926 55015 2927
rect 54949 2894 54950 2926
rect 54944 2862 54950 2894
rect 55014 2894 55015 2926
rect 56309 2926 56375 2927
rect 56309 2894 56310 2926
rect 55014 2862 55020 2894
rect 54944 0 55020 2862
rect 56304 2862 56310 2894
rect 56374 2894 56375 2926
rect 56374 2862 56380 2894
rect 55901 1702 55967 1703
rect 55901 1670 55902 1702
rect 55896 1638 55902 1670
rect 55966 1670 55967 1702
rect 55966 1638 55972 1670
rect 55896 1294 55972 1638
rect 55896 1230 55902 1294
rect 55966 1230 55972 1294
rect 55896 1224 55972 1230
rect 56304 0 56380 2862
rect 56984 0 57060 13062
rect 57256 13062 57262 13126
rect 57326 13062 57332 13126
rect 57256 12582 57332 13062
rect 57256 12550 57262 12582
rect 57261 12518 57262 12550
rect 57326 12550 57332 12582
rect 57326 12518 57327 12550
rect 57261 12517 57327 12518
rect 57392 12038 57468 13470
rect 57528 13262 57604 15102
rect 59845 15102 59846 15134
rect 59910 15134 59916 15166
rect 59976 15166 60052 15172
rect 59910 15102 59911 15134
rect 59845 15101 59911 15102
rect 59976 15102 59982 15166
rect 60046 15102 60052 15166
rect 59845 14350 59911 14351
rect 59845 14318 59846 14350
rect 59840 14286 59846 14318
rect 59910 14318 59911 14350
rect 59910 14286 59916 14318
rect 59840 13670 59916 14286
rect 59840 13606 59846 13670
rect 59910 13606 59916 13670
rect 59840 13600 59916 13606
rect 57528 13230 57534 13262
rect 57533 13198 57534 13230
rect 57598 13230 57604 13262
rect 59840 13534 59916 13540
rect 59840 13470 59846 13534
rect 59910 13470 59916 13534
rect 57598 13198 57599 13230
rect 57533 13197 57599 13198
rect 59301 13126 59367 13127
rect 59301 13094 59302 13126
rect 59296 13062 59302 13094
rect 59366 13094 59367 13126
rect 59366 13062 59372 13094
rect 57533 12310 57599 12311
rect 57533 12278 57534 12310
rect 57392 12006 57398 12038
rect 57397 11974 57398 12006
rect 57462 12006 57468 12038
rect 57528 12246 57534 12278
rect 57598 12278 57599 12310
rect 57598 12246 57604 12278
rect 57462 11974 57463 12006
rect 57397 11973 57463 11974
rect 57261 11902 57327 11903
rect 57261 11870 57262 11902
rect 57256 11838 57262 11870
rect 57326 11870 57327 11902
rect 57326 11838 57332 11870
rect 57256 11086 57332 11838
rect 57528 11766 57604 12246
rect 57528 11702 57534 11766
rect 57598 11702 57604 11766
rect 57528 11696 57604 11702
rect 57256 11022 57262 11086
rect 57326 11022 57332 11086
rect 57256 11016 57332 11022
rect 57533 2926 57599 2927
rect 57533 2894 57534 2926
rect 57528 2862 57534 2894
rect 57598 2894 57599 2926
rect 58621 2926 58687 2927
rect 58621 2894 58622 2926
rect 57598 2862 57604 2894
rect 57397 1702 57463 1703
rect 57397 1670 57398 1702
rect 57392 1638 57398 1670
rect 57462 1670 57463 1702
rect 57462 1638 57468 1670
rect 57392 1294 57468 1638
rect 57392 1230 57398 1294
rect 57462 1230 57468 1294
rect 57392 1224 57468 1230
rect 57528 0 57604 2862
rect 58616 2862 58622 2894
rect 58686 2894 58687 2926
rect 58686 2862 58692 2894
rect 58616 0 58692 2862
rect 59165 1702 59231 1703
rect 59165 1670 59166 1702
rect 59160 1638 59166 1670
rect 59230 1670 59231 1702
rect 59230 1638 59236 1670
rect 59160 1294 59236 1638
rect 59160 1230 59166 1294
rect 59230 1230 59236 1294
rect 59160 1224 59236 1230
rect 59296 0 59372 13062
rect 59573 12310 59639 12311
rect 59573 12278 59574 12310
rect 59568 12246 59574 12278
rect 59638 12278 59639 12310
rect 59638 12246 59644 12278
rect 59568 11766 59644 12246
rect 59840 12038 59916 13470
rect 59976 13262 60052 15102
rect 62424 15166 62500 15172
rect 62424 15102 62430 15166
rect 62494 15102 62500 15166
rect 62560 15166 62636 17006
rect 62560 15134 62566 15166
rect 62293 14350 62359 14351
rect 62293 14318 62294 14350
rect 62288 14286 62294 14318
rect 62358 14318 62359 14350
rect 62358 14286 62364 14318
rect 62288 13670 62364 14286
rect 62288 13606 62294 13670
rect 62358 13606 62364 13670
rect 62288 13600 62364 13606
rect 59976 13230 59982 13262
rect 59981 13198 59982 13230
rect 60046 13230 60052 13262
rect 62288 13534 62364 13540
rect 62288 13470 62294 13534
rect 62358 13470 62364 13534
rect 60046 13198 60047 13230
rect 59981 13197 60047 13198
rect 59976 13126 60052 13132
rect 59976 13062 59982 13126
rect 60046 13062 60052 13126
rect 61885 13126 61951 13127
rect 61885 13094 61886 13126
rect 59976 12582 60052 13062
rect 59976 12550 59982 12582
rect 59981 12518 59982 12550
rect 60046 12550 60052 12582
rect 61880 13062 61886 13094
rect 61950 13094 61951 13126
rect 61950 13062 61956 13094
rect 60046 12518 60047 12550
rect 59981 12517 60047 12518
rect 59840 12006 59846 12038
rect 59845 11974 59846 12006
rect 59910 12006 59916 12038
rect 59910 11974 59911 12006
rect 59845 11973 59911 11974
rect 59709 11902 59775 11903
rect 59709 11870 59710 11902
rect 59568 11702 59574 11766
rect 59638 11702 59644 11766
rect 59568 11696 59644 11702
rect 59704 11838 59710 11870
rect 59774 11870 59775 11902
rect 59774 11838 59780 11870
rect 59704 11086 59780 11838
rect 59704 11022 59710 11086
rect 59774 11022 59780 11086
rect 59704 11016 59780 11022
rect 59709 2926 59775 2927
rect 59709 2894 59710 2926
rect 59704 2862 59710 2894
rect 59774 2894 59775 2926
rect 59774 2862 59780 2894
rect 59704 0 59780 2862
rect 60933 1702 60999 1703
rect 60933 1670 60934 1702
rect 60928 1638 60934 1670
rect 60998 1670 60999 1702
rect 60998 1638 61004 1670
rect 60928 1294 61004 1638
rect 60928 1230 60934 1294
rect 60998 1230 61004 1294
rect 60928 1224 61004 1230
rect 61880 0 61956 13062
rect 62288 12038 62364 13470
rect 62424 13262 62500 15102
rect 62565 15102 62566 15134
rect 62630 15134 62636 15166
rect 64872 17070 64948 17076
rect 64872 17006 64878 17070
rect 64942 17006 64948 17070
rect 64872 15166 64948 17006
rect 67592 17070 67668 17076
rect 67592 17006 67598 17070
rect 67662 17006 67668 17070
rect 64872 15134 64878 15166
rect 62630 15102 62631 15134
rect 62565 15101 62631 15102
rect 64877 15102 64878 15134
rect 64942 15134 64948 15166
rect 65008 15166 65084 15172
rect 64942 15102 64943 15134
rect 64877 15101 64943 15102
rect 65008 15102 65014 15166
rect 65078 15102 65084 15166
rect 64877 14350 64943 14351
rect 64877 14318 64878 14350
rect 64872 14286 64878 14318
rect 64942 14318 64943 14350
rect 64942 14286 64948 14318
rect 64872 13670 64948 14286
rect 64872 13606 64878 13670
rect 64942 13606 64948 13670
rect 64872 13600 64948 13606
rect 62424 13230 62430 13262
rect 62429 13198 62430 13230
rect 62494 13230 62500 13262
rect 64736 13534 64812 13540
rect 64736 13470 64742 13534
rect 64806 13470 64812 13534
rect 62494 13198 62495 13230
rect 62429 13197 62495 13198
rect 62424 13126 62500 13132
rect 62424 13062 62430 13126
rect 62494 13062 62500 13126
rect 64469 13126 64535 13127
rect 64469 13094 64470 13126
rect 62424 12582 62500 13062
rect 62424 12550 62430 12582
rect 62429 12518 62430 12550
rect 62494 12550 62500 12582
rect 64464 13062 64470 13094
rect 64534 13094 64535 13126
rect 64534 13062 64540 13094
rect 62494 12518 62495 12550
rect 62429 12517 62495 12518
rect 62429 12310 62495 12311
rect 62429 12278 62430 12310
rect 62288 12006 62294 12038
rect 62293 11974 62294 12006
rect 62358 12006 62364 12038
rect 62424 12246 62430 12278
rect 62494 12278 62495 12310
rect 62494 12246 62500 12278
rect 62358 11974 62359 12006
rect 62293 11973 62359 11974
rect 62157 11902 62223 11903
rect 62157 11870 62158 11902
rect 62152 11838 62158 11870
rect 62222 11870 62223 11902
rect 62222 11838 62228 11870
rect 62152 11086 62228 11838
rect 62424 11766 62500 12246
rect 62424 11702 62430 11766
rect 62494 11702 62500 11766
rect 62424 11696 62500 11702
rect 62152 11022 62158 11086
rect 62222 11022 62228 11086
rect 62152 11016 62228 11022
rect 62701 1702 62767 1703
rect 62701 1670 62702 1702
rect 62696 1638 62702 1670
rect 62766 1670 62767 1702
rect 64197 1702 64263 1703
rect 64197 1670 64198 1702
rect 62766 1638 62772 1670
rect 62696 1294 62772 1638
rect 62696 1230 62702 1294
rect 62766 1230 62772 1294
rect 62696 1224 62772 1230
rect 64192 1638 64198 1670
rect 64262 1670 64263 1702
rect 64262 1638 64268 1670
rect 64192 1294 64268 1638
rect 64192 1230 64198 1294
rect 64262 1230 64268 1294
rect 64192 1224 64268 1230
rect 64464 0 64540 13062
rect 64736 12038 64812 13470
rect 65008 13262 65084 15102
rect 67456 15166 67532 15172
rect 67456 15102 67462 15166
rect 67526 15102 67532 15166
rect 67592 15166 67668 17006
rect 67592 15134 67598 15166
rect 67189 14350 67255 14351
rect 67189 14318 67190 14350
rect 67184 14286 67190 14318
rect 67254 14318 67255 14350
rect 67254 14286 67260 14318
rect 67184 13670 67260 14286
rect 67184 13606 67190 13670
rect 67254 13606 67260 13670
rect 67184 13600 67260 13606
rect 65008 13230 65014 13262
rect 65013 13198 65014 13230
rect 65078 13230 65084 13262
rect 67320 13534 67396 13540
rect 67320 13470 67326 13534
rect 67390 13470 67396 13534
rect 65078 13198 65079 13230
rect 65013 13197 65079 13198
rect 64872 13126 64948 13132
rect 64872 13062 64878 13126
rect 64942 13062 64948 13126
rect 66917 13126 66983 13127
rect 66917 13094 66918 13126
rect 64872 12582 64948 13062
rect 64872 12550 64878 12582
rect 64877 12518 64878 12550
rect 64942 12550 64948 12582
rect 66912 13062 66918 13094
rect 66982 13094 66983 13126
rect 66982 13062 66988 13094
rect 64942 12518 64943 12550
rect 64877 12517 64943 12518
rect 64877 12310 64943 12311
rect 64877 12278 64878 12310
rect 64736 12006 64742 12038
rect 64741 11974 64742 12006
rect 64806 12006 64812 12038
rect 64872 12246 64878 12278
rect 64942 12278 64943 12310
rect 64942 12246 64948 12278
rect 64806 11974 64807 12006
rect 64741 11973 64807 11974
rect 64741 11902 64807 11903
rect 64741 11870 64742 11902
rect 64736 11838 64742 11870
rect 64806 11870 64807 11902
rect 64806 11838 64812 11870
rect 64736 11086 64812 11838
rect 64872 11766 64948 12246
rect 64872 11702 64878 11766
rect 64942 11702 64948 11766
rect 64872 11696 64948 11702
rect 64736 11022 64742 11086
rect 64806 11022 64812 11086
rect 64736 11016 64812 11022
rect 65829 1702 65895 1703
rect 65829 1670 65830 1702
rect 65824 1638 65830 1670
rect 65894 1670 65895 1702
rect 65894 1638 65900 1670
rect 65824 1294 65900 1638
rect 65824 1230 65830 1294
rect 65894 1230 65900 1294
rect 65824 1224 65900 1230
rect 66912 0 66988 13062
rect 67320 12038 67396 13470
rect 67456 13262 67532 15102
rect 67597 15102 67598 15134
rect 67662 15134 67668 15166
rect 69904 17070 69980 17076
rect 69904 17006 69910 17070
rect 69974 17006 69980 17070
rect 69904 15166 69980 17006
rect 72352 17070 72428 17076
rect 72352 17006 72358 17070
rect 72422 17006 72428 17070
rect 69904 15134 69910 15166
rect 67662 15102 67663 15134
rect 67597 15101 67663 15102
rect 69909 15102 69910 15134
rect 69974 15134 69980 15166
rect 70040 15166 70116 15172
rect 69974 15102 69975 15134
rect 69909 15101 69975 15102
rect 70040 15102 70046 15166
rect 70110 15102 70116 15166
rect 72352 15166 72428 17006
rect 75072 17070 75148 17076
rect 75072 17006 75078 17070
rect 75142 17006 75148 17070
rect 72352 15134 72358 15166
rect 69637 14350 69703 14351
rect 69637 14318 69638 14350
rect 69632 14286 69638 14318
rect 69702 14318 69703 14350
rect 69702 14286 69708 14318
rect 69632 13670 69708 14286
rect 69632 13606 69638 13670
rect 69702 13606 69708 13670
rect 69632 13600 69708 13606
rect 69768 13670 69844 13676
rect 69768 13606 69774 13670
rect 69838 13606 69844 13670
rect 67456 13230 67462 13262
rect 67461 13198 67462 13230
rect 67526 13230 67532 13262
rect 67526 13198 67527 13230
rect 67461 13197 67527 13198
rect 67456 13126 67532 13132
rect 67456 13062 67462 13126
rect 67526 13062 67532 13126
rect 69501 13126 69567 13127
rect 69501 13094 69502 13126
rect 67456 12582 67532 13062
rect 67456 12550 67462 12582
rect 67461 12518 67462 12550
rect 67526 12550 67532 12582
rect 69496 13062 69502 13094
rect 69566 13094 69567 13126
rect 69566 13062 69572 13094
rect 67526 12518 67527 12550
rect 67461 12517 67527 12518
rect 67461 12310 67527 12311
rect 67461 12278 67462 12310
rect 67320 12006 67326 12038
rect 67325 11974 67326 12006
rect 67390 12006 67396 12038
rect 67456 12246 67462 12278
rect 67526 12278 67527 12310
rect 67526 12246 67532 12278
rect 67390 11974 67391 12006
rect 67325 11973 67391 11974
rect 67189 11902 67255 11903
rect 67189 11870 67190 11902
rect 67184 11838 67190 11870
rect 67254 11870 67255 11902
rect 67254 11838 67260 11870
rect 67184 11086 67260 11838
rect 67456 11766 67532 12246
rect 67456 11702 67462 11766
rect 67526 11702 67532 11766
rect 67456 11696 67532 11702
rect 67184 11022 67190 11086
rect 67254 11022 67260 11086
rect 67184 11016 67260 11022
rect 67597 1702 67663 1703
rect 67597 1670 67598 1702
rect 67592 1638 67598 1670
rect 67662 1670 67663 1702
rect 69229 1702 69295 1703
rect 69229 1670 69230 1702
rect 67662 1638 67668 1670
rect 67592 1294 67668 1638
rect 67592 1230 67598 1294
rect 67662 1230 67668 1294
rect 67592 1224 67668 1230
rect 69224 1638 69230 1670
rect 69294 1670 69295 1702
rect 69294 1638 69300 1670
rect 69224 1294 69300 1638
rect 69224 1230 69230 1294
rect 69294 1230 69300 1294
rect 69224 1224 69300 1230
rect 69496 0 69572 13062
rect 69768 12038 69844 13606
rect 69904 13126 69980 13132
rect 69904 13062 69910 13126
rect 69974 13062 69980 13126
rect 69904 12582 69980 13062
rect 70040 12990 70116 15102
rect 72357 15102 72358 15134
rect 72422 15134 72428 15166
rect 72488 15166 72564 15172
rect 72422 15102 72423 15134
rect 72357 15101 72423 15102
rect 72488 15102 72494 15166
rect 72558 15102 72564 15166
rect 72080 14350 72156 14356
rect 72080 14286 72086 14350
rect 72150 14286 72156 14350
rect 72221 14350 72287 14351
rect 72221 14318 72222 14350
rect 72080 13670 72156 14286
rect 72080 13638 72086 13670
rect 72085 13606 72086 13638
rect 72150 13638 72156 13670
rect 72216 14286 72222 14318
rect 72286 14318 72287 14350
rect 72286 14286 72292 14318
rect 72216 13670 72292 14286
rect 72150 13606 72151 13638
rect 72085 13605 72151 13606
rect 72216 13606 72222 13670
rect 72286 13606 72292 13670
rect 72216 13600 72292 13606
rect 72352 13534 72428 13540
rect 72352 13470 72358 13534
rect 72422 13470 72428 13534
rect 71949 13126 72015 13127
rect 71949 13094 71950 13126
rect 70040 12958 70046 12990
rect 70045 12926 70046 12958
rect 70110 12958 70116 12990
rect 71944 13062 71950 13094
rect 72014 13094 72015 13126
rect 72014 13062 72020 13094
rect 70110 12926 70111 12958
rect 70045 12925 70111 12926
rect 69904 12550 69910 12582
rect 69909 12518 69910 12550
rect 69974 12550 69980 12582
rect 69974 12518 69975 12550
rect 69909 12517 69975 12518
rect 69909 12310 69975 12311
rect 69909 12278 69910 12310
rect 69768 12006 69774 12038
rect 69773 11974 69774 12006
rect 69838 12006 69844 12038
rect 69904 12246 69910 12278
rect 69974 12278 69975 12310
rect 69974 12246 69980 12278
rect 69838 11974 69839 12006
rect 69773 11973 69839 11974
rect 69773 11902 69839 11903
rect 69773 11870 69774 11902
rect 69768 11838 69774 11870
rect 69838 11870 69839 11902
rect 69838 11838 69844 11870
rect 69768 11086 69844 11838
rect 69904 11766 69980 12246
rect 69904 11702 69910 11766
rect 69974 11702 69980 11766
rect 69904 11696 69980 11702
rect 69768 11022 69774 11086
rect 69838 11022 69844 11086
rect 69768 11016 69844 11022
rect 71133 1702 71199 1703
rect 71133 1670 71134 1702
rect 71128 1638 71134 1670
rect 71198 1670 71199 1702
rect 71198 1638 71204 1670
rect 71128 1294 71204 1638
rect 71128 1230 71134 1294
rect 71198 1230 71204 1294
rect 71128 1224 71204 1230
rect 71944 0 72020 13062
rect 72352 12038 72428 13470
rect 72488 13262 72564 15102
rect 74936 15166 75012 15172
rect 74936 15102 74942 15166
rect 75006 15102 75012 15166
rect 75072 15166 75148 17006
rect 75072 15134 75078 15166
rect 74805 14350 74871 14351
rect 74805 14318 74806 14350
rect 74800 14286 74806 14318
rect 74870 14318 74871 14350
rect 74870 14286 74876 14318
rect 74800 13670 74876 14286
rect 74800 13606 74806 13670
rect 74870 13606 74876 13670
rect 74800 13600 74876 13606
rect 72488 13230 72494 13262
rect 72493 13198 72494 13230
rect 72558 13230 72564 13262
rect 74800 13534 74876 13540
rect 74800 13470 74806 13534
rect 74870 13470 74876 13534
rect 72558 13198 72559 13230
rect 72493 13197 72559 13198
rect 72488 13126 72564 13132
rect 72488 13062 72494 13126
rect 72558 13062 72564 13126
rect 74397 13126 74463 13127
rect 74397 13094 74398 13126
rect 72488 12582 72564 13062
rect 72488 12550 72494 12582
rect 72493 12518 72494 12550
rect 72558 12550 72564 12582
rect 74392 13062 74398 13094
rect 74462 13094 74463 13126
rect 74462 13062 74468 13094
rect 72558 12518 72559 12550
rect 72493 12517 72559 12518
rect 72493 12310 72559 12311
rect 72493 12278 72494 12310
rect 72352 12006 72358 12038
rect 72357 11974 72358 12006
rect 72422 12006 72428 12038
rect 72488 12246 72494 12278
rect 72558 12278 72559 12310
rect 72558 12246 72564 12278
rect 72422 11974 72423 12006
rect 72357 11973 72423 11974
rect 72221 11902 72287 11903
rect 72221 11870 72222 11902
rect 72216 11838 72222 11870
rect 72286 11870 72287 11902
rect 72286 11838 72292 11870
rect 72216 11086 72292 11838
rect 72488 11766 72564 12246
rect 72488 11702 72494 11766
rect 72558 11702 72564 11766
rect 72488 11696 72564 11702
rect 72216 11022 72222 11086
rect 72286 11022 72292 11086
rect 72216 11016 72292 11022
rect 72629 1702 72695 1703
rect 72629 1670 72630 1702
rect 72624 1638 72630 1670
rect 72694 1670 72695 1702
rect 74261 1702 74327 1703
rect 74261 1670 74262 1702
rect 72694 1638 72700 1670
rect 72624 1294 72700 1638
rect 72624 1230 72630 1294
rect 72694 1230 72700 1294
rect 72624 1224 72700 1230
rect 74256 1638 74262 1670
rect 74326 1670 74327 1702
rect 74326 1638 74332 1670
rect 74256 1294 74332 1638
rect 74256 1230 74262 1294
rect 74326 1230 74332 1294
rect 74256 1224 74332 1230
rect 74392 0 74468 13062
rect 74669 12310 74735 12311
rect 74669 12278 74670 12310
rect 74664 12246 74670 12278
rect 74734 12278 74735 12310
rect 74734 12246 74740 12278
rect 74533 11902 74599 11903
rect 74533 11870 74534 11902
rect 74528 11838 74534 11870
rect 74598 11870 74599 11902
rect 74598 11838 74604 11870
rect 74528 11086 74604 11838
rect 74664 11766 74740 12246
rect 74800 12038 74876 13470
rect 74936 13262 75012 15102
rect 75077 15102 75078 15134
rect 75142 15134 75148 15166
rect 75142 15102 75143 15134
rect 75077 15101 75143 15102
rect 77112 14486 77188 18638
rect 110160 17206 110236 19726
rect 121312 18566 121388 20134
rect 124168 20134 124174 20166
rect 124238 20166 124239 20198
rect 124238 20134 124244 20166
rect 124168 19926 124244 20134
rect 124168 19862 124174 19926
rect 124238 19862 124244 19926
rect 124168 19856 124244 19862
rect 121312 18502 121318 18566
rect 121382 18502 121388 18566
rect 121312 18496 121388 18502
rect 124304 19790 124380 19796
rect 124304 19726 124310 19790
rect 124374 19726 124380 19790
rect 124173 18430 124239 18431
rect 124173 18398 124174 18430
rect 110160 17174 110166 17206
rect 110165 17142 110166 17174
rect 110230 17174 110236 17206
rect 124168 18366 124174 18398
rect 124238 18398 124239 18430
rect 124238 18366 124244 18398
rect 110230 17142 110231 17174
rect 110165 17141 110231 17142
rect 77520 17070 77596 17076
rect 77520 17006 77526 17070
rect 77590 17006 77596 17070
rect 77112 14422 77118 14486
rect 77182 14422 77188 14486
rect 77112 14416 77188 14422
rect 77384 15166 77460 15172
rect 77384 15102 77390 15166
rect 77454 15102 77460 15166
rect 77520 15166 77596 17006
rect 77520 15134 77526 15166
rect 76981 14350 77047 14351
rect 76981 14318 76982 14350
rect 76976 14286 76982 14318
rect 77046 14318 77047 14350
rect 77253 14350 77319 14351
rect 77253 14318 77254 14350
rect 77046 14286 77052 14318
rect 76976 13670 77052 14286
rect 77248 14286 77254 14318
rect 77318 14318 77319 14350
rect 77318 14286 77324 14318
rect 76976 13606 76982 13670
rect 77046 13606 77052 13670
rect 76976 13600 77052 13606
rect 77112 13670 77188 13676
rect 77112 13606 77118 13670
rect 77182 13606 77188 13670
rect 74936 13230 74942 13262
rect 74941 13198 74942 13230
rect 75006 13230 75012 13262
rect 75006 13198 75007 13230
rect 74941 13197 75007 13198
rect 74936 13126 75012 13132
rect 74936 13062 74942 13126
rect 75006 13062 75012 13126
rect 76845 13126 76911 13127
rect 76845 13094 76846 13126
rect 74936 12582 75012 13062
rect 74936 12550 74942 12582
rect 74941 12518 74942 12550
rect 75006 12550 75012 12582
rect 76840 13062 76846 13094
rect 76910 13094 76911 13126
rect 76910 13062 76916 13094
rect 75006 12518 75007 12550
rect 74941 12517 75007 12518
rect 74800 12006 74806 12038
rect 74805 11974 74806 12006
rect 74870 12006 74876 12038
rect 74870 11974 74871 12006
rect 74805 11973 74871 11974
rect 74664 11702 74670 11766
rect 74734 11702 74740 11766
rect 74664 11696 74740 11702
rect 74528 11022 74534 11086
rect 74598 11022 74604 11086
rect 74528 11016 74604 11022
rect 76029 1702 76095 1703
rect 76029 1670 76030 1702
rect 76024 1638 76030 1670
rect 76094 1670 76095 1702
rect 76094 1638 76100 1670
rect 76024 1294 76100 1638
rect 76024 1230 76030 1294
rect 76094 1230 76100 1294
rect 76024 1224 76100 1230
rect 76840 0 76916 13062
rect 76981 12310 77047 12311
rect 76981 12278 76982 12310
rect 76976 12246 76982 12278
rect 77046 12278 77047 12310
rect 77046 12246 77052 12278
rect 76976 11766 77052 12246
rect 77112 12038 77188 13606
rect 77248 13670 77324 14286
rect 77248 13606 77254 13670
rect 77318 13606 77324 13670
rect 77248 13600 77324 13606
rect 77248 13126 77324 13132
rect 77248 13062 77254 13126
rect 77318 13062 77324 13126
rect 77384 13126 77460 15102
rect 77525 15102 77526 15134
rect 77590 15134 77596 15166
rect 79832 17070 79908 17076
rect 79832 17006 79838 17070
rect 79902 17006 79908 17070
rect 79832 15166 79908 17006
rect 82552 17070 82628 17076
rect 82552 17006 82558 17070
rect 82622 17006 82628 17070
rect 79832 15134 79838 15166
rect 77590 15102 77591 15134
rect 77525 15101 77591 15102
rect 79837 15102 79838 15134
rect 79902 15134 79908 15166
rect 79968 15166 80044 15172
rect 79902 15102 79903 15134
rect 79837 15101 79903 15102
rect 79968 15102 79974 15166
rect 80038 15102 80044 15166
rect 79837 14350 79903 14351
rect 79837 14318 79838 14350
rect 79832 14286 79838 14318
rect 79902 14318 79903 14350
rect 79902 14286 79908 14318
rect 79832 13670 79908 14286
rect 79832 13606 79838 13670
rect 79902 13606 79908 13670
rect 79832 13600 79908 13606
rect 79832 13534 79908 13540
rect 79832 13470 79838 13534
rect 79902 13470 79908 13534
rect 77384 13094 77390 13126
rect 77248 12582 77324 13062
rect 77389 13062 77390 13094
rect 77454 13094 77460 13126
rect 79429 13126 79495 13127
rect 79429 13094 79430 13126
rect 77454 13062 77455 13094
rect 77389 13061 77455 13062
rect 79424 13062 79430 13094
rect 79494 13094 79495 13126
rect 79494 13062 79500 13094
rect 77248 12550 77254 12582
rect 77253 12518 77254 12550
rect 77318 12550 77324 12582
rect 77318 12518 77319 12550
rect 77253 12517 77319 12518
rect 77112 12006 77118 12038
rect 77117 11974 77118 12006
rect 77182 12006 77188 12038
rect 77182 11974 77183 12006
rect 77117 11973 77183 11974
rect 77253 11902 77319 11903
rect 77253 11870 77254 11902
rect 76976 11702 76982 11766
rect 77046 11702 77052 11766
rect 76976 11696 77052 11702
rect 77248 11838 77254 11870
rect 77318 11870 77319 11902
rect 77318 11838 77324 11870
rect 77248 11086 77324 11838
rect 77248 11022 77254 11086
rect 77318 11022 77324 11086
rect 77248 11016 77324 11022
rect 77661 1702 77727 1703
rect 77661 1670 77662 1702
rect 77656 1638 77662 1670
rect 77726 1670 77727 1702
rect 79293 1702 79359 1703
rect 79293 1670 79294 1702
rect 77726 1638 77732 1670
rect 77656 1294 77732 1638
rect 77656 1230 77662 1294
rect 77726 1230 77732 1294
rect 77656 1224 77732 1230
rect 79288 1638 79294 1670
rect 79358 1670 79359 1702
rect 79358 1638 79364 1670
rect 79288 1294 79364 1638
rect 79288 1230 79294 1294
rect 79358 1230 79364 1294
rect 79288 1224 79364 1230
rect 79424 0 79500 13062
rect 79832 12038 79908 13470
rect 79968 13262 80044 15102
rect 82416 15166 82492 15172
rect 82416 15102 82422 15166
rect 82486 15102 82492 15166
rect 82552 15166 82628 17006
rect 82552 15134 82558 15166
rect 82285 14350 82351 14351
rect 82285 14318 82286 14350
rect 82280 14286 82286 14318
rect 82350 14318 82351 14350
rect 82350 14286 82356 14318
rect 82280 13670 82356 14286
rect 82280 13606 82286 13670
rect 82350 13606 82356 13670
rect 82280 13600 82356 13606
rect 79968 13230 79974 13262
rect 79973 13198 79974 13230
rect 80038 13230 80044 13262
rect 82280 13534 82356 13540
rect 82280 13470 82286 13534
rect 82350 13470 82356 13534
rect 80038 13198 80039 13230
rect 79973 13197 80039 13198
rect 79968 13126 80044 13132
rect 79968 13062 79974 13126
rect 80038 13062 80044 13126
rect 81877 13126 81943 13127
rect 81877 13094 81878 13126
rect 79968 12582 80044 13062
rect 79968 12550 79974 12582
rect 79973 12518 79974 12550
rect 80038 12550 80044 12582
rect 81872 13062 81878 13094
rect 81942 13094 81943 13126
rect 81942 13062 81948 13094
rect 80038 12518 80039 12550
rect 79973 12517 80039 12518
rect 79973 12310 80039 12311
rect 79973 12278 79974 12310
rect 79832 12006 79838 12038
rect 79837 11974 79838 12006
rect 79902 12006 79908 12038
rect 79968 12246 79974 12278
rect 80038 12278 80039 12310
rect 80038 12246 80044 12278
rect 79902 11974 79903 12006
rect 79837 11973 79903 11974
rect 79701 11902 79767 11903
rect 79701 11870 79702 11902
rect 79696 11838 79702 11870
rect 79766 11870 79767 11902
rect 79766 11838 79772 11870
rect 79696 11086 79772 11838
rect 79968 11766 80044 12246
rect 79968 11702 79974 11766
rect 80038 11702 80044 11766
rect 79968 11696 80044 11702
rect 79696 11022 79702 11086
rect 79766 11022 79772 11086
rect 79696 11016 79772 11022
rect 81197 1702 81263 1703
rect 81197 1670 81198 1702
rect 81192 1638 81198 1670
rect 81262 1670 81263 1702
rect 81262 1638 81268 1670
rect 81192 1294 81268 1638
rect 81192 1230 81198 1294
rect 81262 1230 81268 1294
rect 81192 1224 81268 1230
rect 81872 0 81948 13062
rect 82280 12038 82356 13470
rect 82416 13262 82492 15102
rect 82557 15102 82558 15134
rect 82622 15134 82628 15166
rect 84864 17070 84940 17076
rect 84864 17006 84870 17070
rect 84934 17006 84940 17070
rect 84864 15166 84940 17006
rect 87312 17070 87388 17076
rect 87312 17006 87318 17070
rect 87382 17006 87388 17070
rect 84864 15134 84870 15166
rect 82622 15102 82623 15134
rect 82557 15101 82623 15102
rect 84869 15102 84870 15134
rect 84934 15134 84940 15166
rect 85000 15166 85076 15172
rect 84934 15102 84935 15134
rect 84869 15101 84935 15102
rect 85000 15102 85006 15166
rect 85070 15102 85076 15166
rect 87312 15166 87388 17006
rect 90032 17070 90108 17076
rect 90032 17006 90038 17070
rect 90102 17006 90108 17070
rect 87312 15134 87318 15166
rect 84597 14350 84663 14351
rect 84597 14318 84598 14350
rect 84592 14286 84598 14318
rect 84662 14318 84663 14350
rect 84662 14286 84668 14318
rect 84592 13670 84668 14286
rect 84592 13606 84598 13670
rect 84662 13606 84668 13670
rect 84592 13600 84668 13606
rect 82416 13230 82422 13262
rect 82421 13198 82422 13230
rect 82486 13230 82492 13262
rect 84864 13534 84940 13540
rect 84864 13470 84870 13534
rect 84934 13470 84940 13534
rect 82486 13198 82487 13230
rect 82421 13197 82487 13198
rect 82416 13126 82492 13132
rect 82416 13062 82422 13126
rect 82486 13062 82492 13126
rect 84325 13126 84391 13127
rect 84325 13094 84326 13126
rect 82416 12582 82492 13062
rect 82416 12550 82422 12582
rect 82421 12518 82422 12550
rect 82486 12550 82492 12582
rect 84320 13062 84326 13094
rect 84390 13094 84391 13126
rect 84728 13126 84804 13132
rect 84390 13062 84396 13094
rect 82486 12518 82487 12550
rect 82421 12517 82487 12518
rect 82421 12310 82487 12311
rect 82421 12278 82422 12310
rect 82280 12006 82286 12038
rect 82285 11974 82286 12006
rect 82350 12006 82356 12038
rect 82416 12246 82422 12278
rect 82486 12278 82487 12310
rect 82486 12246 82492 12278
rect 82350 11974 82351 12006
rect 82285 11973 82351 11974
rect 82149 11902 82215 11903
rect 82149 11870 82150 11902
rect 82144 11838 82150 11870
rect 82214 11870 82215 11902
rect 82214 11838 82220 11870
rect 82144 11086 82220 11838
rect 82416 11766 82492 12246
rect 82416 11702 82422 11766
rect 82486 11702 82492 11766
rect 82416 11696 82492 11702
rect 82144 11022 82150 11086
rect 82214 11022 82220 11086
rect 82144 11016 82220 11022
rect 82693 1702 82759 1703
rect 82693 1670 82694 1702
rect 82688 1638 82694 1670
rect 82758 1670 82759 1702
rect 82758 1638 82764 1670
rect 82688 1294 82764 1638
rect 82688 1230 82694 1294
rect 82758 1230 82764 1294
rect 82688 1224 82764 1230
rect 84320 0 84396 13062
rect 84728 13062 84734 13126
rect 84798 13062 84804 13126
rect 84728 12582 84804 13062
rect 84728 12550 84734 12582
rect 84733 12518 84734 12550
rect 84798 12550 84804 12582
rect 84798 12518 84799 12550
rect 84733 12517 84799 12518
rect 84733 12310 84799 12311
rect 84733 12278 84734 12310
rect 84728 12246 84734 12278
rect 84798 12278 84799 12310
rect 84798 12246 84804 12278
rect 84597 11902 84663 11903
rect 84597 11870 84598 11902
rect 84592 11838 84598 11870
rect 84662 11870 84663 11902
rect 84662 11838 84668 11870
rect 84592 11086 84668 11838
rect 84728 11766 84804 12246
rect 84864 12038 84940 13470
rect 85000 13262 85076 15102
rect 87317 15102 87318 15134
rect 87382 15134 87388 15166
rect 87448 15166 87524 15172
rect 87382 15102 87383 15134
rect 87317 15101 87383 15102
rect 87448 15102 87454 15166
rect 87518 15102 87524 15166
rect 87317 14350 87383 14351
rect 87317 14318 87318 14350
rect 87312 14286 87318 14318
rect 87382 14318 87383 14350
rect 87382 14286 87388 14318
rect 87312 13670 87388 14286
rect 87312 13606 87318 13670
rect 87382 13606 87388 13670
rect 87312 13600 87388 13606
rect 85000 13230 85006 13262
rect 85005 13198 85006 13230
rect 85070 13230 85076 13262
rect 87312 13534 87388 13540
rect 87312 13470 87318 13534
rect 87382 13470 87388 13534
rect 85070 13198 85071 13230
rect 85005 13197 85071 13198
rect 86909 13126 86975 13127
rect 86909 13094 86910 13126
rect 84864 12006 84870 12038
rect 84869 11974 84870 12006
rect 84934 12006 84940 12038
rect 86904 13062 86910 13094
rect 86974 13094 86975 13126
rect 86974 13062 86980 13094
rect 84934 11974 84935 12006
rect 84869 11973 84935 11974
rect 84728 11702 84734 11766
rect 84798 11702 84804 11766
rect 84728 11696 84804 11702
rect 84592 11022 84598 11086
rect 84662 11022 84668 11086
rect 84592 11016 84668 11022
rect 84597 1702 84663 1703
rect 84597 1670 84598 1702
rect 84592 1638 84598 1670
rect 84662 1670 84663 1702
rect 86093 1702 86159 1703
rect 86093 1670 86094 1702
rect 84662 1638 84668 1670
rect 84592 1294 84668 1638
rect 84592 1230 84598 1294
rect 84662 1230 84668 1294
rect 84592 1224 84668 1230
rect 86088 1638 86094 1670
rect 86158 1670 86159 1702
rect 86158 1638 86164 1670
rect 86088 1294 86164 1638
rect 86088 1230 86094 1294
rect 86158 1230 86164 1294
rect 86088 1224 86164 1230
rect 86904 0 86980 13062
rect 87045 12310 87111 12311
rect 87045 12278 87046 12310
rect 87040 12246 87046 12278
rect 87110 12278 87111 12310
rect 87110 12246 87116 12278
rect 87040 11766 87116 12246
rect 87312 12038 87388 13470
rect 87448 13262 87524 15102
rect 89896 15166 89972 15172
rect 89896 15102 89902 15166
rect 89966 15102 89972 15166
rect 90032 15166 90108 17006
rect 90032 15134 90038 15166
rect 89629 14350 89695 14351
rect 89629 14318 89630 14350
rect 89624 14286 89630 14318
rect 89694 14318 89695 14350
rect 89694 14286 89700 14318
rect 89624 13670 89700 14286
rect 89624 13606 89630 13670
rect 89694 13606 89700 13670
rect 89624 13600 89700 13606
rect 87448 13230 87454 13262
rect 87453 13198 87454 13230
rect 87518 13230 87524 13262
rect 89760 13534 89836 13540
rect 89760 13470 89766 13534
rect 89830 13470 89836 13534
rect 87518 13198 87519 13230
rect 87453 13197 87519 13198
rect 87448 13126 87524 13132
rect 87448 13062 87454 13126
rect 87518 13062 87524 13126
rect 89085 13126 89151 13127
rect 89085 13094 89086 13126
rect 87448 12582 87524 13062
rect 87448 12550 87454 12582
rect 87453 12518 87454 12550
rect 87518 12550 87524 12582
rect 89080 13062 89086 13094
rect 89150 13094 89151 13126
rect 89150 13062 89156 13094
rect 87518 12518 87519 12550
rect 87453 12517 87519 12518
rect 87312 12006 87318 12038
rect 87317 11974 87318 12006
rect 87382 12006 87388 12038
rect 87382 11974 87383 12006
rect 87317 11973 87383 11974
rect 87181 11902 87247 11903
rect 87181 11870 87182 11902
rect 87040 11702 87046 11766
rect 87110 11702 87116 11766
rect 87040 11696 87116 11702
rect 87176 11838 87182 11870
rect 87246 11870 87247 11902
rect 87246 11838 87252 11870
rect 87176 11086 87252 11838
rect 87176 11022 87182 11086
rect 87246 11022 87252 11086
rect 87176 11016 87252 11022
rect 87725 1702 87791 1703
rect 87725 1670 87726 1702
rect 87720 1638 87726 1670
rect 87790 1670 87791 1702
rect 87790 1638 87796 1670
rect 87720 1294 87796 1638
rect 87720 1230 87726 1294
rect 87790 1230 87796 1294
rect 87720 1224 87796 1230
rect 89080 0 89156 13062
rect 89629 12310 89695 12311
rect 89629 12278 89630 12310
rect 89624 12246 89630 12278
rect 89694 12278 89695 12310
rect 89694 12246 89700 12278
rect 89493 11902 89559 11903
rect 89493 11870 89494 11902
rect 89488 11838 89494 11870
rect 89558 11870 89559 11902
rect 89558 11838 89564 11870
rect 89488 11086 89564 11838
rect 89624 11766 89700 12246
rect 89760 12038 89836 13470
rect 89896 13262 89972 15102
rect 90037 15102 90038 15134
rect 90102 15134 90108 15166
rect 92344 17070 92420 17076
rect 92344 17006 92350 17070
rect 92414 17006 92420 17070
rect 92344 15166 92420 17006
rect 94792 17070 95004 17076
rect 94792 17006 94934 17070
rect 94998 17006 95004 17070
rect 94792 17000 95004 17006
rect 97512 17070 97588 17076
rect 97512 17006 97518 17070
rect 97582 17006 97588 17070
rect 92344 15134 92350 15166
rect 90102 15102 90103 15134
rect 90037 15101 90103 15102
rect 92349 15102 92350 15134
rect 92414 15134 92420 15166
rect 92480 15166 92556 15172
rect 92414 15102 92415 15134
rect 92349 15101 92415 15102
rect 92480 15102 92486 15166
rect 92550 15102 92556 15166
rect 94792 15166 94868 17000
rect 94792 15134 94798 15166
rect 92213 14350 92279 14351
rect 92213 14318 92214 14350
rect 92208 14286 92214 14318
rect 92278 14318 92279 14350
rect 92278 14286 92284 14318
rect 92208 13670 92284 14286
rect 92208 13606 92214 13670
rect 92278 13606 92284 13670
rect 92208 13600 92284 13606
rect 89896 13230 89902 13262
rect 89901 13198 89902 13230
rect 89966 13230 89972 13262
rect 92344 13534 92420 13540
rect 92344 13470 92350 13534
rect 92414 13470 92420 13534
rect 89966 13198 89967 13230
rect 89901 13197 89967 13198
rect 89896 13126 89972 13132
rect 89896 13062 89902 13126
rect 89966 13062 89972 13126
rect 91941 13126 92007 13127
rect 91941 13094 91942 13126
rect 89896 12582 89972 13062
rect 89896 12550 89902 12582
rect 89901 12518 89902 12550
rect 89966 12550 89972 12582
rect 91936 13062 91942 13094
rect 92006 13094 92007 13126
rect 92208 13126 92284 13132
rect 92006 13062 92012 13094
rect 89966 12518 89967 12550
rect 89901 12517 89967 12518
rect 89760 12006 89766 12038
rect 89765 11974 89766 12006
rect 89830 12006 89836 12038
rect 89830 11974 89831 12006
rect 89765 11973 89831 11974
rect 89624 11702 89630 11766
rect 89694 11702 89700 11766
rect 89624 11696 89700 11702
rect 89488 11022 89494 11086
rect 89558 11022 89564 11086
rect 89488 11016 89564 11022
rect 89357 1702 89423 1703
rect 89357 1670 89358 1702
rect 89352 1638 89358 1670
rect 89422 1670 89423 1702
rect 91125 1702 91191 1703
rect 91125 1670 91126 1702
rect 89422 1638 89428 1670
rect 89352 1294 89428 1638
rect 89352 1230 89358 1294
rect 89422 1230 89428 1294
rect 89352 1224 89428 1230
rect 91120 1638 91126 1670
rect 91190 1670 91191 1702
rect 91190 1638 91196 1670
rect 91120 1294 91196 1638
rect 91120 1230 91126 1294
rect 91190 1230 91196 1294
rect 91120 1224 91196 1230
rect 91936 0 92012 13062
rect 92208 13062 92214 13126
rect 92278 13062 92284 13126
rect 92208 12582 92284 13062
rect 92208 12550 92214 12582
rect 92213 12518 92214 12550
rect 92278 12550 92284 12582
rect 92278 12518 92279 12550
rect 92213 12517 92279 12518
rect 92344 12038 92420 13470
rect 92480 13262 92556 15102
rect 94797 15102 94798 15134
rect 94862 15134 94868 15166
rect 94928 15166 95004 15172
rect 94862 15102 94863 15134
rect 94797 15101 94863 15102
rect 94928 15102 94934 15166
rect 94998 15102 95004 15166
rect 94661 14350 94727 14351
rect 94661 14318 94662 14350
rect 94656 14286 94662 14318
rect 94726 14318 94727 14350
rect 94726 14286 94732 14318
rect 94656 13670 94732 14286
rect 94656 13606 94662 13670
rect 94726 13606 94732 13670
rect 94656 13600 94732 13606
rect 92480 13230 92486 13262
rect 92485 13198 92486 13230
rect 92550 13230 92556 13262
rect 94792 13534 94868 13540
rect 94792 13470 94798 13534
rect 94862 13470 94868 13534
rect 92550 13198 92551 13230
rect 92485 13197 92551 13198
rect 94389 13126 94455 13127
rect 94389 13094 94390 13126
rect 94384 13062 94390 13094
rect 94454 13094 94455 13126
rect 94454 13062 94460 13094
rect 92485 12310 92551 12311
rect 92485 12278 92486 12310
rect 92344 12006 92350 12038
rect 92349 11974 92350 12006
rect 92414 12006 92420 12038
rect 92480 12246 92486 12278
rect 92550 12278 92551 12310
rect 92550 12246 92556 12278
rect 92414 11974 92415 12006
rect 92349 11973 92415 11974
rect 92213 11902 92279 11903
rect 92213 11870 92214 11902
rect 92208 11838 92214 11870
rect 92278 11870 92279 11902
rect 92278 11838 92284 11870
rect 92208 11086 92284 11838
rect 92480 11766 92556 12246
rect 92480 11702 92486 11766
rect 92550 11702 92556 11766
rect 92480 11696 92556 11702
rect 92208 11022 92214 11086
rect 92278 11022 92284 11086
rect 92208 11016 92284 11022
rect 92893 1702 92959 1703
rect 92893 1670 92894 1702
rect 92888 1638 92894 1670
rect 92958 1670 92959 1702
rect 92958 1638 92964 1670
rect 92888 1294 92964 1638
rect 92888 1230 92894 1294
rect 92958 1230 92964 1294
rect 92888 1224 92964 1230
rect 94384 0 94460 13062
rect 94792 12038 94868 13470
rect 94928 13262 95004 15102
rect 97376 15166 97452 15172
rect 97376 15102 97382 15166
rect 97446 15102 97452 15166
rect 97512 15166 97588 17006
rect 97512 15134 97518 15166
rect 97245 14350 97311 14351
rect 97245 14318 97246 14350
rect 97240 14286 97246 14318
rect 97310 14318 97311 14350
rect 97310 14286 97316 14318
rect 97240 13670 97316 14286
rect 97240 13606 97246 13670
rect 97310 13606 97316 13670
rect 97240 13600 97316 13606
rect 94928 13230 94934 13262
rect 94933 13198 94934 13230
rect 94998 13230 95004 13262
rect 97240 13534 97316 13540
rect 97240 13470 97246 13534
rect 97310 13470 97316 13534
rect 94998 13198 94999 13230
rect 94933 13197 94999 13198
rect 94928 13126 95004 13132
rect 94928 13062 94934 13126
rect 94998 13062 95004 13126
rect 96837 13126 96903 13127
rect 96837 13094 96838 13126
rect 94928 12582 95004 13062
rect 94928 12550 94934 12582
rect 94933 12518 94934 12550
rect 94998 12550 95004 12582
rect 96832 13062 96838 13094
rect 96902 13094 96903 13126
rect 96902 13062 96908 13094
rect 94998 12518 94999 12550
rect 94933 12517 94999 12518
rect 94933 12310 94999 12311
rect 94933 12278 94934 12310
rect 94792 12006 94798 12038
rect 94797 11974 94798 12006
rect 94862 12006 94868 12038
rect 94928 12246 94934 12278
rect 94998 12278 94999 12310
rect 94998 12246 95004 12278
rect 94862 11974 94863 12006
rect 94797 11973 94863 11974
rect 94661 11902 94727 11903
rect 94661 11870 94662 11902
rect 94656 11838 94662 11870
rect 94726 11870 94727 11902
rect 94726 11838 94732 11870
rect 94656 11086 94732 11838
rect 94928 11766 95004 12246
rect 94928 11702 94934 11766
rect 94998 11702 95004 11766
rect 94928 11696 95004 11702
rect 94656 11022 94662 11086
rect 94726 11022 94732 11086
rect 94656 11016 94732 11022
rect 94661 1702 94727 1703
rect 94661 1670 94662 1702
rect 94656 1638 94662 1670
rect 94726 1670 94727 1702
rect 96157 1702 96223 1703
rect 96157 1670 96158 1702
rect 94726 1638 94732 1670
rect 94656 1294 94732 1638
rect 94656 1230 94662 1294
rect 94726 1230 94732 1294
rect 94656 1224 94732 1230
rect 96152 1638 96158 1670
rect 96222 1670 96223 1702
rect 96222 1638 96228 1670
rect 96152 1294 96228 1638
rect 96152 1230 96158 1294
rect 96222 1230 96228 1294
rect 96152 1224 96228 1230
rect 96832 0 96908 13062
rect 97240 12038 97316 13470
rect 97376 13262 97452 15102
rect 97517 15102 97518 15134
rect 97582 15134 97588 15166
rect 99824 17070 99900 17076
rect 99824 17006 99830 17070
rect 99894 17006 99900 17070
rect 99824 15166 99900 17006
rect 102272 17070 102484 17076
rect 102272 17006 102414 17070
rect 102478 17006 102484 17070
rect 102272 17000 102484 17006
rect 104992 17070 105068 17076
rect 104992 17006 104998 17070
rect 105062 17006 105068 17070
rect 99824 15134 99830 15166
rect 97582 15102 97583 15134
rect 97517 15101 97583 15102
rect 99829 15102 99830 15134
rect 99894 15134 99900 15166
rect 99960 15166 100036 15172
rect 99894 15102 99895 15134
rect 99829 15101 99895 15102
rect 99960 15102 99966 15166
rect 100030 15102 100036 15166
rect 102272 15166 102348 17000
rect 102272 15134 102278 15166
rect 99693 14350 99759 14351
rect 99693 14318 99694 14350
rect 99688 14286 99694 14318
rect 99758 14318 99759 14350
rect 99758 14286 99764 14318
rect 99688 13670 99764 14286
rect 99688 13606 99694 13670
rect 99758 13606 99764 13670
rect 99688 13600 99764 13606
rect 97376 13230 97382 13262
rect 97381 13198 97382 13230
rect 97446 13230 97452 13262
rect 99824 13534 99900 13540
rect 99824 13470 99830 13534
rect 99894 13470 99900 13534
rect 97446 13198 97447 13230
rect 97381 13197 97447 13198
rect 97376 13126 97452 13132
rect 97376 13062 97382 13126
rect 97446 13062 97452 13126
rect 99421 13126 99487 13127
rect 99421 13094 99422 13126
rect 97376 12582 97452 13062
rect 97376 12550 97382 12582
rect 97381 12518 97382 12550
rect 97446 12550 97452 12582
rect 99416 13062 99422 13094
rect 99486 13094 99487 13126
rect 99688 13126 99764 13132
rect 99486 13062 99492 13094
rect 97446 12518 97447 12550
rect 97381 12517 97447 12518
rect 97381 12310 97447 12311
rect 97381 12278 97382 12310
rect 97240 12006 97246 12038
rect 97245 11974 97246 12006
rect 97310 12006 97316 12038
rect 97376 12246 97382 12278
rect 97446 12278 97447 12310
rect 97446 12246 97452 12278
rect 97310 11974 97311 12006
rect 97245 11973 97311 11974
rect 97109 11902 97175 11903
rect 97109 11870 97110 11902
rect 97104 11838 97110 11870
rect 97174 11870 97175 11902
rect 97174 11838 97180 11870
rect 97104 11086 97180 11838
rect 97376 11766 97452 12246
rect 97376 11702 97382 11766
rect 97446 11702 97452 11766
rect 97376 11696 97452 11702
rect 97104 11022 97110 11086
rect 97174 11022 97180 11086
rect 97104 11016 97180 11022
rect 97925 1702 97991 1703
rect 97925 1670 97926 1702
rect 97920 1638 97926 1670
rect 97990 1670 97991 1702
rect 97990 1638 97996 1670
rect 97920 1294 97996 1638
rect 97920 1230 97926 1294
rect 97990 1230 97996 1294
rect 97920 1224 97996 1230
rect 99416 0 99492 13062
rect 99688 13062 99694 13126
rect 99758 13062 99764 13126
rect 99688 12582 99764 13062
rect 99688 12550 99694 12582
rect 99693 12518 99694 12550
rect 99758 12550 99764 12582
rect 99758 12518 99759 12550
rect 99693 12517 99759 12518
rect 99693 12310 99759 12311
rect 99693 12278 99694 12310
rect 99688 12246 99694 12278
rect 99758 12278 99759 12310
rect 99758 12246 99764 12278
rect 99557 11902 99623 11903
rect 99557 11870 99558 11902
rect 99552 11838 99558 11870
rect 99622 11870 99623 11902
rect 99622 11838 99628 11870
rect 99552 11086 99628 11838
rect 99688 11766 99764 12246
rect 99824 12038 99900 13470
rect 99960 13262 100036 15102
rect 102277 15102 102278 15134
rect 102342 15134 102348 15166
rect 102408 15166 102484 15172
rect 102342 15102 102343 15134
rect 102277 15101 102343 15102
rect 102408 15102 102414 15166
rect 102478 15102 102484 15166
rect 102277 14350 102343 14351
rect 102277 14318 102278 14350
rect 102272 14286 102278 14318
rect 102342 14318 102343 14350
rect 102342 14286 102348 14318
rect 102272 13670 102348 14286
rect 102272 13606 102278 13670
rect 102342 13606 102348 13670
rect 102272 13600 102348 13606
rect 99960 13230 99966 13262
rect 99965 13198 99966 13230
rect 100030 13230 100036 13262
rect 102272 13534 102348 13540
rect 102272 13470 102278 13534
rect 102342 13470 102348 13534
rect 100030 13198 100031 13230
rect 99965 13197 100031 13198
rect 101869 13126 101935 13127
rect 101869 13094 101870 13126
rect 99824 12006 99830 12038
rect 99829 11974 99830 12006
rect 99894 12006 99900 12038
rect 101864 13062 101870 13094
rect 101934 13094 101935 13126
rect 101934 13062 101940 13094
rect 99894 11974 99895 12006
rect 99829 11973 99895 11974
rect 99688 11702 99694 11766
rect 99758 11702 99764 11766
rect 99688 11696 99764 11702
rect 99552 11022 99558 11086
rect 99622 11022 99628 11086
rect 99552 11016 99628 11022
rect 99693 1702 99759 1703
rect 99693 1670 99694 1702
rect 99688 1638 99694 1670
rect 99758 1670 99759 1702
rect 101189 1702 101255 1703
rect 101189 1670 101190 1702
rect 99758 1638 99764 1670
rect 99688 1294 99764 1638
rect 99688 1230 99694 1294
rect 99758 1230 99764 1294
rect 99688 1224 99764 1230
rect 101184 1638 101190 1670
rect 101254 1670 101255 1702
rect 101254 1638 101260 1670
rect 101184 1294 101260 1638
rect 101184 1230 101190 1294
rect 101254 1230 101260 1294
rect 101184 1224 101260 1230
rect 101864 0 101940 13062
rect 102005 12310 102071 12311
rect 102005 12278 102006 12310
rect 102000 12246 102006 12278
rect 102070 12278 102071 12310
rect 102070 12246 102076 12278
rect 102000 11766 102076 12246
rect 102272 12038 102348 13470
rect 102408 13262 102484 15102
rect 104856 15166 104932 15172
rect 104856 15102 104862 15166
rect 104926 15102 104932 15166
rect 104992 15166 105068 17006
rect 104992 15134 104998 15166
rect 104725 14350 104791 14351
rect 104725 14318 104726 14350
rect 104720 14286 104726 14318
rect 104790 14318 104791 14350
rect 104790 14286 104796 14318
rect 104720 13670 104796 14286
rect 104720 13606 104726 13670
rect 104790 13606 104796 13670
rect 104720 13600 104796 13606
rect 102408 13230 102414 13262
rect 102413 13198 102414 13230
rect 102478 13230 102484 13262
rect 104720 13534 104796 13540
rect 104720 13470 104726 13534
rect 104790 13470 104796 13534
rect 102478 13198 102479 13230
rect 102413 13197 102479 13198
rect 102408 13126 102484 13132
rect 102408 13062 102414 13126
rect 102478 13062 102484 13126
rect 104317 13126 104383 13127
rect 104317 13094 104318 13126
rect 102408 12582 102484 13062
rect 102408 12550 102414 12582
rect 102413 12518 102414 12550
rect 102478 12550 102484 12582
rect 104312 13062 104318 13094
rect 104382 13094 104383 13126
rect 104382 13062 104388 13094
rect 102478 12518 102479 12550
rect 102413 12517 102479 12518
rect 102272 12006 102278 12038
rect 102277 11974 102278 12006
rect 102342 12006 102348 12038
rect 102342 11974 102343 12006
rect 102277 11973 102343 11974
rect 102141 11902 102207 11903
rect 102141 11870 102142 11902
rect 102000 11702 102006 11766
rect 102070 11702 102076 11766
rect 102000 11696 102076 11702
rect 102136 11838 102142 11870
rect 102206 11870 102207 11902
rect 102206 11838 102212 11870
rect 102136 11086 102212 11838
rect 102136 11022 102142 11086
rect 102206 11022 102212 11086
rect 102136 11016 102212 11022
rect 102957 1702 103023 1703
rect 102957 1670 102958 1702
rect 102952 1638 102958 1670
rect 103022 1670 103023 1702
rect 103022 1638 103028 1670
rect 102952 1294 103028 1638
rect 102952 1230 102958 1294
rect 103022 1230 103028 1294
rect 102952 1224 103028 1230
rect 104312 0 104388 13062
rect 104453 12310 104519 12311
rect 104453 12278 104454 12310
rect 104448 12246 104454 12278
rect 104518 12278 104519 12310
rect 104518 12246 104524 12278
rect 104448 11766 104524 12246
rect 104720 12038 104796 13470
rect 104856 13262 104932 15102
rect 104997 15102 104998 15134
rect 105062 15134 105068 15166
rect 107304 17070 107380 17076
rect 107304 17006 107310 17070
rect 107374 17006 107380 17070
rect 107304 15166 107380 17006
rect 124168 15710 124244 18366
rect 124304 17070 124380 19726
rect 124304 17038 124310 17070
rect 124309 17006 124310 17038
rect 124374 17038 124380 17070
rect 137496 18838 137844 20406
rect 137496 18774 137502 18838
rect 137566 18774 137844 18838
rect 137496 17070 137844 18774
rect 124374 17006 124375 17038
rect 124309 17005 124375 17006
rect 137496 17006 137502 17070
rect 137566 17006 137844 17070
rect 124168 15646 124174 15710
rect 124238 15646 124244 15710
rect 124168 15640 124244 15646
rect 124440 16934 124516 16940
rect 124440 16870 124446 16934
rect 124510 16870 124516 16934
rect 124304 15574 124380 15580
rect 124304 15510 124310 15574
rect 124374 15510 124380 15574
rect 107304 15134 107310 15166
rect 105062 15102 105063 15134
rect 104997 15101 105063 15102
rect 107309 15102 107310 15134
rect 107374 15134 107380 15166
rect 107440 15166 107516 15172
rect 107374 15102 107375 15134
rect 107309 15101 107375 15102
rect 107440 15102 107446 15166
rect 107510 15102 107516 15166
rect 107309 14350 107375 14351
rect 107309 14318 107310 14350
rect 107304 14286 107310 14318
rect 107374 14318 107375 14350
rect 107374 14286 107380 14318
rect 107304 13670 107380 14286
rect 107304 13606 107310 13670
rect 107374 13606 107380 13670
rect 107304 13600 107380 13606
rect 104856 13230 104862 13262
rect 104861 13198 104862 13230
rect 104926 13230 104932 13262
rect 107304 13534 107380 13540
rect 107304 13470 107310 13534
rect 107374 13470 107380 13534
rect 104926 13198 104927 13230
rect 104861 13197 104927 13198
rect 104856 13126 104932 13132
rect 104856 13062 104862 13126
rect 104926 13062 104932 13126
rect 106901 13126 106967 13127
rect 106901 13094 106902 13126
rect 104856 12582 104932 13062
rect 104856 12550 104862 12582
rect 104861 12518 104862 12550
rect 104926 12550 104932 12582
rect 106896 13062 106902 13094
rect 106966 13094 106967 13126
rect 106966 13062 106972 13094
rect 104926 12518 104927 12550
rect 104861 12517 104927 12518
rect 104720 12006 104726 12038
rect 104725 11974 104726 12006
rect 104790 12006 104796 12038
rect 104790 11974 104791 12006
rect 104725 11973 104791 11974
rect 104589 11902 104655 11903
rect 104589 11870 104590 11902
rect 104448 11702 104454 11766
rect 104518 11702 104524 11766
rect 104448 11696 104524 11702
rect 104584 11838 104590 11870
rect 104654 11870 104655 11902
rect 104654 11838 104660 11870
rect 104584 11086 104660 11838
rect 104584 11022 104590 11086
rect 104654 11022 104660 11086
rect 104584 11016 104660 11022
rect 104589 1702 104655 1703
rect 104589 1670 104590 1702
rect 104584 1638 104590 1670
rect 104654 1670 104655 1702
rect 106221 1702 106287 1703
rect 106221 1670 106222 1702
rect 104654 1638 104660 1670
rect 104584 1294 104660 1638
rect 104584 1230 104590 1294
rect 104654 1230 104660 1294
rect 104584 1224 104660 1230
rect 106216 1638 106222 1670
rect 106286 1670 106287 1702
rect 106286 1638 106292 1670
rect 106216 1294 106292 1638
rect 106216 1230 106222 1294
rect 106286 1230 106292 1294
rect 106216 1224 106292 1230
rect 106896 0 106972 13062
rect 107304 12038 107380 13470
rect 107440 13262 107516 15102
rect 124173 14078 124239 14079
rect 124173 14046 124174 14078
rect 107440 13230 107446 13262
rect 107445 13198 107446 13230
rect 107510 13230 107516 13262
rect 124168 14014 124174 14046
rect 124238 14046 124239 14078
rect 124238 14014 124244 14046
rect 107510 13198 107511 13230
rect 107445 13197 107511 13198
rect 107440 13126 107516 13132
rect 107440 13062 107446 13126
rect 107510 13062 107516 13126
rect 107440 12582 107516 13062
rect 107440 12550 107446 12582
rect 107445 12518 107446 12550
rect 107510 12550 107516 12582
rect 107510 12518 107511 12550
rect 107445 12517 107511 12518
rect 107445 12310 107511 12311
rect 107445 12278 107446 12310
rect 107304 12006 107310 12038
rect 107309 11974 107310 12006
rect 107374 12006 107380 12038
rect 107440 12246 107446 12278
rect 107510 12278 107511 12310
rect 107510 12246 107516 12278
rect 107374 11974 107375 12006
rect 107309 11973 107375 11974
rect 107173 11902 107239 11903
rect 107173 11870 107174 11902
rect 107168 11838 107174 11870
rect 107238 11870 107239 11902
rect 107238 11838 107244 11870
rect 107168 11086 107244 11838
rect 107440 11766 107516 12246
rect 107440 11702 107446 11766
rect 107510 11702 107516 11766
rect 107440 11696 107516 11702
rect 124168 11494 124244 14014
rect 124304 12854 124380 15510
rect 124440 14350 124516 16870
rect 124440 14318 124446 14350
rect 124445 14286 124446 14318
rect 124510 14318 124516 14350
rect 137496 15574 137844 17006
rect 137496 15510 137502 15574
rect 137566 15510 137844 15574
rect 124510 14286 124511 14318
rect 124445 14285 124511 14286
rect 137496 13942 137844 15510
rect 137496 13878 137502 13942
rect 137566 13878 137844 13942
rect 124853 13534 124919 13535
rect 124853 13502 124854 13534
rect 124304 12822 124310 12854
rect 124309 12790 124310 12822
rect 124374 12822 124380 12854
rect 124848 13470 124854 13502
rect 124918 13502 124919 13534
rect 124918 13470 124924 13502
rect 124374 12790 124375 12822
rect 124309 12789 124375 12790
rect 124309 12718 124375 12719
rect 124309 12686 124310 12718
rect 124168 11430 124174 11494
rect 124238 11430 124244 11494
rect 124168 11424 124244 11430
rect 124304 12654 124310 12686
rect 124374 12686 124375 12718
rect 124374 12654 124380 12686
rect 109349 11358 109415 11359
rect 109349 11326 109350 11358
rect 109344 11294 109350 11326
rect 109414 11326 109415 11358
rect 124168 11358 124244 11364
rect 109414 11294 109420 11326
rect 107168 11022 107174 11086
rect 107238 11022 107244 11086
rect 109213 11086 109279 11087
rect 109213 11054 109214 11086
rect 107168 11016 107244 11022
rect 109208 11022 109214 11054
rect 109278 11054 109279 11086
rect 109278 11022 109284 11054
rect 109208 10678 109284 11022
rect 109208 10614 109214 10678
rect 109278 10614 109284 10678
rect 109208 10608 109284 10614
rect 109344 9590 109420 11294
rect 109344 9526 109350 9590
rect 109414 9526 109420 9590
rect 109344 9520 109420 9526
rect 124168 11294 124174 11358
rect 124238 11294 124244 11358
rect 124168 8638 124244 11294
rect 124304 9998 124380 12654
rect 124445 11902 124511 11903
rect 124445 11870 124446 11902
rect 124304 9934 124310 9998
rect 124374 9934 124380 9998
rect 124304 9928 124380 9934
rect 124440 11838 124446 11870
rect 124510 11870 124511 11902
rect 124510 11838 124516 11870
rect 124168 8606 124174 8638
rect 124173 8574 124174 8606
rect 124238 8606 124244 8638
rect 124238 8574 124239 8606
rect 124173 8573 124239 8574
rect 107853 1702 107919 1703
rect 107853 1670 107854 1702
rect 107848 1638 107854 1670
rect 107918 1670 107919 1702
rect 109621 1702 109687 1703
rect 109621 1670 109622 1702
rect 107918 1638 107924 1670
rect 107848 1294 107924 1638
rect 107848 1230 107854 1294
rect 107918 1230 107924 1294
rect 107848 1224 107924 1230
rect 109616 1638 109622 1670
rect 109686 1670 109687 1702
rect 111389 1702 111455 1703
rect 111389 1670 111390 1702
rect 109686 1638 109692 1670
rect 109616 1294 109692 1638
rect 109616 1230 109622 1294
rect 109686 1230 109692 1294
rect 109616 1224 109692 1230
rect 111384 1638 111390 1670
rect 111454 1670 111455 1702
rect 112885 1702 112951 1703
rect 112885 1670 112886 1702
rect 111454 1638 111460 1670
rect 111384 1294 111460 1638
rect 111384 1230 111390 1294
rect 111454 1230 111460 1294
rect 111384 1224 111460 1230
rect 112880 1638 112886 1670
rect 112950 1670 112951 1702
rect 114653 1702 114719 1703
rect 114653 1670 114654 1702
rect 112950 1638 112956 1670
rect 112880 1294 112956 1638
rect 112880 1230 112886 1294
rect 112950 1230 112956 1294
rect 112880 1224 112956 1230
rect 114648 1638 114654 1670
rect 114718 1670 114719 1702
rect 116285 1702 116351 1703
rect 116285 1670 116286 1702
rect 114718 1638 114724 1670
rect 114648 1294 114724 1638
rect 114648 1230 114654 1294
rect 114718 1230 114724 1294
rect 114648 1224 114724 1230
rect 116280 1638 116286 1670
rect 116350 1670 116351 1702
rect 118053 1702 118119 1703
rect 118053 1670 118054 1702
rect 116350 1638 116356 1670
rect 116280 1294 116356 1638
rect 116280 1230 116286 1294
rect 116350 1230 116356 1294
rect 116280 1224 116356 1230
rect 118048 1638 118054 1670
rect 118118 1670 118119 1702
rect 119685 1702 119751 1703
rect 119685 1670 119686 1702
rect 118118 1638 118124 1670
rect 118048 1294 118124 1638
rect 118048 1230 118054 1294
rect 118118 1230 118124 1294
rect 118048 1224 118124 1230
rect 119680 1638 119686 1670
rect 119750 1670 119751 1702
rect 121453 1702 121519 1703
rect 121453 1670 121454 1702
rect 119750 1638 119756 1670
rect 119680 1294 119756 1638
rect 119680 1230 119686 1294
rect 119750 1230 119756 1294
rect 119680 1224 119756 1230
rect 121448 1638 121454 1670
rect 121518 1670 121519 1702
rect 122949 1702 123015 1703
rect 122949 1670 122950 1702
rect 121518 1638 121524 1670
rect 121448 1294 121524 1638
rect 121448 1230 121454 1294
rect 121518 1230 121524 1294
rect 121448 1224 121524 1230
rect 122944 1638 122950 1670
rect 123014 1670 123015 1702
rect 123014 1638 123020 1670
rect 122944 1294 123020 1638
rect 122944 1230 122950 1294
rect 123014 1230 123020 1294
rect 122944 1224 123020 1230
rect 124440 0 124516 11838
rect 124581 10814 124647 10815
rect 124581 10782 124582 10814
rect 124576 10750 124582 10782
rect 124646 10782 124647 10814
rect 124646 10750 124652 10782
rect 124576 0 124652 10750
rect 124717 9046 124783 9047
rect 124717 9014 124718 9046
rect 124712 8982 124718 9014
rect 124782 9014 124783 9046
rect 124782 8982 124788 9014
rect 124712 0 124788 8982
rect 124848 0 124924 13470
rect 137496 12038 137844 13878
rect 137496 11974 137502 12038
rect 137566 11974 137844 12038
rect 137496 10542 137844 11974
rect 137496 10478 137502 10542
rect 137566 10478 137844 10542
rect 137496 8774 137844 10478
rect 137496 8710 137502 8774
rect 137566 8710 137844 8774
rect 137496 7142 137844 8710
rect 137496 7078 137502 7142
rect 137566 7078 137844 7142
rect 137496 5510 137844 7078
rect 137496 5446 137502 5510
rect 137566 5446 137844 5510
rect 137496 3878 137844 5446
rect 137496 3814 137502 3878
rect 137566 3814 137844 3878
rect 125125 1702 125191 1703
rect 125125 1670 125126 1702
rect 125120 1638 125126 1670
rect 125190 1670 125191 1702
rect 126349 1702 126415 1703
rect 126349 1670 126350 1702
rect 125190 1638 125196 1670
rect 125120 1294 125196 1638
rect 125120 1230 125126 1294
rect 125190 1230 125196 1294
rect 125120 1224 125196 1230
rect 126344 1638 126350 1670
rect 126414 1670 126415 1702
rect 128117 1702 128183 1703
rect 128117 1670 128118 1702
rect 126414 1638 126420 1670
rect 126344 1294 126420 1638
rect 126344 1230 126350 1294
rect 126414 1230 126420 1294
rect 126344 1224 126420 1230
rect 128112 1638 128118 1670
rect 128182 1670 128183 1702
rect 129885 1702 129951 1703
rect 129885 1670 129886 1702
rect 128182 1638 128188 1670
rect 128112 1294 128188 1638
rect 128112 1230 128118 1294
rect 128182 1230 128188 1294
rect 128112 1224 128188 1230
rect 129880 1638 129886 1670
rect 129950 1670 129951 1702
rect 131381 1702 131447 1703
rect 131381 1670 131382 1702
rect 129950 1638 129956 1670
rect 129880 1294 129956 1638
rect 129880 1230 129886 1294
rect 129950 1230 129956 1294
rect 129880 1224 129956 1230
rect 131376 1638 131382 1670
rect 131446 1670 131447 1702
rect 133149 1702 133215 1703
rect 133149 1670 133150 1702
rect 131446 1638 131452 1670
rect 131376 1294 131452 1638
rect 131376 1230 131382 1294
rect 131446 1230 131452 1294
rect 131376 1224 131452 1230
rect 133144 1638 133150 1670
rect 133214 1670 133215 1702
rect 134781 1702 134847 1703
rect 134781 1670 134782 1702
rect 133214 1638 133220 1670
rect 133144 1294 133220 1638
rect 133144 1230 133150 1294
rect 133214 1230 133220 1294
rect 133144 1224 133220 1230
rect 134776 1638 134782 1670
rect 134846 1670 134847 1702
rect 136549 1702 136615 1703
rect 136549 1670 136550 1702
rect 134846 1638 134852 1670
rect 134776 1294 134852 1638
rect 134776 1230 134782 1294
rect 134846 1230 134852 1294
rect 134776 1224 134852 1230
rect 136544 1638 136550 1670
rect 136614 1670 136615 1702
rect 136614 1638 136620 1670
rect 136544 1294 136620 1638
rect 136544 1230 136550 1294
rect 136614 1230 136620 1294
rect 136544 1224 136620 1230
rect 137496 1294 137844 3814
rect 137496 1230 137502 1294
rect 137566 1230 137638 1294
rect 137702 1230 137774 1294
rect 137838 1230 137844 1294
rect 137496 1158 137844 1230
rect 137496 1094 137502 1158
rect 137566 1094 137638 1158
rect 137702 1094 137774 1158
rect 137838 1094 137844 1158
rect 137496 1022 137844 1094
rect 137496 958 137502 1022
rect 137566 958 137638 1022
rect 137702 958 137774 1022
rect 137838 958 137844 1022
rect 137496 952 137844 958
rect 138176 130494 138524 133150
rect 138176 130430 138182 130494
rect 138246 130430 138524 130494
rect 138176 123422 138524 130430
rect 138176 123358 138182 123422
rect 138246 123358 138524 123422
rect 138176 114854 138524 123358
rect 138176 114790 138182 114854
rect 138246 114790 138524 114854
rect 138176 614 138524 114790
rect 138176 550 138182 614
rect 138246 550 138318 614
rect 138382 550 138454 614
rect 138518 550 138524 614
rect 138176 478 138524 550
rect 138176 414 138182 478
rect 138246 414 138318 478
rect 138382 414 138454 478
rect 138518 414 138524 478
rect 138176 342 138524 414
rect 138176 278 138182 342
rect 138246 278 138318 342
rect 138382 278 138454 342
rect 138518 278 138524 342
rect 138176 272 138524 278
use contact_39  contact_39_5
timestamp 1624857261
transform 1 0 408 0 1 413
box 0 0 192 192
use contact_39  contact_39_9
timestamp 1624857261
transform 1 0 544 0 1 549
box 0 0 192 192
use contact_39  contact_39_13
timestamp 1624857261
transform 1 0 272 0 1 549
box 0 0 192 192
use contact_39  contact_39_23
timestamp 1624857261
transform 1 0 408 0 1 549
box 0 0 192 192
use contact_39  contact_39_26
timestamp 1624857261
transform 1 0 272 0 1 277
box 0 0 192 192
use contact_39  contact_39_28
timestamp 1624857261
transform 1 0 544 0 1 413
box 0 0 192 192
use contact_39  contact_39_29
timestamp 1624857261
transform 1 0 408 0 1 277
box 0 0 192 192
use contact_39  contact_39_31
timestamp 1624857261
transform 1 0 544 0 1 277
box 0 0 192 192
use contact_39  contact_39_35
timestamp 1624857261
transform 1 0 272 0 1 413
box 0 0 192 192
use contact_33  contact_33_2303
timestamp 1624857261
transform 1 0 19312 0 1 549
box 0 0 1 1
use contact_39  contact_39_42
timestamp 1624857261
transform 1 0 952 0 1 1093
box 0 0 192 192
use contact_39  contact_39_48
timestamp 1624857261
transform 1 0 1088 0 1 1093
box 0 0 192 192
use contact_39  contact_39_60
timestamp 1624857261
transform 1 0 952 0 1 957
box 0 0 192 192
use contact_39  contact_39_70
timestamp 1624857261
transform 1 0 1088 0 1 957
box 0 0 192 192
use contact_39  contact_39_41
timestamp 1624857261
transform 1 0 1224 0 1 957
box 0 0 192 192
use contact_39  contact_39_64
timestamp 1624857261
transform 1 0 1224 0 1 1093
box 0 0 192 192
use contact_39  contact_39_63
timestamp 1624857261
transform 1 0 1088 0 1 1229
box 0 0 192 192
use contact_39  contact_39_65
timestamp 1624857261
transform 1 0 952 0 1 1229
box 0 0 192 192
use contact_39  contact_39_57
timestamp 1624857261
transform 1 0 1224 0 1 1229
box 0 0 192 192
use contact_33  contact_33_5294
timestamp 1624857261
transform 1 0 2040 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5290
timestamp 1624857261
transform 1 0 3808 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5284
timestamp 1624857261
transform 1 0 5440 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5282
timestamp 1624857261
transform 1 0 7208 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5278
timestamp 1624857261
transform 1 0 8704 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5274
timestamp 1624857261
transform 1 0 10472 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5270
timestamp 1624857261
transform 1 0 12104 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5266
timestamp 1624857261
transform 1 0 13872 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5242
timestamp 1624857261
transform 1 0 15640 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5236
timestamp 1624857261
transform 1 0 17136 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5228
timestamp 1624857261
transform 1 0 19040 0 1 1229
box 0 0 1 1
use contact_33  contact_33_5200
timestamp 1624857261
transform 1 0 20536 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4904
timestamp 1624857261
transform 1 0 22168 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4326
timestamp 1624857261
transform 1 0 23936 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4322
timestamp 1624857261
transform 1 0 25704 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4314
timestamp 1624857261
transform 1 0 27200 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4310
timestamp 1624857261
transform 1 0 28832 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4284
timestamp 1624857261
transform 1 0 30464 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4266
timestamp 1624857261
transform 1 0 32232 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4258
timestamp 1624857261
transform 1 0 34272 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4230
timestamp 1624857261
transform 1 0 35632 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4210
timestamp 1624857261
transform 1 0 37264 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4200
timestamp 1624857261
transform 1 0 39032 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4178
timestamp 1624857261
transform 1 0 40664 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4160
timestamp 1624857261
transform 1 0 42432 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4140
timestamp 1624857261
transform 1 0 44064 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4122
timestamp 1624857261
transform 1 0 45696 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4102
timestamp 1624857261
transform 1 0 47464 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4088
timestamp 1624857261
transform 1 0 48960 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4064
timestamp 1624857261
transform 1 0 50728 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4048
timestamp 1624857261
transform 1 0 52496 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4036
timestamp 1624857261
transform 1 0 54128 0 1 1229
box 0 0 1 1
use contact_33  contact_33_4012
timestamp 1624857261
transform 1 0 55896 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3986
timestamp 1624857261
transform 1 0 57392 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3974
timestamp 1624857261
transform 1 0 59160 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3958
timestamp 1624857261
transform 1 0 60928 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3936
timestamp 1624857261
transform 1 0 62696 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3920
timestamp 1624857261
transform 1 0 64192 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3900
timestamp 1624857261
transform 1 0 65824 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3882
timestamp 1624857261
transform 1 0 67592 0 1 1229
box 0 0 1 1
use contact_38  contact_38_3
timestamp 1624857261
transform 1 0 1730 0 1 1628
box 0 0 192 192
use contact_7  contact_7_317
timestamp 1624857261
transform 1 0 2129 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1573
timestamp 1624857261
transform 1 0 2133 0 1 1691
box 0 0 1 1
use contact_19  contact_19_933
timestamp 1624857261
transform 1 0 2130 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1573
timestamp 1624857261
transform 1 0 2137 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5295
timestamp 1624857261
transform 1 0 2040 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1571
timestamp 1624857261
transform 1 0 2805 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1572
timestamp 1624857261
transform 1 0 2469 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1571
timestamp 1624857261
transform 1 0 2809 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1572
timestamp 1624857261
transform 1 0 2473 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1570
timestamp 1624857261
transform 1 0 3141 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1570
timestamp 1624857261
transform 1 0 3145 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1569
timestamp 1624857261
transform 1 0 3477 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1569
timestamp 1624857261
transform 1 0 3481 0 1 1683
box 0 0 1 1
use contact_7  contact_7_316
timestamp 1624857261
transform 1 0 3809 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1568
timestamp 1624857261
transform 1 0 3813 0 1 1691
box 0 0 1 1
use contact_19  contact_19_932
timestamp 1624857261
transform 1 0 3810 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1568
timestamp 1624857261
transform 1 0 3817 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5291
timestamp 1624857261
transform 1 0 3808 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1566
timestamp 1624857261
transform 1 0 4485 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1567
timestamp 1624857261
transform 1 0 4149 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1566
timestamp 1624857261
transform 1 0 4489 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1567
timestamp 1624857261
transform 1 0 4153 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1565
timestamp 1624857261
transform 1 0 4821 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1565
timestamp 1624857261
transform 1 0 4825 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1564
timestamp 1624857261
transform 1 0 5157 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1564
timestamp 1624857261
transform 1 0 5161 0 1 1683
box 0 0 1 1
use contact_7  contact_7_315
timestamp 1624857261
transform 1 0 5489 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1563
timestamp 1624857261
transform 1 0 5493 0 1 1691
box 0 0 1 1
use contact_19  contact_19_931
timestamp 1624857261
transform 1 0 5490 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1563
timestamp 1624857261
transform 1 0 5497 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5285
timestamp 1624857261
transform 1 0 5440 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1561
timestamp 1624857261
transform 1 0 6165 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1562
timestamp 1624857261
transform 1 0 5829 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1561
timestamp 1624857261
transform 1 0 6169 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1562
timestamp 1624857261
transform 1 0 5833 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1560
timestamp 1624857261
transform 1 0 6501 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1560
timestamp 1624857261
transform 1 0 6505 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1559
timestamp 1624857261
transform 1 0 6837 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1559
timestamp 1624857261
transform 1 0 6841 0 1 1683
box 0 0 1 1
use contact_7  contact_7_314
timestamp 1624857261
transform 1 0 7169 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1558
timestamp 1624857261
transform 1 0 7173 0 1 1691
box 0 0 1 1
use contact_19  contact_19_930
timestamp 1624857261
transform 1 0 7170 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1558
timestamp 1624857261
transform 1 0 7177 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5283
timestamp 1624857261
transform 1 0 7208 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1556
timestamp 1624857261
transform 1 0 7845 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1557
timestamp 1624857261
transform 1 0 7509 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1556
timestamp 1624857261
transform 1 0 7849 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1557
timestamp 1624857261
transform 1 0 7513 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1555
timestamp 1624857261
transform 1 0 8181 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1555
timestamp 1624857261
transform 1 0 8185 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1554
timestamp 1624857261
transform 1 0 8517 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1554
timestamp 1624857261
transform 1 0 8521 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5279
timestamp 1624857261
transform 1 0 8704 0 1 1637
box 0 0 1 1
use contact_7  contact_7_313
timestamp 1624857261
transform 1 0 8849 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1553
timestamp 1624857261
transform 1 0 8853 0 1 1691
box 0 0 1 1
use contact_19  contact_19_929
timestamp 1624857261
transform 1 0 8850 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1553
timestamp 1624857261
transform 1 0 8857 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1551
timestamp 1624857261
transform 1 0 9525 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1552
timestamp 1624857261
transform 1 0 9189 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1551
timestamp 1624857261
transform 1 0 9529 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1552
timestamp 1624857261
transform 1 0 9193 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1550
timestamp 1624857261
transform 1 0 9861 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1550
timestamp 1624857261
transform 1 0 9865 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1549
timestamp 1624857261
transform 1 0 10197 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1549
timestamp 1624857261
transform 1 0 10201 0 1 1683
box 0 0 1 1
use contact_7  contact_7_312
timestamp 1624857261
transform 1 0 10529 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1548
timestamp 1624857261
transform 1 0 10533 0 1 1691
box 0 0 1 1
use contact_19  contact_19_928
timestamp 1624857261
transform 1 0 10530 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1548
timestamp 1624857261
transform 1 0 10537 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5275
timestamp 1624857261
transform 1 0 10472 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1546
timestamp 1624857261
transform 1 0 11205 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1547
timestamp 1624857261
transform 1 0 10869 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1546
timestamp 1624857261
transform 1 0 11209 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1547
timestamp 1624857261
transform 1 0 10873 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1545
timestamp 1624857261
transform 1 0 11541 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1545
timestamp 1624857261
transform 1 0 11545 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1544
timestamp 1624857261
transform 1 0 11877 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1544
timestamp 1624857261
transform 1 0 11881 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5271
timestamp 1624857261
transform 1 0 12104 0 1 1637
box 0 0 1 1
use contact_7  contact_7_311
timestamp 1624857261
transform 1 0 12209 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1543
timestamp 1624857261
transform 1 0 12213 0 1 1691
box 0 0 1 1
use contact_19  contact_19_927
timestamp 1624857261
transform 1 0 12210 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1543
timestamp 1624857261
transform 1 0 12217 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1541
timestamp 1624857261
transform 1 0 12885 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1542
timestamp 1624857261
transform 1 0 12549 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1541
timestamp 1624857261
transform 1 0 12889 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1542
timestamp 1624857261
transform 1 0 12553 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1540
timestamp 1624857261
transform 1 0 13221 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1540
timestamp 1624857261
transform 1 0 13225 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1539
timestamp 1624857261
transform 1 0 13557 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1539
timestamp 1624857261
transform 1 0 13561 0 1 1683
box 0 0 1 1
use contact_7  contact_7_310
timestamp 1624857261
transform 1 0 13889 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1537
timestamp 1624857261
transform 1 0 14229 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1538
timestamp 1624857261
transform 1 0 13893 0 1 1691
box 0 0 1 1
use contact_19  contact_19_926
timestamp 1624857261
transform 1 0 13890 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1538
timestamp 1624857261
transform 1 0 13897 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5267
timestamp 1624857261
transform 1 0 13872 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1536
timestamp 1624857261
transform 1 0 14565 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1536
timestamp 1624857261
transform 1 0 14569 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1537
timestamp 1624857261
transform 1 0 14233 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1535
timestamp 1624857261
transform 1 0 14901 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1535
timestamp 1624857261
transform 1 0 14905 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1534
timestamp 1624857261
transform 1 0 15237 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1534
timestamp 1624857261
transform 1 0 15241 0 1 1683
box 0 0 1 1
use contact_7  contact_7_309
timestamp 1624857261
transform 1 0 15569 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1532
timestamp 1624857261
transform 1 0 15909 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1533
timestamp 1624857261
transform 1 0 15573 0 1 1691
box 0 0 1 1
use contact_19  contact_19_925
timestamp 1624857261
transform 1 0 15570 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1532
timestamp 1624857261
transform 1 0 15913 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1533
timestamp 1624857261
transform 1 0 15577 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5243
timestamp 1624857261
transform 1 0 15640 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1531
timestamp 1624857261
transform 1 0 16245 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1531
timestamp 1624857261
transform 1 0 16249 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1530
timestamp 1624857261
transform 1 0 16581 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1530
timestamp 1624857261
transform 1 0 16585 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1529
timestamp 1624857261
transform 1 0 16917 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1529
timestamp 1624857261
transform 1 0 16921 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5237
timestamp 1624857261
transform 1 0 17136 0 1 1637
box 0 0 1 1
use contact_7  contact_7_308
timestamp 1624857261
transform 1 0 17249 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1527
timestamp 1624857261
transform 1 0 17589 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1528
timestamp 1624857261
transform 1 0 17253 0 1 1691
box 0 0 1 1
use contact_19  contact_19_924
timestamp 1624857261
transform 1 0 17250 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1527
timestamp 1624857261
transform 1 0 17593 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1528
timestamp 1624857261
transform 1 0 17257 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1526
timestamp 1624857261
transform 1 0 17925 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1526
timestamp 1624857261
transform 1 0 17929 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1525
timestamp 1624857261
transform 1 0 18261 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1525
timestamp 1624857261
transform 1 0 18265 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1524
timestamp 1624857261
transform 1 0 18597 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1524
timestamp 1624857261
transform 1 0 18601 0 1 1683
box 0 0 1 1
use contact_7  contact_7_307
timestamp 1624857261
transform 1 0 18929 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1522
timestamp 1624857261
transform 1 0 19269 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1523
timestamp 1624857261
transform 1 0 18933 0 1 1691
box 0 0 1 1
use contact_19  contact_19_923
timestamp 1624857261
transform 1 0 18930 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1522
timestamp 1624857261
transform 1 0 19273 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1523
timestamp 1624857261
transform 1 0 18937 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5229
timestamp 1624857261
transform 1 0 19040 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1521
timestamp 1624857261
transform 1 0 19605 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1521
timestamp 1624857261
transform 1 0 19609 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1520
timestamp 1624857261
transform 1 0 19941 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1520
timestamp 1624857261
transform 1 0 19945 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1519
timestamp 1624857261
transform 1 0 20277 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1519
timestamp 1624857261
transform 1 0 20281 0 1 1683
box 0 0 1 1
use contact_33  contact_33_5201
timestamp 1624857261
transform 1 0 20536 0 1 1637
box 0 0 1 1
use contact_7  contact_7_306
timestamp 1624857261
transform 1 0 20609 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1517
timestamp 1624857261
transform 1 0 20949 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1518
timestamp 1624857261
transform 1 0 20613 0 1 1691
box 0 0 1 1
use contact_19  contact_19_922
timestamp 1624857261
transform 1 0 20610 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1517
timestamp 1624857261
transform 1 0 20953 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1518
timestamp 1624857261
transform 1 0 20617 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1516
timestamp 1624857261
transform 1 0 21285 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1516
timestamp 1624857261
transform 1 0 21289 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1515
timestamp 1624857261
transform 1 0 21621 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1515
timestamp 1624857261
transform 1 0 21625 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1514
timestamp 1624857261
transform 1 0 21957 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1514
timestamp 1624857261
transform 1 0 21961 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4905
timestamp 1624857261
transform 1 0 22168 0 1 1637
box 0 0 1 1
use contact_7  contact_7_305
timestamp 1624857261
transform 1 0 22289 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1512
timestamp 1624857261
transform 1 0 22629 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1513
timestamp 1624857261
transform 1 0 22293 0 1 1691
box 0 0 1 1
use contact_19  contact_19_921
timestamp 1624857261
transform 1 0 22290 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1512
timestamp 1624857261
transform 1 0 22633 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1513
timestamp 1624857261
transform 1 0 22297 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1511
timestamp 1624857261
transform 1 0 22965 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1511
timestamp 1624857261
transform 1 0 22969 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1510
timestamp 1624857261
transform 1 0 23301 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1510
timestamp 1624857261
transform 1 0 23305 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1509
timestamp 1624857261
transform 1 0 23637 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1509
timestamp 1624857261
transform 1 0 23641 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4327
timestamp 1624857261
transform 1 0 23936 0 1 1637
box 0 0 1 1
use contact_7  contact_7_304
timestamp 1624857261
transform 1 0 23969 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1507
timestamp 1624857261
transform 1 0 24309 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1508
timestamp 1624857261
transform 1 0 23973 0 1 1691
box 0 0 1 1
use contact_19  contact_19_920
timestamp 1624857261
transform 1 0 23970 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1507
timestamp 1624857261
transform 1 0 24313 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1508
timestamp 1624857261
transform 1 0 23977 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1506
timestamp 1624857261
transform 1 0 24645 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1506
timestamp 1624857261
transform 1 0 24649 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1505
timestamp 1624857261
transform 1 0 24981 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1505
timestamp 1624857261
transform 1 0 24985 0 1 1683
box 0 0 1 1
use contact_7  contact_7_303
timestamp 1624857261
transform 1 0 25649 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1504
timestamp 1624857261
transform 1 0 25317 0 1 1691
box 0 0 1 1
use contact_19  contact_19_919
timestamp 1624857261
transform 1 0 25650 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1504
timestamp 1624857261
transform 1 0 25321 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1502
timestamp 1624857261
transform 1 0 25989 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1503
timestamp 1624857261
transform 1 0 25653 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1502
timestamp 1624857261
transform 1 0 25993 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1503
timestamp 1624857261
transform 1 0 25657 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4323
timestamp 1624857261
transform 1 0 25704 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1501
timestamp 1624857261
transform 1 0 26325 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1501
timestamp 1624857261
transform 1 0 26329 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1500
timestamp 1624857261
transform 1 0 26661 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1500
timestamp 1624857261
transform 1 0 26665 0 1 1683
box 0 0 1 1
use contact_7  contact_7_302
timestamp 1624857261
transform 1 0 27329 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1498
timestamp 1624857261
transform 1 0 27333 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1499
timestamp 1624857261
transform 1 0 26997 0 1 1691
box 0 0 1 1
use contact_19  contact_19_918
timestamp 1624857261
transform 1 0 27330 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1498
timestamp 1624857261
transform 1 0 27337 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1499
timestamp 1624857261
transform 1 0 27001 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4315
timestamp 1624857261
transform 1 0 27200 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1497
timestamp 1624857261
transform 1 0 27669 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1497
timestamp 1624857261
transform 1 0 27673 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1496
timestamp 1624857261
transform 1 0 28005 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1496
timestamp 1624857261
transform 1 0 28009 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1495
timestamp 1624857261
transform 1 0 28341 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1495
timestamp 1624857261
transform 1 0 28345 0 1 1683
box 0 0 1 1
use contact_7  contact_7_301
timestamp 1624857261
transform 1 0 29009 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1493
timestamp 1624857261
transform 1 0 29013 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1494
timestamp 1624857261
transform 1 0 28677 0 1 1691
box 0 0 1 1
use contact_19  contact_19_917
timestamp 1624857261
transform 1 0 29010 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1493
timestamp 1624857261
transform 1 0 29017 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1494
timestamp 1624857261
transform 1 0 28681 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4311
timestamp 1624857261
transform 1 0 28832 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1492
timestamp 1624857261
transform 1 0 29349 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1492
timestamp 1624857261
transform 1 0 29353 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1491
timestamp 1624857261
transform 1 0 29685 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1491
timestamp 1624857261
transform 1 0 29689 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1490
timestamp 1624857261
transform 1 0 30021 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1490
timestamp 1624857261
transform 1 0 30025 0 1 1683
box 0 0 1 1
use contact_7  contact_7_300
timestamp 1624857261
transform 1 0 30689 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1488
timestamp 1624857261
transform 1 0 30693 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1489
timestamp 1624857261
transform 1 0 30357 0 1 1691
box 0 0 1 1
use contact_19  contact_19_916
timestamp 1624857261
transform 1 0 30690 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1488
timestamp 1624857261
transform 1 0 30697 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1489
timestamp 1624857261
transform 1 0 30361 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4285
timestamp 1624857261
transform 1 0 30464 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1487
timestamp 1624857261
transform 1 0 31029 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1487
timestamp 1624857261
transform 1 0 31033 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1486
timestamp 1624857261
transform 1 0 31365 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1486
timestamp 1624857261
transform 1 0 31369 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1485
timestamp 1624857261
transform 1 0 31701 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1485
timestamp 1624857261
transform 1 0 31705 0 1 1683
box 0 0 1 1
use contact_7  contact_7_299
timestamp 1624857261
transform 1 0 32369 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1483
timestamp 1624857261
transform 1 0 32373 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1484
timestamp 1624857261
transform 1 0 32037 0 1 1691
box 0 0 1 1
use contact_19  contact_19_915
timestamp 1624857261
transform 1 0 32370 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1483
timestamp 1624857261
transform 1 0 32377 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1484
timestamp 1624857261
transform 1 0 32041 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4267
timestamp 1624857261
transform 1 0 32232 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1482
timestamp 1624857261
transform 1 0 32709 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1482
timestamp 1624857261
transform 1 0 32713 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1481
timestamp 1624857261
transform 1 0 33045 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1481
timestamp 1624857261
transform 1 0 33049 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1480
timestamp 1624857261
transform 1 0 33381 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1480
timestamp 1624857261
transform 1 0 33385 0 1 1683
box 0 0 1 1
use contact_7  contact_7_298
timestamp 1624857261
transform 1 0 34049 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1478
timestamp 1624857261
transform 1 0 34053 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1479
timestamp 1624857261
transform 1 0 33717 0 1 1691
box 0 0 1 1
use contact_19  contact_19_914
timestamp 1624857261
transform 1 0 34050 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1478
timestamp 1624857261
transform 1 0 34057 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1479
timestamp 1624857261
transform 1 0 33721 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1477
timestamp 1624857261
transform 1 0 34389 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1477
timestamp 1624857261
transform 1 0 34393 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4259
timestamp 1624857261
transform 1 0 34272 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1476
timestamp 1624857261
transform 1 0 34725 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1476
timestamp 1624857261
transform 1 0 34729 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1475
timestamp 1624857261
transform 1 0 35061 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1475
timestamp 1624857261
transform 1 0 35065 0 1 1683
box 0 0 1 1
use contact_7  contact_7_297
timestamp 1624857261
transform 1 0 35729 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1473
timestamp 1624857261
transform 1 0 35733 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1474
timestamp 1624857261
transform 1 0 35397 0 1 1691
box 0 0 1 1
use contact_19  contact_19_913
timestamp 1624857261
transform 1 0 35730 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1473
timestamp 1624857261
transform 1 0 35737 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1474
timestamp 1624857261
transform 1 0 35401 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4231
timestamp 1624857261
transform 1 0 35632 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1472
timestamp 1624857261
transform 1 0 36069 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1472
timestamp 1624857261
transform 1 0 36073 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1471
timestamp 1624857261
transform 1 0 36405 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1471
timestamp 1624857261
transform 1 0 36409 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1470
timestamp 1624857261
transform 1 0 36741 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1470
timestamp 1624857261
transform 1 0 36745 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4222
timestamp 1624857261
transform 1 0 36720 0 1 1773
box 0 0 1 1
use contact_7  contact_7_296
timestamp 1624857261
transform 1 0 37409 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1468
timestamp 1624857261
transform 1 0 37413 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1469
timestamp 1624857261
transform 1 0 37077 0 1 1691
box 0 0 1 1
use contact_19  contact_19_912
timestamp 1624857261
transform 1 0 37410 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1468
timestamp 1624857261
transform 1 0 37417 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1469
timestamp 1624857261
transform 1 0 37081 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4211
timestamp 1624857261
transform 1 0 37264 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1467
timestamp 1624857261
transform 1 0 37749 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1467
timestamp 1624857261
transform 1 0 37753 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1466
timestamp 1624857261
transform 1 0 38085 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1466
timestamp 1624857261
transform 1 0 38089 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1464
timestamp 1624857261
transform 1 0 38757 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1465
timestamp 1624857261
transform 1 0 38421 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1464
timestamp 1624857261
transform 1 0 38761 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1465
timestamp 1624857261
transform 1 0 38425 0 1 1683
box 0 0 1 1
use contact_7  contact_7_295
timestamp 1624857261
transform 1 0 39089 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1463
timestamp 1624857261
transform 1 0 39093 0 1 1691
box 0 0 1 1
use contact_19  contact_19_911
timestamp 1624857261
transform 1 0 39090 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1463
timestamp 1624857261
transform 1 0 39097 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4201
timestamp 1624857261
transform 1 0 39032 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1462
timestamp 1624857261
transform 1 0 39429 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1462
timestamp 1624857261
transform 1 0 39433 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1461
timestamp 1624857261
transform 1 0 39765 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1461
timestamp 1624857261
transform 1 0 39769 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1459
timestamp 1624857261
transform 1 0 40437 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1460
timestamp 1624857261
transform 1 0 40101 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1459
timestamp 1624857261
transform 1 0 40441 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1460
timestamp 1624857261
transform 1 0 40105 0 1 1683
box 0 0 1 1
use contact_7  contact_7_294
timestamp 1624857261
transform 1 0 40769 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1458
timestamp 1624857261
transform 1 0 40773 0 1 1691
box 0 0 1 1
use contact_19  contact_19_910
timestamp 1624857261
transform 1 0 40770 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1458
timestamp 1624857261
transform 1 0 40777 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4179
timestamp 1624857261
transform 1 0 40664 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1457
timestamp 1624857261
transform 1 0 41109 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1457
timestamp 1624857261
transform 1 0 41113 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1456
timestamp 1624857261
transform 1 0 41445 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1456
timestamp 1624857261
transform 1 0 41449 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1454
timestamp 1624857261
transform 1 0 42117 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1455
timestamp 1624857261
transform 1 0 41781 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1454
timestamp 1624857261
transform 1 0 42121 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1455
timestamp 1624857261
transform 1 0 41785 0 1 1683
box 0 0 1 1
use contact_7  contact_7_293
timestamp 1624857261
transform 1 0 42449 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1453
timestamp 1624857261
transform 1 0 42453 0 1 1691
box 0 0 1 1
use contact_19  contact_19_909
timestamp 1624857261
transform 1 0 42450 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1453
timestamp 1624857261
transform 1 0 42457 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4161
timestamp 1624857261
transform 1 0 42432 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1452
timestamp 1624857261
transform 1 0 42789 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1452
timestamp 1624857261
transform 1 0 42793 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1451
timestamp 1624857261
transform 1 0 43125 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1451
timestamp 1624857261
transform 1 0 43129 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1449
timestamp 1624857261
transform 1 0 43797 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1450
timestamp 1624857261
transform 1 0 43461 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1449
timestamp 1624857261
transform 1 0 43801 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1450
timestamp 1624857261
transform 1 0 43465 0 1 1683
box 0 0 1 1
use contact_7  contact_7_292
timestamp 1624857261
transform 1 0 44129 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1448
timestamp 1624857261
transform 1 0 44133 0 1 1691
box 0 0 1 1
use contact_19  contact_19_908
timestamp 1624857261
transform 1 0 44130 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1448
timestamp 1624857261
transform 1 0 44137 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4141
timestamp 1624857261
transform 1 0 44064 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1447
timestamp 1624857261
transform 1 0 44469 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1447
timestamp 1624857261
transform 1 0 44473 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1446
timestamp 1624857261
transform 1 0 44805 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1446
timestamp 1624857261
transform 1 0 44809 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1444
timestamp 1624857261
transform 1 0 45477 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1445
timestamp 1624857261
transform 1 0 45141 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1444
timestamp 1624857261
transform 1 0 45481 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1445
timestamp 1624857261
transform 1 0 45145 0 1 1683
box 0 0 1 1
use contact_7  contact_7_291
timestamp 1624857261
transform 1 0 45809 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1443
timestamp 1624857261
transform 1 0 45813 0 1 1691
box 0 0 1 1
use contact_19  contact_19_907
timestamp 1624857261
transform 1 0 45810 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1443
timestamp 1624857261
transform 1 0 45817 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4123
timestamp 1624857261
transform 1 0 45696 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1442
timestamp 1624857261
transform 1 0 46149 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1442
timestamp 1624857261
transform 1 0 46153 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1441
timestamp 1624857261
transform 1 0 46485 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1441
timestamp 1624857261
transform 1 0 46489 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1439
timestamp 1624857261
transform 1 0 47157 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1440
timestamp 1624857261
transform 1 0 46821 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1439
timestamp 1624857261
transform 1 0 47161 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1440
timestamp 1624857261
transform 1 0 46825 0 1 1683
box 0 0 1 1
use contact_7  contact_7_290
timestamp 1624857261
transform 1 0 47489 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1438
timestamp 1624857261
transform 1 0 47493 0 1 1691
box 0 0 1 1
use contact_19  contact_19_906
timestamp 1624857261
transform 1 0 47490 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1438
timestamp 1624857261
transform 1 0 47497 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4103
timestamp 1624857261
transform 1 0 47464 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1437
timestamp 1624857261
transform 1 0 47829 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1437
timestamp 1624857261
transform 1 0 47833 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1436
timestamp 1624857261
transform 1 0 48165 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1436
timestamp 1624857261
transform 1 0 48169 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1434
timestamp 1624857261
transform 1 0 48837 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1435
timestamp 1624857261
transform 1 0 48501 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1434
timestamp 1624857261
transform 1 0 48841 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1435
timestamp 1624857261
transform 1 0 48505 0 1 1683
box 0 0 1 1
use contact_7  contact_7_289
timestamp 1624857261
transform 1 0 49169 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1433
timestamp 1624857261
transform 1 0 49173 0 1 1691
box 0 0 1 1
use contact_19  contact_19_905
timestamp 1624857261
transform 1 0 49170 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1433
timestamp 1624857261
transform 1 0 49177 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4089
timestamp 1624857261
transform 1 0 48960 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1432
timestamp 1624857261
transform 1 0 49509 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1432
timestamp 1624857261
transform 1 0 49513 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1430
timestamp 1624857261
transform 1 0 50181 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1431
timestamp 1624857261
transform 1 0 49845 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1430
timestamp 1624857261
transform 1 0 50185 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1431
timestamp 1624857261
transform 1 0 49849 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1429
timestamp 1624857261
transform 1 0 50517 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1429
timestamp 1624857261
transform 1 0 50521 0 1 1683
box 0 0 1 1
use contact_7  contact_7_288
timestamp 1624857261
transform 1 0 50849 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1428
timestamp 1624857261
transform 1 0 50853 0 1 1691
box 0 0 1 1
use contact_19  contact_19_904
timestamp 1624857261
transform 1 0 50850 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1428
timestamp 1624857261
transform 1 0 50857 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4065
timestamp 1624857261
transform 1 0 50728 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1427
timestamp 1624857261
transform 1 0 51189 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1427
timestamp 1624857261
transform 1 0 51193 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1425
timestamp 1624857261
transform 1 0 51861 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1426
timestamp 1624857261
transform 1 0 51525 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1425
timestamp 1624857261
transform 1 0 51865 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1426
timestamp 1624857261
transform 1 0 51529 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1424
timestamp 1624857261
transform 1 0 52197 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1424
timestamp 1624857261
transform 1 0 52201 0 1 1683
box 0 0 1 1
use contact_7  contact_7_287
timestamp 1624857261
transform 1 0 52529 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1423
timestamp 1624857261
transform 1 0 52533 0 1 1691
box 0 0 1 1
use contact_19  contact_19_903
timestamp 1624857261
transform 1 0 52530 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1423
timestamp 1624857261
transform 1 0 52537 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4049
timestamp 1624857261
transform 1 0 52496 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1422
timestamp 1624857261
transform 1 0 52869 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1422
timestamp 1624857261
transform 1 0 52873 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1420
timestamp 1624857261
transform 1 0 53541 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1421
timestamp 1624857261
transform 1 0 53205 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1420
timestamp 1624857261
transform 1 0 53545 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1421
timestamp 1624857261
transform 1 0 53209 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1419
timestamp 1624857261
transform 1 0 53877 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1419
timestamp 1624857261
transform 1 0 53881 0 1 1683
box 0 0 1 1
use contact_7  contact_7_286
timestamp 1624857261
transform 1 0 54209 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1418
timestamp 1624857261
transform 1 0 54213 0 1 1691
box 0 0 1 1
use contact_19  contact_19_902
timestamp 1624857261
transform 1 0 54210 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1418
timestamp 1624857261
transform 1 0 54217 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4037
timestamp 1624857261
transform 1 0 54128 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1417
timestamp 1624857261
transform 1 0 54549 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1417
timestamp 1624857261
transform 1 0 54553 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1415
timestamp 1624857261
transform 1 0 55221 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1416
timestamp 1624857261
transform 1 0 54885 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1415
timestamp 1624857261
transform 1 0 55225 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1416
timestamp 1624857261
transform 1 0 54889 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1414
timestamp 1624857261
transform 1 0 55557 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1414
timestamp 1624857261
transform 1 0 55561 0 1 1683
box 0 0 1 1
use contact_7  contact_7_285
timestamp 1624857261
transform 1 0 55889 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1413
timestamp 1624857261
transform 1 0 55893 0 1 1691
box 0 0 1 1
use contact_19  contact_19_901
timestamp 1624857261
transform 1 0 55890 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1413
timestamp 1624857261
transform 1 0 55897 0 1 1683
box 0 0 1 1
use contact_33  contact_33_4013
timestamp 1624857261
transform 1 0 55896 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1412
timestamp 1624857261
transform 1 0 56229 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1412
timestamp 1624857261
transform 1 0 56233 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1410
timestamp 1624857261
transform 1 0 56901 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1411
timestamp 1624857261
transform 1 0 56565 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1410
timestamp 1624857261
transform 1 0 56905 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1411
timestamp 1624857261
transform 1 0 56569 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1409
timestamp 1624857261
transform 1 0 57237 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1409
timestamp 1624857261
transform 1 0 57241 0 1 1683
box 0 0 1 1
use contact_7  contact_7_284
timestamp 1624857261
transform 1 0 57569 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1408
timestamp 1624857261
transform 1 0 57573 0 1 1691
box 0 0 1 1
use contact_19  contact_19_900
timestamp 1624857261
transform 1 0 57570 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1408
timestamp 1624857261
transform 1 0 57577 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3987
timestamp 1624857261
transform 1 0 57392 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1407
timestamp 1624857261
transform 1 0 57909 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1407
timestamp 1624857261
transform 1 0 57913 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1405
timestamp 1624857261
transform 1 0 58581 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1406
timestamp 1624857261
transform 1 0 58245 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1405
timestamp 1624857261
transform 1 0 58585 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1406
timestamp 1624857261
transform 1 0 58249 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1404
timestamp 1624857261
transform 1 0 58917 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1404
timestamp 1624857261
transform 1 0 58921 0 1 1683
box 0 0 1 1
use contact_7  contact_7_283
timestamp 1624857261
transform 1 0 59249 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1403
timestamp 1624857261
transform 1 0 59253 0 1 1691
box 0 0 1 1
use contact_19  contact_19_899
timestamp 1624857261
transform 1 0 59250 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1403
timestamp 1624857261
transform 1 0 59257 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3975
timestamp 1624857261
transform 1 0 59160 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1402
timestamp 1624857261
transform 1 0 59589 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1402
timestamp 1624857261
transform 1 0 59593 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1400
timestamp 1624857261
transform 1 0 60261 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1401
timestamp 1624857261
transform 1 0 59925 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1400
timestamp 1624857261
transform 1 0 60265 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1401
timestamp 1624857261
transform 1 0 59929 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1399
timestamp 1624857261
transform 1 0 60597 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1399
timestamp 1624857261
transform 1 0 60601 0 1 1683
box 0 0 1 1
use contact_7  contact_7_282
timestamp 1624857261
transform 1 0 60929 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1398
timestamp 1624857261
transform 1 0 60933 0 1 1691
box 0 0 1 1
use contact_19  contact_19_898
timestamp 1624857261
transform 1 0 60930 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1398
timestamp 1624857261
transform 1 0 60937 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3959
timestamp 1624857261
transform 1 0 60928 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1396
timestamp 1624857261
transform 1 0 61605 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1397
timestamp 1624857261
transform 1 0 61269 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1397
timestamp 1624857261
transform 1 0 61273 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1395
timestamp 1624857261
transform 1 0 61941 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1395
timestamp 1624857261
transform 1 0 61945 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1396
timestamp 1624857261
transform 1 0 61609 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1394
timestamp 1624857261
transform 1 0 62277 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1394
timestamp 1624857261
transform 1 0 62281 0 1 1683
box 0 0 1 1
use contact_7  contact_7_281
timestamp 1624857261
transform 1 0 62609 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1393
timestamp 1624857261
transform 1 0 62613 0 1 1691
box 0 0 1 1
use contact_19  contact_19_897
timestamp 1624857261
transform 1 0 62610 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1393
timestamp 1624857261
transform 1 0 62617 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3937
timestamp 1624857261
transform 1 0 62696 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1391
timestamp 1624857261
transform 1 0 63285 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1392
timestamp 1624857261
transform 1 0 62949 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1391
timestamp 1624857261
transform 1 0 63289 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1392
timestamp 1624857261
transform 1 0 62953 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1390
timestamp 1624857261
transform 1 0 63621 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1390
timestamp 1624857261
transform 1 0 63625 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1389
timestamp 1624857261
transform 1 0 63957 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1389
timestamp 1624857261
transform 1 0 63961 0 1 1683
box 0 0 1 1
use contact_7  contact_7_280
timestamp 1624857261
transform 1 0 64289 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1388
timestamp 1624857261
transform 1 0 64293 0 1 1691
box 0 0 1 1
use contact_19  contact_19_896
timestamp 1624857261
transform 1 0 64290 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1388
timestamp 1624857261
transform 1 0 64297 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3921
timestamp 1624857261
transform 1 0 64192 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1386
timestamp 1624857261
transform 1 0 64965 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1387
timestamp 1624857261
transform 1 0 64629 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1386
timestamp 1624857261
transform 1 0 64969 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1387
timestamp 1624857261
transform 1 0 64633 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1385
timestamp 1624857261
transform 1 0 65301 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1385
timestamp 1624857261
transform 1 0 65305 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1384
timestamp 1624857261
transform 1 0 65637 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1384
timestamp 1624857261
transform 1 0 65641 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3901
timestamp 1624857261
transform 1 0 65824 0 1 1637
box 0 0 1 1
use contact_7  contact_7_279
timestamp 1624857261
transform 1 0 65969 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1383
timestamp 1624857261
transform 1 0 65973 0 1 1691
box 0 0 1 1
use contact_19  contact_19_895
timestamp 1624857261
transform 1 0 65970 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1383
timestamp 1624857261
transform 1 0 65977 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1381
timestamp 1624857261
transform 1 0 66645 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1382
timestamp 1624857261
transform 1 0 66309 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1381
timestamp 1624857261
transform 1 0 66649 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1382
timestamp 1624857261
transform 1 0 66313 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1380
timestamp 1624857261
transform 1 0 66981 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1380
timestamp 1624857261
transform 1 0 66985 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1379
timestamp 1624857261
transform 1 0 67317 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1379
timestamp 1624857261
transform 1 0 67321 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3883
timestamp 1624857261
transform 1 0 67592 0 1 1637
box 0 0 1 1
use contact_7  contact_7_155
timestamp 1624857261
transform 1 0 1793 0 1 2023
box 0 0 1 1
use contact_14  contact_14_770
timestamp 1624857261
transform 1 0 1797 0 1 2363
box 0 0 1 1
use contact_14  contact_14_771
timestamp 1624857261
transform 1 0 1797 0 1 2027
box 0 0 1 1
use contact_19  contact_19_770
timestamp 1624857261
transform 1 0 1794 0 1 2364
box 0 0 1 1
use contact_19  contact_19_771
timestamp 1624857261
transform 1 0 1794 0 1 2028
box 0 0 1 1
use contact_13  contact_13_770
timestamp 1624857261
transform 1 0 1801 0 1 2355
box 0 0 1 1
use contact_13  contact_13_771
timestamp 1624857261
transform 1 0 1801 0 1 2019
box 0 0 1 1
use contact_14  contact_14_768
timestamp 1624857261
transform 1 0 1797 0 1 3035
box 0 0 1 1
use contact_14  contact_14_769
timestamp 1624857261
transform 1 0 1797 0 1 2699
box 0 0 1 1
use contact_19  contact_19_768
timestamp 1624857261
transform 1 0 1794 0 1 3036
box 0 0 1 1
use contact_19  contact_19_769
timestamp 1624857261
transform 1 0 1794 0 1 2700
box 0 0 1 1
use contact_13  contact_13_768
timestamp 1624857261
transform 1 0 1801 0 1 3027
box 0 0 1 1
use contact_13  contact_13_769
timestamp 1624857261
transform 1 0 1801 0 1 2691
box 0 0 1 1
use wmask_dff  wmask_dff_0
timestamp 1624857261
transform 1 0 18742 0 1 2396
box -36 -49 4708 1467
use col_addr_dff  col_addr_dff_1
timestamp 1624857261
transform 1 0 16406 0 1 2396
box -36 -49 1204 1467
use contact_33  contact_33_5456
timestamp 1624857261
transform 1 0 16592 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5455
timestamp 1624857261
transform 1 0 17680 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5454
timestamp 1624857261
transform 1 0 18768 0 1 2861
box 0 0 1 1
use contact_7  contact_7_375
timestamp 1624857261
transform 1 0 16543 0 1 2923
box 0 0 1 1
use contact_7  contact_7_374
timestamp 1624857261
transform 1 0 17711 0 1 2923
box 0 0 1 1
use contact_7  contact_7_365
timestamp 1624857261
transform 1 0 18879 0 1 2923
box 0 0 1 1
use contact_32  contact_32_2
timestamp 1624857261
transform 1 0 15289 0 1 2667
box 0 0 1 1
use contact_33  contact_33_5488
timestamp 1624857261
transform 1 0 23664 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5453
timestamp 1624857261
transform 1 0 20128 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5452
timestamp 1624857261
transform 1 0 21080 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5451
timestamp 1624857261
transform 1 0 22304 0 1 2861
box 0 0 1 1
use contact_33  contact_33_2304
timestamp 1624857261
transform 1 0 19312 0 1 2317
box 0 0 1 1
use contact_7  contact_7_439
timestamp 1624857261
transform 1 0 23551 0 1 2923
box 0 0 1 1
use contact_7  contact_7_364
timestamp 1624857261
transform 1 0 20047 0 1 2923
box 0 0 1 1
use contact_7  contact_7_363
timestamp 1624857261
transform 1 0 21215 0 1 2923
box 0 0 1 1
use contact_7  contact_7_362
timestamp 1624857261
transform 1 0 22383 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5487
timestamp 1624857261
transform 1 0 24752 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5486
timestamp 1624857261
transform 1 0 25976 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5485
timestamp 1624857261
transform 1 0 27064 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5484
timestamp 1624857261
transform 1 0 28152 0 1 2861
box 0 0 1 1
use contact_7  contact_7_438
timestamp 1624857261
transform 1 0 24719 0 1 2923
box 0 0 1 1
use contact_7  contact_7_437
timestamp 1624857261
transform 1 0 25887 0 1 2923
box 0 0 1 1
use contact_7  contact_7_436
timestamp 1624857261
transform 1 0 27055 0 1 2923
box 0 0 1 1
use contact_7  contact_7_435
timestamp 1624857261
transform 1 0 28223 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5483
timestamp 1624857261
transform 1 0 29240 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5482
timestamp 1624857261
transform 1 0 30600 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5481
timestamp 1624857261
transform 1 0 31824 0 1 2861
box 0 0 1 1
use contact_33  contact_33_5480
timestamp 1624857261
transform 1 0 32912 0 1 2861
box 0 0 1 1
use contact_7  contact_7_434
timestamp 1624857261
transform 1 0 29391 0 1 2923
box 0 0 1 1
use contact_7  contact_7_433
timestamp 1624857261
transform 1 0 30559 0 1 2923
box 0 0 1 1
use contact_7  contact_7_432
timestamp 1624857261
transform 1 0 31727 0 1 2923
box 0 0 1 1
use contact_7  contact_7_431
timestamp 1624857261
transform 1 0 32895 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5479
timestamp 1624857261
transform 1 0 34000 0 1 2861
box 0 0 1 1
use contact_7  contact_7_430
timestamp 1624857261
transform 1 0 34063 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5478
timestamp 1624857261
transform 1 0 35088 0 1 2861
box 0 0 1 1
use contact_7  contact_7_429
timestamp 1624857261
transform 1 0 35231 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5477
timestamp 1624857261
transform 1 0 36448 0 1 2861
box 0 0 1 1
use contact_7  contact_7_428
timestamp 1624857261
transform 1 0 36399 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5476
timestamp 1624857261
transform 1 0 37536 0 1 2861
box 0 0 1 1
use contact_7  contact_7_427
timestamp 1624857261
transform 1 0 37567 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5475
timestamp 1624857261
transform 1 0 38624 0 1 2861
box 0 0 1 1
use contact_7  contact_7_426
timestamp 1624857261
transform 1 0 38735 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5474
timestamp 1624857261
transform 1 0 39984 0 1 2861
box 0 0 1 1
use contact_7  contact_7_425
timestamp 1624857261
transform 1 0 39903 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5473
timestamp 1624857261
transform 1 0 41208 0 1 2861
box 0 0 1 1
use contact_7  contact_7_424
timestamp 1624857261
transform 1 0 41071 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5472
timestamp 1624857261
transform 1 0 42296 0 1 2861
box 0 0 1 1
use contact_7  contact_7_423
timestamp 1624857261
transform 1 0 42239 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5471
timestamp 1624857261
transform 1 0 43384 0 1 2861
box 0 0 1 1
use contact_7  contact_7_422
timestamp 1624857261
transform 1 0 43407 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5470
timestamp 1624857261
transform 1 0 44472 0 1 2861
box 0 0 1 1
use contact_7  contact_7_421
timestamp 1624857261
transform 1 0 44575 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5469
timestamp 1624857261
transform 1 0 45832 0 1 2861
box 0 0 1 1
use contact_7  contact_7_420
timestamp 1624857261
transform 1 0 45743 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5468
timestamp 1624857261
transform 1 0 46920 0 1 2861
box 0 0 1 1
use contact_7  contact_7_419
timestamp 1624857261
transform 1 0 46911 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5467
timestamp 1624857261
transform 1 0 48144 0 1 2861
box 0 0 1 1
use contact_7  contact_7_418
timestamp 1624857261
transform 1 0 48079 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5466
timestamp 1624857261
transform 1 0 49232 0 1 2861
box 0 0 1 1
use contact_7  contact_7_417
timestamp 1624857261
transform 1 0 49247 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5465
timestamp 1624857261
transform 1 0 50320 0 1 2861
box 0 0 1 1
use contact_7  contact_7_416
timestamp 1624857261
transform 1 0 50415 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5464
timestamp 1624857261
transform 1 0 51680 0 1 2861
box 0 0 1 1
use contact_7  contact_7_415
timestamp 1624857261
transform 1 0 51583 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5463
timestamp 1624857261
transform 1 0 52768 0 1 2861
box 0 0 1 1
use contact_7  contact_7_414
timestamp 1624857261
transform 1 0 52751 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5462
timestamp 1624857261
transform 1 0 53856 0 1 2861
box 0 0 1 1
use contact_7  contact_7_413
timestamp 1624857261
transform 1 0 53919 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5461
timestamp 1624857261
transform 1 0 54944 0 1 2861
box 0 0 1 1
use contact_7  contact_7_412
timestamp 1624857261
transform 1 0 55087 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5460
timestamp 1624857261
transform 1 0 56304 0 1 2861
box 0 0 1 1
use contact_7  contact_7_411
timestamp 1624857261
transform 1 0 56255 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5459
timestamp 1624857261
transform 1 0 57528 0 1 2861
box 0 0 1 1
use contact_7  contact_7_410
timestamp 1624857261
transform 1 0 57423 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5458
timestamp 1624857261
transform 1 0 58616 0 1 2861
box 0 0 1 1
use contact_7  contact_7_409
timestamp 1624857261
transform 1 0 58591 0 1 2923
box 0 0 1 1
use contact_33  contact_33_5457
timestamp 1624857261
transform 1 0 59704 0 1 2861
box 0 0 1 1
use contact_7  contact_7_408
timestamp 1624857261
transform 1 0 59759 0 1 2923
box 0 0 1 1
use data_dff  data_dff_0
timestamp 1624857261
transform 1 0 23414 0 1 2396
box -36 -49 37412 1467
use contact_33  contact_33_5345
timestamp 1624857261
transform 1 0 1224 0 1 3813
box 0 0 1 1
use contact_13  contact_13_767
timestamp 1624857261
transform 1 0 1801 0 1 3363
box 0 0 1 1
use contact_13  contact_13_766
timestamp 1624857261
transform 1 0 1801 0 1 3699
box 0 0 1 1
use contact_19  contact_19_767
timestamp 1624857261
transform 1 0 1794 0 1 3372
box 0 0 1 1
use contact_19  contact_19_766
timestamp 1624857261
transform 1 0 1794 0 1 3708
box 0 0 1 1
use contact_14  contact_14_767
timestamp 1624857261
transform 1 0 1797 0 1 3371
box 0 0 1 1
use contact_14  contact_14_766
timestamp 1624857261
transform 1 0 1797 0 1 3707
box 0 0 1 1
use contact_7  contact_7_154
timestamp 1624857261
transform 1 0 1793 0 1 3703
box 0 0 1 1
use contact_13  contact_13_765
timestamp 1624857261
transform 1 0 1801 0 1 4035
box 0 0 1 1
use contact_13  contact_13_764
timestamp 1624857261
transform 1 0 1801 0 1 4371
box 0 0 1 1
use contact_19  contact_19_765
timestamp 1624857261
transform 1 0 1794 0 1 4044
box 0 0 1 1
use contact_19  contact_19_764
timestamp 1624857261
transform 1 0 1794 0 1 4380
box 0 0 1 1
use contact_14  contact_14_765
timestamp 1624857261
transform 1 0 1797 0 1 4043
box 0 0 1 1
use contact_14  contact_14_764
timestamp 1624857261
transform 1 0 1797 0 1 4379
box 0 0 1 1
use contact_13  contact_13_763
timestamp 1624857261
transform 1 0 1801 0 1 4707
box 0 0 1 1
use contact_19  contact_19_763
timestamp 1624857261
transform 1 0 1794 0 1 4716
box 0 0 1 1
use contact_14  contact_14_763
timestamp 1624857261
transform 1 0 1797 0 1 4715
box 0 0 1 1
use contact_33  contact_33_5252
timestamp 1624857261
transform 1 0 16864 0 1 3813
box 0 0 1 1
use contact_33  contact_33_4223
timestamp 1624857261
transform 1 0 36720 0 1 3677
box 0 0 1 1
use contact_33  contact_33_5333
timestamp 1624857261
transform 1 0 1224 0 1 6941
box 0 0 1 1
use contact_33  contact_33_5332
timestamp 1624857261
transform 1 0 1224 0 1 5445
box 0 0 1 1
use contact_33  contact_33_5323
timestamp 1624857261
transform 1 0 1224 0 1 8845
box 0 0 1 1
use contact_33  contact_33_2350
timestamp 1624857261
transform 1 0 544 0 1 7621
box 0 0 1 1
use contact_14  contact_14_762
timestamp 1624857261
transform 1 0 1797 0 1 5051
box 0 0 1 1
use contact_19  contact_19_762
timestamp 1624857261
transform 1 0 1794 0 1 5052
box 0 0 1 1
use contact_13  contact_13_762
timestamp 1624857261
transform 1 0 1801 0 1 5043
box 0 0 1 1
use contact_7  contact_7_153
timestamp 1624857261
transform 1 0 1793 0 1 5383
box 0 0 1 1
use contact_14  contact_14_761
timestamp 1624857261
transform 1 0 1797 0 1 5387
box 0 0 1 1
use contact_19  contact_19_761
timestamp 1624857261
transform 1 0 1794 0 1 5388
box 0 0 1 1
use contact_13  contact_13_761
timestamp 1624857261
transform 1 0 1801 0 1 5379
box 0 0 1 1
use contact_14  contact_14_760
timestamp 1624857261
transform 1 0 1797 0 1 5723
box 0 0 1 1
use contact_19  contact_19_760
timestamp 1624857261
transform 1 0 1794 0 1 5724
box 0 0 1 1
use contact_13  contact_13_760
timestamp 1624857261
transform 1 0 1801 0 1 5715
box 0 0 1 1
use contact_14  contact_14_759
timestamp 1624857261
transform 1 0 1797 0 1 6059
box 0 0 1 1
use contact_19  contact_19_759
timestamp 1624857261
transform 1 0 1794 0 1 6060
box 0 0 1 1
use contact_13  contact_13_759
timestamp 1624857261
transform 1 0 1801 0 1 6051
box 0 0 1 1
use contact_14  contact_14_758
timestamp 1624857261
transform 1 0 1797 0 1 6395
box 0 0 1 1
use contact_19  contact_19_758
timestamp 1624857261
transform 1 0 1794 0 1 6396
box 0 0 1 1
use contact_13  contact_13_758
timestamp 1624857261
transform 1 0 1801 0 1 6387
box 0 0 1 1
use contact_14  contact_14_757
timestamp 1624857261
transform 1 0 1797 0 1 6731
box 0 0 1 1
use contact_19  contact_19_757
timestamp 1624857261
transform 1 0 1794 0 1 6732
box 0 0 1 1
use contact_13  contact_13_757
timestamp 1624857261
transform 1 0 1801 0 1 6723
box 0 0 1 1
use contact_7  contact_7_152
timestamp 1624857261
transform 1 0 1793 0 1 7063
box 0 0 1 1
use contact_14  contact_14_756
timestamp 1624857261
transform 1 0 1797 0 1 7067
box 0 0 1 1
use contact_19  contact_19_756
timestamp 1624857261
transform 1 0 1794 0 1 7068
box 0 0 1 1
use contact_13  contact_13_756
timestamp 1624857261
transform 1 0 1801 0 1 7059
box 0 0 1 1
use contact_14  contact_14_755
timestamp 1624857261
transform 1 0 1797 0 1 7403
box 0 0 1 1
use contact_19  contact_19_755
timestamp 1624857261
transform 1 0 1794 0 1 7404
box 0 0 1 1
use contact_13  contact_13_755
timestamp 1624857261
transform 1 0 1801 0 1 7395
box 0 0 1 1
use contact_14  contact_14_754
timestamp 1624857261
transform 1 0 1797 0 1 7739
box 0 0 1 1
use contact_19  contact_19_754
timestamp 1624857261
transform 1 0 1794 0 1 7740
box 0 0 1 1
use contact_13  contact_13_753
timestamp 1624857261
transform 1 0 1801 0 1 8067
box 0 0 1 1
use contact_13  contact_13_754
timestamp 1624857261
transform 1 0 1801 0 1 7731
box 0 0 1 1
use contact_14  contact_14_752
timestamp 1624857261
transform 1 0 1797 0 1 8411
box 0 0 1 1
use contact_14  contact_14_753
timestamp 1624857261
transform 1 0 1797 0 1 8075
box 0 0 1 1
use contact_19  contact_19_752
timestamp 1624857261
transform 1 0 1794 0 1 8412
box 0 0 1 1
use contact_19  contact_19_753
timestamp 1624857261
transform 1 0 1794 0 1 8076
box 0 0 1 1
use contact_13  contact_13_752
timestamp 1624857261
transform 1 0 1801 0 1 8403
box 0 0 1 1
use contact_7  contact_7_442
timestamp 1624857261
transform 1 0 2753 0 1 8147
box 0 0 1 1
use contact_7  contact_7_151
timestamp 1624857261
transform 1 0 1793 0 1 8743
box 0 0 1 1
use contact_14  contact_14_751
timestamp 1624857261
transform 1 0 1797 0 1 8747
box 0 0 1 1
use contact_19  contact_19_751
timestamp 1624857261
transform 1 0 1794 0 1 8748
box 0 0 1 1
use contact_13  contact_13_751
timestamp 1624857261
transform 1 0 1801 0 1 8739
box 0 0 1 1
use contact_14  contact_14_750
timestamp 1624857261
transform 1 0 1797 0 1 9083
box 0 0 1 1
use contact_19  contact_19_750
timestamp 1624857261
transform 1 0 1794 0 1 9084
box 0 0 1 1
use contact_13  contact_13_750
timestamp 1624857261
transform 1 0 1801 0 1 9075
box 0 0 1 1
use contact_14  contact_14_749
timestamp 1624857261
transform 1 0 1797 0 1 9419
box 0 0 1 1
use contact_19  contact_19_749
timestamp 1624857261
transform 1 0 1794 0 1 9420
box 0 0 1 1
use contact_13  contact_13_749
timestamp 1624857261
transform 1 0 1801 0 1 9411
box 0 0 1 1
use contact_7  contact_7_440
timestamp 1624857261
transform 1 0 5974 0 1 8252
box 0 0 1 1
use contact_33  contact_33_5255
timestamp 1624857261
transform 1 0 15096 0 1 9117
box 0 0 1 1
use contact_33  contact_33_2329
timestamp 1624857261
transform 1 0 15232 0 1 7621
box 0 0 1 1
use contact_33  contact_33_5253
timestamp 1624857261
transform 1 0 16864 0 1 8981
box 0 0 1 1
use cr_4  cr_4_0
timestamp 1624857261
transform 1 0 15406 0 1 9422
box 3208 -3962 52705 1462
use contact_33  contact_33_2351
timestamp 1624857261
transform 1 0 544 0 1 10205
box 0 0 1 1
use contact_33  contact_33_5371
timestamp 1624857261
transform 1 0 1224 0 1 10341
box 0 0 1 1
use contact_13  contact_13_748
timestamp 1624857261
transform 1 0 1801 0 1 9747
box 0 0 1 1
use contact_19  contact_19_748
timestamp 1624857261
transform 1 0 1794 0 1 9756
box 0 0 1 1
use contact_14  contact_14_748
timestamp 1624857261
transform 1 0 1797 0 1 9755
box 0 0 1 1
use contact_7  contact_7_441
timestamp 1624857261
transform 1 0 2753 0 1 9847
box 0 0 1 1
use contact_13  contact_13_747
timestamp 1624857261
transform 1 0 1801 0 1 10083
box 0 0 1 1
use contact_19  contact_19_747
timestamp 1624857261
transform 1 0 1794 0 1 10092
box 0 0 1 1
use contact_14  contact_14_747
timestamp 1624857261
transform 1 0 1797 0 1 10091
box 0 0 1 1
use contact_13  contact_13_746
timestamp 1624857261
transform 1 0 1801 0 1 10419
box 0 0 1 1
use contact_19  contact_19_746
timestamp 1624857261
transform 1 0 1794 0 1 10428
box 0 0 1 1
use contact_14  contact_14_746
timestamp 1624857261
transform 1 0 1797 0 1 10427
box 0 0 1 1
use contact_7  contact_7_150
timestamp 1624857261
transform 1 0 1793 0 1 10423
box 0 0 1 1
use contact_13  contact_13_745
timestamp 1624857261
transform 1 0 1801 0 1 10755
box 0 0 1 1
use contact_33  contact_33_2330
timestamp 1624857261
transform 1 0 15232 0 1 10341
box 0 0 1 1
use contact_33  contact_33_2332
timestamp 1624857261
transform 1 0 15232 0 1 10477
box 0 0 1 1
use contact_33  contact_33_1524
timestamp 1624857261
transform 1 0 29240 0 1 9525
box 0 0 1 1
use contact_33  contact_33_4313
timestamp 1624857261
transform 1 0 29512 0 1 10613
box 0 0 1 1
use contact_13  contact_13_744
timestamp 1624857261
transform 1 0 1801 0 1 11091
box 0 0 1 1
use contact_19  contact_19_745
timestamp 1624857261
transform 1 0 1794 0 1 10764
box 0 0 1 1
use contact_19  contact_19_744
timestamp 1624857261
transform 1 0 1794 0 1 11100
box 0 0 1 1
use contact_14  contact_14_745
timestamp 1624857261
transform 1 0 1797 0 1 10763
box 0 0 1 1
use contact_14  contact_14_744
timestamp 1624857261
transform 1 0 1797 0 1 11099
box 0 0 1 1
use contact_13  contact_13_743
timestamp 1624857261
transform 1 0 1801 0 1 11427
box 0 0 1 1
use contact_19  contact_19_743
timestamp 1624857261
transform 1 0 1794 0 1 11436
box 0 0 1 1
use contact_14  contact_14_743
timestamp 1624857261
transform 1 0 1797 0 1 11435
box 0 0 1 1
use contact_13  contact_13_742
timestamp 1624857261
transform 1 0 1801 0 1 11763
box 0 0 1 1
use contact_19  contact_19_742
timestamp 1624857261
transform 1 0 1794 0 1 11772
box 0 0 1 1
use contact_14  contact_14_742
timestamp 1624857261
transform 1 0 1797 0 1 11771
box 0 0 1 1
use contact_33  contact_33_5251
timestamp 1624857261
transform 1 0 15096 0 1 11973
box 0 0 1 1
use contact_33  contact_33_5254
timestamp 1624857261
transform 1 0 15096 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1901
timestamp 1624857261
transform 1 0 22168 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1357
timestamp 1624857261
transform 1 0 29784 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1523
timestamp 1624857261
transform 1 0 29240 0 1 11293
box 0 0 1 1
use contact_33  contact_33_4299
timestamp 1624857261
transform 1 0 29920 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4300
timestamp 1624857261
transform 1 0 29648 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4301
timestamp 1624857261
transform 1 0 29648 0 1 11837
box 0 0 1 1
use contact_33  contact_33_4312
timestamp 1624857261
transform 1 0 29512 0 1 11021
box 0 0 1 1
use contact_33  contact_33_1345
timestamp 1624857261
transform 1 0 32232 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4273
timestamp 1624857261
transform 1 0 32368 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4274
timestamp 1624857261
transform 1 0 32096 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4275
timestamp 1624857261
transform 1 0 32096 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1333
timestamp 1624857261
transform 1 0 34816 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4245
timestamp 1624857261
transform 1 0 34680 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4246
timestamp 1624857261
transform 1 0 34680 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4247
timestamp 1624857261
transform 1 0 34680 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1321
timestamp 1624857261
transform 1 0 37400 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4217
timestamp 1624857261
transform 1 0 37264 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4218
timestamp 1624857261
transform 1 0 37264 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4219
timestamp 1624857261
transform 1 0 37264 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1309
timestamp 1624857261
transform 1 0 39848 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4189
timestamp 1624857261
transform 1 0 39712 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4190
timestamp 1624857261
transform 1 0 39712 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4191
timestamp 1624857261
transform 1 0 39712 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1297
timestamp 1624857261
transform 1 0 42160 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4167
timestamp 1624857261
transform 1 0 42432 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4168
timestamp 1624857261
transform 1 0 42296 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4169
timestamp 1624857261
transform 1 0 42296 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1285
timestamp 1624857261
transform 1 0 44608 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4135
timestamp 1624857261
transform 1 0 44880 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4136
timestamp 1624857261
transform 1 0 44744 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4137
timestamp 1624857261
transform 1 0 44744 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1273
timestamp 1624857261
transform 1 0 47192 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4113
timestamp 1624857261
transform 1 0 47328 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4114
timestamp 1624857261
transform 1 0 47056 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4115
timestamp 1624857261
transform 1 0 47056 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1261
timestamp 1624857261
transform 1 0 49504 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4079
timestamp 1624857261
transform 1 0 49640 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4080
timestamp 1624857261
transform 1 0 49776 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4081
timestamp 1624857261
transform 1 0 49776 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1249
timestamp 1624857261
transform 1 0 52360 0 1 11701
box 0 0 1 1
use contact_33  contact_33_4057
timestamp 1624857261
transform 1 0 52224 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4058
timestamp 1624857261
transform 1 0 52224 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4059
timestamp 1624857261
transform 1 0 52224 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1238
timestamp 1624857261
transform 1 0 54400 0 1 11429
box 0 0 1 1
use contact_33  contact_33_4027
timestamp 1624857261
transform 1 0 54808 0 1 11973
box 0 0 1 1
use contact_33  contact_33_4028
timestamp 1624857261
transform 1 0 54808 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4029
timestamp 1624857261
transform 1 0 54808 0 1 11837
box 0 0 1 1
use contact_33  contact_33_4000
timestamp 1624857261
transform 1 0 57256 0 1 11021
box 0 0 1 1
use contact_33  contact_33_4001
timestamp 1624857261
transform 1 0 57256 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1225
timestamp 1624857261
transform 1 0 57528 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3999
timestamp 1624857261
transform 1 0 57392 0 1 11973
box 0 0 1 1
use contact_33  contact_33_1213
timestamp 1624857261
transform 1 0 59568 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3970
timestamp 1624857261
transform 1 0 59704 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3971
timestamp 1624857261
transform 1 0 59704 0 1 11837
box 0 0 1 1
use contact_33  contact_33_3969
timestamp 1624857261
transform 1 0 59840 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3945
timestamp 1624857261
transform 1 0 62288 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3946
timestamp 1624857261
transform 1 0 62152 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3947
timestamp 1624857261
transform 1 0 62152 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1201
timestamp 1624857261
transform 1 0 62424 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3913
timestamp 1624857261
transform 1 0 64736 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3914
timestamp 1624857261
transform 1 0 64736 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3915
timestamp 1624857261
transform 1 0 64736 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1189
timestamp 1624857261
transform 1 0 64872 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3892
timestamp 1624857261
transform 1 0 67184 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3893
timestamp 1624857261
transform 1 0 67184 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1177
timestamp 1624857261
transform 1 0 67456 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3891
timestamp 1624857261
transform 1 0 67320 0 1 11973
box 0 0 1 1
use contact_33  contact_33_5334
timestamp 1624857261
transform 1 0 1224 0 1 12109
box 0 0 1 1
use contact_13  contact_13_741
timestamp 1624857261
transform 1 0 1801 0 1 12099
box 0 0 1 1
use contact_19  contact_19_741
timestamp 1624857261
transform 1 0 1794 0 1 12108
box 0 0 1 1
use contact_14  contact_14_741
timestamp 1624857261
transform 1 0 1797 0 1 12107
box 0 0 1 1
use contact_7  contact_7_149
timestamp 1624857261
transform 1 0 1793 0 1 12103
box 0 0 1 1
use contact_13  contact_13_740
timestamp 1624857261
transform 1 0 1801 0 1 12435
box 0 0 1 1
use contact_19  contact_19_740
timestamp 1624857261
transform 1 0 1794 0 1 12444
box 0 0 1 1
use contact_14  contact_14_740
timestamp 1624857261
transform 1 0 1797 0 1 12443
box 0 0 1 1
use contact_13  contact_13_739
timestamp 1624857261
transform 1 0 1801 0 1 12771
box 0 0 1 1
use contact_19  contact_19_739
timestamp 1624857261
transform 1 0 1794 0 1 12780
box 0 0 1 1
use contact_14  contact_14_739
timestamp 1624857261
transform 1 0 1797 0 1 12779
box 0 0 1 1
use contact_13  contact_13_738
timestamp 1624857261
transform 1 0 1801 0 1 13107
box 0 0 1 1
use contact_19  contact_19_738
timestamp 1624857261
transform 1 0 1794 0 1 13116
box 0 0 1 1
use contact_14  contact_14_738
timestamp 1624857261
transform 1 0 1797 0 1 13115
box 0 0 1 1
use contact_7  contact_7_490
timestamp 1624857261
transform 1 0 15205 0 1 12532
box 0 0 1 1
use contact_33  contact_33_2331
timestamp 1624857261
transform 1 0 15232 0 1 13197
box 0 0 1 1
use contact_33  contact_33_4901
timestamp 1624857261
transform 1 0 22304 0 1 13061
box 0 0 1 1
use contact_7  contact_7_489
timestamp 1624857261
transform 1 0 27574 0 1 12532
box 0 0 1 1
use contact_7  contact_7_407
timestamp 1624857261
transform 1 0 29557 0 1 13196
box 0 0 1 1
use contact_19  contact_19_997
timestamp 1624857261
transform 1 0 29558 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1358
timestamp 1624857261
transform 1 0 29784 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5414
timestamp 1624857261
transform 1 0 28968 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1352
timestamp 1624857261
transform 1 0 30056 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1355
timestamp 1624857261
transform 1 0 30056 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1356
timestamp 1624857261
transform 1 0 30056 0 1 12517
box 0 0 1 1
use contact_7  contact_7_406
timestamp 1624857261
transform 1 0 32053 0 1 13196
box 0 0 1 1
use contact_19  contact_19_996
timestamp 1624857261
transform 1 0 32054 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1340
timestamp 1624857261
transform 1 0 32504 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1343
timestamp 1624857261
transform 1 0 32504 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1344
timestamp 1624857261
transform 1 0 32504 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1346
timestamp 1624857261
transform 1 0 32232 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5413
timestamp 1624857261
transform 1 0 31960 0 1 13061
box 0 0 1 1
use contact_7  contact_7_405
timestamp 1624857261
transform 1 0 34549 0 1 13196
box 0 0 1 1
use contact_19  contact_19_995
timestamp 1624857261
transform 1 0 34550 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1328
timestamp 1624857261
transform 1 0 34952 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1331
timestamp 1624857261
transform 1 0 34816 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1332
timestamp 1624857261
transform 1 0 34816 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1334
timestamp 1624857261
transform 1 0 34816 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5412
timestamp 1624857261
transform 1 0 34408 0 1 13061
box 0 0 1 1
use contact_7  contact_7_404
timestamp 1624857261
transform 1 0 37045 0 1 13196
box 0 0 1 1
use contact_19  contact_19_994
timestamp 1624857261
transform 1 0 37046 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1319
timestamp 1624857261
transform 1 0 37400 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1320
timestamp 1624857261
transform 1 0 37400 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1322
timestamp 1624857261
transform 1 0 37400 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5411
timestamp 1624857261
transform 1 0 36992 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1316
timestamp 1624857261
transform 1 0 37536 0 1 13197
box 0 0 1 1
use contact_7  contact_7_403
timestamp 1624857261
transform 1 0 39541 0 1 13196
box 0 0 1 1
use contact_19  contact_19_993
timestamp 1624857261
transform 1 0 39542 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1307
timestamp 1624857261
transform 1 0 39848 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1308
timestamp 1624857261
transform 1 0 39848 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1310
timestamp 1624857261
transform 1 0 39848 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5410
timestamp 1624857261
transform 1 0 39440 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1306
timestamp 1624857261
transform 1 0 39984 0 1 13197
box 0 0 1 1
use contact_7  contact_7_402
timestamp 1624857261
transform 1 0 42037 0 1 13196
box 0 0 1 1
use contact_19  contact_19_992
timestamp 1624857261
transform 1 0 42038 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1295
timestamp 1624857261
transform 1 0 42296 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1296
timestamp 1624857261
transform 1 0 42296 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1298
timestamp 1624857261
transform 1 0 42160 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5409
timestamp 1624857261
transform 1 0 41752 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1292
timestamp 1624857261
transform 1 0 42568 0 1 13197
box 0 0 1 1
use contact_7  contact_7_401
timestamp 1624857261
transform 1 0 44533 0 1 13196
box 0 0 1 1
use contact_19  contact_19_991
timestamp 1624857261
transform 1 0 44534 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1286
timestamp 1624857261
transform 1 0 44608 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5408
timestamp 1624857261
transform 1 0 44200 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1282
timestamp 1624857261
transform 1 0 45016 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1283
timestamp 1624857261
transform 1 0 45016 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1284
timestamp 1624857261
transform 1 0 45016 0 1 12517
box 0 0 1 1
use contact_7  contact_7_400
timestamp 1624857261
transform 1 0 47029 0 1 13196
box 0 0 1 1
use contact_19  contact_19_990
timestamp 1624857261
transform 1 0 47030 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1274
timestamp 1624857261
transform 1 0 47192 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5407
timestamp 1624857261
transform 1 0 46512 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1270
timestamp 1624857261
transform 1 0 47464 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1271
timestamp 1624857261
transform 1 0 47464 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1272
timestamp 1624857261
transform 1 0 47464 0 1 12517
box 0 0 1 1
use contact_7  contact_7_399
timestamp 1624857261
transform 1 0 49525 0 1 13196
box 0 0 1 1
use contact_19  contact_19_989
timestamp 1624857261
transform 1 0 49526 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1259
timestamp 1624857261
transform 1 0 49776 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1260
timestamp 1624857261
transform 1 0 49776 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1262
timestamp 1624857261
transform 1 0 49504 0 1 12245
box 0 0 1 1
use contact_33  contact_33_1258
timestamp 1624857261
transform 1 0 50184 0 1 13061
box 0 0 1 1
use contact_7  contact_7_398
timestamp 1624857261
transform 1 0 52021 0 1 13196
box 0 0 1 1
use contact_19  contact_19_988
timestamp 1624857261
transform 1 0 52022 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1246
timestamp 1624857261
transform 1 0 52360 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1247
timestamp 1624857261
transform 1 0 52360 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1248
timestamp 1624857261
transform 1 0 52360 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1250
timestamp 1624857261
transform 1 0 52360 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5405
timestamp 1624857261
transform 1 0 51952 0 1 13061
box 0 0 1 1
use contact_7  contact_7_397
timestamp 1624857261
transform 1 0 54517 0 1 13196
box 0 0 1 1
use contact_19  contact_19_987
timestamp 1624857261
transform 1 0 54518 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1237
timestamp 1624857261
transform 1 0 54400 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5404
timestamp 1624857261
transform 1 0 54536 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1234
timestamp 1624857261
transform 1 0 54944 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1235
timestamp 1624857261
transform 1 0 54944 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1236
timestamp 1624857261
transform 1 0 54944 0 1 12517
box 0 0 1 1
use contact_7  contact_7_396
timestamp 1624857261
transform 1 0 57013 0 1 13196
box 0 0 1 1
use contact_19  contact_19_986
timestamp 1624857261
transform 1 0 57014 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1223
timestamp 1624857261
transform 1 0 57256 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1224
timestamp 1624857261
transform 1 0 57256 0 1 12517
box 0 0 1 1
use contact_33  contact_33_5403
timestamp 1624857261
transform 1 0 56984 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1222
timestamp 1624857261
transform 1 0 57528 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1226
timestamp 1624857261
transform 1 0 57528 0 1 12245
box 0 0 1 1
use contact_7  contact_7_395
timestamp 1624857261
transform 1 0 59509 0 1 13196
box 0 0 1 1
use contact_19  contact_19_985
timestamp 1624857261
transform 1 0 59510 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1214
timestamp 1624857261
transform 1 0 59568 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5402
timestamp 1624857261
transform 1 0 59296 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1210
timestamp 1624857261
transform 1 0 59976 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1211
timestamp 1624857261
transform 1 0 59976 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1212
timestamp 1624857261
transform 1 0 59976 0 1 12517
box 0 0 1 1
use contact_7  contact_7_394
timestamp 1624857261
transform 1 0 62005 0 1 13196
box 0 0 1 1
use contact_19  contact_19_984
timestamp 1624857261
transform 1 0 62006 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5401
timestamp 1624857261
transform 1 0 61880 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1198
timestamp 1624857261
transform 1 0 62424 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1199
timestamp 1624857261
transform 1 0 62424 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1200
timestamp 1624857261
transform 1 0 62424 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1202
timestamp 1624857261
transform 1 0 62424 0 1 12245
box 0 0 1 1
use contact_7  contact_7_393
timestamp 1624857261
transform 1 0 64501 0 1 13196
box 0 0 1 1
use contact_19  contact_19_983
timestamp 1624857261
transform 1 0 64502 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5400
timestamp 1624857261
transform 1 0 64464 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1186
timestamp 1624857261
transform 1 0 65008 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1187
timestamp 1624857261
transform 1 0 64872 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1188
timestamp 1624857261
transform 1 0 64872 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1190
timestamp 1624857261
transform 1 0 64872 0 1 12245
box 0 0 1 1
use contact_7  contact_7_392
timestamp 1624857261
transform 1 0 66997 0 1 13196
box 0 0 1 1
use contact_19  contact_19_982
timestamp 1624857261
transform 1 0 66998 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5399
timestamp 1624857261
transform 1 0 66912 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1174
timestamp 1624857261
transform 1 0 67456 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1175
timestamp 1624857261
transform 1 0 67456 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1176
timestamp 1624857261
transform 1 0 67456 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1178
timestamp 1624857261
transform 1 0 67456 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5305
timestamp 1624857261
transform 1 0 1224 0 1 13877
box 0 0 1 1
use contact_13  contact_13_737
timestamp 1624857261
transform 1 0 1801 0 1 13443
box 0 0 1 1
use contact_19  contact_19_737
timestamp 1624857261
transform 1 0 1794 0 1 13452
box 0 0 1 1
use contact_14  contact_14_737
timestamp 1624857261
transform 1 0 1797 0 1 13451
box 0 0 1 1
use contact_13  contact_13_736
timestamp 1624857261
transform 1 0 1801 0 1 13779
box 0 0 1 1
use contact_19  contact_19_736
timestamp 1624857261
transform 1 0 1794 0 1 13788
box 0 0 1 1
use contact_14  contact_14_736
timestamp 1624857261
transform 1 0 1797 0 1 13787
box 0 0 1 1
use contact_7  contact_7_148
timestamp 1624857261
transform 1 0 1793 0 1 13783
box 0 0 1 1
use contact_13  contact_13_735
timestamp 1624857261
transform 1 0 1801 0 1 14115
box 0 0 1 1
use contact_19  contact_19_735
timestamp 1624857261
transform 1 0 1794 0 1 14124
box 0 0 1 1
use contact_14  contact_14_735
timestamp 1624857261
transform 1 0 1797 0 1 14123
box 0 0 1 1
use contact_13  contact_13_734
timestamp 1624857261
transform 1 0 1801 0 1 14451
box 0 0 1 1
use contact_19  contact_19_734
timestamp 1624857261
transform 1 0 1794 0 1 14460
box 0 0 1 1
use contact_14  contact_14_734
timestamp 1624857261
transform 1 0 1797 0 1 14459
box 0 0 1 1
use contact_33  contact_33_5306
timestamp 1624857261
transform 1 0 3128 0 1 13333
box 0 0 1 1
use contact_33  contact_33_5307
timestamp 1624857261
transform 1 0 3128 0 1 13741
box 0 0 1 1
use contact_7  contact_7_488
timestamp 1624857261
transform 1 0 15205 0 1 13946
box 0 0 1 1
use contact_33  contact_33_2328
timestamp 1624857261
transform 1 0 15232 0 1 13333
box 0 0 1 1
use contact_33  contact_33_1902
timestamp 1624857261
transform 1 0 22168 0 1 14285
box 0 0 1 1
use contact_7  contact_7_487
timestamp 1624857261
transform 1 0 27698 0 1 13946
box 0 0 1 1
use contact_33  contact_33_4294
timestamp 1624857261
transform 1 0 29920 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4295
timestamp 1624857261
transform 1 0 29920 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4298
timestamp 1624857261
transform 1 0 29920 0 1 13469
box 0 0 1 1
use contact_33  contact_33_4270
timestamp 1624857261
transform 1 0 32368 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4271
timestamp 1624857261
transform 1 0 32368 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4272
timestamp 1624857261
transform 1 0 32368 0 1 13469
box 0 0 1 1
use contact_33  contact_33_4242
timestamp 1624857261
transform 1 0 34816 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4243
timestamp 1624857261
transform 1 0 34816 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4244
timestamp 1624857261
transform 1 0 34680 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4214
timestamp 1624857261
transform 1 0 37400 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4215
timestamp 1624857261
transform 1 0 37400 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4216
timestamp 1624857261
transform 1 0 37264 0 1 13469
box 0 0 1 1
use contact_33  contact_33_4184
timestamp 1624857261
transform 1 0 39848 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4185
timestamp 1624857261
transform 1 0 39848 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4188
timestamp 1624857261
transform 1 0 39712 0 1 13469
box 0 0 1 1
use contact_33  contact_33_4164
timestamp 1624857261
transform 1 0 42160 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4165
timestamp 1624857261
transform 1 0 42160 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4166
timestamp 1624857261
transform 1 0 42432 0 1 13469
box 0 0 1 1
use contact_33  contact_33_4132
timestamp 1624857261
transform 1 0 44880 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4133
timestamp 1624857261
transform 1 0 44880 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4134
timestamp 1624857261
transform 1 0 44880 0 1 13469
box 0 0 1 1
use contact_33  contact_33_4108
timestamp 1624857261
transform 1 0 47192 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4109
timestamp 1624857261
transform 1 0 47192 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4112
timestamp 1624857261
transform 1 0 47328 0 1 13469
box 0 0 1 1
use contact_33  contact_33_4074
timestamp 1624857261
transform 1 0 49776 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4075
timestamp 1624857261
transform 1 0 49776 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4078
timestamp 1624857261
transform 1 0 49640 0 1 13605
box 0 0 1 1
use contact_33  contact_33_5406
timestamp 1624857261
transform 1 0 49912 0 1 13333
box 0 0 1 1
use contact_33  contact_33_4054
timestamp 1624857261
transform 1 0 52224 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4055
timestamp 1624857261
transform 1 0 52224 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4056
timestamp 1624857261
transform 1 0 52224 0 1 13469
box 0 0 1 1
use contact_33  contact_33_4024
timestamp 1624857261
transform 1 0 54808 0 1 13605
box 0 0 1 1
use contact_33  contact_33_4025
timestamp 1624857261
transform 1 0 54808 0 1 14285
box 0 0 1 1
use contact_33  contact_33_4026
timestamp 1624857261
transform 1 0 54808 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3994
timestamp 1624857261
transform 1 0 57392 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3995
timestamp 1624857261
transform 1 0 57392 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3998
timestamp 1624857261
transform 1 0 57392 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3966
timestamp 1624857261
transform 1 0 59840 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3967
timestamp 1624857261
transform 1 0 59840 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3968
timestamp 1624857261
transform 1 0 59840 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3942
timestamp 1624857261
transform 1 0 62288 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3943
timestamp 1624857261
transform 1 0 62288 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3944
timestamp 1624857261
transform 1 0 62288 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3912
timestamp 1624857261
transform 1 0 64736 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3908
timestamp 1624857261
transform 1 0 64872 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3909
timestamp 1624857261
transform 1 0 64872 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3886
timestamp 1624857261
transform 1 0 67184 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3887
timestamp 1624857261
transform 1 0 67184 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3890
timestamp 1624857261
transform 1 0 67320 0 1 13469
box 0 0 1 1
use contact_33  contact_33_2345
timestamp 1624857261
transform 1 0 544 0 1 14693
box 0 0 1 1
use contact_33  contact_33_5319
timestamp 1624857261
transform 1 0 1224 0 1 15509
box 0 0 1 1
use contact_13  contact_13_733
timestamp 1624857261
transform 1 0 1801 0 1 14787
box 0 0 1 1
use contact_19  contact_19_733
timestamp 1624857261
transform 1 0 1794 0 1 14796
box 0 0 1 1
use contact_14  contact_14_733
timestamp 1624857261
transform 1 0 1797 0 1 14795
box 0 0 1 1
use contact_13  contact_13_732
timestamp 1624857261
transform 1 0 1801 0 1 15123
box 0 0 1 1
use contact_19  contact_19_732
timestamp 1624857261
transform 1 0 1794 0 1 15132
box 0 0 1 1
use contact_14  contact_14_732
timestamp 1624857261
transform 1 0 1797 0 1 15131
box 0 0 1 1
use contact_13  contact_13_731
timestamp 1624857261
transform 1 0 1801 0 1 15459
box 0 0 1 1
use contact_19  contact_19_731
timestamp 1624857261
transform 1 0 1794 0 1 15468
box 0 0 1 1
use contact_14  contact_14_731
timestamp 1624857261
transform 1 0 1797 0 1 15467
box 0 0 1 1
use contact_7  contact_7_147
timestamp 1624857261
transform 1 0 1793 0 1 15463
box 0 0 1 1
use contact_33  contact_33_5321
timestamp 1624857261
transform 1 0 3128 0 1 15509
box 0 0 1 1
use contact_33  contact_33_5249
timestamp 1624857261
transform 1 0 15096 0 1 14693
box 0 0 1 1
use contact_33  contact_33_5250
timestamp 1624857261
transform 1 0 15096 0 1 14557
box 0 0 1 1
use contact_7  contact_7_486
timestamp 1624857261
transform 1 0 15205 0 1 15360
box 0 0 1 1
use contact_33  contact_33_2284
timestamp 1624857261
transform 1 0 21080 0 1 14557
box 0 0 1 1
use contact_7  contact_7_485
timestamp 1624857261
transform 1 0 27450 0 1 15360
box 0 0 1 1
use contact_33  contact_33_1350
timestamp 1624857261
transform 1 0 29920 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1351
timestamp 1624857261
transform 1 0 30056 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1339
timestamp 1624857261
transform 1 0 32504 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1336
timestamp 1624857261
transform 1 0 32640 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1327
timestamp 1624857261
transform 1 0 34952 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1324
timestamp 1624857261
transform 1 0 35088 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1314
timestamp 1624857261
transform 1 0 37400 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1315
timestamp 1624857261
transform 1 0 37536 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1300
timestamp 1624857261
transform 1 0 40120 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1305
timestamp 1624857261
transform 1 0 39984 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1290
timestamp 1624857261
transform 1 0 42432 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1291
timestamp 1624857261
transform 1 0 42568 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1276
timestamp 1624857261
transform 1 0 44880 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1281
timestamp 1624857261
transform 1 0 45016 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1266
timestamp 1624857261
transform 1 0 47600 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1269
timestamp 1624857261
transform 1 0 47464 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1254
timestamp 1624857261
transform 1 0 49912 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1257
timestamp 1624857261
transform 1 0 50184 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1245
timestamp 1624857261
transform 1 0 52360 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1242
timestamp 1624857261
transform 1 0 52496 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1228
timestamp 1624857261
transform 1 0 55080 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1233
timestamp 1624857261
transform 1 0 54944 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1216
timestamp 1624857261
transform 1 0 57392 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1221
timestamp 1624857261
transform 1 0 57528 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1204
timestamp 1624857261
transform 1 0 59840 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1209
timestamp 1624857261
transform 1 0 59976 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1194
timestamp 1624857261
transform 1 0 62560 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1197
timestamp 1624857261
transform 1 0 62424 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1182
timestamp 1624857261
transform 1 0 64872 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1185
timestamp 1624857261
transform 1 0 65008 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1168
timestamp 1624857261
transform 1 0 67592 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1173
timestamp 1624857261
transform 1 0 67456 0 1 15101
box 0 0 1 1
use contact_13  contact_13_730
timestamp 1624857261
transform 1 0 1801 0 1 15795
box 0 0 1 1
use contact_19  contact_19_730
timestamp 1624857261
transform 1 0 1794 0 1 15804
box 0 0 1 1
use contact_14  contact_14_730
timestamp 1624857261
transform 1 0 1797 0 1 15803
box 0 0 1 1
use contact_13  contact_13_729
timestamp 1624857261
transform 1 0 1801 0 1 16131
box 0 0 1 1
use contact_19  contact_19_729
timestamp 1624857261
transform 1 0 1794 0 1 16140
box 0 0 1 1
use contact_14  contact_14_729
timestamp 1624857261
transform 1 0 1797 0 1 16139
box 0 0 1 1
use contact_13  contact_13_728
timestamp 1624857261
transform 1 0 1801 0 1 16467
box 0 0 1 1
use contact_19  contact_19_728
timestamp 1624857261
transform 1 0 1794 0 1 16476
box 0 0 1 1
use contact_14  contact_14_728
timestamp 1624857261
transform 1 0 1797 0 1 16475
box 0 0 1 1
use contact_13  contact_13_727
timestamp 1624857261
transform 1 0 1801 0 1 16803
box 0 0 1 1
use contact_19  contact_19_727
timestamp 1624857261
transform 1 0 1794 0 1 16812
box 0 0 1 1
use contact_14  contact_14_727
timestamp 1624857261
transform 1 0 1797 0 1 16811
box 0 0 1 1
use contact_33  contact_33_5320
timestamp 1624857261
transform 1 0 3128 0 1 16053
box 0 0 1 1
use contact_33  contact_33_2326
timestamp 1624857261
transform 1 0 15232 0 1 16189
box 0 0 1 1
use contact_33  contact_33_2327
timestamp 1624857261
transform 1 0 15232 0 1 16053
box 0 0 1 1
use contact_33  contact_33_4900
timestamp 1624857261
transform 1 0 22304 0 1 15781
box 0 0 1 1
use contact_33  contact_33_4899
timestamp 1624857261
transform 1 0 23392 0 1 15781
box 0 0 1 1
use contact_33  contact_33_5356
timestamp 1624857261
transform 1 0 1224 0 1 17005
box 0 0 1 1
use contact_13  contact_13_726
timestamp 1624857261
transform 1 0 1801 0 1 17139
box 0 0 1 1
use contact_19  contact_19_726
timestamp 1624857261
transform 1 0 1794 0 1 17148
box 0 0 1 1
use contact_14  contact_14_726
timestamp 1624857261
transform 1 0 1797 0 1 17147
box 0 0 1 1
use contact_7  contact_7_146
timestamp 1624857261
transform 1 0 1793 0 1 17143
box 0 0 1 1
use contact_13  contact_13_725
timestamp 1624857261
transform 1 0 1801 0 1 17475
box 0 0 1 1
use contact_19  contact_19_725
timestamp 1624857261
transform 1 0 1794 0 1 17484
box 0 0 1 1
use contact_14  contact_14_725
timestamp 1624857261
transform 1 0 1797 0 1 17483
box 0 0 1 1
use contact_13  contact_13_724
timestamp 1624857261
transform 1 0 1801 0 1 17811
box 0 0 1 1
use contact_19  contact_19_724
timestamp 1624857261
transform 1 0 1794 0 1 17820
box 0 0 1 1
use contact_14  contact_14_724
timestamp 1624857261
transform 1 0 1797 0 1 17819
box 0 0 1 1
use contact_33  contact_33_5494
timestamp 1624857261
transform 1 0 2535 0 1 17893
box 0 0 1 1
use contact_13  contact_13_723
timestamp 1624857261
transform 1 0 1801 0 1 18147
box 0 0 1 1
use contact_19  contact_19_723
timestamp 1624857261
transform 1 0 1794 0 1 18156
box 0 0 1 1
use contact_14  contact_14_723
timestamp 1624857261
transform 1 0 1797 0 1 18155
box 0 0 1 1
use contact_33  contact_33_2344
timestamp 1624857261
transform 1 0 3808 0 1 17549
box 0 0 1 1
use contact_33  contact_33_5248
timestamp 1624857261
transform 1 0 15096 0 1 17413
box 0 0 1 1
use contact_7  contact_7_484
timestamp 1624857261
transform 1 0 15205 0 1 18188
box 0 0 1 1
use contact_33  contact_33_5247
timestamp 1624857261
transform 1 0 17544 0 1 17549
box 0 0 1 1
use contact_33  contact_33_2283
timestamp 1624857261
transform 1 0 21080 0 1 17141
box 0 0 1 1
use contact_33  contact_33_2282
timestamp 1624857261
transform 1 0 21760 0 1 17277
box 0 0 1 1
use contact_7  contact_7_483
timestamp 1624857261
transform 1 0 23747 0 1 18188
box 0 0 1 1
use contact_33  contact_33_1349
timestamp 1624857261
transform 1 0 29920 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1335
timestamp 1624857261
transform 1 0 32640 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1323
timestamp 1624857261
transform 1 0 35088 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1313
timestamp 1624857261
transform 1 0 37400 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1299
timestamp 1624857261
transform 1 0 40120 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1289
timestamp 1624857261
transform 1 0 42432 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1275
timestamp 1624857261
transform 1 0 44880 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1265
timestamp 1624857261
transform 1 0 47600 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1253
timestamp 1624857261
transform 1 0 49912 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1241
timestamp 1624857261
transform 1 0 52496 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1227
timestamp 1624857261
transform 1 0 55080 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1215
timestamp 1624857261
transform 1 0 57392 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1203
timestamp 1624857261
transform 1 0 59976 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1193
timestamp 1624857261
transform 1 0 62560 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1181
timestamp 1624857261
transform 1 0 64872 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1167
timestamp 1624857261
transform 1 0 67592 0 1 17005
box 0 0 1 1
use contact_14  contact_14_722
timestamp 1624857261
transform 1 0 1797 0 1 18491
box 0 0 1 1
use contact_19  contact_19_722
timestamp 1624857261
transform 1 0 1794 0 1 18492
box 0 0 1 1
use contact_13  contact_13_722
timestamp 1624857261
transform 1 0 1801 0 1 18483
box 0 0 1 1
use cr_3  cr_3_0
timestamp 1624857261
transform 1 0 15406 0 1 9422
box 2083 -3939 6102 5492
use control_logic_rw  control_logic_rw_0
timestamp 1624857261
transform 1 0 2616 0 1 7620
box -75 -49 11650 18431
use contact_33  contact_33_5346
timestamp 1624857261
transform 1 0 1224 0 1 18909
box 0 0 1 1
use contact_33  contact_33_2346
timestamp 1624857261
transform 1 0 544 0 1 20269
box 0 0 1 1
use contact_33  contact_33_5379
timestamp 1624857261
transform 1 0 1224 0 1 20405
box 0 0 1 1
use contact_33  contact_33_5327
timestamp 1624857261
transform 1 0 1224 0 1 22309
box 0 0 1 1
use contact_33  contact_33_5365
timestamp 1624857261
transform 1 0 1224 0 1 23941
box 0 0 1 1
use contact_33  contact_33_2347
timestamp 1624857261
transform 1 0 544 0 1 25845
box 0 0 1 1
use contact_33  contact_33_5340
timestamp 1624857261
transform 1 0 1224 0 1 25573
box 0 0 1 1
use contact_33  contact_33_5335
timestamp 1624857261
transform 1 0 1224 0 1 27341
box 0 0 1 1
use contact_33  contact_33_5359
timestamp 1624857261
transform 1 0 1224 0 1 28837
box 0 0 1 1
use contact_33  contact_33_5368
timestamp 1624857261
transform 1 0 1224 0 1 30605
box 0 0 1 1
use contact_33  contact_33_5315
timestamp 1624857261
transform 1 0 1224 0 1 32373
box 0 0 1 1
use contact_33  contact_33_5344
timestamp 1624857261
transform 1 0 1224 0 1 34005
box 0 0 1 1
use contact_33  contact_33_5353
timestamp 1624857261
transform 1 0 1224 0 1 35773
box 0 0 1 1
use contact_7  contact_7_145
timestamp 1624857261
transform 1 0 1793 0 1 18823
box 0 0 1 1
use contact_14  contact_14_721
timestamp 1624857261
transform 1 0 1797 0 1 18827
box 0 0 1 1
use contact_19  contact_19_721
timestamp 1624857261
transform 1 0 1794 0 1 18828
box 0 0 1 1
use contact_13  contact_13_721
timestamp 1624857261
transform 1 0 1801 0 1 18819
box 0 0 1 1
use contact_14  contact_14_720
timestamp 1624857261
transform 1 0 1797 0 1 19163
box 0 0 1 1
use contact_19  contact_19_720
timestamp 1624857261
transform 1 0 1794 0 1 19164
box 0 0 1 1
use contact_13  contact_13_720
timestamp 1624857261
transform 1 0 1801 0 1 19155
box 0 0 1 1
use contact_14  contact_14_719
timestamp 1624857261
transform 1 0 1797 0 1 19499
box 0 0 1 1
use contact_19  contact_19_719
timestamp 1624857261
transform 1 0 1794 0 1 19500
box 0 0 1 1
use contact_13  contact_13_719
timestamp 1624857261
transform 1 0 1801 0 1 19491
box 0 0 1 1
use contact_14  contact_14_717
timestamp 1624857261
transform 1 0 1797 0 1 20171
box 0 0 1 1
use contact_14  contact_14_718
timestamp 1624857261
transform 1 0 1797 0 1 19835
box 0 0 1 1
use contact_19  contact_19_717
timestamp 1624857261
transform 1 0 1794 0 1 20172
box 0 0 1 1
use contact_19  contact_19_718
timestamp 1624857261
transform 1 0 1794 0 1 19836
box 0 0 1 1
use contact_13  contact_13_717
timestamp 1624857261
transform 1 0 1801 0 1 20163
box 0 0 1 1
use contact_13  contact_13_718
timestamp 1624857261
transform 1 0 1801 0 1 19827
box 0 0 1 1
use contact_7  contact_7_144
timestamp 1624857261
transform 1 0 1793 0 1 20503
box 0 0 1 1
use contact_14  contact_14_716
timestamp 1624857261
transform 1 0 1797 0 1 20507
box 0 0 1 1
use contact_19  contact_19_716
timestamp 1624857261
transform 1 0 1794 0 1 20508
box 0 0 1 1
use contact_13  contact_13_716
timestamp 1624857261
transform 1 0 1801 0 1 20499
box 0 0 1 1
use contact_14  contact_14_715
timestamp 1624857261
transform 1 0 1797 0 1 20843
box 0 0 1 1
use contact_19  contact_19_715
timestamp 1624857261
transform 1 0 1794 0 1 20844
box 0 0 1 1
use contact_13  contact_13_715
timestamp 1624857261
transform 1 0 1801 0 1 20835
box 0 0 1 1
use contact_14  contact_14_714
timestamp 1624857261
transform 1 0 1797 0 1 21179
box 0 0 1 1
use contact_19  contact_19_714
timestamp 1624857261
transform 1 0 1794 0 1 21180
box 0 0 1 1
use contact_13  contact_13_714
timestamp 1624857261
transform 1 0 1801 0 1 21171
box 0 0 1 1
use contact_14  contact_14_713
timestamp 1624857261
transform 1 0 1797 0 1 21515
box 0 0 1 1
use contact_19  contact_19_713
timestamp 1624857261
transform 1 0 1794 0 1 21516
box 0 0 1 1
use contact_13  contact_13_713
timestamp 1624857261
transform 1 0 1801 0 1 21507
box 0 0 1 1
use contact_14  contact_14_712
timestamp 1624857261
transform 1 0 1797 0 1 21851
box 0 0 1 1
use contact_19  contact_19_712
timestamp 1624857261
transform 1 0 1794 0 1 21852
box 0 0 1 1
use contact_13  contact_13_712
timestamp 1624857261
transform 1 0 1801 0 1 21843
box 0 0 1 1
use contact_7  contact_7_143
timestamp 1624857261
transform 1 0 1793 0 1 22183
box 0 0 1 1
use contact_14  contact_14_711
timestamp 1624857261
transform 1 0 1797 0 1 22187
box 0 0 1 1
use contact_19  contact_19_711
timestamp 1624857261
transform 1 0 1794 0 1 22188
box 0 0 1 1
use contact_13  contact_13_711
timestamp 1624857261
transform 1 0 1801 0 1 22179
box 0 0 1 1
use contact_14  contact_14_710
timestamp 1624857261
transform 1 0 1797 0 1 22523
box 0 0 1 1
use contact_19  contact_19_710
timestamp 1624857261
transform 1 0 1794 0 1 22524
box 0 0 1 1
use contact_13  contact_13_710
timestamp 1624857261
transform 1 0 1801 0 1 22515
box 0 0 1 1
use contact_14  contact_14_709
timestamp 1624857261
transform 1 0 1797 0 1 22859
box 0 0 1 1
use contact_19  contact_19_709
timestamp 1624857261
transform 1 0 1794 0 1 22860
box 0 0 1 1
use contact_13  contact_13_709
timestamp 1624857261
transform 1 0 1801 0 1 22851
box 0 0 1 1
use contact_14  contact_14_708
timestamp 1624857261
transform 1 0 1797 0 1 23195
box 0 0 1 1
use contact_19  contact_19_708
timestamp 1624857261
transform 1 0 1794 0 1 23196
box 0 0 1 1
use contact_13  contact_13_708
timestamp 1624857261
transform 1 0 1801 0 1 23187
box 0 0 1 1
use contact_14  contact_14_707
timestamp 1624857261
transform 1 0 1797 0 1 23531
box 0 0 1 1
use contact_19  contact_19_707
timestamp 1624857261
transform 1 0 1794 0 1 23532
box 0 0 1 1
use contact_13  contact_13_707
timestamp 1624857261
transform 1 0 1801 0 1 23523
box 0 0 1 1
use contact_7  contact_7_142
timestamp 1624857261
transform 1 0 1793 0 1 23863
box 0 0 1 1
use contact_14  contact_14_706
timestamp 1624857261
transform 1 0 1797 0 1 23867
box 0 0 1 1
use contact_19  contact_19_706
timestamp 1624857261
transform 1 0 1794 0 1 23868
box 0 0 1 1
use contact_13  contact_13_706
timestamp 1624857261
transform 1 0 1801 0 1 23859
box 0 0 1 1
use contact_33  contact_33_5367
timestamp 1624857261
transform 1 0 2312 0 1 23941
box 0 0 1 1
use contact_14  contact_14_705
timestamp 1624857261
transform 1 0 1797 0 1 24203
box 0 0 1 1
use contact_19  contact_19_705
timestamp 1624857261
transform 1 0 1794 0 1 24204
box 0 0 1 1
use contact_13  contact_13_705
timestamp 1624857261
transform 1 0 1801 0 1 24195
box 0 0 1 1
use contact_14  contact_14_704
timestamp 1624857261
transform 1 0 1797 0 1 24539
box 0 0 1 1
use contact_19  contact_19_704
timestamp 1624857261
transform 1 0 1794 0 1 24540
box 0 0 1 1
use contact_13  contact_13_704
timestamp 1624857261
transform 1 0 1801 0 1 24531
box 0 0 1 1
use contact_33  contact_33_5366
timestamp 1624857261
transform 1 0 2312 0 1 24485
box 0 0 1 1
use contact_14  contact_14_703
timestamp 1624857261
transform 1 0 1797 0 1 24875
box 0 0 1 1
use contact_19  contact_19_703
timestamp 1624857261
transform 1 0 1794 0 1 24876
box 0 0 1 1
use contact_13  contact_13_703
timestamp 1624857261
transform 1 0 1801 0 1 24867
box 0 0 1 1
use contact_14  contact_14_702
timestamp 1624857261
transform 1 0 1797 0 1 25211
box 0 0 1 1
use contact_19  contact_19_702
timestamp 1624857261
transform 1 0 1794 0 1 25212
box 0 0 1 1
use contact_13  contact_13_702
timestamp 1624857261
transform 1 0 1801 0 1 25203
box 0 0 1 1
use contact_7  contact_7_476
timestamp 1624857261
transform 1 0 2540 0 1 25296
box 0 0 1 1
use contact_33  contact_33_5493
timestamp 1624857261
transform 1 0 2535 0 1 25300
box 0 0 1 1
use contact_7  contact_7_141
timestamp 1624857261
transform 1 0 1793 0 1 25543
box 0 0 1 1
use contact_14  contact_14_701
timestamp 1624857261
transform 1 0 1797 0 1 25547
box 0 0 1 1
use contact_19  contact_19_701
timestamp 1624857261
transform 1 0 1794 0 1 25548
box 0 0 1 1
use contact_13  contact_13_700
timestamp 1624857261
transform 1 0 1801 0 1 25875
box 0 0 1 1
use contact_13  contact_13_701
timestamp 1624857261
transform 1 0 1801 0 1 25539
box 0 0 1 1
use contact_14  contact_14_699
timestamp 1624857261
transform 1 0 1797 0 1 26219
box 0 0 1 1
use contact_14  contact_14_700
timestamp 1624857261
transform 1 0 1797 0 1 25883
box 0 0 1 1
use contact_19  contact_19_699
timestamp 1624857261
transform 1 0 1794 0 1 26220
box 0 0 1 1
use contact_19  contact_19_700
timestamp 1624857261
transform 1 0 1794 0 1 25884
box 0 0 1 1
use contact_13  contact_13_699
timestamp 1624857261
transform 1 0 1801 0 1 26211
box 0 0 1 1
use contact_14  contact_14_698
timestamp 1624857261
transform 1 0 1797 0 1 26555
box 0 0 1 1
use contact_19  contact_19_698
timestamp 1624857261
transform 1 0 1794 0 1 26556
box 0 0 1 1
use contact_13  contact_13_698
timestamp 1624857261
transform 1 0 1801 0 1 26547
box 0 0 1 1
use contact_14  contact_14_697
timestamp 1624857261
transform 1 0 1797 0 1 26891
box 0 0 1 1
use contact_19  contact_19_697
timestamp 1624857261
transform 1 0 1794 0 1 26892
box 0 0 1 1
use contact_13  contact_13_697
timestamp 1624857261
transform 1 0 1801 0 1 26883
box 0 0 1 1
use contact_7  contact_7_140
timestamp 1624857261
transform 1 0 1793 0 1 27223
box 0 0 1 1
use contact_14  contact_14_696
timestamp 1624857261
transform 1 0 1797 0 1 27227
box 0 0 1 1
use contact_19  contact_19_696
timestamp 1624857261
transform 1 0 1794 0 1 27228
box 0 0 1 1
use contact_13  contact_13_696
timestamp 1624857261
transform 1 0 1801 0 1 27219
box 0 0 1 1
use contact_14  contact_14_695
timestamp 1624857261
transform 1 0 1797 0 1 27563
box 0 0 1 1
use contact_19  contact_19_695
timestamp 1624857261
transform 1 0 1794 0 1 27564
box 0 0 1 1
use contact_13  contact_13_695
timestamp 1624857261
transform 1 0 1801 0 1 27555
box 0 0 1 1
use contact_14  contact_14_694
timestamp 1624857261
transform 1 0 1797 0 1 27899
box 0 0 1 1
use contact_19  contact_19_694
timestamp 1624857261
transform 1 0 1794 0 1 27900
box 0 0 1 1
use contact_13  contact_13_694
timestamp 1624857261
transform 1 0 1801 0 1 27891
box 0 0 1 1
use contact_14  contact_14_693
timestamp 1624857261
transform 1 0 1797 0 1 28235
box 0 0 1 1
use contact_19  contact_19_693
timestamp 1624857261
transform 1 0 1794 0 1 28236
box 0 0 1 1
use contact_13  contact_13_693
timestamp 1624857261
transform 1 0 1801 0 1 28227
box 0 0 1 1
use contact_14  contact_14_692
timestamp 1624857261
transform 1 0 1797 0 1 28571
box 0 0 1 1
use contact_19  contact_19_692
timestamp 1624857261
transform 1 0 1794 0 1 28572
box 0 0 1 1
use contact_13  contact_13_692
timestamp 1624857261
transform 1 0 1801 0 1 28563
box 0 0 1 1
use contact_7  contact_7_139
timestamp 1624857261
transform 1 0 1793 0 1 28903
box 0 0 1 1
use contact_14  contact_14_691
timestamp 1624857261
transform 1 0 1797 0 1 28907
box 0 0 1 1
use contact_19  contact_19_691
timestamp 1624857261
transform 1 0 1794 0 1 28908
box 0 0 1 1
use contact_13  contact_13_691
timestamp 1624857261
transform 1 0 1801 0 1 28899
box 0 0 1 1
use contact_14  contact_14_690
timestamp 1624857261
transform 1 0 1797 0 1 29243
box 0 0 1 1
use contact_19  contact_19_690
timestamp 1624857261
transform 1 0 1794 0 1 29244
box 0 0 1 1
use contact_13  contact_13_690
timestamp 1624857261
transform 1 0 1801 0 1 29235
box 0 0 1 1
use contact_14  contact_14_689
timestamp 1624857261
transform 1 0 1797 0 1 29579
box 0 0 1 1
use contact_19  contact_19_689
timestamp 1624857261
transform 1 0 1794 0 1 29580
box 0 0 1 1
use contact_13  contact_13_689
timestamp 1624857261
transform 1 0 1801 0 1 29571
box 0 0 1 1
use contact_14  contact_14_688
timestamp 1624857261
transform 1 0 1797 0 1 29915
box 0 0 1 1
use contact_19  contact_19_688
timestamp 1624857261
transform 1 0 1794 0 1 29916
box 0 0 1 1
use contact_13  contact_13_688
timestamp 1624857261
transform 1 0 1801 0 1 29907
box 0 0 1 1
use contact_14  contact_14_687
timestamp 1624857261
transform 1 0 1797 0 1 30251
box 0 0 1 1
use contact_19  contact_19_687
timestamp 1624857261
transform 1 0 1794 0 1 30252
box 0 0 1 1
use contact_13  contact_13_687
timestamp 1624857261
transform 1 0 1801 0 1 30243
box 0 0 1 1
use contact_7  contact_7_138
timestamp 1624857261
transform 1 0 1793 0 1 30583
box 0 0 1 1
use contact_14  contact_14_686
timestamp 1624857261
transform 1 0 1797 0 1 30587
box 0 0 1 1
use contact_19  contact_19_686
timestamp 1624857261
transform 1 0 1794 0 1 30588
box 0 0 1 1
use contact_13  contact_13_686
timestamp 1624857261
transform 1 0 1801 0 1 30579
box 0 0 1 1
use contact_14  contact_14_685
timestamp 1624857261
transform 1 0 1797 0 1 30923
box 0 0 1 1
use contact_19  contact_19_685
timestamp 1624857261
transform 1 0 1794 0 1 30924
box 0 0 1 1
use contact_13  contact_13_685
timestamp 1624857261
transform 1 0 1801 0 1 30915
box 0 0 1 1
use contact_14  contact_14_684
timestamp 1624857261
transform 1 0 1797 0 1 31259
box 0 0 1 1
use contact_19  contact_19_684
timestamp 1624857261
transform 1 0 1794 0 1 31260
box 0 0 1 1
use contact_13  contact_13_684
timestamp 1624857261
transform 1 0 1801 0 1 31251
box 0 0 1 1
use contact_14  contact_14_683
timestamp 1624857261
transform 1 0 1797 0 1 31595
box 0 0 1 1
use contact_19  contact_19_683
timestamp 1624857261
transform 1 0 1794 0 1 31596
box 0 0 1 1
use contact_13  contact_13_682
timestamp 1624857261
transform 1 0 1801 0 1 31923
box 0 0 1 1
use contact_13  contact_13_683
timestamp 1624857261
transform 1 0 1801 0 1 31587
box 0 0 1 1
use contact_7  contact_7_137
timestamp 1624857261
transform 1 0 1793 0 1 32263
box 0 0 1 1
use contact_14  contact_14_681
timestamp 1624857261
transform 1 0 1797 0 1 32267
box 0 0 1 1
use contact_14  contact_14_682
timestamp 1624857261
transform 1 0 1797 0 1 31931
box 0 0 1 1
use contact_19  contact_19_681
timestamp 1624857261
transform 1 0 1794 0 1 32268
box 0 0 1 1
use contact_19  contact_19_682
timestamp 1624857261
transform 1 0 1794 0 1 31932
box 0 0 1 1
use contact_13  contact_13_681
timestamp 1624857261
transform 1 0 1801 0 1 32259
box 0 0 1 1
use contact_14  contact_14_680
timestamp 1624857261
transform 1 0 1797 0 1 32603
box 0 0 1 1
use contact_19  contact_19_680
timestamp 1624857261
transform 1 0 1794 0 1 32604
box 0 0 1 1
use contact_13  contact_13_680
timestamp 1624857261
transform 1 0 1801 0 1 32595
box 0 0 1 1
use contact_14  contact_14_679
timestamp 1624857261
transform 1 0 1797 0 1 32939
box 0 0 1 1
use contact_19  contact_19_679
timestamp 1624857261
transform 1 0 1794 0 1 32940
box 0 0 1 1
use contact_13  contact_13_679
timestamp 1624857261
transform 1 0 1801 0 1 32931
box 0 0 1 1
use contact_14  contact_14_678
timestamp 1624857261
transform 1 0 1797 0 1 33275
box 0 0 1 1
use contact_19  contact_19_678
timestamp 1624857261
transform 1 0 1794 0 1 33276
box 0 0 1 1
use contact_13  contact_13_678
timestamp 1624857261
transform 1 0 1801 0 1 33267
box 0 0 1 1
use contact_14  contact_14_677
timestamp 1624857261
transform 1 0 1797 0 1 33611
box 0 0 1 1
use contact_19  contact_19_677
timestamp 1624857261
transform 1 0 1794 0 1 33612
box 0 0 1 1
use contact_13  contact_13_677
timestamp 1624857261
transform 1 0 1801 0 1 33603
box 0 0 1 1
use contact_7  contact_7_136
timestamp 1624857261
transform 1 0 1793 0 1 33943
box 0 0 1 1
use contact_14  contact_14_676
timestamp 1624857261
transform 1 0 1797 0 1 33947
box 0 0 1 1
use contact_19  contact_19_676
timestamp 1624857261
transform 1 0 1794 0 1 33948
box 0 0 1 1
use contact_13  contact_13_676
timestamp 1624857261
transform 1 0 1801 0 1 33939
box 0 0 1 1
use contact_14  contact_14_675
timestamp 1624857261
transform 1 0 1797 0 1 34283
box 0 0 1 1
use contact_19  contact_19_675
timestamp 1624857261
transform 1 0 1794 0 1 34284
box 0 0 1 1
use contact_13  contact_13_675
timestamp 1624857261
transform 1 0 1801 0 1 34275
box 0 0 1 1
use contact_14  contact_14_674
timestamp 1624857261
transform 1 0 1797 0 1 34619
box 0 0 1 1
use contact_19  contact_19_674
timestamp 1624857261
transform 1 0 1794 0 1 34620
box 0 0 1 1
use contact_13  contact_13_674
timestamp 1624857261
transform 1 0 1801 0 1 34611
box 0 0 1 1
use contact_14  contact_14_673
timestamp 1624857261
transform 1 0 1797 0 1 34955
box 0 0 1 1
use contact_19  contact_19_673
timestamp 1624857261
transform 1 0 1794 0 1 34956
box 0 0 1 1
use contact_13  contact_13_673
timestamp 1624857261
transform 1 0 1801 0 1 34947
box 0 0 1 1
use contact_14  contact_14_672
timestamp 1624857261
transform 1 0 1797 0 1 35291
box 0 0 1 1
use contact_19  contact_19_672
timestamp 1624857261
transform 1 0 1794 0 1 35292
box 0 0 1 1
use contact_13  contact_13_672
timestamp 1624857261
transform 1 0 1801 0 1 35283
box 0 0 1 1
use contact_7  contact_7_135
timestamp 1624857261
transform 1 0 1793 0 1 35623
box 0 0 1 1
use contact_14  contact_14_671
timestamp 1624857261
transform 1 0 1797 0 1 35627
box 0 0 1 1
use contact_19  contact_19_671
timestamp 1624857261
transform 1 0 1794 0 1 35628
box 0 0 1 1
use contact_13  contact_13_671
timestamp 1624857261
transform 1 0 1801 0 1 35619
box 0 0 1 1
use contact_14  contact_14_670
timestamp 1624857261
transform 1 0 1797 0 1 35963
box 0 0 1 1
use contact_19  contact_19_670
timestamp 1624857261
transform 1 0 1794 0 1 35964
box 0 0 1 1
use contact_13  contact_13_670
timestamp 1624857261
transform 1 0 1801 0 1 35955
box 0 0 1 1
use contact_14  contact_14_669
timestamp 1624857261
transform 1 0 1797 0 1 36299
box 0 0 1 1
use contact_19  contact_19_669
timestamp 1624857261
transform 1 0 1794 0 1 36300
box 0 0 1 1
use contact_13  contact_13_669
timestamp 1624857261
transform 1 0 1801 0 1 36291
box 0 0 1 1
use contact_14  contact_14_668
timestamp 1624857261
transform 1 0 1797 0 1 36635
box 0 0 1 1
use contact_19  contact_19_668
timestamp 1624857261
transform 1 0 1794 0 1 36636
box 0 0 1 1
use contact_13  contact_13_668
timestamp 1624857261
transform 1 0 1801 0 1 36627
box 0 0 1 1
use contact_14  contact_14_667
timestamp 1624857261
transform 1 0 1797 0 1 36971
box 0 0 1 1
use contact_19  contact_19_667
timestamp 1624857261
transform 1 0 1794 0 1 36972
box 0 0 1 1
use contact_13  contact_13_667
timestamp 1624857261
transform 1 0 1801 0 1 36963
box 0 0 1 1
use contact_33  contact_33_5329
timestamp 1624857261
transform 1 0 3128 0 1 22173
box 0 0 1 1
use contact_33  contact_33_5328
timestamp 1624857261
transform 1 0 3128 0 1 21765
box 0 0 1 1
use contact_33  contact_33_2349
timestamp 1624857261
transform 1 0 3808 0 1 23261
box 0 0 1 1
use contact_33  contact_33_2348
timestamp 1624857261
transform 1 0 3808 0 1 25845
box 0 0 1 1
use contact_33  contact_33_2343
timestamp 1624857261
transform 1 0 3944 0 1 20269
box 0 0 1 1
use contact_33  contact_33_2335
timestamp 1624857261
transform 1 0 14552 0 1 29381
box 0 0 1 1
use contact_7  contact_7_474
timestamp 1624857261
transform 1 0 15152 0 1 29924
box 0 0 1 1
use contact_7  contact_7_373
timestamp 1624857261
transform 1 0 14207 0 1 29853
box 0 0 1 1
use contact_33  contact_33_5262
timestamp 1624857261
transform 1 0 14688 0 1 30741
box 0 0 1 1
use contact_7  contact_7_472
timestamp 1624857261
transform 1 0 15152 0 1 31482
box 0 0 1 1
use contact_7  contact_7_372
timestamp 1624857261
transform 1 0 14207 0 1 31553
box 0 0 1 1
use contact_33  contact_33_2336
timestamp 1624857261
transform 1 0 14552 0 1 32101
box 0 0 1 1
use contact_33  contact_33_2337
timestamp 1624857261
transform 1 0 14552 0 1 32237
box 0 0 1 1
use contact_7  contact_7_470
timestamp 1624857261
transform 1 0 15152 0 1 32752
box 0 0 1 1
use contact_7  contact_7_371
timestamp 1624857261
transform 1 0 14207 0 1 32681
box 0 0 1 1
use contact_33  contact_33_5263
timestamp 1624857261
transform 1 0 14688 0 1 33461
box 0 0 1 1
use contact_33  contact_33_5261
timestamp 1624857261
transform 1 0 14688 0 1 33597
box 0 0 1 1
use contact_7  contact_7_468
timestamp 1624857261
transform 1 0 15152 0 1 34310
box 0 0 1 1
use contact_7  contact_7_370
timestamp 1624857261
transform 1 0 14207 0 1 34381
box 0 0 1 1
use contact_33  contact_33_2339
timestamp 1624857261
transform 1 0 14824 0 1 35093
box 0 0 1 1
use contact_33  contact_33_2338
timestamp 1624857261
transform 1 0 14552 0 1 34821
box 0 0 1 1
use contact_7  contact_7_369
timestamp 1624857261
transform 1 0 14207 0 1 35509
box 0 0 1 1
use contact_7  contact_7_466
timestamp 1624857261
transform 1 0 15152 0 1 35580
box 0 0 1 1
use contact_33  contact_33_5260
timestamp 1624857261
transform 1 0 14688 0 1 36317
box 0 0 1 1
use contact_33  contact_33_5256
timestamp 1624857261
transform 1 0 14552 0 1 36453
box 0 0 1 1
use contact_7  contact_7_464
timestamp 1624857261
transform 1 0 15152 0 1 37138
box 0 0 1 1
use contact_7  contact_7_368
timestamp 1624857261
transform 1 0 14207 0 1 37209
box 0 0 1 1
use row_addr_dff  row_addr_dff_1
timestamp 1624857261
transform 1 0 14070 0 1 29326
box -36 -49 1204 9951
use contact_33  contact_33_2325
timestamp 1624857261
transform 1 0 15232 0 1 18773
box 0 0 1 1
use contact_32  contact_32_3
timestamp 1624857261
transform 1 0 15289 0 1 29597
box 0 0 1 1
use contact_7  contact_7_473
timestamp 1624857261
transform 1 0 15406 0 1 29924
box 0 0 1 1
use contact_19  contact_19_1013
timestamp 1624857261
transform 1 0 15407 0 1 29929
box 0 0 1 1
use contact_7  contact_7_471
timestamp 1624857261
transform 1 0 15486 0 1 31482
box 0 0 1 1
use contact_19  contact_19_1012
timestamp 1624857261
transform 1 0 15487 0 1 31487
box 0 0 1 1
use contact_7  contact_7_469
timestamp 1624857261
transform 1 0 15566 0 1 32752
box 0 0 1 1
use contact_19  contact_19_1011
timestamp 1624857261
transform 1 0 15567 0 1 32757
box 0 0 1 1
use contact_7  contact_7_467
timestamp 1624857261
transform 1 0 15646 0 1 34310
box 0 0 1 1
use contact_19  contact_19_1010
timestamp 1624857261
transform 1 0 15647 0 1 34315
box 0 0 1 1
use contact_7  contact_7_465
timestamp 1624857261
transform 1 0 15726 0 1 35580
box 0 0 1 1
use contact_19  contact_19_1009
timestamp 1624857261
transform 1 0 15727 0 1 35585
box 0 0 1 1
use contact_7  contact_7_463
timestamp 1624857261
transform 1 0 15806 0 1 37138
box 0 0 1 1
use contact_19  contact_19_1008
timestamp 1624857261
transform 1 0 15807 0 1 37143
box 0 0 1 1
use contact_33  contact_33_5246
timestamp 1624857261
transform 1 0 17544 0 1 20133
box 0 0 1 1
use contact_33  contact_33_2334
timestamp 1624857261
transform 1 0 16592 0 1 29245
box 0 0 1 1
use contact_33  contact_33_2333
timestamp 1624857261
transform 1 0 16592 0 1 26661
box 0 0 1 1
use contact_33  contact_33_2324
timestamp 1624857261
transform 1 0 17136 0 1 19045
box 0 0 1 1
use contact_33  contact_33_2323
timestamp 1624857261
transform 1 0 17136 0 1 20133
box 0 0 1 1
use contact_33  contact_33_2306
timestamp 1624857261
transform 1 0 18632 0 1 21085
box 0 0 1 1
use contact_33  contact_33_2305
timestamp 1624857261
transform 1 0 18632 0 1 22445
box 0 0 1 1
use contact_33  contact_33_2311
timestamp 1624857261
transform 1 0 18360 0 1 23125
box 0 0 1 1
use contact_33  contact_33_2312
timestamp 1624857261
transform 1 0 18360 0 1 22717
box 0 0 1 1
use contact_33  contact_33_2319
timestamp 1624857261
transform 1 0 18224 0 1 22717
box 0 0 1 1
use contact_33  contact_33_2320
timestamp 1624857261
transform 1 0 18224 0 1 23261
box 0 0 1 1
use contact_33  contact_33_5230
timestamp 1624857261
transform 1 0 18632 0 1 23261
box 0 0 1 1
use contact_33  contact_33_5231
timestamp 1624857261
transform 1 0 18632 0 1 22717
box 0 0 1 1
use contact_33  contact_33_2321
timestamp 1624857261
transform 1 0 18224 0 1 24077
box 0 0 1 1
use contact_33  contact_33_2322
timestamp 1624857261
transform 1 0 18224 0 1 23533
box 0 0 1 1
use contact_33  contact_33_5234
timestamp 1624857261
transform 1 0 18496 0 1 23533
box 0 0 1 1
use contact_33  contact_33_5235
timestamp 1624857261
transform 1 0 18496 0 1 24077
box 0 0 1 1
use contact_33  contact_33_2313
timestamp 1624857261
transform 1 0 18224 0 1 24893
box 0 0 1 1
use contact_33  contact_33_2314
timestamp 1624857261
transform 1 0 18224 0 1 24213
box 0 0 1 1
use contact_33  contact_33_5241
timestamp 1624857261
transform 1 0 18496 0 1 26389
box 0 0 1 1
use contact_33  contact_33_2317
timestamp 1624857261
transform 1 0 18088 0 1 27205
box 0 0 1 1
use contact_33  contact_33_2318
timestamp 1624857261
transform 1 0 18088 0 1 26661
box 0 0 1 1
use contact_33  contact_33_5240
timestamp 1624857261
transform 1 0 18496 0 1 27205
box 0 0 1 1
use contact_33  contact_33_2310
timestamp 1624857261
transform 1 0 18088 0 1 27477
box 0 0 1 1
use contact_33  contact_33_2309
timestamp 1624857261
transform 1 0 18088 0 1 28021
box 0 0 1 1
use contact_33  contact_33_2315
timestamp 1624857261
transform 1 0 18088 0 1 28157
box 0 0 1 1
use contact_33  contact_33_2316
timestamp 1624857261
transform 1 0 18088 0 1 28837
box 0 0 1 1
use contact_33  contact_33_5258
timestamp 1624857261
transform 1 0 18496 0 1 28973
box 0 0 1 1
use contact_33  contact_33_5259
timestamp 1624857261
transform 1 0 18496 0 1 30605
box 0 0 1 1
use contact_33  contact_33_2301
timestamp 1624857261
transform 1 0 19312 0 1 20269
box 0 0 1 1
use contact_33  contact_33_5215
timestamp 1624857261
transform 1 0 19856 0 1 20269
box 0 0 1 1
use contact_33  contact_33_5218
timestamp 1624857261
transform 1 0 18904 0 1 20269
box 0 0 1 1
use contact_33  contact_33_2302
timestamp 1624857261
transform 1 0 19312 0 1 20949
box 0 0 1 1
use contact_33  contact_33_5204
timestamp 1624857261
transform 1 0 19856 0 1 21085
box 0 0 1 1
use contact_33  contact_33_5214
timestamp 1624857261
transform 1 0 19856 0 1 20949
box 0 0 1 1
use contact_33  contact_33_5219
timestamp 1624857261
transform 1 0 18904 0 1 20949
box 0 0 1 1
use contact_33  contact_33_5205
timestamp 1624857261
transform 1 0 19856 0 1 22445
box 0 0 1 1
use contact_33  contact_33_2287
timestamp 1624857261
transform 1 0 19312 0 1 22717
box 0 0 1 1
use contact_33  contact_33_5208
timestamp 1624857261
transform 1 0 19720 0 1 22717
box 0 0 1 1
use contact_33  contact_33_2288
timestamp 1624857261
transform 1 0 19312 0 1 23261
box 0 0 1 1
use contact_33  contact_33_5209
timestamp 1624857261
transform 1 0 19720 0 1 23261
box 0 0 1 1
use contact_33  contact_33_2295
timestamp 1624857261
transform 1 0 19312 0 1 23397
box 0 0 1 1
use contact_33  contact_33_5216
timestamp 1624857261
transform 1 0 19856 0 1 23397
box 0 0 1 1
use contact_33  contact_33_2294
timestamp 1624857261
transform 1 0 19312 0 1 24213
box 0 0 1 1
use contact_33  contact_33_2296
timestamp 1624857261
transform 1 0 19312 0 1 24077
box 0 0 1 1
use contact_33  contact_33_5217
timestamp 1624857261
transform 1 0 19856 0 1 24077
box 0 0 1 1
use contact_33  contact_33_5223
timestamp 1624857261
transform 1 0 18904 0 1 24213
box 0 0 1 1
use contact_33  contact_33_2286
timestamp 1624857261
transform 1 0 19584 0 1 25029
box 0 0 1 1
use contact_33  contact_33_2293
timestamp 1624857261
transform 1 0 19312 0 1 24893
box 0 0 1 1
use contact_33  contact_33_2297
timestamp 1624857261
transform 1 0 19448 0 1 25029
box 0 0 1 1
use contact_33  contact_33_5210
timestamp 1624857261
transform 1 0 19720 0 1 25029
box 0 0 1 1
use contact_33  contact_33_5222
timestamp 1624857261
transform 1 0 18904 0 1 24893
box 0 0 1 1
use contact_33  contact_33_2285
timestamp 1624857261
transform 1 0 19584 0 1 25301
box 0 0 1 1
use contact_33  contact_33_2298
timestamp 1624857261
transform 1 0 19448 0 1 26389
box 0 0 1 1
use contact_33  contact_33_2300
timestamp 1624857261
transform 1 0 19312 0 1 26661
box 0 0 1 1
use contact_33  contact_33_5211
timestamp 1624857261
transform 1 0 19720 0 1 26389
box 0 0 1 1
use contact_33  contact_33_5213
timestamp 1624857261
transform 1 0 19856 0 1 26661
box 0 0 1 1
use contact_33  contact_33_5232
timestamp 1624857261
transform 1 0 18904 0 1 26661
box 0 0 1 1
use contact_33  contact_33_5233
timestamp 1624857261
transform 1 0 18904 0 1 27069
box 0 0 1 1
use contact_33  contact_33_2289
timestamp 1624857261
transform 1 0 19448 0 1 27341
box 0 0 1 1
use contact_33  contact_33_2299
timestamp 1624857261
transform 1 0 19312 0 1 27205
box 0 0 1 1
use contact_33  contact_33_2307
timestamp 1624857261
transform 1 0 19312 0 1 27341
box 0 0 1 1
use contact_33  contact_33_5206
timestamp 1624857261
transform 1 0 19720 0 1 27341
box 0 0 1 1
use contact_33  contact_33_5212
timestamp 1624857261
transform 1 0 19856 0 1 27205
box 0 0 1 1
use contact_33  contact_33_5221
timestamp 1624857261
transform 1 0 19040 0 1 27477
box 0 0 1 1
use contact_33  contact_33_2308
timestamp 1624857261
transform 1 0 19312 0 1 27613
box 0 0 1 1
use contact_33  contact_33_2290
timestamp 1624857261
transform 1 0 19448 0 1 28021
box 0 0 1 1
use contact_33  contact_33_2292
timestamp 1624857261
transform 1 0 19448 0 1 28157
box 0 0 1 1
use contact_33  contact_33_5207
timestamp 1624857261
transform 1 0 19720 0 1 28021
box 0 0 1 1
use contact_33  contact_33_5220
timestamp 1624857261
transform 1 0 19040 0 1 28021
box 0 0 1 1
use contact_33  contact_33_5224
timestamp 1624857261
transform 1 0 18904 0 1 28157
box 0 0 1 1
use contact_33  contact_33_2291
timestamp 1624857261
transform 1 0 19448 0 1 28837
box 0 0 1 1
use contact_33  contact_33_5225
timestamp 1624857261
transform 1 0 18904 0 1 28837
box 0 0 1 1
use contact_33  contact_33_2281
timestamp 1624857261
transform 1 0 21760 0 1 20133
box 0 0 1 1
use contact_33  contact_33_1905
timestamp 1624857261
transform 1 0 21896 0 1 20269
box 0 0 1 1
use contact_33  contact_33_5088
timestamp 1624857261
transform 1 0 22304 0 1 20269
box 0 0 1 1
use contact_33  contact_33_2031
timestamp 1624857261
transform 1 0 21760 0 1 20677
box 0 0 1 1
use contact_33  contact_33_1906
timestamp 1624857261
transform 1 0 21896 0 1 20541
box 0 0 1 1
use contact_33  contact_33_5089
timestamp 1624857261
transform 1 0 22304 0 1 20541
box 0 0 1 1
use contact_33  contact_33_2032
timestamp 1624857261
transform 1 0 21760 0 1 20949
box 0 0 1 1
use contact_33  contact_33_2177
timestamp 1624857261
transform 1 0 21896 0 1 21085
box 0 0 1 1
use contact_33  contact_33_5108
timestamp 1624857261
transform 1 0 22440 0 1 21085
box 0 0 1 1
use contact_33  contact_33_5110
timestamp 1624857261
transform 1 0 22304 0 1 21085
box 0 0 1 1
use contact_33  contact_33_2176
timestamp 1624857261
transform 1 0 21896 0 1 21493
box 0 0 1 1
use contact_33  contact_33_2178
timestamp 1624857261
transform 1 0 21896 0 1 21357
box 0 0 1 1
use contact_33  contact_33_5109
timestamp 1624857261
transform 1 0 22440 0 1 21357
box 0 0 1 1
use contact_33  contact_33_5111
timestamp 1624857261
transform 1 0 22304 0 1 21357
box 0 0 1 1
use contact_33  contact_33_5113
timestamp 1624857261
transform 1 0 22304 0 1 21493
box 0 0 1 1
use contact_33  contact_33_2249
timestamp 1624857261
transform 1 0 21760 0 1 21901
box 0 0 1 1
use contact_33  contact_33_2175
timestamp 1624857261
transform 1 0 21896 0 1 21765
box 0 0 1 1
use contact_33  contact_33_5112
timestamp 1624857261
transform 1 0 22304 0 1 21765
box 0 0 1 1
use contact_33  contact_33_2250
timestamp 1624857261
transform 1 0 21760 0 1 22173
box 0 0 1 1
use contact_33  contact_33_2252
timestamp 1624857261
transform 1 0 21760 0 1 22309
box 0 0 1 1
use contact_33  contact_33_4946
timestamp 1624857261
transform 1 0 22440 0 1 22309
box 0 0 1 1
use contact_33  contact_33_2097
timestamp 1624857261
transform 1 0 21760 0 1 22717
box 0 0 1 1
use contact_33  contact_33_2251
timestamp 1624857261
transform 1 0 21760 0 1 22581
box 0 0 1 1
use contact_33  contact_33_4947
timestamp 1624857261
transform 1 0 22440 0 1 22581
box 0 0 1 1
use contact_33  contact_33_2098
timestamp 1624857261
transform 1 0 21760 0 1 22989
box 0 0 1 1
use contact_33  contact_33_5102
timestamp 1624857261
transform 1 0 22168 0 1 22989
box 0 0 1 1
use contact_33  contact_33_5103
timestamp 1624857261
transform 1 0 22168 0 1 23261
box 0 0 1 1
use contact_33  contact_33_4804
timestamp 1624857261
transform 1 0 22576 0 1 23261
box 0 0 1 1
use contact_33  contact_33_4805
timestamp 1624857261
transform 1 0 22576 0 1 22989
box 0 0 1 1
use contact_33  contact_33_4758
timestamp 1624857261
transform 1 0 22576 0 1 23805
box 0 0 1 1
use contact_33  contact_33_4759
timestamp 1624857261
transform 1 0 22576 0 1 24077
box 0 0 1 1
use contact_33  contact_33_5170
timestamp 1624857261
transform 1 0 22304 0 1 24077
box 0 0 1 1
use contact_33  contact_33_5171
timestamp 1624857261
transform 1 0 22304 0 1 23805
box 0 0 1 1
use contact_33  contact_33_2115
timestamp 1624857261
transform 1 0 21760 0 1 24485
box 0 0 1 1
use contact_33  contact_33_2116
timestamp 1624857261
transform 1 0 21760 0 1 24213
box 0 0 1 1
use contact_33  contact_33_5118
timestamp 1624857261
transform 1 0 22304 0 1 24213
box 0 0 1 1
use contact_33  contact_33_5119
timestamp 1624857261
transform 1 0 22304 0 1 24485
box 0 0 1 1
use contact_33  contact_33_1925
timestamp 1624857261
transform 1 0 21896 0 1 24893
box 0 0 1 1
use contact_33  contact_33_1926
timestamp 1624857261
transform 1 0 21896 0 1 24621
box 0 0 1 1
use contact_33  contact_33_5116
timestamp 1624857261
transform 1 0 22168 0 1 24893
box 0 0 1 1
use contact_33  contact_33_5117
timestamp 1624857261
transform 1 0 22168 0 1 24621
box 0 0 1 1
use contact_33  contact_33_1921
timestamp 1624857261
transform 1 0 21760 0 1 25029
box 0 0 1 1
use contact_33  contact_33_1922
timestamp 1624857261
transform 1 0 21760 0 1 25301
box 0 0 1 1
use contact_33  contact_33_2207
timestamp 1624857261
transform 1 0 21896 0 1 25437
box 0 0 1 1
use contact_33  contact_33_5008
timestamp 1624857261
transform 1 0 22168 0 1 25029
box 0 0 1 1
use contact_33  contact_33_5009
timestamp 1624857261
transform 1 0 22168 0 1 25301
box 0 0 1 1
use contact_33  contact_33_4914
timestamp 1624857261
transform 1 0 22440 0 1 25437
box 0 0 1 1
use contact_33  contact_33_2208
timestamp 1624857261
transform 1 0 21896 0 1 25709
box 0 0 1 1
use contact_33  contact_33_2210
timestamp 1624857261
transform 1 0 21896 0 1 25845
box 0 0 1 1
use contact_33  contact_33_4908
timestamp 1624857261
transform 1 0 22576 0 1 25845
box 0 0 1 1
use contact_33  contact_33_4915
timestamp 1624857261
transform 1 0 22440 0 1 25709
box 0 0 1 1
use contact_33  contact_33_1928
timestamp 1624857261
transform 1 0 21760 0 1 26253
box 0 0 1 1
use contact_33  contact_33_2209
timestamp 1624857261
transform 1 0 21896 0 1 26117
box 0 0 1 1
use contact_33  contact_33_4909
timestamp 1624857261
transform 1 0 22440 0 1 25981
box 0 0 1 1
use contact_33  contact_33_1927
timestamp 1624857261
transform 1 0 21760 0 1 26525
box 0 0 1 1
use contact_33  contact_33_2077
timestamp 1624857261
transform 1 0 21896 0 1 26661
box 0 0 1 1
use contact_33  contact_33_2078
timestamp 1624857261
transform 1 0 21896 0 1 26933
box 0 0 1 1
use contact_33  contact_33_5195
timestamp 1624857261
transform 1 0 22304 0 1 26933
box 0 0 1 1
use contact_33  contact_33_5194
timestamp 1624857261
transform 1 0 22304 0 1 27205
box 0 0 1 1
use contact_33  contact_33_5126
timestamp 1624857261
transform 1 0 22304 0 1 27749
box 0 0 1 1
use contact_33  contact_33_1933
timestamp 1624857261
transform 1 0 21760 0 1 28157
box 0 0 1 1
use contact_33  contact_33_5127
timestamp 1624857261
transform 1 0 22304 0 1 28021
box 0 0 1 1
use contact_33  contact_33_1934
timestamp 1624857261
transform 1 0 21760 0 1 28429
box 0 0 1 1
use contact_33  contact_33_1987
timestamp 1624857261
transform 1 0 21760 0 1 28565
box 0 0 1 1
use contact_33  contact_33_4979
timestamp 1624857261
transform 1 0 22168 0 1 28565
box 0 0 1 1
use contact_33  contact_33_4932
timestamp 1624857261
transform 1 0 22440 0 1 28565
box 0 0 1 1
use contact_33  contact_33_1988
timestamp 1624857261
transform 1 0 21760 0 1 28837
box 0 0 1 1
use contact_33  contact_33_1986
timestamp 1624857261
transform 1 0 21896 0 1 28973
box 0 0 1 1
use contact_33  contact_33_4978
timestamp 1624857261
transform 1 0 22168 0 1 28837
box 0 0 1 1
use contact_33  contact_33_4933
timestamp 1624857261
transform 1 0 22440 0 1 28837
box 0 0 1 1
use contact_33  contact_33_1913
timestamp 1624857261
transform 1 0 21760 0 1 29381
box 0 0 1 1
use contact_33  contact_33_1985
timestamp 1624857261
transform 1 0 21896 0 1 29245
box 0 0 1 1
use contact_33  contact_33_4814
timestamp 1624857261
transform 1 0 22576 0 1 29381
box 0 0 1 1
use contact_33  contact_33_1914
timestamp 1624857261
transform 1 0 21760 0 1 29653
box 0 0 1 1
use contact_33  contact_33_1916
timestamp 1624857261
transform 1 0 21760 0 1 29789
box 0 0 1 1
use contact_33  contact_33_4815
timestamp 1624857261
transform 1 0 22576 0 1 29653
box 0 0 1 1
use contact_33  contact_33_1915
timestamp 1624857261
transform 1 0 21760 0 1 30061
box 0 0 1 1
use contact_33  contact_33_2201
timestamp 1624857261
transform 1 0 21896 0 1 30197
box 0 0 1 1
use contact_33  contact_33_4911
timestamp 1624857261
transform 1 0 22440 0 1 30197
box 0 0 1 1
use contact_33  contact_33_2203
timestamp 1624857261
transform 1 0 21760 0 1 30877
box 0 0 1 1
use contact_33  contact_33_2204
timestamp 1624857261
transform 1 0 21760 0 1 30605
box 0 0 1 1
use contact_33  contact_33_2202
timestamp 1624857261
transform 1 0 21896 0 1 30469
box 0 0 1 1
use contact_33  contact_33_4749
timestamp 1624857261
transform 1 0 22576 0 1 30877
box 0 0 1 1
use contact_33  contact_33_4910
timestamp 1624857261
transform 1 0 22440 0 1 30469
box 0 0 1 1
use contact_33  contact_33_4748
timestamp 1624857261
transform 1 0 22576 0 1 31149
box 0 0 1 1
use contact_33  contact_33_2187
timestamp 1624857261
transform 1 0 21760 0 1 31421
box 0 0 1 1
use contact_33  contact_33_2188
timestamp 1624857261
transform 1 0 21760 0 1 31693
box 0 0 1 1
use contact_33  contact_33_4894
timestamp 1624857261
transform 1 0 22576 0 1 31693
box 0 0 1 1
use contact_33  contact_33_1961
timestamp 1624857261
transform 1 0 21896 0 1 32101
box 0 0 1 1
use contact_33  contact_33_4895
timestamp 1624857261
transform 1 0 22576 0 1 31965
box 0 0 1 1
use contact_33  contact_33_1962
timestamp 1624857261
transform 1 0 21896 0 1 32373
box 0 0 1 1
use contact_33  contact_33_1964
timestamp 1624857261
transform 1 0 21896 0 1 32509
box 0 0 1 1
use contact_33  contact_33_5003
timestamp 1624857261
transform 1 0 22440 0 1 32509
box 0 0 1 1
use contact_33  contact_33_5005
timestamp 1624857261
transform 1 0 22304 0 1 32509
box 0 0 1 1
use contact_33  contact_33_2169
timestamp 1624857261
transform 1 0 21760 0 1 32917
box 0 0 1 1
use contact_33  contact_33_1963
timestamp 1624857261
transform 1 0 21896 0 1 32781
box 0 0 1 1
use contact_33  contact_33_5044
timestamp 1624857261
transform 1 0 22168 0 1 32917
box 0 0 1 1
use contact_33  contact_33_4869
timestamp 1624857261
transform 1 0 22576 0 1 32917
box 0 0 1 1
use contact_33  contact_33_5002
timestamp 1624857261
transform 1 0 22440 0 1 32781
box 0 0 1 1
use contact_33  contact_33_5004
timestamp 1624857261
transform 1 0 22304 0 1 32781
box 0 0 1 1
use contact_33  contact_33_2170
timestamp 1624857261
transform 1 0 21760 0 1 33189
box 0 0 1 1
use contact_33  contact_33_2168
timestamp 1624857261
transform 1 0 21896 0 1 33325
box 0 0 1 1
use contact_33  contact_33_5045
timestamp 1624857261
transform 1 0 22168 0 1 33189
box 0 0 1 1
use contact_33  contact_33_4868
timestamp 1624857261
transform 1 0 22576 0 1 33189
box 0 0 1 1
use contact_33  contact_33_1981
timestamp 1624857261
transform 1 0 21760 0 1 33733
box 0 0 1 1
use contact_33  contact_33_2167
timestamp 1624857261
transform 1 0 21896 0 1 33597
box 0 0 1 1
use contact_33  contact_33_5190
timestamp 1624857261
transform 1 0 22168 0 1 33733
box 0 0 1 1
use contact_33  contact_33_1982
timestamp 1624857261
transform 1 0 21760 0 1 34005
box 0 0 1 1
use contact_33  contact_33_2275
timestamp 1624857261
transform 1 0 21896 0 1 34141
box 0 0 1 1
use contact_33  contact_33_5191
timestamp 1624857261
transform 1 0 22168 0 1 34005
box 0 0 1 1
use contact_33  contact_33_5046
timestamp 1624857261
transform 1 0 22440 0 1 34141
box 0 0 1 1
use contact_33  contact_33_2274
timestamp 1624857261
transform 1 0 21896 0 1 34549
box 0 0 1 1
use contact_33  contact_33_2276
timestamp 1624857261
transform 1 0 21896 0 1 34413
box 0 0 1 1
use contact_33  contact_33_5047
timestamp 1624857261
transform 1 0 22440 0 1 34413
box 0 0 1 1
use contact_33  contact_33_1980
timestamp 1624857261
transform 1 0 21760 0 1 34957
box 0 0 1 1
use contact_33  contact_33_2273
timestamp 1624857261
transform 1 0 21896 0 1 34821
box 0 0 1 1
use contact_33  contact_33_4848
timestamp 1624857261
transform 1 0 22576 0 1 34821
box 0 0 1 1
use contact_33  contact_33_1979
timestamp 1624857261
transform 1 0 21760 0 1 35229
box 0 0 1 1
use contact_33  contact_33_2117
timestamp 1624857261
transform 1 0 21896 0 1 35365
box 0 0 1 1
use contact_33  contact_33_4849
timestamp 1624857261
transform 1 0 22576 0 1 35229
box 0 0 1 1
use contact_33  contact_33_2118
timestamp 1624857261
transform 1 0 21896 0 1 35637
box 0 0 1 1
use contact_33  contact_33_2271
timestamp 1624857261
transform 1 0 21896 0 1 36045
box 0 0 1 1
use contact_33  contact_33_5094
timestamp 1624857261
transform 1 0 22168 0 1 36045
box 0 0 1 1
use contact_33  contact_33_4716
timestamp 1624857261
transform 1 0 22576 0 1 36045
box 0 0 1 1
use contact_33  contact_33_2272
timestamp 1624857261
transform 1 0 21896 0 1 36317
box 0 0 1 1
use contact_33  contact_33_5095
timestamp 1624857261
transform 1 0 22168 0 1 36317
box 0 0 1 1
use contact_33  contact_33_5096
timestamp 1624857261
transform 1 0 22168 0 1 36725
box 0 0 1 1
use contact_33  contact_33_5097
timestamp 1624857261
transform 1 0 22168 0 1 36453
box 0 0 1 1
use contact_33  contact_33_4717
timestamp 1624857261
transform 1 0 22576 0 1 36317
box 0 0 1 1
use contact_33  contact_33_2029
timestamp 1624857261
transform 1 0 21896 0 1 37133
box 0 0 1 1
use contact_33  contact_33_2030
timestamp 1624857261
transform 1 0 21896 0 1 36861
box 0 0 1 1
use contact_33  contact_33_4898
timestamp 1624857261
transform 1 0 23392 0 1 19589
box 0 0 1 1
use contact_33  contact_33_4478
timestamp 1624857261
transform 1 0 23528 0 1 19725
box 0 0 1 1
use contact_33  contact_33_1555
timestamp 1624857261
transform 1 0 22984 0 1 20269
box 0 0 1 1
use contact_33  contact_33_4845
timestamp 1624857261
transform 1 0 22712 0 1 20269
box 0 0 1 1
use contact_33  contact_33_4481
timestamp 1624857261
transform 1 0 23392 0 1 20269
box 0 0 1 1
use contact_33  contact_33_4479
timestamp 1624857261
transform 1 0 23528 0 1 20133
box 0 0 1 1
use contact_33  contact_33_1556
timestamp 1624857261
transform 1 0 22984 0 1 20541
box 0 0 1 1
use contact_33  contact_33_1565
timestamp 1624857261
transform 1 0 22984 0 1 20677
box 0 0 1 1
use contact_33  contact_33_4785
timestamp 1624857261
transform 1 0 22712 0 1 20677
box 0 0 1 1
use contact_33  contact_33_4844
timestamp 1624857261
transform 1 0 22712 0 1 20541
box 0 0 1 1
use contact_33  contact_33_4480
timestamp 1624857261
transform 1 0 23392 0 1 20541
box 0 0 1 1
use contact_33  contact_33_4382
timestamp 1624857261
transform 1 0 23528 0 1 20677
box 0 0 1 1
use contact_33  contact_33_1564
timestamp 1624857261
transform 1 0 22984 0 1 21085
box 0 0 1 1
use contact_33  contact_33_1566
timestamp 1624857261
transform 1 0 22984 0 1 20949
box 0 0 1 1
use contact_33  contact_33_4784
timestamp 1624857261
transform 1 0 22712 0 1 20949
box 0 0 1 1
use contact_33  contact_33_4536
timestamp 1624857261
transform 1 0 23392 0 1 21085
box 0 0 1 1
use contact_33  contact_33_4383
timestamp 1624857261
transform 1 0 23528 0 1 20949
box 0 0 1 1
use contact_33  contact_33_1563
timestamp 1624857261
transform 1 0 22984 0 1 21357
box 0 0 1 1
use contact_33  contact_33_1550
timestamp 1624857261
transform 1 0 23120 0 1 21493
box 0 0 1 1
use contact_33  contact_33_4535
timestamp 1624857261
transform 1 0 23392 0 1 21493
box 0 0 1 1
use contact_33  contact_33_4537
timestamp 1624857261
transform 1 0 23392 0 1 21357
box 0 0 1 1
use contact_33  contact_33_1549
timestamp 1624857261
transform 1 0 23120 0 1 21765
box 0 0 1 1
use contact_33  contact_33_4534
timestamp 1624857261
transform 1 0 23392 0 1 21765
box 0 0 1 1
use contact_33  contact_33_1710
timestamp 1624857261
transform 1 0 23120 0 1 22989
box 0 0 1 1
use contact_33  contact_33_4469
timestamp 1624857261
transform 1 0 23528 0 1 22989
box 0 0 1 1
use contact_33  contact_33_1875
timestamp 1624857261
transform 1 0 22984 0 1 23397
box 0 0 1 1
use contact_33  contact_33_1709
timestamp 1624857261
transform 1 0 23120 0 1 23261
box 0 0 1 1
use contact_33  contact_33_4638
timestamp 1624857261
transform 1 0 23392 0 1 23397
box 0 0 1 1
use contact_33  contact_33_4468
timestamp 1624857261
transform 1 0 23528 0 1 23261
box 0 0 1 1
use contact_33  contact_33_1876
timestamp 1624857261
transform 1 0 22984 0 1 23669
box 0 0 1 1
use contact_33  contact_33_1878
timestamp 1624857261
transform 1 0 22984 0 1 23805
box 0 0 1 1
use contact_33  contact_33_4637
timestamp 1624857261
transform 1 0 23392 0 1 23805
box 0 0 1 1
use contact_33  contact_33_4639
timestamp 1624857261
transform 1 0 23392 0 1 23669
box 0 0 1 1
use contact_33  contact_33_1877
timestamp 1624857261
transform 1 0 22984 0 1 24077
box 0 0 1 1
use contact_33  contact_33_1626
timestamp 1624857261
transform 1 0 23120 0 1 24213
box 0 0 1 1
use contact_33  contact_33_4636
timestamp 1624857261
transform 1 0 23392 0 1 24077
box 0 0 1 1
use contact_33  contact_33_4378
timestamp 1624857261
transform 1 0 23528 0 1 24213
box 0 0 1 1
use contact_33  contact_33_1596
timestamp 1624857261
transform 1 0 23120 0 1 24621
box 0 0 1 1
use contact_33  contact_33_1625
timestamp 1624857261
transform 1 0 23120 0 1 24485
box 0 0 1 1
use contact_33  contact_33_4404
timestamp 1624857261
transform 1 0 23392 0 1 24621
box 0 0 1 1
use contact_33  contact_33_4379
timestamp 1624857261
transform 1 0 23528 0 1 24485
box 0 0 1 1
use contact_33  contact_33_1811
timestamp 1624857261
transform 1 0 22984 0 1 25029
box 0 0 1 1
use contact_33  contact_33_4833
timestamp 1624857261
transform 1 0 22712 0 1 25029
box 0 0 1 1
use contact_33  contact_33_1595
timestamp 1624857261
transform 1 0 23120 0 1 24893
box 0 0 1 1
use contact_33  contact_33_4405
timestamp 1624857261
transform 1 0 23392 0 1 24893
box 0 0 1 1
use contact_33  contact_33_4520
timestamp 1624857261
transform 1 0 23528 0 1 25029
box 0 0 1 1
use contact_33  contact_33_1812
timestamp 1624857261
transform 1 0 22984 0 1 25301
box 0 0 1 1
use contact_33  contact_33_4832
timestamp 1624857261
transform 1 0 22712 0 1 25301
box 0 0 1 1
use contact_33  contact_33_1810
timestamp 1624857261
transform 1 0 23120 0 1 25437
box 0 0 1 1
use contact_33  contact_33_4521
timestamp 1624857261
transform 1 0 23528 0 1 25301
box 0 0 1 1
use contact_33  contact_33_4523
timestamp 1624857261
transform 1 0 23528 0 1 25437
box 0 0 1 1
use contact_33  contact_33_1539
timestamp 1624857261
transform 1 0 22984 0 1 25845
box 0 0 1 1
use contact_33  contact_33_1809
timestamp 1624857261
transform 1 0 23120 0 1 25709
box 0 0 1 1
use contact_33  contact_33_4447
timestamp 1624857261
transform 1 0 23392 0 1 25845
box 0 0 1 1
use contact_33  contact_33_4522
timestamp 1624857261
transform 1 0 23528 0 1 25709
box 0 0 1 1
use contact_33  contact_33_1540
timestamp 1624857261
transform 1 0 22984 0 1 26117
box 0 0 1 1
use contact_33  contact_33_4729
timestamp 1624857261
transform 1 0 22712 0 1 26253
box 0 0 1 1
use contact_33  contact_33_4446
timestamp 1624857261
transform 1 0 23392 0 1 26117
box 0 0 1 1
use contact_33  contact_33_4728
timestamp 1624857261
transform 1 0 22712 0 1 26525
box 0 0 1 1
use contact_33  contact_33_1634
timestamp 1624857261
transform 1 0 23120 0 1 27341
box 0 0 1 1
use contact_33  contact_33_4433
timestamp 1624857261
transform 1 0 23528 0 1 27341
box 0 0 1 1
use contact_33  contact_33_1843
timestamp 1624857261
transform 1 0 22984 0 1 27749
box 0 0 1 1
use contact_33  contact_33_4840
timestamp 1624857261
transform 1 0 22712 0 1 27749
box 0 0 1 1
use contact_33  contact_33_1633
timestamp 1624857261
transform 1 0 23120 0 1 27613
box 0 0 1 1
use contact_33  contact_33_4670
timestamp 1624857261
transform 1 0 23392 0 1 27749
box 0 0 1 1
use contact_33  contact_33_4432
timestamp 1624857261
transform 1 0 23528 0 1 27613
box 0 0 1 1
use contact_33  contact_33_1844
timestamp 1624857261
transform 1 0 22984 0 1 28021
box 0 0 1 1
use contact_33  contact_33_1846
timestamp 1624857261
transform 1 0 22984 0 1 28157
box 0 0 1 1
use contact_33  contact_33_4841
timestamp 1624857261
transform 1 0 22712 0 1 28021
box 0 0 1 1
use contact_33  contact_33_4671
timestamp 1624857261
transform 1 0 23392 0 1 28021
box 0 0 1 1
use contact_33  contact_33_4673
timestamp 1624857261
transform 1 0 23392 0 1 28157
box 0 0 1 1
use contact_33  contact_33_1733
timestamp 1624857261
transform 1 0 22984 0 1 28565
box 0 0 1 1
use contact_33  contact_33_1845
timestamp 1624857261
transform 1 0 22984 0 1 28429
box 0 0 1 1
use contact_33  contact_33_4672
timestamp 1624857261
transform 1 0 23392 0 1 28429
box 0 0 1 1
use contact_33  contact_33_4502
timestamp 1624857261
transform 1 0 23528 0 1 28565
box 0 0 1 1
use contact_33  contact_33_1734
timestamp 1624857261
transform 1 0 22984 0 1 28837
box 0 0 1 1
use contact_33  contact_33_1777
timestamp 1624857261
transform 1 0 22984 0 1 28973
box 0 0 1 1
use contact_33  contact_33_4889
timestamp 1624857261
transform 1 0 22712 0 1 28973
box 0 0 1 1
use contact_33  contact_33_4505
timestamp 1624857261
transform 1 0 23392 0 1 28973
box 0 0 1 1
use contact_33  contact_33_4503
timestamp 1624857261
transform 1 0 23528 0 1 28837
box 0 0 1 1
use contact_33  contact_33_1776
timestamp 1624857261
transform 1 0 22984 0 1 29381
box 0 0 1 1
use contact_33  contact_33_1778
timestamp 1624857261
transform 1 0 22984 0 1 29245
box 0 0 1 1
use contact_33  contact_33_4888
timestamp 1624857261
transform 1 0 22712 0 1 29245
box 0 0 1 1
use contact_33  contact_33_4399
timestamp 1624857261
transform 1 0 23392 0 1 29381
box 0 0 1 1
use contact_33  contact_33_4504
timestamp 1624857261
transform 1 0 23392 0 1 29245
box 0 0 1 1
use contact_33  contact_33_1775
timestamp 1624857261
transform 1 0 22984 0 1 29653
box 0 0 1 1
use contact_33  contact_33_1599
timestamp 1624857261
transform 1 0 23120 0 1 29789
box 0 0 1 1
use contact_33  contact_33_4398
timestamp 1624857261
transform 1 0 23392 0 1 29653
box 0 0 1 1
use contact_33  contact_33_4430
timestamp 1624857261
transform 1 0 23392 0 1 29789
box 0 0 1 1
use contact_33  contact_33_4745
timestamp 1624857261
transform 1 0 22712 0 1 30197
box 0 0 1 1
use contact_33  contact_33_1600
timestamp 1624857261
transform 1 0 23120 0 1 30061
box 0 0 1 1
use contact_33  contact_33_4431
timestamp 1624857261
transform 1 0 23392 0 1 30061
box 0 0 1 1
use contact_33  contact_33_4744
timestamp 1624857261
transform 1 0 22712 0 1 30469
box 0 0 1 1
use contact_33  contact_33_1851
timestamp 1624857261
transform 1 0 22984 0 1 31285
box 0 0 1 1
use contact_33  contact_33_4572
timestamp 1624857261
transform 1 0 23392 0 1 31285
box 0 0 1 1
use contact_33  contact_33_1852
timestamp 1624857261
transform 1 0 22984 0 1 31557
box 0 0 1 1
use contact_33  contact_33_1850
timestamp 1624857261
transform 1 0 23120 0 1 31693
box 0 0 1 1
use contact_33  contact_33_4573
timestamp 1624857261
transform 1 0 23392 0 1 31557
box 0 0 1 1
use contact_33  contact_33_4571
timestamp 1624857261
transform 1 0 23528 0 1 31693
box 0 0 1 1
use contact_33  contact_33_1767
timestamp 1624857261
transform 1 0 22984 0 1 32101
box 0 0 1 1
use contact_33  contact_33_1849
timestamp 1624857261
transform 1 0 23120 0 1 31965
box 0 0 1 1
use contact_33  contact_33_4330
timestamp 1624857261
transform 1 0 23392 0 1 32101
box 0 0 1 1
use contact_33  contact_33_4570
timestamp 1624857261
transform 1 0 23528 0 1 31965
box 0 0 1 1
use contact_33  contact_33_1766
timestamp 1624857261
transform 1 0 22984 0 1 32509
box 0 0 1 1
use contact_33  contact_33_1768
timestamp 1624857261
transform 1 0 22984 0 1 32373
box 0 0 1 1
use contact_33  contact_33_4331
timestamp 1624857261
transform 1 0 23392 0 1 32373
box 0 0 1 1
use contact_33  contact_33_4524
timestamp 1624857261
transform 1 0 23528 0 1 32509
box 0 0 1 1
use contact_33  contact_33_1747
timestamp 1624857261
transform 1 0 22984 0 1 32917
box 0 0 1 1
use contact_33  contact_33_1765
timestamp 1624857261
transform 1 0 22984 0 1 32781
box 0 0 1 1
use contact_33  contact_33_4525
timestamp 1624857261
transform 1 0 23528 0 1 32781
box 0 0 1 1
use contact_33  contact_33_4527
timestamp 1624857261
transform 1 0 23528 0 1 32917
box 0 0 1 1
use contact_33  contact_33_1748
timestamp 1624857261
transform 1 0 22984 0 1 33189
box 0 0 1 1
use contact_33  contact_33_1750
timestamp 1624857261
transform 1 0 23120 0 1 33325
box 0 0 1 1
use contact_33  contact_33_4373
timestamp 1624857261
transform 1 0 23392 0 1 33325
box 0 0 1 1
use contact_33  contact_33_4526
timestamp 1624857261
transform 1 0 23528 0 1 33189
box 0 0 1 1
use contact_33  contact_33_1724
timestamp 1624857261
transform 1 0 22984 0 1 33733
box 0 0 1 1
use contact_33  contact_33_4769
timestamp 1624857261
transform 1 0 22712 0 1 33733
box 0 0 1 1
use contact_33  contact_33_1749
timestamp 1624857261
transform 1 0 23120 0 1 33597
box 0 0 1 1
use contact_33  contact_33_4372
timestamp 1624857261
transform 1 0 23392 0 1 33597
box 0 0 1 1
use contact_33  contact_33_4416
timestamp 1624857261
transform 1 0 23528 0 1 33733
box 0 0 1 1
use contact_33  contact_33_1723
timestamp 1624857261
transform 1 0 22984 0 1 34005
box 0 0 1 1
use contact_33  contact_33_4768
timestamp 1624857261
transform 1 0 22712 0 1 34005
box 0 0 1 1
use contact_33  contact_33_1651
timestamp 1624857261
transform 1 0 23120 0 1 34141
box 0 0 1 1
use contact_33  contact_33_4424
timestamp 1624857261
transform 1 0 23392 0 1 34141
box 0 0 1 1
use contact_33  contact_33_4417
timestamp 1624857261
transform 1 0 23528 0 1 34005
box 0 0 1 1
use contact_33  contact_33_1652
timestamp 1624857261
transform 1 0 23120 0 1 34413
box 0 0 1 1
use contact_33  contact_33_4425
timestamp 1624857261
transform 1 0 23392 0 1 34413
box 0 0 1 1
use contact_33  contact_33_4733
timestamp 1624857261
transform 1 0 22712 0 1 35637
box 0 0 1 1
use contact_33  contact_33_1758
timestamp 1624857261
transform 1 0 23120 0 1 35637
box 0 0 1 1
use contact_33  contact_33_4695
timestamp 1624857261
transform 1 0 23392 0 1 35637
box 0 0 1 1
use contact_33  contact_33_1621
timestamp 1624857261
transform 1 0 22984 0 1 36045
box 0 0 1 1
use contact_33  contact_33_4732
timestamp 1624857261
transform 1 0 22712 0 1 35909
box 0 0 1 1
use contact_33  contact_33_1757
timestamp 1624857261
transform 1 0 23120 0 1 35909
box 0 0 1 1
use contact_33  contact_33_4694
timestamp 1624857261
transform 1 0 23392 0 1 35909
box 0 0 1 1
use contact_33  contact_33_4353
timestamp 1624857261
transform 1 0 23528 0 1 36045
box 0 0 1 1
use contact_33  contact_33_1622
timestamp 1624857261
transform 1 0 22984 0 1 36317
box 0 0 1 1
use contact_33  contact_33_1631
timestamp 1624857261
transform 1 0 22984 0 1 36453
box 0 0 1 1
use contact_33  contact_33_4722
timestamp 1624857261
transform 1 0 22712 0 1 36453
box 0 0 1 1
use contact_33  contact_33_4338
timestamp 1624857261
transform 1 0 23392 0 1 36453
box 0 0 1 1
use contact_33  contact_33_4352
timestamp 1624857261
transform 1 0 23528 0 1 36317
box 0 0 1 1
use contact_33  contact_33_1630
timestamp 1624857261
transform 1 0 22984 0 1 36861
box 0 0 1 1
use contact_33  contact_33_1632
timestamp 1624857261
transform 1 0 22984 0 1 36725
box 0 0 1 1
use contact_33  contact_33_4723
timestamp 1624857261
transform 1 0 22712 0 1 36725
box 0 0 1 1
use contact_33  contact_33_4337
timestamp 1624857261
transform 1 0 23392 0 1 36861
box 0 0 1 1
use contact_33  contact_33_4339
timestamp 1624857261
transform 1 0 23392 0 1 36725
box 0 0 1 1
use contact_33  contact_33_1629
timestamp 1624857261
transform 1 0 22984 0 1 37133
box 0 0 1 1
use contact_33  contact_33_4336
timestamp 1624857261
transform 1 0 23392 0 1 37133
box 0 0 1 1
use contact_33  contact_33_4477
timestamp 1624857261
transform 1 0 24208 0 1 20133
box 0 0 1 1
use contact_33  contact_33_4476
timestamp 1624857261
transform 1 0 24208 0 1 19725
box 0 0 1 1
use contact_33  contact_33_4318
timestamp 1624857261
transform 1 0 27880 0 1 19317
box 0 0 1 1
use contact_33  contact_33_1522
timestamp 1624857261
transform 1 0 28288 0 1 19589
box 0 0 1 1
use contact_33  contact_33_4319
timestamp 1624857261
transform 1 0 27880 0 1 19589
box 0 0 1 1
use contact_33  contact_33_1521
timestamp 1624857261
transform 1 0 28288 0 1 19997
box 0 0 1 1
use contact_33  contact_33_1379
timestamp 1624857261
transform 1 0 28288 0 1 22037
box 0 0 1 1
use contact_33  contact_33_1443
timestamp 1624857261
transform 1 0 28424 0 1 22037
box 0 0 1 1
use contact_33  contact_33_1444
timestamp 1624857261
transform 1 0 28424 0 1 21765
box 0 0 1 1
use contact_33  contact_33_1359
timestamp 1624857261
transform 1 0 28560 0 1 22717
box 0 0 1 1
use contact_33  contact_33_1360
timestamp 1624857261
transform 1 0 28560 0 1 22309
box 0 0 1 1
use contact_33  contact_33_1380
timestamp 1624857261
transform 1 0 28288 0 1 22309
box 0 0 1 1
use contact_33  contact_33_1489
timestamp 1624857261
transform 1 0 28424 0 1 23941
box 0 0 1 1
use contact_33  contact_33_1490
timestamp 1624857261
transform 1 0 28424 0 1 23669
box 0 0 1 1
use contact_33  contact_33_1519
timestamp 1624857261
transform 1 0 28560 0 1 25437
box 0 0 1 1
use contact_33  contact_33_1520
timestamp 1624857261
transform 1 0 28560 0 1 25845
box 0 0 1 1
use contact_33  contact_33_1399
timestamp 1624857261
transform 1 0 28288 0 1 26389
box 0 0 1 1
use contact_33  contact_33_1400
timestamp 1624857261
transform 1 0 28288 0 1 26661
box 0 0 1 1
use contact_33  contact_33_1435
timestamp 1624857261
transform 1 0 28560 0 1 26797
box 0 0 1 1
use contact_33  contact_33_1436
timestamp 1624857261
transform 1 0 28560 0 1 27069
box 0 0 1 1
use contact_33  contact_33_1501
timestamp 1624857261
transform 1 0 28424 0 1 27341
box 0 0 1 1
use contact_33  contact_33_1502
timestamp 1624857261
transform 1 0 28424 0 1 27069
box 0 0 1 1
use contact_33  contact_33_1451
timestamp 1624857261
transform 1 0 28288 0 1 27885
box 0 0 1 1
use contact_33  contact_33_1452
timestamp 1624857261
transform 1 0 28288 0 1 27613
box 0 0 1 1
use contact_33  contact_33_1499
timestamp 1624857261
transform 1 0 28288 0 1 30197
box 0 0 1 1
use contact_33  contact_33_1500
timestamp 1624857261
transform 1 0 28288 0 1 29925
box 0 0 1 1
use contact_33  contact_33_1385
timestamp 1624857261
transform 1 0 28288 0 1 30741
box 0 0 1 1
use contact_33  contact_33_1431
timestamp 1624857261
transform 1 0 28288 0 1 30605
box 0 0 1 1
use contact_33  contact_33_1432
timestamp 1624857261
transform 1 0 28288 0 1 30333
box 0 0 1 1
use contact_33  contact_33_1386
timestamp 1624857261
transform 1 0 28288 0 1 31013
box 0 0 1 1
use contact_33  contact_33_1391
timestamp 1624857261
transform 1 0 28288 0 1 34141
box 0 0 1 1
use contact_33  contact_33_1392
timestamp 1624857261
transform 1 0 28288 0 1 33869
box 0 0 1 1
use contact_33  contact_33_1419
timestamp 1624857261
transform 1 0 28560 0 1 35773
box 0 0 1 1
use contact_33  contact_33_1420
timestamp 1624857261
transform 1 0 28560 0 1 35501
box 0 0 1 1
use contact_33  contact_33_4307
timestamp 1624857261
transform 1 0 29104 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4306
timestamp 1624857261
transform 1 0 29104 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4291
timestamp 1624857261
transform 1 0 30464 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4290
timestamp 1624857261
transform 1 0 30464 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4279
timestamp 1624857261
transform 1 0 32232 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4278
timestamp 1624857261
transform 1 0 32232 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4277
timestamp 1624857261
transform 1 0 32776 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4276
timestamp 1624857261
transform 1 0 32776 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4263
timestamp 1624857261
transform 1 0 32912 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4262
timestamp 1624857261
transform 1 0 32912 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4253
timestamp 1624857261
transform 1 0 34136 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4252
timestamp 1624857261
transform 1 0 34136 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4249
timestamp 1624857261
transform 1 0 34680 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4248
timestamp 1624857261
transform 1 0 34680 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4235
timestamp 1624857261
transform 1 0 35496 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4234
timestamp 1624857261
transform 1 0 35496 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4233
timestamp 1624857261
transform 1 0 35904 0 1 18909
box 0 0 1 1
use contact_33  contact_33_4232
timestamp 1624857261
transform 1 0 35904 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4225
timestamp 1624857261
transform 1 0 36720 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4224
timestamp 1624857261
transform 1 0 36720 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4207
timestamp 1624857261
transform 1 0 38488 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4206
timestamp 1624857261
transform 1 0 38488 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4199
timestamp 1624857261
transform 1 0 39168 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4198
timestamp 1624857261
transform 1 0 39168 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4195
timestamp 1624857261
transform 1 0 39576 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4194
timestamp 1624857261
transform 1 0 39576 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4175
timestamp 1624857261
transform 1 0 40936 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4174
timestamp 1624857261
transform 1 0 40936 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4173
timestamp 1624857261
transform 1 0 41616 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4172
timestamp 1624857261
transform 1 0 41616 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4157
timestamp 1624857261
transform 1 0 42840 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4156
timestamp 1624857261
transform 1 0 42840 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4151
timestamp 1624857261
transform 1 0 43384 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4150
timestamp 1624857261
transform 1 0 43384 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4147
timestamp 1624857261
transform 1 0 44064 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4146
timestamp 1624857261
transform 1 0 44064 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4127
timestamp 1624857261
transform 1 0 45696 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4126
timestamp 1624857261
transform 1 0 45696 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4121
timestamp 1624857261
transform 1 0 46648 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4120
timestamp 1624857261
transform 1 0 46648 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4117
timestamp 1624857261
transform 1 0 47192 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4116
timestamp 1624857261
transform 1 0 47192 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4099
timestamp 1624857261
transform 1 0 47872 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4098
timestamp 1624857261
transform 1 0 47872 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4095
timestamp 1624857261
transform 1 0 48416 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4094
timestamp 1624857261
transform 1 0 48416 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4093
timestamp 1624857261
transform 1 0 49096 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4092
timestamp 1624857261
transform 1 0 49096 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4083
timestamp 1624857261
transform 1 0 49640 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4082
timestamp 1624857261
transform 1 0 49640 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4071
timestamp 1624857261
transform 1 0 50456 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4070
timestamp 1624857261
transform 1 0 50456 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4063
timestamp 1624857261
transform 1 0 52088 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4062
timestamp 1624857261
transform 1 0 52088 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4045
timestamp 1624857261
transform 1 0 52904 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4044
timestamp 1624857261
transform 1 0 52904 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4039
timestamp 1624857261
transform 1 0 54128 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4038
timestamp 1624857261
transform 1 0 54128 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4031
timestamp 1624857261
transform 1 0 54672 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4030
timestamp 1624857261
transform 1 0 54672 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4019
timestamp 1624857261
transform 1 0 55352 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4018
timestamp 1624857261
transform 1 0 55352 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4015
timestamp 1624857261
transform 1 0 55896 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4014
timestamp 1624857261
transform 1 0 55896 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4007
timestamp 1624857261
transform 1 0 56712 0 1 19181
box 0 0 1 1
use contact_33  contact_33_4006
timestamp 1624857261
transform 1 0 56712 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4003
timestamp 1624857261
transform 1 0 57120 0 1 18773
box 0 0 1 1
use contact_33  contact_33_4002
timestamp 1624857261
transform 1 0 57120 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3997
timestamp 1624857261
transform 1 0 57664 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3996
timestamp 1624857261
transform 1 0 57664 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3983
timestamp 1624857261
transform 1 0 58344 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3982
timestamp 1624857261
transform 1 0 58344 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3981
timestamp 1624857261
transform 1 0 59160 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3980
timestamp 1624857261
transform 1 0 59160 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3973
timestamp 1624857261
transform 1 0 59704 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3972
timestamp 1624857261
transform 1 0 59704 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3963
timestamp 1624857261
transform 1 0 60520 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3962
timestamp 1624857261
transform 1 0 60520 0 1 19317
box 0 0 1 1
use contact_33  contact_33_3953
timestamp 1624857261
transform 1 0 61608 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3952
timestamp 1624857261
transform 1 0 61608 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3951
timestamp 1624857261
transform 1 0 62152 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3950
timestamp 1624857261
transform 1 0 62152 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3935
timestamp 1624857261
transform 1 0 62832 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3934
timestamp 1624857261
transform 1 0 62832 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3931
timestamp 1624857261
transform 1 0 63376 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3930
timestamp 1624857261
transform 1 0 63376 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3925
timestamp 1624857261
transform 1 0 64192 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3924
timestamp 1624857261
transform 1 0 64192 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3919
timestamp 1624857261
transform 1 0 64600 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3918
timestamp 1624857261
transform 1 0 64600 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3903
timestamp 1624857261
transform 1 0 65824 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3902
timestamp 1624857261
transform 1 0 65824 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3895
timestamp 1624857261
transform 1 0 67184 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3894
timestamp 1624857261
transform 1 0 67184 0 1 19181
box 0 0 1 1
use contact_33  contact_33_5339
timestamp 1624857261
transform 1 0 1224 0 1 37405
box 0 0 1 1
use contact_7  contact_7_134
timestamp 1624857261
transform 1 0 1793 0 1 37303
box 0 0 1 1
use contact_14  contact_14_666
timestamp 1624857261
transform 1 0 1797 0 1 37307
box 0 0 1 1
use contact_19  contact_19_666
timestamp 1624857261
transform 1 0 1794 0 1 37308
box 0 0 1 1
use contact_13  contact_13_666
timestamp 1624857261
transform 1 0 1801 0 1 37299
box 0 0 1 1
use contact_14  contact_14_664
timestamp 1624857261
transform 1 0 1797 0 1 37979
box 0 0 1 1
use contact_14  contact_14_665
timestamp 1624857261
transform 1 0 1797 0 1 37643
box 0 0 1 1
use contact_19  contact_19_664
timestamp 1624857261
transform 1 0 1794 0 1 37980
box 0 0 1 1
use contact_19  contact_19_665
timestamp 1624857261
transform 1 0 1794 0 1 37644
box 0 0 1 1
use contact_13  contact_13_664
timestamp 1624857261
transform 1 0 1801 0 1 37971
box 0 0 1 1
use contact_13  contact_13_665
timestamp 1624857261
transform 1 0 1801 0 1 37635
box 0 0 1 1
use contact_14  contact_14_663
timestamp 1624857261
transform 1 0 1797 0 1 38315
box 0 0 1 1
use contact_19  contact_19_663
timestamp 1624857261
transform 1 0 1794 0 1 38316
box 0 0 1 1
use contact_13  contact_13_663
timestamp 1624857261
transform 1 0 1801 0 1 38307
box 0 0 1 1
use contact_14  contact_14_662
timestamp 1624857261
transform 1 0 1797 0 1 38651
box 0 0 1 1
use contact_19  contact_19_662
timestamp 1624857261
transform 1 0 1794 0 1 38652
box 0 0 1 1
use contact_13  contact_13_662
timestamp 1624857261
transform 1 0 1801 0 1 38643
box 0 0 1 1
use contact_33  contact_33_2342
timestamp 1624857261
transform 1 0 14688 0 1 37813
box 0 0 1 1
use contact_33  contact_33_2340
timestamp 1624857261
transform 1 0 14824 0 1 37677
box 0 0 1 1
use contact_7  contact_7_462
timestamp 1624857261
transform 1 0 15152 0 1 38408
box 0 0 1 1
use contact_7  contact_7_367
timestamp 1624857261
transform 1 0 14207 0 1 38337
box 0 0 1 1
use contact_19  contact_19_1007
timestamp 1624857261
transform 1 0 15887 0 1 38413
box 0 0 1 1
use contact_7  contact_7_461
timestamp 1624857261
transform 1 0 15886 0 1 38408
box 0 0 1 1
use contact_33  contact_33_1942
timestamp 1624857261
transform 1 0 21760 0 1 37269
box 0 0 1 1
use contact_33  contact_33_1941
timestamp 1624857261
transform 1 0 21760 0 1 37541
box 0 0 1 1
use contact_33  contact_33_5086
timestamp 1624857261
transform 1 0 22440 0 1 37269
box 0 0 1 1
use contact_33  contact_33_5087
timestamp 1624857261
transform 1 0 22440 0 1 37541
box 0 0 1 1
use contact_33  contact_33_5152
timestamp 1624857261
transform 1 0 22168 0 1 37541
box 0 0 1 1
use contact_33  contact_33_5153
timestamp 1624857261
transform 1 0 22168 0 1 37269
box 0 0 1 1
use contact_33  contact_33_1577
timestamp 1624857261
transform 1 0 23120 0 1 37541
box 0 0 1 1
use contact_33  contact_33_1578
timestamp 1624857261
transform 1 0 23120 0 1 37269
box 0 0 1 1
use contact_33  contact_33_1989
timestamp 1624857261
transform 1 0 21896 0 1 37677
box 0 0 1 1
use contact_33  contact_33_1639
timestamp 1624857261
transform 1 0 22984 0 1 37677
box 0 0 1 1
use contact_33  contact_33_1990
timestamp 1624857261
transform 1 0 21896 0 1 37949
box 0 0 1 1
use contact_33  contact_33_1992
timestamp 1624857261
transform 1 0 21896 0 1 38085
box 0 0 1 1
use contact_33  contact_33_5150
timestamp 1624857261
transform 1 0 22168 0 1 38085
box 0 0 1 1
use contact_33  contact_33_4855
timestamp 1624857261
transform 1 0 22712 0 1 38085
box 0 0 1 1
use contact_33  contact_33_1640
timestamp 1624857261
transform 1 0 22984 0 1 37949
box 0 0 1 1
use contact_33  contact_33_1642
timestamp 1624857261
transform 1 0 22984 0 1 38085
box 0 0 1 1
use contact_33  contact_33_1991
timestamp 1624857261
transform 1 0 21896 0 1 38357
box 0 0 1 1
use contact_33  contact_33_2009
timestamp 1624857261
transform 1 0 21896 0 1 38493
box 0 0 1 1
use contact_33  contact_33_5151
timestamp 1624857261
transform 1 0 22168 0 1 38357
box 0 0 1 1
use contact_33  contact_33_4854
timestamp 1624857261
transform 1 0 22712 0 1 38357
box 0 0 1 1
use contact_33  contact_33_1641
timestamp 1624857261
transform 1 0 22984 0 1 38357
box 0 0 1 1
use contact_33  contact_33_2010
timestamp 1624857261
transform 1 0 21896 0 1 38765
box 0 0 1 1
use contact_33  contact_33_4627
timestamp 1624857261
transform 1 0 23392 0 1 38085
box 0 0 1 1
use contact_33  contact_33_4626
timestamp 1624857261
transform 1 0 23392 0 1 38357
box 0 0 1 1
use contact_33  contact_33_4625
timestamp 1624857261
transform 1 0 23392 0 1 37949
box 0 0 1 1
use contact_33  contact_33_4624
timestamp 1624857261
transform 1 0 23392 0 1 37677
box 0 0 1 1
use contact_33  contact_33_4333
timestamp 1624857261
transform 1 0 23528 0 1 37541
box 0 0 1 1
use contact_33  contact_33_4332
timestamp 1624857261
transform 1 0 23528 0 1 37269
box 0 0 1 1
use contact_33  contact_33_1511
timestamp 1624857261
transform 1 0 28288 0 1 38629
box 0 0 1 1
use contact_33  contact_33_5318
timestamp 1624857261
transform 1 0 1224 0 1 39037
box 0 0 1 1
use contact_7  contact_7_133
timestamp 1624857261
transform 1 0 1793 0 1 38983
box 0 0 1 1
use contact_14  contact_14_661
timestamp 1624857261
transform 1 0 1797 0 1 38987
box 0 0 1 1
use contact_19  contact_19_661
timestamp 1624857261
transform 1 0 1794 0 1 38988
box 0 0 1 1
use contact_13  contact_13_661
timestamp 1624857261
transform 1 0 1801 0 1 38979
box 0 0 1 1
use contact_14  contact_14_660
timestamp 1624857261
transform 1 0 1797 0 1 39323
box 0 0 1 1
use contact_19  contact_19_660
timestamp 1624857261
transform 1 0 1794 0 1 39324
box 0 0 1 1
use contact_13  contact_13_660
timestamp 1624857261
transform 1 0 1801 0 1 39315
box 0 0 1 1
use contact_14  contact_14_658
timestamp 1624857261
transform 1 0 1797 0 1 39995
box 0 0 1 1
use contact_14  contact_14_659
timestamp 1624857261
transform 1 0 1797 0 1 39659
box 0 0 1 1
use contact_19  contact_19_658
timestamp 1624857261
transform 1 0 1794 0 1 39996
box 0 0 1 1
use contact_19  contact_19_659
timestamp 1624857261
transform 1 0 1794 0 1 39660
box 0 0 1 1
use contact_13  contact_13_658
timestamp 1624857261
transform 1 0 1801 0 1 39987
box 0 0 1 1
use contact_13  contact_13_659
timestamp 1624857261
transform 1 0 1801 0 1 39651
box 0 0 1 1
use contact_33  contact_33_5257
timestamp 1624857261
transform 1 0 14552 0 1 39173
box 0 0 1 1
use contact_7  contact_7_460
timestamp 1624857261
transform 1 0 15152 0 1 39966
box 0 0 1 1
use contact_7  contact_7_366
timestamp 1624857261
transform 1 0 14207 0 1 40037
box 0 0 1 1
use contact_19  contact_19_1006
timestamp 1624857261
transform 1 0 15967 0 1 39971
box 0 0 1 1
use contact_7  contact_7_459
timestamp 1624857261
transform 1 0 15966 0 1 39966
box 0 0 1 1
use contact_33  contact_33_2134
timestamp 1624857261
transform 1 0 21760 0 1 39581
box 0 0 1 1
use contact_33  contact_33_2133
timestamp 1624857261
transform 1 0 21760 0 1 39309
box 0 0 1 1
use contact_33  contact_33_2043
timestamp 1624857261
transform 1 0 21896 0 1 38901
box 0 0 1 1
use contact_33  contact_33_2044
timestamp 1624857261
transform 1 0 21896 0 1 39173
box 0 0 1 1
use contact_33  contact_33_5186
timestamp 1624857261
transform 1 0 22440 0 1 38901
box 0 0 1 1
use contact_33  contact_33_5187
timestamp 1624857261
transform 1 0 22440 0 1 39173
box 0 0 1 1
use contact_33  contact_33_5188
timestamp 1624857261
transform 1 0 22304 0 1 38901
box 0 0 1 1
use contact_33  contact_33_5189
timestamp 1624857261
transform 1 0 22304 0 1 39173
box 0 0 1 1
use contact_33  contact_33_4721
timestamp 1624857261
transform 1 0 22576 0 1 39581
box 0 0 1 1
use contact_33  contact_33_1740
timestamp 1624857261
transform 1 0 23120 0 1 39581
box 0 0 1 1
use contact_33  contact_33_4720
timestamp 1624857261
transform 1 0 22576 0 1 39853
box 0 0 1 1
use contact_33  contact_33_1739
timestamp 1624857261
transform 1 0 23120 0 1 39853
box 0 0 1 1
use contact_33  contact_33_1879
timestamp 1624857261
transform 1 0 22984 0 1 39989
box 0 0 1 1
use contact_33  contact_33_1880
timestamp 1624857261
transform 1 0 22984 0 1 40261
box 0 0 1 1
use contact_33  contact_33_4665
timestamp 1624857261
transform 1 0 23528 0 1 39581
box 0 0 1 1
use contact_33  contact_33_4664
timestamp 1624857261
transform 1 0 23528 0 1 39853
box 0 0 1 1
use contact_33  contact_33_4539
timestamp 1624857261
transform 1 0 23392 0 1 39989
box 0 0 1 1
use contact_33  contact_33_4538
timestamp 1624857261
transform 1 0 23392 0 1 40261
box 0 0 1 1
use contact_33  contact_33_1512
timestamp 1624857261
transform 1 0 28288 0 1 38901
box 0 0 1 1
use contact_33  contact_33_1510
timestamp 1624857261
transform 1 0 28288 0 1 39037
box 0 0 1 1
use contact_33  contact_33_1509
timestamp 1624857261
transform 1 0 28288 0 1 39309
box 0 0 1 1
use contact_33  contact_33_1374
timestamp 1624857261
transform 1 0 28424 0 1 39445
box 0 0 1 1
use contact_33  contact_33_1373
timestamp 1624857261
transform 1 0 28424 0 1 39717
box 0 0 1 1
use contact_33  contact_33_5347
timestamp 1624857261
transform 1 0 1224 0 1 40669
box 0 0 1 1
use contact_7  contact_7_132
timestamp 1624857261
transform 1 0 1793 0 1 40663
box 0 0 1 1
use contact_14  contact_14_656
timestamp 1624857261
transform 1 0 1797 0 1 40667
box 0 0 1 1
use contact_14  contact_14_657
timestamp 1624857261
transform 1 0 1797 0 1 40331
box 0 0 1 1
use contact_19  contact_19_656
timestamp 1624857261
transform 1 0 1794 0 1 40668
box 0 0 1 1
use contact_19  contact_19_657
timestamp 1624857261
transform 1 0 1794 0 1 40332
box 0 0 1 1
use contact_13  contact_13_656
timestamp 1624857261
transform 1 0 1801 0 1 40659
box 0 0 1 1
use contact_13  contact_13_657
timestamp 1624857261
transform 1 0 1801 0 1 40323
box 0 0 1 1
use contact_14  contact_14_655
timestamp 1624857261
transform 1 0 1797 0 1 41003
box 0 0 1 1
use contact_19  contact_19_655
timestamp 1624857261
transform 1 0 1794 0 1 41004
box 0 0 1 1
use contact_13  contact_13_655
timestamp 1624857261
transform 1 0 1801 0 1 40995
box 0 0 1 1
use contact_14  contact_14_654
timestamp 1624857261
transform 1 0 1797 0 1 41339
box 0 0 1 1
use contact_19  contact_19_654
timestamp 1624857261
transform 1 0 1794 0 1 41340
box 0 0 1 1
use contact_13  contact_13_654
timestamp 1624857261
transform 1 0 1801 0 1 41331
box 0 0 1 1
use contact_14  contact_14_653
timestamp 1624857261
transform 1 0 1797 0 1 41675
box 0 0 1 1
use contact_19  contact_19_653
timestamp 1624857261
transform 1 0 1794 0 1 41676
box 0 0 1 1
use contact_13  contact_13_653
timestamp 1624857261
transform 1 0 1801 0 1 41667
box 0 0 1 1
use contact_33  contact_33_2341
timestamp 1624857261
transform 1 0 14688 0 1 40533
box 0 0 1 1
use contact_33  contact_33_2270
timestamp 1624857261
transform 1 0 21760 0 1 41621
box 0 0 1 1
use contact_33  contact_33_2268
timestamp 1624857261
transform 1 0 21760 0 1 41485
box 0 0 1 1
use contact_33  contact_33_2267
timestamp 1624857261
transform 1 0 21760 0 1 41213
box 0 0 1 1
use contact_33  contact_33_2016
timestamp 1624857261
transform 1 0 21760 0 1 40805
box 0 0 1 1
use contact_33  contact_33_2015
timestamp 1624857261
transform 1 0 21760 0 1 41077
box 0 0 1 1
use contact_33  contact_33_4724
timestamp 1624857261
transform 1 0 22576 0 1 40669
box 0 0 1 1
use contact_33  contact_33_4725
timestamp 1624857261
transform 1 0 22576 0 1 40397
box 0 0 1 1
use contact_33  contact_33_1881
timestamp 1624857261
transform 1 0 23120 0 1 40669
box 0 0 1 1
use contact_33  contact_33_1882
timestamp 1624857261
transform 1 0 23120 0 1 40397
box 0 0 1 1
use contact_33  contact_33_4936
timestamp 1624857261
transform 1 0 22168 0 1 41077
box 0 0 1 1
use contact_33  contact_33_4937
timestamp 1624857261
transform 1 0 22168 0 1 40805
box 0 0 1 1
use contact_33  contact_33_1761
timestamp 1624857261
transform 1 0 22984 0 1 41077
box 0 0 1 1
use contact_33  contact_33_1762
timestamp 1624857261
transform 1 0 22984 0 1 40805
box 0 0 1 1
use contact_33  contact_33_4762
timestamp 1624857261
transform 1 0 22712 0 1 40805
box 0 0 1 1
use contact_33  contact_33_4763
timestamp 1624857261
transform 1 0 22712 0 1 41077
box 0 0 1 1
use contact_33  contact_33_1729
timestamp 1624857261
transform 1 0 23120 0 1 41213
box 0 0 1 1
use contact_33  contact_33_1730
timestamp 1624857261
transform 1 0 23120 0 1 41485
box 0 0 1 1
use contact_33  contact_33_5163
timestamp 1624857261
transform 1 0 22168 0 1 41621
box 0 0 1 1
use contact_33  contact_33_5156
timestamp 1624857261
transform 1 0 22440 0 1 41621
box 0 0 1 1
use contact_33  contact_33_1732
timestamp 1624857261
transform 1 0 23120 0 1 41621
box 0 0 1 1
use contact_33  contact_33_4599
timestamp 1624857261
transform 1 0 23528 0 1 40805
box 0 0 1 1
use contact_33  contact_33_4598
timestamp 1624857261
transform 1 0 23528 0 1 41077
box 0 0 1 1
use contact_33  contact_33_4597
timestamp 1624857261
transform 1 0 23528 0 1 40669
box 0 0 1 1
use contact_33  contact_33_4596
timestamp 1624857261
transform 1 0 23528 0 1 40397
box 0 0 1 1
use contact_33  contact_33_4488
timestamp 1624857261
transform 1 0 23528 0 1 41621
box 0 0 1 1
use contact_33  contact_33_4421
timestamp 1624857261
transform 1 0 23392 0 1 41213
box 0 0 1 1
use contact_33  contact_33_4420
timestamp 1624857261
transform 1 0 23392 0 1 41485
box 0 0 1 1
use contact_14  contact_14_652
timestamp 1624857261
transform 1 0 1797 0 1 42011
box 0 0 1 1
use contact_19  contact_19_652
timestamp 1624857261
transform 1 0 1794 0 1 42012
box 0 0 1 1
use contact_13  contact_13_652
timestamp 1624857261
transform 1 0 1801 0 1 42003
box 0 0 1 1
use contact_33  contact_33_5374
timestamp 1624857261
transform 1 0 1224 0 1 42437
box 0 0 1 1
use contact_7  contact_7_131
timestamp 1624857261
transform 1 0 1793 0 1 42343
box 0 0 1 1
use contact_14  contact_14_651
timestamp 1624857261
transform 1 0 1797 0 1 42347
box 0 0 1 1
use contact_19  contact_19_651
timestamp 1624857261
transform 1 0 1794 0 1 42348
box 0 0 1 1
use contact_13  contact_13_651
timestamp 1624857261
transform 1 0 1801 0 1 42339
box 0 0 1 1
use contact_14  contact_14_650
timestamp 1624857261
transform 1 0 1797 0 1 42683
box 0 0 1 1
use contact_19  contact_19_650
timestamp 1624857261
transform 1 0 1794 0 1 42684
box 0 0 1 1
use contact_13  contact_13_650
timestamp 1624857261
transform 1 0 1801 0 1 42675
box 0 0 1 1
use contact_14  contact_14_649
timestamp 1624857261
transform 1 0 1797 0 1 43019
box 0 0 1 1
use contact_19  contact_19_649
timestamp 1624857261
transform 1 0 1794 0 1 43020
box 0 0 1 1
use contact_13  contact_13_649
timestamp 1624857261
transform 1 0 1801 0 1 43011
box 0 0 1 1
use contact_14  contact_14_648
timestamp 1624857261
transform 1 0 1797 0 1 43355
box 0 0 1 1
use contact_19  contact_19_648
timestamp 1624857261
transform 1 0 1794 0 1 43356
box 0 0 1 1
use contact_13  contact_13_648
timestamp 1624857261
transform 1 0 1801 0 1 43347
box 0 0 1 1
use contact_33  contact_33_2269
timestamp 1624857261
transform 1 0 21760 0 1 41893
box 0 0 1 1
use contact_33  contact_33_2092
timestamp 1624857261
transform 1 0 21760 0 1 42709
box 0 0 1 1
use contact_33  contact_33_2091
timestamp 1624857261
transform 1 0 21760 0 1 42437
box 0 0 1 1
use contact_33  contact_33_2090
timestamp 1624857261
transform 1 0 21760 0 1 42845
box 0 0 1 1
use contact_33  contact_33_2089
timestamp 1624857261
transform 1 0 21760 0 1 43117
box 0 0 1 1
use contact_33  contact_33_2038
timestamp 1624857261
transform 1 0 21896 0 1 42029
box 0 0 1 1
use contact_33  contact_33_5162
timestamp 1624857261
transform 1 0 22168 0 1 41893
box 0 0 1 1
use contact_33  contact_33_5157
timestamp 1624857261
transform 1 0 22440 0 1 41893
box 0 0 1 1
use contact_33  contact_33_1646
timestamp 1624857261
transform 1 0 23120 0 1 42029
box 0 0 1 1
use contact_33  contact_33_1731
timestamp 1624857261
transform 1 0 23120 0 1 41893
box 0 0 1 1
use contact_33  contact_33_2037
timestamp 1624857261
transform 1 0 21896 0 1 42301
box 0 0 1 1
use contact_33  contact_33_1527
timestamp 1624857261
transform 1 0 23120 0 1 42437
box 0 0 1 1
use contact_33  contact_33_1645
timestamp 1624857261
transform 1 0 23120 0 1 42301
box 0 0 1 1
use contact_33  contact_33_5114
timestamp 1624857261
transform 1 0 22440 0 1 42845
box 0 0 1 1
use contact_33  contact_33_5115
timestamp 1624857261
transform 1 0 22440 0 1 43117
box 0 0 1 1
use contact_33  contact_33_1528
timestamp 1624857261
transform 1 0 23120 0 1 42709
box 0 0 1 1
use contact_33  contact_33_1909
timestamp 1624857261
transform 1 0 21896 0 1 43253
box 0 0 1 1
use contact_33  contact_33_4924
timestamp 1624857261
transform 1 0 22576 0 1 43253
box 0 0 1 1
use contact_33  contact_33_4491
timestamp 1624857261
transform 1 0 23392 0 1 42029
box 0 0 1 1
use contact_33  contact_33_4490
timestamp 1624857261
transform 1 0 23392 0 1 42301
box 0 0 1 1
use contact_33  contact_33_4489
timestamp 1624857261
transform 1 0 23528 0 1 41893
box 0 0 1 1
use contact_33  contact_33_4451
timestamp 1624857261
transform 1 0 23392 0 1 42437
box 0 0 1 1
use contact_33  contact_33_4450
timestamp 1624857261
transform 1 0 23392 0 1 42709
box 0 0 1 1
use contact_33  contact_33_1368
timestamp 1624857261
transform 1 0 28288 0 1 43253
box 0 0 1 1
use contact_33  contact_33_1367
timestamp 1624857261
transform 1 0 28288 0 1 42981
box 0 0 1 1
use contact_33  contact_33_1362
timestamp 1624857261
transform 1 0 28288 0 1 42573
box 0 0 1 1
use contact_33  contact_33_1361
timestamp 1624857261
transform 1 0 28288 0 1 42845
box 0 0 1 1
use contact_14  contact_14_647
timestamp 1624857261
transform 1 0 1797 0 1 43691
box 0 0 1 1
use contact_19  contact_19_647
timestamp 1624857261
transform 1 0 1794 0 1 43692
box 0 0 1 1
use contact_13  contact_13_647
timestamp 1624857261
transform 1 0 1801 0 1 43683
box 0 0 1 1
use contact_33  contact_33_5302
timestamp 1624857261
transform 1 0 1224 0 1 44069
box 0 0 1 1
use contact_7  contact_7_130
timestamp 1624857261
transform 1 0 1793 0 1 44023
box 0 0 1 1
use contact_14  contact_14_646
timestamp 1624857261
transform 1 0 1797 0 1 44027
box 0 0 1 1
use contact_19  contact_19_646
timestamp 1624857261
transform 1 0 1794 0 1 44028
box 0 0 1 1
use contact_13  contact_13_646
timestamp 1624857261
transform 1 0 1801 0 1 44019
box 0 0 1 1
use contact_14  contact_14_645
timestamp 1624857261
transform 1 0 1797 0 1 44363
box 0 0 1 1
use contact_19  contact_19_645
timestamp 1624857261
transform 1 0 1794 0 1 44364
box 0 0 1 1
use contact_13  contact_13_645
timestamp 1624857261
transform 1 0 1801 0 1 44355
box 0 0 1 1
use contact_14  contact_14_644
timestamp 1624857261
transform 1 0 1797 0 1 44699
box 0 0 1 1
use contact_19  contact_19_644
timestamp 1624857261
transform 1 0 1794 0 1 44700
box 0 0 1 1
use contact_13  contact_13_644
timestamp 1624857261
transform 1 0 1801 0 1 44691
box 0 0 1 1
use contact_33  contact_33_2024
timestamp 1624857261
transform 1 0 21760 0 1 44749
box 0 0 1 1
use contact_33  contact_33_1910
timestamp 1624857261
transform 1 0 21896 0 1 43525
box 0 0 1 1
use contact_33  contact_33_4925
timestamp 1624857261
transform 1 0 22440 0 1 43525
box 0 0 1 1
use contact_33  contact_33_5130
timestamp 1624857261
transform 1 0 22168 0 1 43525
box 0 0 1 1
use contact_33  contact_33_4852
timestamp 1624857261
transform 1 0 22576 0 1 43525
box 0 0 1 1
use contact_33  contact_33_1638
timestamp 1624857261
transform 1 0 22984 0 1 43525
box 0 0 1 1
use contact_33  contact_33_5131
timestamp 1624857261
transform 1 0 22168 0 1 43797
box 0 0 1 1
use contact_33  contact_33_4853
timestamp 1624857261
transform 1 0 22576 0 1 43797
box 0 0 1 1
use contact_33  contact_33_1592
timestamp 1624857261
transform 1 0 22984 0 1 43933
box 0 0 1 1
use contact_33  contact_33_1637
timestamp 1624857261
transform 1 0 22984 0 1 43797
box 0 0 1 1
use contact_33  contact_33_5198
timestamp 1624857261
transform 1 0 22304 0 1 44341
box 0 0 1 1
use contact_33  contact_33_4800
timestamp 1624857261
transform 1 0 22712 0 1 44341
box 0 0 1 1
use contact_33  contact_33_1542
timestamp 1624857261
transform 1 0 23120 0 1 44341
box 0 0 1 1
use contact_33  contact_33_1591
timestamp 1624857261
transform 1 0 22984 0 1 44205
box 0 0 1 1
use contact_33  contact_33_5197
timestamp 1624857261
transform 1 0 22168 0 1 44749
box 0 0 1 1
use contact_33  contact_33_5199
timestamp 1624857261
transform 1 0 22304 0 1 44613
box 0 0 1 1
use contact_33  contact_33_4801
timestamp 1624857261
transform 1 0 22712 0 1 44613
box 0 0 1 1
use contact_33  contact_33_4884
timestamp 1624857261
transform 1 0 22576 0 1 44749
box 0 0 1 1
use contact_33  contact_33_1541
timestamp 1624857261
transform 1 0 23120 0 1 44613
box 0 0 1 1
use contact_33  contact_33_1547
timestamp 1624857261
transform 1 0 22984 0 1 44749
box 0 0 1 1
use contact_33  contact_33_4377
timestamp 1624857261
transform 1 0 23392 0 1 44341
box 0 0 1 1
use contact_33  contact_33_4376
timestamp 1624857261
transform 1 0 23392 0 1 44613
box 0 0 1 1
use contact_33  contact_33_4375
timestamp 1624857261
transform 1 0 23392 0 1 44205
box 0 0 1 1
use contact_33  contact_33_4374
timestamp 1624857261
transform 1 0 23392 0 1 43933
box 0 0 1 1
use contact_33  contact_33_4367
timestamp 1624857261
transform 1 0 23528 0 1 44749
box 0 0 1 1
use contact_33  contact_33_4335
timestamp 1624857261
transform 1 0 23392 0 1 43525
box 0 0 1 1
use contact_33  contact_33_4334
timestamp 1624857261
transform 1 0 23392 0 1 43797
box 0 0 1 1
use contact_14  contact_14_643
timestamp 1624857261
transform 1 0 1797 0 1 45035
box 0 0 1 1
use contact_19  contact_19_643
timestamp 1624857261
transform 1 0 1794 0 1 45036
box 0 0 1 1
use contact_13  contact_13_643
timestamp 1624857261
transform 1 0 1801 0 1 45027
box 0 0 1 1
use contact_33  contact_33_5364
timestamp 1624857261
transform 1 0 1224 0 1 45565
box 0 0 1 1
use contact_14  contact_14_642
timestamp 1624857261
transform 1 0 1797 0 1 45371
box 0 0 1 1
use contact_19  contact_19_642
timestamp 1624857261
transform 1 0 1794 0 1 45372
box 0 0 1 1
use contact_13  contact_13_642
timestamp 1624857261
transform 1 0 1801 0 1 45363
box 0 0 1 1
use contact_7  contact_7_129
timestamp 1624857261
transform 1 0 1793 0 1 45703
box 0 0 1 1
use contact_14  contact_14_640
timestamp 1624857261
transform 1 0 1797 0 1 46043
box 0 0 1 1
use contact_14  contact_14_641
timestamp 1624857261
transform 1 0 1797 0 1 45707
box 0 0 1 1
use contact_19  contact_19_640
timestamp 1624857261
transform 1 0 1794 0 1 46044
box 0 0 1 1
use contact_19  contact_19_641
timestamp 1624857261
transform 1 0 1794 0 1 45708
box 0 0 1 1
use contact_13  contact_13_640
timestamp 1624857261
transform 1 0 1801 0 1 46035
box 0 0 1 1
use contact_13  contact_13_641
timestamp 1624857261
transform 1 0 1801 0 1 45699
box 0 0 1 1
use contact_14  contact_14_639
timestamp 1624857261
transform 1 0 1797 0 1 46379
box 0 0 1 1
use contact_19  contact_19_639
timestamp 1624857261
transform 1 0 1794 0 1 46380
box 0 0 1 1
use contact_13  contact_13_639
timestamp 1624857261
transform 1 0 1801 0 1 46371
box 0 0 1 1
use contact_33  contact_33_2023
timestamp 1624857261
transform 1 0 21760 0 1 45021
box 0 0 1 1
use contact_33  contact_33_2012
timestamp 1624857261
transform 1 0 21760 0 1 45973
box 0 0 1 1
use contact_33  contact_33_2011
timestamp 1624857261
transform 1 0 21760 0 1 46245
box 0 0 1 1
use contact_33  contact_33_2141
timestamp 1624857261
transform 1 0 21896 0 1 45157
box 0 0 1 1
use contact_33  contact_33_5196
timestamp 1624857261
transform 1 0 22168 0 1 45021
box 0 0 1 1
use contact_33  contact_33_4885
timestamp 1624857261
transform 1 0 22576 0 1 45021
box 0 0 1 1
use contact_33  contact_33_4887
timestamp 1624857261
transform 1 0 22576 0 1 45157
box 0 0 1 1
use contact_33  contact_33_1548
timestamp 1624857261
transform 1 0 22984 0 1 45021
box 0 0 1 1
use contact_33  contact_33_1585
timestamp 1624857261
transform 1 0 22984 0 1 45157
box 0 0 1 1
use contact_33  contact_33_2142
timestamp 1624857261
transform 1 0 21896 0 1 45429
box 0 0 1 1
use contact_33  contact_33_2144
timestamp 1624857261
transform 1 0 21896 0 1 45565
box 0 0 1 1
use contact_33  contact_33_4919
timestamp 1624857261
transform 1 0 22304 0 1 45565
box 0 0 1 1
use contact_33  contact_33_4886
timestamp 1624857261
transform 1 0 22576 0 1 45429
box 0 0 1 1
use contact_33  contact_33_1586
timestamp 1624857261
transform 1 0 22984 0 1 45429
box 0 0 1 1
use contact_33  contact_33_1609
timestamp 1624857261
transform 1 0 23120 0 1 45565
box 0 0 1 1
use contact_33  contact_33_2143
timestamp 1624857261
transform 1 0 21896 0 1 45837
box 0 0 1 1
use contact_33  contact_33_4918
timestamp 1624857261
transform 1 0 22304 0 1 45837
box 0 0 1 1
use contact_33  contact_33_1610
timestamp 1624857261
transform 1 0 23120 0 1 45837
box 0 0 1 1
use contact_33  contact_33_5026
timestamp 1624857261
transform 1 0 22168 0 1 45973
box 0 0 1 1
use contact_33  contact_33_5027
timestamp 1624857261
transform 1 0 22168 0 1 46245
box 0 0 1 1
use contact_33  contact_33_1607
timestamp 1624857261
transform 1 0 23120 0 1 46245
box 0 0 1 1
use contact_33  contact_33_1608
timestamp 1624857261
transform 1 0 23120 0 1 45973
box 0 0 1 1
use contact_33  contact_33_1965
timestamp 1624857261
transform 1 0 21896 0 1 46381
box 0 0 1 1
use contact_33  contact_33_1601
timestamp 1624857261
transform 1 0 22984 0 1 46381
box 0 0 1 1
use contact_33  contact_33_4591
timestamp 1624857261
transform 1 0 23392 0 1 46381
box 0 0 1 1
use contact_33  contact_33_4589
timestamp 1624857261
transform 1 0 23528 0 1 46245
box 0 0 1 1
use contact_33  contact_33_4588
timestamp 1624857261
transform 1 0 23528 0 1 45973
box 0 0 1 1
use contact_33  contact_33_4413
timestamp 1624857261
transform 1 0 23392 0 1 45429
box 0 0 1 1
use contact_33  contact_33_4412
timestamp 1624857261
transform 1 0 23392 0 1 45157
box 0 0 1 1
use contact_33  contact_33_4411
timestamp 1624857261
transform 1 0 23392 0 1 45565
box 0 0 1 1
use contact_33  contact_33_4410
timestamp 1624857261
transform 1 0 23392 0 1 45837
box 0 0 1 1
use contact_33  contact_33_4366
timestamp 1624857261
transform 1 0 23528 0 1 45021
box 0 0 1 1
use contact_33  contact_33_1478
timestamp 1624857261
transform 1 0 28288 0 1 45973
box 0 0 1 1
use contact_33  contact_33_1477
timestamp 1624857261
transform 1 0 28288 0 1 46381
box 0 0 1 1
use contact_14  contact_14_638
timestamp 1624857261
transform 1 0 1797 0 1 46715
box 0 0 1 1
use contact_19  contact_19_638
timestamp 1624857261
transform 1 0 1794 0 1 46716
box 0 0 1 1
use contact_13  contact_13_638
timestamp 1624857261
transform 1 0 1801 0 1 46707
box 0 0 1 1
use contact_14  contact_14_637
timestamp 1624857261
transform 1 0 1797 0 1 47051
box 0 0 1 1
use contact_19  contact_19_637
timestamp 1624857261
transform 1 0 1794 0 1 47052
box 0 0 1 1
use contact_13  contact_13_637
timestamp 1624857261
transform 1 0 1801 0 1 47043
box 0 0 1 1
use contact_33  contact_33_5363
timestamp 1624857261
transform 1 0 1224 0 1 47333
box 0 0 1 1
use contact_7  contact_7_128
timestamp 1624857261
transform 1 0 1793 0 1 47383
box 0 0 1 1
use contact_14  contact_14_636
timestamp 1624857261
transform 1 0 1797 0 1 47387
box 0 0 1 1
use contact_19  contact_19_636
timestamp 1624857261
transform 1 0 1794 0 1 47388
box 0 0 1 1
use contact_13  contact_13_636
timestamp 1624857261
transform 1 0 1801 0 1 47379
box 0 0 1 1
use contact_14  contact_14_635
timestamp 1624857261
transform 1 0 1797 0 1 47723
box 0 0 1 1
use contact_19  contact_19_635
timestamp 1624857261
transform 1 0 1794 0 1 47724
box 0 0 1 1
use contact_13  contact_13_635
timestamp 1624857261
transform 1 0 1801 0 1 47715
box 0 0 1 1
use contact_33  contact_33_2266
timestamp 1624857261
transform 1 0 21760 0 1 47061
box 0 0 1 1
use contact_33  contact_33_2265
timestamp 1624857261
transform 1 0 21760 0 1 46789
box 0 0 1 1
use contact_33  contact_33_2264
timestamp 1624857261
transform 1 0 21760 0 1 47197
box 0 0 1 1
use contact_33  contact_33_2263
timestamp 1624857261
transform 1 0 21760 0 1 47469
box 0 0 1 1
use contact_33  contact_33_5143
timestamp 1624857261
transform 1 0 22440 0 1 47061
box 0 0 1 1
use contact_33  contact_33_5142
timestamp 1624857261
transform 1 0 22440 0 1 46789
box 0 0 1 1
use contact_33  contact_33_4831
timestamp 1624857261
transform 1 0 22712 0 1 47469
box 0 0 1 1
use contact_33  contact_33_4830
timestamp 1624857261
transform 1 0 22712 0 1 47741
box 0 0 1 1
use contact_33  contact_33_1966
timestamp 1624857261
transform 1 0 21896 0 1 46653
box 0 0 1 1
use contact_33  contact_33_1716
timestamp 1624857261
transform 1 0 22984 0 1 47877
box 0 0 1 1
use contact_33  contact_33_1602
timestamp 1624857261
transform 1 0 22984 0 1 46653
box 0 0 1 1
use contact_33  contact_33_4590
timestamp 1624857261
transform 1 0 23392 0 1 46653
box 0 0 1 1
use contact_33  contact_33_4553
timestamp 1624857261
transform 1 0 23392 0 1 47877
box 0 0 1 1
use contact_33  contact_33_1424
timestamp 1624857261
transform 1 0 28288 0 1 46925
box 0 0 1 1
use contact_33  contact_33_1423
timestamp 1624857261
transform 1 0 28288 0 1 47197
box 0 0 1 1
use contact_14  contact_14_634
timestamp 1624857261
transform 1 0 1797 0 1 48059
box 0 0 1 1
use contact_19  contact_19_634
timestamp 1624857261
transform 1 0 1794 0 1 48060
box 0 0 1 1
use contact_13  contact_13_634
timestamp 1624857261
transform 1 0 1801 0 1 48051
box 0 0 1 1
use contact_14  contact_14_632
timestamp 1624857261
transform 1 0 1797 0 1 48731
box 0 0 1 1
use contact_14  contact_14_633
timestamp 1624857261
transform 1 0 1797 0 1 48395
box 0 0 1 1
use contact_19  contact_19_632
timestamp 1624857261
transform 1 0 1794 0 1 48732
box 0 0 1 1
use contact_19  contact_19_633
timestamp 1624857261
transform 1 0 1794 0 1 48396
box 0 0 1 1
use contact_13  contact_13_632
timestamp 1624857261
transform 1 0 1801 0 1 48723
box 0 0 1 1
use contact_13  contact_13_633
timestamp 1624857261
transform 1 0 1801 0 1 48387
box 0 0 1 1
use contact_33  contact_33_5380
timestamp 1624857261
transform 1 0 1224 0 1 49101
box 0 0 1 1
use contact_7  contact_7_127
timestamp 1624857261
transform 1 0 1793 0 1 49063
box 0 0 1 1
use contact_14  contact_14_631
timestamp 1624857261
transform 1 0 1797 0 1 49067
box 0 0 1 1
use contact_19  contact_19_631
timestamp 1624857261
transform 1 0 1794 0 1 49068
box 0 0 1 1
use contact_13  contact_13_631
timestamp 1624857261
transform 1 0 1801 0 1 49059
box 0 0 1 1
use contact_14  contact_14_630
timestamp 1624857261
transform 1 0 1797 0 1 49403
box 0 0 1 1
use contact_19  contact_19_630
timestamp 1624857261
transform 1 0 1794 0 1 49404
box 0 0 1 1
use contact_13  contact_13_630
timestamp 1624857261
transform 1 0 1801 0 1 49395
box 0 0 1 1
use contact_33  contact_33_2166
timestamp 1624857261
transform 1 0 21760 0 1 48285
box 0 0 1 1
use contact_33  contact_33_2165
timestamp 1624857261
transform 1 0 21760 0 1 48013
box 0 0 1 1
use contact_33  contact_33_1912
timestamp 1624857261
transform 1 0 21760 0 1 49101
box 0 0 1 1
use contact_33  contact_33_1911
timestamp 1624857261
transform 1 0 21760 0 1 49373
box 0 0 1 1
use contact_33  contact_33_4954
timestamp 1624857261
transform 1 0 22304 0 1 48285
box 0 0 1 1
use contact_33  contact_33_1571
timestamp 1624857261
transform 1 0 23120 0 1 48285
box 0 0 1 1
use contact_33  contact_33_1715
timestamp 1624857261
transform 1 0 22984 0 1 48149
box 0 0 1 1
use contact_33  contact_33_1946
timestamp 1624857261
transform 1 0 21896 0 1 48693
box 0 0 1 1
use contact_33  contact_33_4955
timestamp 1624857261
transform 1 0 22304 0 1 48557
box 0 0 1 1
use contact_33  contact_33_4867
timestamp 1624857261
transform 1 0 22712 0 1 48693
box 0 0 1 1
use contact_33  contact_33_1570
timestamp 1624857261
transform 1 0 23120 0 1 48693
box 0 0 1 1
use contact_33  contact_33_1572
timestamp 1624857261
transform 1 0 23120 0 1 48557
box 0 0 1 1
use contact_33  contact_33_1945
timestamp 1624857261
transform 1 0 21896 0 1 48965
box 0 0 1 1
use contact_33  contact_33_4866
timestamp 1624857261
transform 1 0 22712 0 1 48965
box 0 0 1 1
use contact_33  contact_33_1569
timestamp 1624857261
transform 1 0 23120 0 1 48965
box 0 0 1 1
use contact_33  contact_33_4742
timestamp 1624857261
transform 1 0 22576 0 1 49373
box 0 0 1 1
use contact_33  contact_33_4743
timestamp 1624857261
transform 1 0 22576 0 1 49101
box 0 0 1 1
use contact_33  contact_33_1681
timestamp 1624857261
transform 1 0 22984 0 1 49101
box 0 0 1 1
use contact_33  contact_33_1682
timestamp 1624857261
transform 1 0 22984 0 1 49373
box 0 0 1 1
use contact_33  contact_33_2235
timestamp 1624857261
transform 1 0 21896 0 1 49509
box 0 0 1 1
use contact_33  contact_33_5165
timestamp 1624857261
transform 1 0 22168 0 1 49509
box 0 0 1 1
use contact_33  contact_33_4719
timestamp 1624857261
transform 1 0 22576 0 1 49509
box 0 0 1 1
use contact_33  contact_33_1684
timestamp 1624857261
transform 1 0 22984 0 1 49509
box 0 0 1 1
use contact_33  contact_33_4681
timestamp 1624857261
transform 1 0 23528 0 1 49101
box 0 0 1 1
use contact_33  contact_33_4680
timestamp 1624857261
transform 1 0 23528 0 1 49373
box 0 0 1 1
use contact_33  contact_33_4679
timestamp 1624857261
transform 1 0 23392 0 1 48965
box 0 0 1 1
use contact_33  contact_33_4678
timestamp 1624857261
transform 1 0 23392 0 1 48693
box 0 0 1 1
use contact_33  contact_33_4552
timestamp 1624857261
transform 1 0 23392 0 1 48149
box 0 0 1 1
use contact_33  contact_33_4513
timestamp 1624857261
transform 1 0 23528 0 1 49509
box 0 0 1 1
use contact_33  contact_33_4495
timestamp 1624857261
transform 1 0 23392 0 1 48557
box 0 0 1 1
use contact_33  contact_33_4494
timestamp 1624857261
transform 1 0 23392 0 1 48285
box 0 0 1 1
use contact_14  contact_14_629
timestamp 1624857261
transform 1 0 1797 0 1 49739
box 0 0 1 1
use contact_19  contact_19_629
timestamp 1624857261
transform 1 0 1794 0 1 49740
box 0 0 1 1
use contact_13  contact_13_629
timestamp 1624857261
transform 1 0 1801 0 1 49731
box 0 0 1 1
use contact_14  contact_14_628
timestamp 1624857261
transform 1 0 1797 0 1 50075
box 0 0 1 1
use contact_19  contact_19_628
timestamp 1624857261
transform 1 0 1794 0 1 50076
box 0 0 1 1
use contact_13  contact_13_628
timestamp 1624857261
transform 1 0 1801 0 1 50067
box 0 0 1 1
use contact_14  contact_14_627
timestamp 1624857261
transform 1 0 1797 0 1 50411
box 0 0 1 1
use contact_19  contact_19_627
timestamp 1624857261
transform 1 0 1794 0 1 50412
box 0 0 1 1
use contact_13  contact_13_627
timestamp 1624857261
transform 1 0 1801 0 1 50403
box 0 0 1 1
use contact_33  contact_33_5310
timestamp 1624857261
transform 1 0 1224 0 1 50869
box 0 0 1 1
use contact_7  contact_7_126
timestamp 1624857261
transform 1 0 1793 0 1 50743
box 0 0 1 1
use contact_14  contact_14_626
timestamp 1624857261
transform 1 0 1797 0 1 50747
box 0 0 1 1
use contact_19  contact_19_626
timestamp 1624857261
transform 1 0 1794 0 1 50748
box 0 0 1 1
use contact_13  contact_13_625
timestamp 1624857261
transform 1 0 1801 0 1 51075
box 0 0 1 1
use contact_13  contact_13_626
timestamp 1624857261
transform 1 0 1801 0 1 50739
box 0 0 1 1
use contact_33  contact_33_2206
timestamp 1624857261
transform 1 0 21760 0 1 50325
box 0 0 1 1
use contact_33  contact_33_2205
timestamp 1624857261
transform 1 0 21760 0 1 50597
box 0 0 1 1
use contact_33  contact_33_2236
timestamp 1624857261
transform 1 0 21896 0 1 49781
box 0 0 1 1
use contact_33  contact_33_5164
timestamp 1624857261
transform 1 0 22168 0 1 49781
box 0 0 1 1
use contact_33  contact_33_4718
timestamp 1624857261
transform 1 0 22576 0 1 49781
box 0 0 1 1
use contact_33  contact_33_1683
timestamp 1624857261
transform 1 0 22984 0 1 49781
box 0 0 1 1
use contact_33  contact_33_2238
timestamp 1624857261
transform 1 0 21896 0 1 49917
box 0 0 1 1
use contact_33  contact_33_5017
timestamp 1624857261
transform 1 0 22440 0 1 49917
box 0 0 1 1
use contact_33  contact_33_1543
timestamp 1624857261
transform 1 0 23120 0 1 49917
box 0 0 1 1
use contact_33  contact_33_2237
timestamp 1624857261
transform 1 0 21896 0 1 50189
box 0 0 1 1
use contact_33  contact_33_5159
timestamp 1624857261
transform 1 0 22168 0 1 50325
box 0 0 1 1
use contact_33  contact_33_4863
timestamp 1624857261
transform 1 0 22576 0 1 50325
box 0 0 1 1
use contact_33  contact_33_5016
timestamp 1624857261
transform 1 0 22440 0 1 50189
box 0 0 1 1
use contact_33  contact_33_1643
timestamp 1624857261
transform 1 0 22984 0 1 50325
box 0 0 1 1
use contact_33  contact_33_1544
timestamp 1624857261
transform 1 0 23120 0 1 50189
box 0 0 1 1
use contact_33  contact_33_1938
timestamp 1624857261
transform 1 0 21896 0 1 50733
box 0 0 1 1
use contact_33  contact_33_5024
timestamp 1624857261
transform 1 0 22304 0 1 50733
box 0 0 1 1
use contact_33  contact_33_5158
timestamp 1624857261
transform 1 0 22168 0 1 50597
box 0 0 1 1
use contact_33  contact_33_4862
timestamp 1624857261
transform 1 0 22576 0 1 50597
box 0 0 1 1
use contact_33  contact_33_5022
timestamp 1624857261
transform 1 0 22440 0 1 50733
box 0 0 1 1
use contact_33  contact_33_1644
timestamp 1624857261
transform 1 0 22984 0 1 50597
box 0 0 1 1
use contact_33  contact_33_1823
timestamp 1624857261
transform 1 0 22984 0 1 50733
box 0 0 1 1
use contact_33  contact_33_1937
timestamp 1624857261
transform 1 0 21896 0 1 51005
box 0 0 1 1
use contact_33  contact_33_5025
timestamp 1624857261
transform 1 0 22304 0 1 51005
box 0 0 1 1
use contact_33  contact_33_5023
timestamp 1624857261
transform 1 0 22440 0 1 51005
box 0 0 1 1
use contact_33  contact_33_1824
timestamp 1624857261
transform 1 0 22984 0 1 51005
box 0 0 1 1
use contact_33  contact_33_4611
timestamp 1624857261
transform 1 0 23392 0 1 50733
box 0 0 1 1
use contact_33  contact_33_4610
timestamp 1624857261
transform 1 0 23392 0 1 51005
box 0 0 1 1
use contact_33  contact_33_4609
timestamp 1624857261
transform 1 0 23528 0 1 50597
box 0 0 1 1
use contact_33  contact_33_4608
timestamp 1624857261
transform 1 0 23528 0 1 50325
box 0 0 1 1
use contact_33  contact_33_4512
timestamp 1624857261
transform 1 0 23528 0 1 49781
box 0 0 1 1
use contact_33  contact_33_4435
timestamp 1624857261
transform 1 0 23528 0 1 50189
box 0 0 1 1
use contact_33  contact_33_4434
timestamp 1624857261
transform 1 0 23528 0 1 49917
box 0 0 1 1
use contact_14  contact_14_624
timestamp 1624857261
transform 1 0 1797 0 1 51419
box 0 0 1 1
use contact_14  contact_14_625
timestamp 1624857261
transform 1 0 1797 0 1 51083
box 0 0 1 1
use contact_19  contact_19_624
timestamp 1624857261
transform 1 0 1794 0 1 51420
box 0 0 1 1
use contact_19  contact_19_625
timestamp 1624857261
transform 1 0 1794 0 1 51084
box 0 0 1 1
use contact_13  contact_13_624
timestamp 1624857261
transform 1 0 1801 0 1 51411
box 0 0 1 1
use contact_14  contact_14_623
timestamp 1624857261
transform 1 0 1797 0 1 51755
box 0 0 1 1
use contact_19  contact_19_623
timestamp 1624857261
transform 1 0 1794 0 1 51756
box 0 0 1 1
use contact_13  contact_13_623
timestamp 1624857261
transform 1 0 1801 0 1 51747
box 0 0 1 1
use contact_14  contact_14_622
timestamp 1624857261
transform 1 0 1797 0 1 52091
box 0 0 1 1
use contact_19  contact_19_622
timestamp 1624857261
transform 1 0 1794 0 1 52092
box 0 0 1 1
use contact_13  contact_13_622
timestamp 1624857261
transform 1 0 1801 0 1 52083
box 0 0 1 1
use contact_33  contact_33_5381
timestamp 1624857261
transform 1 0 1224 0 1 52501
box 0 0 1 1
use contact_7  contact_7_125
timestamp 1624857261
transform 1 0 1793 0 1 52423
box 0 0 1 1
use contact_14  contact_14_621
timestamp 1624857261
transform 1 0 1797 0 1 52427
box 0 0 1 1
use contact_19  contact_19_621
timestamp 1624857261
transform 1 0 1794 0 1 52428
box 0 0 1 1
use contact_13  contact_13_621
timestamp 1624857261
transform 1 0 1801 0 1 52419
box 0 0 1 1
use contact_33  contact_33_2080
timestamp 1624857261
transform 1 0 21760 0 1 51413
box 0 0 1 1
use contact_33  contact_33_2079
timestamp 1624857261
transform 1 0 21760 0 1 51141
box 0 0 1 1
use contact_33  contact_33_5175
timestamp 1624857261
transform 1 0 22168 0 1 51413
box 0 0 1 1
use contact_33  contact_33_2136
timestamp 1624857261
transform 1 0 21896 0 1 51957
box 0 0 1 1
use contact_33  contact_33_5174
timestamp 1624857261
transform 1 0 22168 0 1 51685
box 0 0 1 1
use contact_33  contact_33_1583
timestamp 1624857261
transform 1 0 22984 0 1 51821
box 0 0 1 1
use contact_33  contact_33_2135
timestamp 1624857261
transform 1 0 21896 0 1 52229
box 0 0 1 1
use contact_33  contact_33_5192
timestamp 1624857261
transform 1 0 22168 0 1 52229
box 0 0 1 1
use contact_33  contact_33_1584
timestamp 1624857261
transform 1 0 22984 0 1 52093
box 0 0 1 1
use contact_33  contact_33_1673
timestamp 1624857261
transform 1 0 22984 0 1 52229
box 0 0 1 1
use contact_33  contact_33_4865
timestamp 1624857261
transform 1 0 22712 0 1 52229
box 0 0 1 1
use contact_33  contact_33_5193
timestamp 1624857261
transform 1 0 22168 0 1 52501
box 0 0 1 1
use contact_33  contact_33_1674
timestamp 1624857261
transform 1 0 22984 0 1 52501
box 0 0 1 1
use contact_33  contact_33_4864
timestamp 1624857261
transform 1 0 22712 0 1 52501
box 0 0 1 1
use contact_33  contact_33_4581
timestamp 1624857261
transform 1 0 23392 0 1 52229
box 0 0 1 1
use contact_33  contact_33_4580
timestamp 1624857261
transform 1 0 23392 0 1 52501
box 0 0 1 1
use contact_33  contact_33_4579
timestamp 1624857261
transform 1 0 23392 0 1 52093
box 0 0 1 1
use contact_33  contact_33_4578
timestamp 1624857261
transform 1 0 23392 0 1 51821
box 0 0 1 1
use contact_33  contact_33_1514
timestamp 1624857261
transform 1 0 28560 0 1 51549
box 0 0 1 1
use contact_33  contact_33_1513
timestamp 1624857261
transform 1 0 28560 0 1 51277
box 0 0 1 1
use contact_33  contact_33_1398
timestamp 1624857261
transform 1 0 28424 0 1 51821
box 0 0 1 1
use contact_33  contact_33_1397
timestamp 1624857261
transform 1 0 28424 0 1 51549
box 0 0 1 1
use contact_14  contact_14_620
timestamp 1624857261
transform 1 0 1797 0 1 52763
box 0 0 1 1
use contact_19  contact_19_620
timestamp 1624857261
transform 1 0 1794 0 1 52764
box 0 0 1 1
use contact_13  contact_13_620
timestamp 1624857261
transform 1 0 1801 0 1 52755
box 0 0 1 1
use contact_14  contact_14_619
timestamp 1624857261
transform 1 0 1797 0 1 53099
box 0 0 1 1
use contact_19  contact_19_619
timestamp 1624857261
transform 1 0 1794 0 1 53100
box 0 0 1 1
use contact_13  contact_13_619
timestamp 1624857261
transform 1 0 1801 0 1 53091
box 0 0 1 1
use contact_14  contact_14_618
timestamp 1624857261
transform 1 0 1797 0 1 53435
box 0 0 1 1
use contact_19  contact_19_618
timestamp 1624857261
transform 1 0 1794 0 1 53436
box 0 0 1 1
use contact_13  contact_13_618
timestamp 1624857261
transform 1 0 1801 0 1 53427
box 0 0 1 1
use contact_7  contact_7_124
timestamp 1624857261
transform 1 0 1793 0 1 54103
box 0 0 1 1
use contact_14  contact_14_616
timestamp 1624857261
transform 1 0 1797 0 1 54107
box 0 0 1 1
use contact_14  contact_14_617
timestamp 1624857261
transform 1 0 1797 0 1 53771
box 0 0 1 1
use contact_19  contact_19_616
timestamp 1624857261
transform 1 0 1794 0 1 54108
box 0 0 1 1
use contact_19  contact_19_617
timestamp 1624857261
transform 1 0 1794 0 1 53772
box 0 0 1 1
use contact_13  contact_13_616
timestamp 1624857261
transform 1 0 1801 0 1 54099
box 0 0 1 1
use contact_13  contact_13_617
timestamp 1624857261
transform 1 0 1801 0 1 53763
box 0 0 1 1
use contact_33  contact_33_5375
timestamp 1624857261
transform 1 0 1224 0 1 54133
box 0 0 1 1
use contact_33  contact_33_2022
timestamp 1624857261
transform 1 0 21760 0 1 53725
box 0 0 1 1
use contact_33  contact_33_2021
timestamp 1624857261
transform 1 0 21760 0 1 53453
box 0 0 1 1
use contact_33  contact_33_2014
timestamp 1624857261
transform 1 0 21760 0 1 52637
box 0 0 1 1
use contact_33  contact_33_2013
timestamp 1624857261
transform 1 0 21760 0 1 52909
box 0 0 1 1
use contact_33  contact_33_5036
timestamp 1624857261
transform 1 0 22440 0 1 52637
box 0 0 1 1
use contact_33  contact_33_5037
timestamp 1624857261
transform 1 0 22440 0 1 52909
box 0 0 1 1
use contact_33  contact_33_1671
timestamp 1624857261
transform 1 0 23120 0 1 52909
box 0 0 1 1
use contact_33  contact_33_1672
timestamp 1624857261
transform 1 0 23120 0 1 52637
box 0 0 1 1
use contact_33  contact_33_4802
timestamp 1624857261
transform 1 0 22712 0 1 53045
box 0 0 1 1
use contact_33  contact_33_1725
timestamp 1624857261
transform 1 0 22984 0 1 53045
box 0 0 1 1
use contact_33  contact_33_5058
timestamp 1624857261
transform 1 0 22168 0 1 53453
box 0 0 1 1
use contact_33  contact_33_4803
timestamp 1624857261
transform 1 0 22712 0 1 53317
box 0 0 1 1
use contact_33  contact_33_4822
timestamp 1624857261
transform 1 0 22576 0 1 53453
box 0 0 1 1
use contact_33  contact_33_1726
timestamp 1624857261
transform 1 0 22984 0 1 53317
box 0 0 1 1
use contact_33  contact_33_1728
timestamp 1624857261
transform 1 0 23120 0 1 53453
box 0 0 1 1
use contact_33  contact_33_2159
timestamp 1624857261
transform 1 0 21896 0 1 53861
box 0 0 1 1
use contact_33  contact_33_5059
timestamp 1624857261
transform 1 0 22168 0 1 53725
box 0 0 1 1
use contact_33  contact_33_5061
timestamp 1624857261
transform 1 0 22168 0 1 53861
box 0 0 1 1
use contact_33  contact_33_4823
timestamp 1624857261
transform 1 0 22576 0 1 53725
box 0 0 1 1
use contact_33  contact_33_1660
timestamp 1624857261
transform 1 0 22984 0 1 53861
box 0 0 1 1
use contact_33  contact_33_1727
timestamp 1624857261
transform 1 0 23120 0 1 53725
box 0 0 1 1
use contact_33  contact_33_2160
timestamp 1624857261
transform 1 0 21896 0 1 54133
box 0 0 1 1
use contact_33  contact_33_5060
timestamp 1624857261
transform 1 0 22168 0 1 54133
box 0 0 1 1
use contact_33  contact_33_1659
timestamp 1624857261
transform 1 0 22984 0 1 54133
box 0 0 1 1
use contact_33  contact_33_4517
timestamp 1624857261
transform 1 0 23528 0 1 52637
box 0 0 1 1
use contact_33  contact_33_4516
timestamp 1624857261
transform 1 0 23528 0 1 52909
box 0 0 1 1
use contact_33  contact_33_4455
timestamp 1624857261
transform 1 0 23392 0 1 53317
box 0 0 1 1
use contact_33  contact_33_4454
timestamp 1624857261
transform 1 0 23392 0 1 53045
box 0 0 1 1
use contact_33  contact_33_4453
timestamp 1624857261
transform 1 0 23528 0 1 53453
box 0 0 1 1
use contact_33  contact_33_4452
timestamp 1624857261
transform 1 0 23528 0 1 53725
box 0 0 1 1
use contact_33  contact_33_4341
timestamp 1624857261
transform 1 0 23392 0 1 54133
box 0 0 1 1
use contact_33  contact_33_4340
timestamp 1624857261
transform 1 0 23392 0 1 53861
box 0 0 1 1
use contact_14  contact_14_615
timestamp 1624857261
transform 1 0 1797 0 1 54443
box 0 0 1 1
use contact_19  contact_19_615
timestamp 1624857261
transform 1 0 1794 0 1 54444
box 0 0 1 1
use contact_13  contact_13_615
timestamp 1624857261
transform 1 0 1801 0 1 54435
box 0 0 1 1
use contact_14  contact_14_614
timestamp 1624857261
transform 1 0 1797 0 1 54779
box 0 0 1 1
use contact_19  contact_19_614
timestamp 1624857261
transform 1 0 1794 0 1 54780
box 0 0 1 1
use contact_13  contact_13_614
timestamp 1624857261
transform 1 0 1801 0 1 54771
box 0 0 1 1
use contact_14  contact_14_612
timestamp 1624857261
transform 1 0 1797 0 1 55451
box 0 0 1 1
use contact_14  contact_14_613
timestamp 1624857261
transform 1 0 1797 0 1 55115
box 0 0 1 1
use contact_19  contact_19_612
timestamp 1624857261
transform 1 0 1794 0 1 55452
box 0 0 1 1
use contact_19  contact_19_613
timestamp 1624857261
transform 1 0 1794 0 1 55116
box 0 0 1 1
use contact_13  contact_13_612
timestamp 1624857261
transform 1 0 1801 0 1 55443
box 0 0 1 1
use contact_13  contact_13_613
timestamp 1624857261
transform 1 0 1801 0 1 55107
box 0 0 1 1
use contact_33  contact_33_2039
timestamp 1624857261
transform 1 0 21760 0 1 55493
box 0 0 1 1
use contact_33  contact_33_2006
timestamp 1624857261
transform 1 0 21760 0 1 54949
box 0 0 1 1
use contact_33  contact_33_2005
timestamp 1624857261
transform 1 0 21760 0 1 54677
box 0 0 1 1
use contact_33  contact_33_2157
timestamp 1624857261
transform 1 0 21896 0 1 54541
box 0 0 1 1
use contact_33  contact_33_2158
timestamp 1624857261
transform 1 0 21896 0 1 54269
box 0 0 1 1
use contact_33  contact_33_5012
timestamp 1624857261
transform 1 0 22440 0 1 54541
box 0 0 1 1
use contact_33  contact_33_5013
timestamp 1624857261
transform 1 0 22440 0 1 54269
box 0 0 1 1
use contact_33  contact_33_5014
timestamp 1624857261
transform 1 0 22304 0 1 54541
box 0 0 1 1
use contact_33  contact_33_5015
timestamp 1624857261
transform 1 0 22304 0 1 54269
box 0 0 1 1
use contact_33  contact_33_1559
timestamp 1624857261
transform 1 0 22984 0 1 54541
box 0 0 1 1
use contact_33  contact_33_1560
timestamp 1624857261
transform 1 0 22984 0 1 54269
box 0 0 1 1
use contact_33  contact_33_5132
timestamp 1624857261
transform 1 0 22168 0 1 54677
box 0 0 1 1
use contact_33  contact_33_5133
timestamp 1624857261
transform 1 0 22168 0 1 54949
box 0 0 1 1
use contact_33  contact_33_1647
timestamp 1624857261
transform 1 0 22984 0 1 54677
box 0 0 1 1
use contact_33  contact_33_1648
timestamp 1624857261
transform 1 0 22984 0 1 54949
box 0 0 1 1
use contact_33  contact_33_2004
timestamp 1624857261
transform 1 0 21896 0 1 55085
box 0 0 1 1
use contact_33  contact_33_2003
timestamp 1624857261
transform 1 0 21896 0 1 55357
box 0 0 1 1
use contact_33  contact_33_4842
timestamp 1624857261
transform 1 0 22576 0 1 55493
box 0 0 1 1
use contact_33  contact_33_4699
timestamp 1624857261
transform 1 0 23528 0 1 54541
box 0 0 1 1
use contact_33  contact_33_4698
timestamp 1624857261
transform 1 0 23528 0 1 54269
box 0 0 1 1
use contact_33  contact_33_4697
timestamp 1624857261
transform 1 0 23528 0 1 54677
box 0 0 1 1
use contact_33  contact_33_4696
timestamp 1624857261
transform 1 0 23528 0 1 54949
box 0 0 1 1
use contact_33  contact_33_1493
timestamp 1624857261
transform 1 0 28560 0 1 55629
box 0 0 1 1
use contact_33  contact_33_1396
timestamp 1624857261
transform 1 0 28288 0 1 54677
box 0 0 1 1
use contact_33  contact_33_1395
timestamp 1624857261
transform 1 0 28288 0 1 54405
box 0 0 1 1
use contact_33  contact_33_1370
timestamp 1624857261
transform 1 0 28560 0 1 55493
box 0 0 1 1
use contact_33  contact_33_1369
timestamp 1624857261
transform 1 0 28560 0 1 55221
box 0 0 1 1
use contact_33  contact_33_5317
timestamp 1624857261
transform 1 0 1224 0 1 55765
box 0 0 1 1
use contact_7  contact_7_123
timestamp 1624857261
transform 1 0 1793 0 1 55783
box 0 0 1 1
use contact_14  contact_14_610
timestamp 1624857261
transform 1 0 1797 0 1 56123
box 0 0 1 1
use contact_14  contact_14_611
timestamp 1624857261
transform 1 0 1797 0 1 55787
box 0 0 1 1
use contact_19  contact_19_610
timestamp 1624857261
transform 1 0 1794 0 1 56124
box 0 0 1 1
use contact_19  contact_19_611
timestamp 1624857261
transform 1 0 1794 0 1 55788
box 0 0 1 1
use contact_13  contact_13_610
timestamp 1624857261
transform 1 0 1801 0 1 56115
box 0 0 1 1
use contact_13  contact_13_611
timestamp 1624857261
transform 1 0 1801 0 1 55779
box 0 0 1 1
use contact_14  contact_14_609
timestamp 1624857261
transform 1 0 1797 0 1 56459
box 0 0 1 1
use contact_19  contact_19_609
timestamp 1624857261
transform 1 0 1794 0 1 56460
box 0 0 1 1
use contact_13  contact_13_609
timestamp 1624857261
transform 1 0 1801 0 1 56451
box 0 0 1 1
use contact_14  contact_14_608
timestamp 1624857261
transform 1 0 1797 0 1 56795
box 0 0 1 1
use contact_19  contact_19_608
timestamp 1624857261
transform 1 0 1794 0 1 56796
box 0 0 1 1
use contact_13  contact_13_608
timestamp 1624857261
transform 1 0 1801 0 1 56787
box 0 0 1 1
use contact_33  contact_33_5309
timestamp 1624857261
transform 1 0 1224 0 1 57397
box 0 0 1 1
use contact_14  contact_14_607
timestamp 1624857261
transform 1 0 1797 0 1 57131
box 0 0 1 1
use contact_19  contact_19_607
timestamp 1624857261
transform 1 0 1794 0 1 57132
box 0 0 1 1
use contact_13  contact_13_607
timestamp 1624857261
transform 1 0 1801 0 1 57123
box 0 0 1 1
use contact_7  contact_7_122
timestamp 1624857261
transform 1 0 1793 0 1 57463
box 0 0 1 1
use contact_14  contact_14_606
timestamp 1624857261
transform 1 0 1797 0 1 57467
box 0 0 1 1
use contact_19  contact_19_606
timestamp 1624857261
transform 1 0 1794 0 1 57468
box 0 0 1 1
use contact_13  contact_13_606
timestamp 1624857261
transform 1 0 1801 0 1 57459
box 0 0 1 1
use contact_33  contact_33_2042
timestamp 1624857261
transform 1 0 21896 0 1 56173
box 0 0 1 1
use contact_33  contact_33_2041
timestamp 1624857261
transform 1 0 21896 0 1 55901
box 0 0 1 1
use contact_33  contact_33_2040
timestamp 1624857261
transform 1 0 21760 0 1 55765
box 0 0 1 1
use contact_33  contact_33_1978
timestamp 1624857261
transform 1 0 21896 0 1 57397
box 0 0 1 1
use contact_33  contact_33_1977
timestamp 1624857261
transform 1 0 21896 0 1 57669
box 0 0 1 1
use contact_33  contact_33_4843
timestamp 1624857261
transform 1 0 22576 0 1 55765
box 0 0 1 1
use contact_33  contact_33_5070
timestamp 1624857261
transform 1 0 22440 0 1 56445
box 0 0 1 1
use contact_33  contact_33_5071
timestamp 1624857261
transform 1 0 22440 0 1 56173
box 0 0 1 1
use contact_33  contact_33_1679
timestamp 1624857261
transform 1 0 22984 0 1 56173
box 0 0 1 1
use contact_33  contact_33_1680
timestamp 1624857261
transform 1 0 22984 0 1 56445
box 0 0 1 1
use contact_33  contact_33_4846
timestamp 1624857261
transform 1 0 22712 0 1 56445
box 0 0 1 1
use contact_33  contact_33_4847
timestamp 1624857261
transform 1 0 22712 0 1 56173
box 0 0 1 1
use contact_33  contact_33_4444
timestamp 1624857261
transform 1 0 23392 0 1 56445
box 0 0 1 1
use contact_33  contact_33_4445
timestamp 1624857261
transform 1 0 23392 0 1 56173
box 0 0 1 1
use contact_33  contact_33_4994
timestamp 1624857261
transform 1 0 22440 0 1 56853
box 0 0 1 1
use contact_33  contact_33_4995
timestamp 1624857261
transform 1 0 22440 0 1 56581
box 0 0 1 1
use contact_33  contact_33_1677
timestamp 1624857261
transform 1 0 22984 0 1 56853
box 0 0 1 1
use contact_33  contact_33_1678
timestamp 1624857261
transform 1 0 22984 0 1 56581
box 0 0 1 1
use contact_33  contact_33_4540
timestamp 1624857261
transform 1 0 23528 0 1 56581
box 0 0 1 1
use contact_33  contact_33_4541
timestamp 1624857261
transform 1 0 23528 0 1 56853
box 0 0 1 1
use contact_33  contact_33_1707
timestamp 1624857261
transform 1 0 23120 0 1 56989
box 0 0 1 1
use contact_33  contact_33_1708
timestamp 1624857261
transform 1 0 23120 0 1 57261
box 0 0 1 1
use contact_33  contact_33_4542
timestamp 1624857261
transform 1 0 23528 0 1 57261
box 0 0 1 1
use contact_33  contact_33_4543
timestamp 1624857261
transform 1 0 23528 0 1 56989
box 0 0 1 1
use contact_33  contact_33_4712
timestamp 1624857261
transform 1 0 22712 0 1 57669
box 0 0 1 1
use contact_33  contact_33_4713
timestamp 1624857261
transform 1 0 22712 0 1 57397
box 0 0 1 1
use contact_33  contact_33_1705
timestamp 1624857261
transform 1 0 23120 0 1 57669
box 0 0 1 1
use contact_33  contact_33_1706
timestamp 1624857261
transform 1 0 23120 0 1 57397
box 0 0 1 1
use contact_33  contact_33_4642
timestamp 1624857261
transform 1 0 23392 0 1 57397
box 0 0 1 1
use contact_33  contact_33_4643
timestamp 1624857261
transform 1 0 23392 0 1 57669
box 0 0 1 1
use contact_33  contact_33_1494
timestamp 1624857261
transform 1 0 28560 0 1 55901
box 0 0 1 1
use contact_14  contact_14_604
timestamp 1624857261
transform 1 0 1797 0 1 58139
box 0 0 1 1
use contact_14  contact_14_605
timestamp 1624857261
transform 1 0 1797 0 1 57803
box 0 0 1 1
use contact_19  contact_19_604
timestamp 1624857261
transform 1 0 1794 0 1 58140
box 0 0 1 1
use contact_19  contact_19_605
timestamp 1624857261
transform 1 0 1794 0 1 57804
box 0 0 1 1
use contact_13  contact_13_604
timestamp 1624857261
transform 1 0 1801 0 1 58131
box 0 0 1 1
use contact_13  contact_13_605
timestamp 1624857261
transform 1 0 1801 0 1 57795
box 0 0 1 1
use contact_14  contact_14_603
timestamp 1624857261
transform 1 0 1797 0 1 58475
box 0 0 1 1
use contact_19  contact_19_603
timestamp 1624857261
transform 1 0 1794 0 1 58476
box 0 0 1 1
use contact_13  contact_13_603
timestamp 1624857261
transform 1 0 1801 0 1 58467
box 0 0 1 1
use contact_14  contact_14_602
timestamp 1624857261
transform 1 0 1797 0 1 58811
box 0 0 1 1
use contact_19  contact_19_602
timestamp 1624857261
transform 1 0 1794 0 1 58812
box 0 0 1 1
use contact_13  contact_13_602
timestamp 1624857261
transform 1 0 1801 0 1 58803
box 0 0 1 1
use contact_33  contact_33_5313
timestamp 1624857261
transform 1 0 1224 0 1 59165
box 0 0 1 1
use contact_7  contact_7_121
timestamp 1624857261
transform 1 0 1793 0 1 59143
box 0 0 1 1
use contact_14  contact_14_600
timestamp 1624857261
transform 1 0 1797 0 1 59483
box 0 0 1 1
use contact_14  contact_14_601
timestamp 1624857261
transform 1 0 1797 0 1 59147
box 0 0 1 1
use contact_19  contact_19_600
timestamp 1624857261
transform 1 0 1794 0 1 59484
box 0 0 1 1
use contact_19  contact_19_601
timestamp 1624857261
transform 1 0 1794 0 1 59148
box 0 0 1 1
use contact_13  contact_13_600
timestamp 1624857261
transform 1 0 1801 0 1 59475
box 0 0 1 1
use contact_13  contact_13_601
timestamp 1624857261
transform 1 0 1801 0 1 59139
box 0 0 1 1
use contact_33  contact_33_2045
timestamp 1624857261
transform 1 0 21760 0 1 57805
box 0 0 1 1
use contact_33  contact_33_2046
timestamp 1624857261
transform 1 0 21760 0 1 58077
box 0 0 1 1
use contact_33  contact_33_2069
timestamp 1624857261
transform 1 0 21896 0 1 58213
box 0 0 1 1
use contact_33  contact_33_5051
timestamp 1624857261
transform 1 0 22168 0 1 58213
box 0 0 1 1
use contact_33  contact_33_2068
timestamp 1624857261
transform 1 0 21896 0 1 58621
box 0 0 1 1
use contact_33  contact_33_2070
timestamp 1624857261
transform 1 0 21896 0 1 58485
box 0 0 1 1
use contact_33  contact_33_5050
timestamp 1624857261
transform 1 0 22168 0 1 58485
box 0 0 1 1
use contact_33  contact_33_4981
timestamp 1624857261
transform 1 0 22304 0 1 58621
box 0 0 1 1
use contact_33  contact_33_1959
timestamp 1624857261
transform 1 0 21760 0 1 59029
box 0 0 1 1
use contact_33  contact_33_2067
timestamp 1624857261
transform 1 0 21896 0 1 58893
box 0 0 1 1
use contact_33  contact_33_4980
timestamp 1624857261
transform 1 0 22304 0 1 58893
box 0 0 1 1
use contact_33  contact_33_1960
timestamp 1624857261
transform 1 0 21760 0 1 59301
box 0 0 1 1
use contact_33  contact_33_2083
timestamp 1624857261
transform 1 0 21896 0 1 59437
box 0 0 1 1
use contact_33  contact_33_2084
timestamp 1624857261
transform 1 0 21896 0 1 59709
box 0 0 1 1
use contact_33  contact_33_5078
timestamp 1624857261
transform 1 0 22304 0 1 59437
box 0 0 1 1
use contact_33  contact_33_5079
timestamp 1624857261
transform 1 0 22304 0 1 59709
box 0 0 1 1
use contact_33  contact_33_4906
timestamp 1624857261
transform 1 0 22440 0 1 58077
box 0 0 1 1
use contact_33  contact_33_4907
timestamp 1624857261
transform 1 0 22440 0 1 57805
box 0 0 1 1
use contact_33  contact_33_1763
timestamp 1624857261
transform 1 0 22984 0 1 57805
box 0 0 1 1
use contact_33  contact_33_1764
timestamp 1624857261
transform 1 0 22984 0 1 58077
box 0 0 1 1
use contact_33  contact_33_4640
timestamp 1624857261
transform 1 0 23528 0 1 58077
box 0 0 1 1
use contact_33  contact_33_4641
timestamp 1624857261
transform 1 0 23528 0 1 57805
box 0 0 1 1
use contact_33  contact_33_4882
timestamp 1624857261
transform 1 0 22712 0 1 58213
box 0 0 1 1
use contact_33  contact_33_4883
timestamp 1624857261
transform 1 0 22712 0 1 58485
box 0 0 1 1
use contact_33  contact_33_1855
timestamp 1624857261
transform 1 0 22984 0 1 58213
box 0 0 1 1
use contact_33  contact_33_1856
timestamp 1624857261
transform 1 0 22984 0 1 58485
box 0 0 1 1
use contact_33  contact_33_4442
timestamp 1624857261
transform 1 0 23392 0 1 58213
box 0 0 1 1
use contact_33  contact_33_4443
timestamp 1624857261
transform 1 0 23392 0 1 58485
box 0 0 1 1
use contact_33  contact_33_1567
timestamp 1624857261
transform 1 0 22984 0 1 59029
box 0 0 1 1
use contact_33  contact_33_1853
timestamp 1624857261
transform 1 0 22984 0 1 58893
box 0 0 1 1
use contact_33  contact_33_1854
timestamp 1624857261
transform 1 0 22984 0 1 58621
box 0 0 1 1
use contact_33  contact_33_4440
timestamp 1624857261
transform 1 0 23392 0 1 58893
box 0 0 1 1
use contact_33  contact_33_4441
timestamp 1624857261
transform 1 0 23392 0 1 58621
box 0 0 1 1
use contact_33  contact_33_4486
timestamp 1624857261
transform 1 0 23528 0 1 59029
box 0 0 1 1
use contact_33  contact_33_1568
timestamp 1624857261
transform 1 0 22984 0 1 59301
box 0 0 1 1
use contact_33  contact_33_4487
timestamp 1624857261
transform 1 0 23528 0 1 59301
box 0 0 1 1
use contact_33  contact_33_1487
timestamp 1624857261
transform 1 0 28288 0 1 59573
box 0 0 1 1
use contact_33  contact_33_1426
timestamp 1624857261
transform 1 0 28560 0 1 58621
box 0 0 1 1
use contact_33  contact_33_1425
timestamp 1624857261
transform 1 0 28560 0 1 58349
box 0 0 1 1
use contact_14  contact_14_598
timestamp 1624857261
transform 1 0 1797 0 1 60155
box 0 0 1 1
use contact_14  contact_14_599
timestamp 1624857261
transform 1 0 1797 0 1 59819
box 0 0 1 1
use contact_19  contact_19_598
timestamp 1624857261
transform 1 0 1794 0 1 60156
box 0 0 1 1
use contact_19  contact_19_599
timestamp 1624857261
transform 1 0 1794 0 1 59820
box 0 0 1 1
use contact_13  contact_13_598
timestamp 1624857261
transform 1 0 1801 0 1 60147
box 0 0 1 1
use contact_13  contact_13_599
timestamp 1624857261
transform 1 0 1801 0 1 59811
box 0 0 1 1
use contact_14  contact_14_597
timestamp 1624857261
transform 1 0 1797 0 1 60491
box 0 0 1 1
use contact_19  contact_19_597
timestamp 1624857261
transform 1 0 1794 0 1 60492
box 0 0 1 1
use contact_13  contact_13_597
timestamp 1624857261
transform 1 0 1801 0 1 60483
box 0 0 1 1
use contact_33  contact_33_5358
timestamp 1624857261
transform 1 0 1224 0 1 60933
box 0 0 1 1
use contact_7  contact_7_120
timestamp 1624857261
transform 1 0 1793 0 1 60823
box 0 0 1 1
use contact_14  contact_14_596
timestamp 1624857261
transform 1 0 1797 0 1 60827
box 0 0 1 1
use contact_19  contact_19_596
timestamp 1624857261
transform 1 0 1794 0 1 60828
box 0 0 1 1
use contact_13  contact_13_596
timestamp 1624857261
transform 1 0 1801 0 1 60819
box 0 0 1 1
use contact_14  contact_14_594
timestamp 1624857261
transform 1 0 1797 0 1 61499
box 0 0 1 1
use contact_14  contact_14_595
timestamp 1624857261
transform 1 0 1797 0 1 61163
box 0 0 1 1
use contact_19  contact_19_594
timestamp 1624857261
transform 1 0 1794 0 1 61500
box 0 0 1 1
use contact_19  contact_19_595
timestamp 1624857261
transform 1 0 1794 0 1 61164
box 0 0 1 1
use contact_13  contact_13_594
timestamp 1624857261
transform 1 0 1801 0 1 61491
box 0 0 1 1
use contact_13  contact_13_595
timestamp 1624857261
transform 1 0 1801 0 1 61155
box 0 0 1 1
use contact_33  contact_33_5161
timestamp 1624857261
transform 1 0 22168 0 1 60117
box 0 0 1 1
use contact_33  contact_33_5160
timestamp 1624857261
transform 1 0 22168 0 1 60389
box 0 0 1 1
use contact_33  contact_33_4941
timestamp 1624857261
transform 1 0 22304 0 1 61613
box 0 0 1 1
use contact_33  contact_33_4940
timestamp 1624857261
transform 1 0 22304 0 1 61341
box 0 0 1 1
use contact_33  contact_33_2100
timestamp 1624857261
transform 1 0 21896 0 1 61613
box 0 0 1 1
use contact_33  contact_33_2099
timestamp 1624857261
transform 1 0 21896 0 1 61341
box 0 0 1 1
use contact_33  contact_33_2082
timestamp 1624857261
transform 1 0 21896 0 1 59845
box 0 0 1 1
use contact_33  contact_33_2081
timestamp 1624857261
transform 1 0 21896 0 1 60117
box 0 0 1 1
use contact_33  contact_33_1888
timestamp 1624857261
transform 1 0 23120 0 1 60117
box 0 0 1 1
use contact_33  contact_33_4630
timestamp 1624857261
transform 1 0 23528 0 1 60117
box 0 0 1 1
use contact_33  contact_33_1562
timestamp 1624857261
transform 1 0 23120 0 1 60525
box 0 0 1 1
use contact_33  contact_33_1887
timestamp 1624857261
transform 1 0 23120 0 1 60389
box 0 0 1 1
use contact_33  contact_33_4629
timestamp 1624857261
transform 1 0 23392 0 1 60525
box 0 0 1 1
use contact_33  contact_33_4631
timestamp 1624857261
transform 1 0 23528 0 1 60389
box 0 0 1 1
use contact_33  contact_33_4879
timestamp 1624857261
transform 1 0 22712 0 1 60933
box 0 0 1 1
use contact_33  contact_33_4934
timestamp 1624857261
transform 1 0 22440 0 1 60661
box 0 0 1 1
use contact_33  contact_33_4935
timestamp 1624857261
transform 1 0 22440 0 1 60933
box 0 0 1 1
use contact_33  contact_33_1552
timestamp 1624857261
transform 1 0 22984 0 1 60933
box 0 0 1 1
use contact_33  contact_33_1561
timestamp 1624857261
transform 1 0 23120 0 1 60797
box 0 0 1 1
use contact_33  contact_33_4576
timestamp 1624857261
transform 1 0 23528 0 1 60933
box 0 0 1 1
use contact_33  contact_33_4628
timestamp 1624857261
transform 1 0 23392 0 1 60797
box 0 0 1 1
use contact_33  contact_33_4878
timestamp 1624857261
transform 1 0 22712 0 1 61205
box 0 0 1 1
use contact_33  contact_33_4938
timestamp 1624857261
transform 1 0 22440 0 1 61341
box 0 0 1 1
use contact_33  contact_33_1532
timestamp 1624857261
transform 1 0 22984 0 1 61341
box 0 0 1 1
use contact_33  contact_33_1551
timestamp 1624857261
transform 1 0 22984 0 1 61205
box 0 0 1 1
use contact_33  contact_33_4575
timestamp 1624857261
transform 1 0 23528 0 1 61341
box 0 0 1 1
use contact_33  contact_33_4577
timestamp 1624857261
transform 1 0 23528 0 1 61205
box 0 0 1 1
use contact_33  contact_33_4939
timestamp 1624857261
transform 1 0 22440 0 1 61613
box 0 0 1 1
use contact_33  contact_33_1531
timestamp 1624857261
transform 1 0 22984 0 1 61613
box 0 0 1 1
use contact_33  contact_33_4574
timestamp 1624857261
transform 1 0 23528 0 1 61613
box 0 0 1 1
use contact_33  contact_33_1488
timestamp 1624857261
transform 1 0 28288 0 1 59981
box 0 0 1 1
use contact_33  contact_33_1474
timestamp 1624857261
transform 1 0 28560 0 1 59981
box 0 0 1 1
use contact_33  contact_33_1473
timestamp 1624857261
transform 1 0 28560 0 1 60253
box 0 0 1 1
use contact_14  contact_14_592
timestamp 1624857261
transform 1 0 1797 0 1 62171
box 0 0 1 1
use contact_14  contact_14_593
timestamp 1624857261
transform 1 0 1797 0 1 61835
box 0 0 1 1
use contact_19  contact_19_592
timestamp 1624857261
transform 1 0 1794 0 1 62172
box 0 0 1 1
use contact_19  contact_19_593
timestamp 1624857261
transform 1 0 1794 0 1 61836
box 0 0 1 1
use contact_13  contact_13_592
timestamp 1624857261
transform 1 0 1801 0 1 62163
box 0 0 1 1
use contact_13  contact_13_593
timestamp 1624857261
transform 1 0 1801 0 1 61827
box 0 0 1 1
use contact_33  contact_33_5311
timestamp 1624857261
transform 1 0 1224 0 1 62565
box 0 0 1 1
use contact_7  contact_7_119
timestamp 1624857261
transform 1 0 1793 0 1 62503
box 0 0 1 1
use contact_14  contact_14_591
timestamp 1624857261
transform 1 0 1797 0 1 62507
box 0 0 1 1
use contact_19  contact_19_591
timestamp 1624857261
transform 1 0 1794 0 1 62508
box 0 0 1 1
use contact_13  contact_13_591
timestamp 1624857261
transform 1 0 1801 0 1 62499
box 0 0 1 1
use contact_14  contact_14_590
timestamp 1624857261
transform 1 0 1797 0 1 62843
box 0 0 1 1
use contact_19  contact_19_590
timestamp 1624857261
transform 1 0 1794 0 1 62844
box 0 0 1 1
use contact_13  contact_13_590
timestamp 1624857261
transform 1 0 1801 0 1 62835
box 0 0 1 1
use contact_14  contact_14_588
timestamp 1624857261
transform 1 0 1797 0 1 63515
box 0 0 1 1
use contact_14  contact_14_589
timestamp 1624857261
transform 1 0 1797 0 1 63179
box 0 0 1 1
use contact_19  contact_19_588
timestamp 1624857261
transform 1 0 1794 0 1 63516
box 0 0 1 1
use contact_19  contact_19_589
timestamp 1624857261
transform 1 0 1794 0 1 63180
box 0 0 1 1
use contact_13  contact_13_588
timestamp 1624857261
transform 1 0 1801 0 1 63507
box 0 0 1 1
use contact_13  contact_13_589
timestamp 1624857261
transform 1 0 1801 0 1 63171
box 0 0 1 1
use contact_33  contact_33_2256
timestamp 1624857261
transform 1 0 21760 0 1 62157
box 0 0 1 1
use contact_33  contact_33_2257
timestamp 1624857261
transform 1 0 21896 0 1 61749
box 0 0 1 1
use contact_33  contact_33_2258
timestamp 1624857261
transform 1 0 21896 0 1 62021
box 0 0 1 1
use contact_33  contact_33_4953
timestamp 1624857261
transform 1 0 22168 0 1 62157
box 0 0 1 1
use contact_33  contact_33_2086
timestamp 1624857261
transform 1 0 21760 0 1 62565
box 0 0 1 1
use contact_33  contact_33_2255
timestamp 1624857261
transform 1 0 21760 0 1 62429
box 0 0 1 1
use contact_33  contact_33_4952
timestamp 1624857261
transform 1 0 22168 0 1 62429
box 0 0 1 1
use contact_33  contact_33_1943
timestamp 1624857261
transform 1 0 21896 0 1 63245
box 0 0 1 1
use contact_33  contact_33_1944
timestamp 1624857261
transform 1 0 21896 0 1 62973
box 0 0 1 1
use contact_33  contact_33_2085
timestamp 1624857261
transform 1 0 21760 0 1 62837
box 0 0 1 1
use contact_33  contact_33_1995
timestamp 1624857261
transform 1 0 21760 0 1 63381
box 0 0 1 1
use contact_33  contact_33_1996
timestamp 1624857261
transform 1 0 21760 0 1 63653
box 0 0 1 1
use contact_33  contact_33_5080
timestamp 1624857261
transform 1 0 22304 0 1 63381
box 0 0 1 1
use contact_33  contact_33_5081
timestamp 1624857261
transform 1 0 22304 0 1 63653
box 0 0 1 1
use contact_33  contact_33_4950
timestamp 1624857261
transform 1 0 22440 0 1 61749
box 0 0 1 1
use contact_33  contact_33_4951
timestamp 1624857261
transform 1 0 22440 0 1 62021
box 0 0 1 1
use contact_33  contact_33_1613
timestamp 1624857261
transform 1 0 22984 0 1 61749
box 0 0 1 1
use contact_33  contact_33_1614
timestamp 1624857261
transform 1 0 22984 0 1 62021
box 0 0 1 1
use contact_33  contact_33_1693
timestamp 1624857261
transform 1 0 22984 0 1 62157
box 0 0 1 1
use contact_33  contact_33_4560
timestamp 1624857261
transform 1 0 23392 0 1 61749
box 0 0 1 1
use contact_33  contact_33_4561
timestamp 1624857261
transform 1 0 23392 0 1 62021
box 0 0 1 1
use contact_33  contact_33_4582
timestamp 1624857261
transform 1 0 23528 0 1 62157
box 0 0 1 1
use contact_33  contact_33_4795
timestamp 1624857261
transform 1 0 22576 0 1 62565
box 0 0 1 1
use contact_33  contact_33_1692
timestamp 1624857261
transform 1 0 22984 0 1 62565
box 0 0 1 1
use contact_33  contact_33_1694
timestamp 1624857261
transform 1 0 22984 0 1 62429
box 0 0 1 1
use contact_33  contact_33_4583
timestamp 1624857261
transform 1 0 23528 0 1 62429
box 0 0 1 1
use contact_33  contact_33_4606
timestamp 1624857261
transform 1 0 23392 0 1 62565
box 0 0 1 1
use contact_33  contact_33_4794
timestamp 1624857261
transform 1 0 22576 0 1 62837
box 0 0 1 1
use contact_33  contact_33_1553
timestamp 1624857261
transform 1 0 23120 0 1 62973
box 0 0 1 1
use contact_33  contact_33_1691
timestamp 1624857261
transform 1 0 22984 0 1 62837
box 0 0 1 1
use contact_33  contact_33_4605
timestamp 1624857261
transform 1 0 23392 0 1 62973
box 0 0 1 1
use contact_33  contact_33_4607
timestamp 1624857261
transform 1 0 23392 0 1 62837
box 0 0 1 1
use contact_33  contact_33_1554
timestamp 1624857261
transform 1 0 23120 0 1 63245
box 0 0 1 1
use contact_33  contact_33_4604
timestamp 1624857261
transform 1 0 23392 0 1 63245
box 0 0 1 1
use contact_33  contact_33_1496
timestamp 1624857261
transform 1 0 28288 0 1 63381
box 0 0 1 1
use contact_33  contact_33_1495
timestamp 1624857261
transform 1 0 28288 0 1 63109
box 0 0 1 1
use contact_33  contact_33_1498
timestamp 1624857261
transform 1 0 28560 0 1 63517
box 0 0 1 1
use contact_14  contact_14_587
timestamp 1624857261
transform 1 0 1797 0 1 63851
box 0 0 1 1
use contact_19  contact_19_587
timestamp 1624857261
transform 1 0 1794 0 1 63852
box 0 0 1 1
use contact_13  contact_13_587
timestamp 1624857261
transform 1 0 1801 0 1 63843
box 0 0 1 1
use contact_33  contact_33_5298
timestamp 1624857261
transform 1 0 1224 0 1 64333
box 0 0 1 1
use contact_7  contact_7_118
timestamp 1624857261
transform 1 0 1793 0 1 64183
box 0 0 1 1
use contact_14  contact_14_585
timestamp 1624857261
transform 1 0 1797 0 1 64523
box 0 0 1 1
use contact_14  contact_14_586
timestamp 1624857261
transform 1 0 1797 0 1 64187
box 0 0 1 1
use contact_19  contact_19_585
timestamp 1624857261
transform 1 0 1794 0 1 64524
box 0 0 1 1
use contact_19  contact_19_586
timestamp 1624857261
transform 1 0 1794 0 1 64188
box 0 0 1 1
use contact_13  contact_13_585
timestamp 1624857261
transform 1 0 1801 0 1 64515
box 0 0 1 1
use contact_13  contact_13_586
timestamp 1624857261
transform 1 0 1801 0 1 64179
box 0 0 1 1
use contact_14  contact_14_584
timestamp 1624857261
transform 1 0 1797 0 1 64859
box 0 0 1 1
use contact_19  contact_19_584
timestamp 1624857261
transform 1 0 1794 0 1 64860
box 0 0 1 1
use contact_13  contact_13_584
timestamp 1624857261
transform 1 0 1801 0 1 64851
box 0 0 1 1
use contact_14  contact_14_583
timestamp 1624857261
transform 1 0 1797 0 1 65195
box 0 0 1 1
use contact_19  contact_19_583
timestamp 1624857261
transform 1 0 1794 0 1 65196
box 0 0 1 1
use contact_13  contact_13_583
timestamp 1624857261
transform 1 0 1801 0 1 65187
box 0 0 1 1
use contact_14  contact_14_582
timestamp 1624857261
transform 1 0 1797 0 1 65531
box 0 0 1 1
use contact_19  contact_19_582
timestamp 1624857261
transform 1 0 1794 0 1 65532
box 0 0 1 1
use contact_13  contact_13_582
timestamp 1624857261
transform 1 0 1801 0 1 65523
box 0 0 1 1
use contact_33  contact_33_1997
timestamp 1624857261
transform 1 0 21896 0 1 64061
box 0 0 1 1
use contact_33  contact_33_1998
timestamp 1624857261
transform 1 0 21896 0 1 63789
box 0 0 1 1
use contact_33  contact_33_5184
timestamp 1624857261
transform 1 0 22168 0 1 64061
box 0 0 1 1
use contact_33  contact_33_5185
timestamp 1624857261
transform 1 0 22168 0 1 64333
box 0 0 1 1
use contact_33  contact_33_5020
timestamp 1624857261
transform 1 0 22304 0 1 64877
box 0 0 1 1
use contact_33  contact_33_2253
timestamp 1624857261
transform 1 0 21896 0 1 65557
box 0 0 1 1
use contact_33  contact_33_2254
timestamp 1624857261
transform 1 0 21896 0 1 65285
box 0 0 1 1
use contact_33  contact_33_5021
timestamp 1624857261
transform 1 0 22304 0 1 65149
box 0 0 1 1
use contact_33  contact_33_2036
timestamp 1624857261
transform 1 0 21760 0 1 65693
box 0 0 1 1
use contact_33  contact_33_4948
timestamp 1624857261
transform 1 0 22304 0 1 65693
box 0 0 1 1
use contact_33  contact_33_4766
timestamp 1624857261
transform 1 0 22576 0 1 64061
box 0 0 1 1
use contact_33  contact_33_4767
timestamp 1624857261
transform 1 0 22576 0 1 64333
box 0 0 1 1
use contact_33  contact_33_1685
timestamp 1624857261
transform 1 0 22984 0 1 64469
box 0 0 1 1
use contact_33  contact_33_4700
timestamp 1624857261
transform 1 0 23528 0 1 64469
box 0 0 1 1
use contact_33  contact_33_5018
timestamp 1624857261
transform 1 0 22440 0 1 64877
box 0 0 1 1
use contact_33  contact_33_1686
timestamp 1624857261
transform 1 0 22984 0 1 64741
box 0 0 1 1
use contact_33  contact_33_1688
timestamp 1624857261
transform 1 0 23120 0 1 64877
box 0 0 1 1
use contact_33  contact_33_4701
timestamp 1624857261
transform 1 0 23528 0 1 64741
box 0 0 1 1
use contact_33  contact_33_4703
timestamp 1624857261
transform 1 0 23392 0 1 64877
box 0 0 1 1
use contact_33  contact_33_4770
timestamp 1624857261
transform 1 0 22576 0 1 65285
box 0 0 1 1
use contact_33  contact_33_5019
timestamp 1624857261
transform 1 0 22440 0 1 65149
box 0 0 1 1
use contact_33  contact_33_1579
timestamp 1624857261
transform 1 0 22984 0 1 65285
box 0 0 1 1
use contact_33  contact_33_1687
timestamp 1624857261
transform 1 0 23120 0 1 65149
box 0 0 1 1
use contact_33  contact_33_4646
timestamp 1624857261
transform 1 0 23528 0 1 65285
box 0 0 1 1
use contact_33  contact_33_4702
timestamp 1624857261
transform 1 0 23392 0 1 65149
box 0 0 1 1
use contact_33  contact_33_4771
timestamp 1624857261
transform 1 0 22576 0 1 65557
box 0 0 1 1
use contact_33  contact_33_1580
timestamp 1624857261
transform 1 0 22984 0 1 65557
box 0 0 1 1
use contact_33  contact_33_1865
timestamp 1624857261
transform 1 0 23120 0 1 65693
box 0 0 1 1
use contact_33  contact_33_4645
timestamp 1624857261
transform 1 0 23528 0 1 65693
box 0 0 1 1
use contact_33  contact_33_4647
timestamp 1624857261
transform 1 0 23528 0 1 65557
box 0 0 1 1
use contact_33  contact_33_1497
timestamp 1624857261
transform 1 0 28560 0 1 63789
box 0 0 1 1
use contact_33  contact_33_5338
timestamp 1624857261
transform 1 0 1224 0 1 65829
box 0 0 1 1
use contact_7  contact_7_117
timestamp 1624857261
transform 1 0 1793 0 1 65863
box 0 0 1 1
use contact_14  contact_14_580
timestamp 1624857261
transform 1 0 1797 0 1 66203
box 0 0 1 1
use contact_14  contact_14_581
timestamp 1624857261
transform 1 0 1797 0 1 65867
box 0 0 1 1
use contact_19  contact_19_580
timestamp 1624857261
transform 1 0 1794 0 1 66204
box 0 0 1 1
use contact_19  contact_19_581
timestamp 1624857261
transform 1 0 1794 0 1 65868
box 0 0 1 1
use contact_13  contact_13_580
timestamp 1624857261
transform 1 0 1801 0 1 66195
box 0 0 1 1
use contact_13  contact_13_581
timestamp 1624857261
transform 1 0 1801 0 1 65859
box 0 0 1 1
use contact_14  contact_14_579
timestamp 1624857261
transform 1 0 1797 0 1 66539
box 0 0 1 1
use contact_19  contact_19_579
timestamp 1624857261
transform 1 0 1794 0 1 66540
box 0 0 1 1
use contact_13  contact_13_579
timestamp 1624857261
transform 1 0 1801 0 1 66531
box 0 0 1 1
use contact_14  contact_14_578
timestamp 1624857261
transform 1 0 1797 0 1 66875
box 0 0 1 1
use contact_19  contact_19_578
timestamp 1624857261
transform 1 0 1794 0 1 66876
box 0 0 1 1
use contact_13  contact_13_578
timestamp 1624857261
transform 1 0 1801 0 1 66867
box 0 0 1 1
use contact_33  contact_33_4949
timestamp 1624857261
transform 1 0 22304 0 1 65965
box 0 0 1 1
use contact_33  contact_33_2132
timestamp 1624857261
transform 1 0 21760 0 1 66509
box 0 0 1 1
use contact_33  contact_33_2131
timestamp 1624857261
transform 1 0 21760 0 1 66781
box 0 0 1 1
use contact_33  contact_33_2130
timestamp 1624857261
transform 1 0 21896 0 1 66373
box 0 0 1 1
use contact_33  contact_33_2129
timestamp 1624857261
transform 1 0 21896 0 1 66101
box 0 0 1 1
use contact_33  contact_33_2101
timestamp 1624857261
transform 1 0 21896 0 1 66917
box 0 0 1 1
use contact_33  contact_33_2035
timestamp 1624857261
transform 1 0 21760 0 1 65965
box 0 0 1 1
use contact_33  contact_33_4912
timestamp 1624857261
transform 1 0 22440 0 1 66101
box 0 0 1 1
use contact_33  contact_33_1864
timestamp 1624857261
transform 1 0 23120 0 1 66101
box 0 0 1 1
use contact_33  contact_33_1866
timestamp 1624857261
transform 1 0 23120 0 1 65965
box 0 0 1 1
use contact_33  contact_33_4592
timestamp 1624857261
transform 1 0 23392 0 1 66101
box 0 0 1 1
use contact_33  contact_33_4644
timestamp 1624857261
transform 1 0 23528 0 1 65965
box 0 0 1 1
use contact_33  contact_33_4781
timestamp 1624857261
transform 1 0 22576 0 1 66509
box 0 0 1 1
use contact_33  contact_33_4913
timestamp 1624857261
transform 1 0 22440 0 1 66373
box 0 0 1 1
use contact_33  contact_33_1603
timestamp 1624857261
transform 1 0 22984 0 1 66509
box 0 0 1 1
use contact_33  contact_33_1863
timestamp 1624857261
transform 1 0 23120 0 1 66373
box 0 0 1 1
use contact_33  contact_33_4593
timestamp 1624857261
transform 1 0 23392 0 1 66373
box 0 0 1 1
use contact_33  contact_33_4595
timestamp 1624857261
transform 1 0 23528 0 1 66509
box 0 0 1 1
use contact_33  contact_33_4780
timestamp 1624857261
transform 1 0 22576 0 1 66781
box 0 0 1 1
use contact_33  contact_33_1604
timestamp 1624857261
transform 1 0 22984 0 1 66781
box 0 0 1 1
use contact_33  contact_33_1606
timestamp 1624857261
transform 1 0 22984 0 1 66917
box 0 0 1 1
use contact_33  contact_33_4359
timestamp 1624857261
transform 1 0 23528 0 1 66917
box 0 0 1 1
use contact_33  contact_33_4594
timestamp 1624857261
transform 1 0 23528 0 1 66781
box 0 0 1 1
use contact_33  contact_33_5377
timestamp 1624857261
transform 1 0 1224 0 1 67597
box 0 0 1 1
use contact_13  contact_13_577
timestamp 1624857261
transform 1 0 1801 0 1 67203
box 0 0 1 1
use contact_19  contact_19_577
timestamp 1624857261
transform 1 0 1794 0 1 67212
box 0 0 1 1
use contact_14  contact_14_577
timestamp 1624857261
transform 1 0 1797 0 1 67211
box 0 0 1 1
use contact_13  contact_13_576
timestamp 1624857261
transform 1 0 1801 0 1 67539
box 0 0 1 1
use contact_19  contact_19_576
timestamp 1624857261
transform 1 0 1794 0 1 67548
box 0 0 1 1
use contact_14  contact_14_576
timestamp 1624857261
transform 1 0 1797 0 1 67547
box 0 0 1 1
use contact_7  contact_7_116
timestamp 1624857261
transform 1 0 1793 0 1 67543
box 0 0 1 1
use contact_13  contact_13_575
timestamp 1624857261
transform 1 0 1801 0 1 67875
box 0 0 1 1
use contact_19  contact_19_575
timestamp 1624857261
transform 1 0 1794 0 1 67884
box 0 0 1 1
use contact_14  contact_14_575
timestamp 1624857261
transform 1 0 1797 0 1 67883
box 0 0 1 1
use contact_13  contact_13_574
timestamp 1624857261
transform 1 0 1801 0 1 68211
box 0 0 1 1
use contact_19  contact_19_574
timestamp 1624857261
transform 1 0 1794 0 1 68220
box 0 0 1 1
use contact_14  contact_14_574
timestamp 1624857261
transform 1 0 1797 0 1 68219
box 0 0 1 1
use contact_33  contact_33_2102
timestamp 1624857261
transform 1 0 21896 0 1 67189
box 0 0 1 1
use contact_33  contact_33_2217
timestamp 1624857261
transform 1 0 21760 0 1 68005
box 0 0 1 1
use contact_33  contact_33_2218
timestamp 1624857261
transform 1 0 21760 0 1 67733
box 0 0 1 1
use contact_33  contact_33_2219
timestamp 1624857261
transform 1 0 21760 0 1 67325
box 0 0 1 1
use contact_33  contact_33_2220
timestamp 1624857261
transform 1 0 21760 0 1 67597
box 0 0 1 1
use contact_33  contact_33_1605
timestamp 1624857261
transform 1 0 22984 0 1 67189
box 0 0 1 1
use contact_33  contact_33_4730
timestamp 1624857261
transform 1 0 22576 0 1 67597
box 0 0 1 1
use contact_33  contact_33_4731
timestamp 1624857261
transform 1 0 22576 0 1 67325
box 0 0 1 1
use contact_33  contact_33_4734
timestamp 1624857261
transform 1 0 22576 0 1 68005
box 0 0 1 1
use contact_33  contact_33_4735
timestamp 1624857261
transform 1 0 22576 0 1 68277
box 0 0 1 1
use contact_33  contact_33_5062
timestamp 1624857261
transform 1 0 22168 0 1 68005
box 0 0 1 1
use contact_33  contact_33_5063
timestamp 1624857261
transform 1 0 22168 0 1 68277
box 0 0 1 1
use contact_33  contact_33_4358
timestamp 1624857261
transform 1 0 23528 0 1 67189
box 0 0 1 1
use contact_33  contact_33_1406
timestamp 1624857261
transform 1 0 28424 0 1 68277
box 0 0 1 1
use contact_33  contact_33_5312
timestamp 1624857261
transform 1 0 1224 0 1 69229
box 0 0 1 1
use contact_13  contact_13_573
timestamp 1624857261
transform 1 0 1801 0 1 68547
box 0 0 1 1
use contact_19  contact_19_573
timestamp 1624857261
transform 1 0 1794 0 1 68556
box 0 0 1 1
use contact_14  contact_14_573
timestamp 1624857261
transform 1 0 1797 0 1 68555
box 0 0 1 1
use contact_13  contact_13_572
timestamp 1624857261
transform 1 0 1801 0 1 68883
box 0 0 1 1
use contact_19  contact_19_572
timestamp 1624857261
transform 1 0 1794 0 1 68892
box 0 0 1 1
use contact_14  contact_14_572
timestamp 1624857261
transform 1 0 1797 0 1 68891
box 0 0 1 1
use contact_13  contact_13_571
timestamp 1624857261
transform 1 0 1801 0 1 69219
box 0 0 1 1
use contact_19  contact_19_571
timestamp 1624857261
transform 1 0 1794 0 1 69228
box 0 0 1 1
use contact_14  contact_14_571
timestamp 1624857261
transform 1 0 1797 0 1 69227
box 0 0 1 1
use contact_7  contact_7_115
timestamp 1624857261
transform 1 0 1793 0 1 69223
box 0 0 1 1
use contact_13  contact_13_570
timestamp 1624857261
transform 1 0 1801 0 1 69555
box 0 0 1 1
use contact_19  contact_19_570
timestamp 1624857261
transform 1 0 1794 0 1 69564
box 0 0 1 1
use contact_14  contact_14_570
timestamp 1624857261
transform 1 0 1797 0 1 69563
box 0 0 1 1
use contact_33  contact_33_2173
timestamp 1624857261
transform 1 0 21896 0 1 69501
box 0 0 1 1
use contact_33  contact_33_2174
timestamp 1624857261
transform 1 0 21896 0 1 69229
box 0 0 1 1
use contact_33  contact_33_2189
timestamp 1624857261
transform 1 0 21896 0 1 68821
box 0 0 1 1
use contact_33  contact_33_2190
timestamp 1624857261
transform 1 0 21896 0 1 68549
box 0 0 1 1
use contact_33  contact_33_1711
timestamp 1624857261
transform 1 0 23120 0 1 68413
box 0 0 1 1
use contact_33  contact_33_4711
timestamp 1624857261
transform 1 0 22576 0 1 68821
box 0 0 1 1
use contact_33  contact_33_1714
timestamp 1624857261
transform 1 0 23120 0 1 68821
box 0 0 1 1
use contact_33  contact_33_1712
timestamp 1624857261
transform 1 0 23120 0 1 68685
box 0 0 1 1
use contact_33  contact_33_5121
timestamp 1624857261
transform 1 0 22440 0 1 69229
box 0 0 1 1
use contact_33  contact_33_4710
timestamp 1624857261
transform 1 0 22576 0 1 69093
box 0 0 1 1
use contact_33  contact_33_1713
timestamp 1624857261
transform 1 0 23120 0 1 69093
box 0 0 1 1
use contact_33  contact_33_1701
timestamp 1624857261
transform 1 0 22984 0 1 69229
box 0 0 1 1
use contact_33  contact_33_5176
timestamp 1624857261
transform 1 0 22168 0 1 69637
box 0 0 1 1
use contact_33  contact_33_5120
timestamp 1624857261
transform 1 0 22440 0 1 69501
box 0 0 1 1
use contact_33  contact_33_4828
timestamp 1624857261
transform 1 0 22576 0 1 69637
box 0 0 1 1
use contact_33  contact_33_1702
timestamp 1624857261
transform 1 0 22984 0 1 69501
box 0 0 1 1
use contact_33  contact_33_1700
timestamp 1624857261
transform 1 0 22984 0 1 69637
box 0 0 1 1
use contact_33  contact_33_4458
timestamp 1624857261
transform 1 0 23528 0 1 68821
box 0 0 1 1
use contact_33  contact_33_4459
timestamp 1624857261
transform 1 0 23528 0 1 69093
box 0 0 1 1
use contact_33  contact_33_4461
timestamp 1624857261
transform 1 0 23392 0 1 69637
box 0 0 1 1
use contact_33  contact_33_4462
timestamp 1624857261
transform 1 0 23392 0 1 69229
box 0 0 1 1
use contact_33  contact_33_4463
timestamp 1624857261
transform 1 0 23392 0 1 69501
box 0 0 1 1
use contact_33  contact_33_4688
timestamp 1624857261
transform 1 0 23392 0 1 68685
box 0 0 1 1
use contact_33  contact_33_4689
timestamp 1624857261
transform 1 0 23392 0 1 68413
box 0 0 1 1
use contact_33  contact_33_1405
timestamp 1624857261
transform 1 0 28424 0 1 68685
box 0 0 1 1
use contact_33  contact_33_1409
timestamp 1624857261
transform 1 0 28288 0 1 68957
box 0 0 1 1
use contact_33  contact_33_1410
timestamp 1624857261
transform 1 0 28288 0 1 68685
box 0 0 1 1
use contact_33  contact_33_5324
timestamp 1624857261
transform 1 0 1224 0 1 70997
box 0 0 1 1
use contact_13  contact_13_569
timestamp 1624857261
transform 1 0 1801 0 1 69891
box 0 0 1 1
use contact_19  contact_19_569
timestamp 1624857261
transform 1 0 1794 0 1 69900
box 0 0 1 1
use contact_14  contact_14_569
timestamp 1624857261
transform 1 0 1797 0 1 69899
box 0 0 1 1
use contact_13  contact_13_568
timestamp 1624857261
transform 1 0 1801 0 1 70227
box 0 0 1 1
use contact_19  contact_19_568
timestamp 1624857261
transform 1 0 1794 0 1 70236
box 0 0 1 1
use contact_14  contact_14_568
timestamp 1624857261
transform 1 0 1797 0 1 70235
box 0 0 1 1
use contact_13  contact_13_567
timestamp 1624857261
transform 1 0 1801 0 1 70563
box 0 0 1 1
use contact_19  contact_19_567
timestamp 1624857261
transform 1 0 1794 0 1 70572
box 0 0 1 1
use contact_14  contact_14_567
timestamp 1624857261
transform 1 0 1797 0 1 70571
box 0 0 1 1
use contact_13  contact_13_566
timestamp 1624857261
transform 1 0 1801 0 1 70899
box 0 0 1 1
use contact_19  contact_19_566
timestamp 1624857261
transform 1 0 1794 0 1 70908
box 0 0 1 1
use contact_14  contact_14_566
timestamp 1624857261
transform 1 0 1797 0 1 70907
box 0 0 1 1
use contact_7  contact_7_114
timestamp 1624857261
transform 1 0 1793 0 1 70903
box 0 0 1 1
use contact_33  contact_33_1947
timestamp 1624857261
transform 1 0 21896 0 1 70045
box 0 0 1 1
use contact_33  contact_33_1948
timestamp 1624857261
transform 1 0 21896 0 1 70317
box 0 0 1 1
use contact_33  contact_33_2222
timestamp 1624857261
transform 1 0 21760 0 1 70861
box 0 0 1 1
use contact_33  contact_33_2223
timestamp 1624857261
transform 1 0 21896 0 1 70453
box 0 0 1 1
use contact_33  contact_33_2224
timestamp 1624857261
transform 1 0 21896 0 1 70725
box 0 0 1 1
use contact_33  contact_33_5177
timestamp 1624857261
transform 1 0 22168 0 1 69909
box 0 0 1 1
use contact_33  contact_33_4829
timestamp 1624857261
transform 1 0 22576 0 1 69909
box 0 0 1 1
use contact_33  contact_33_1699
timestamp 1624857261
transform 1 0 22984 0 1 69909
box 0 0 1 1
use contact_33  contact_33_5129
timestamp 1624857261
transform 1 0 22440 0 1 70317
box 0 0 1 1
use contact_33  contact_33_5128
timestamp 1624857261
transform 1 0 22440 0 1 70045
box 0 0 1 1
use contact_33  contact_33_1842
timestamp 1624857261
transform 1 0 23120 0 1 70317
box 0 0 1 1
use contact_33  contact_33_1841
timestamp 1624857261
transform 1 0 23120 0 1 70045
box 0 0 1 1
use contact_33  contact_33_4813
timestamp 1624857261
transform 1 0 22712 0 1 70725
box 0 0 1 1
use contact_33  contact_33_4812
timestamp 1624857261
transform 1 0 22712 0 1 70453
box 0 0 1 1
use contact_33  contact_33_1840
timestamp 1624857261
transform 1 0 23120 0 1 70453
box 0 0 1 1
use contact_33  contact_33_1839
timestamp 1624857261
transform 1 0 23120 0 1 70725
box 0 0 1 1
use contact_33  contact_33_5054
timestamp 1624857261
transform 1 0 22168 0 1 70861
box 0 0 1 1
use contact_33  contact_33_4811
timestamp 1624857261
transform 1 0 22576 0 1 70861
box 0 0 1 1
use contact_33  contact_33_1871
timestamp 1624857261
transform 1 0 22984 0 1 70861
box 0 0 1 1
use contact_33  contact_33_4368
timestamp 1624857261
transform 1 0 24208 0 1 70317
box 0 0 1 1
use contact_33  contact_33_4369
timestamp 1624857261
transform 1 0 24208 0 1 70045
box 0 0 1 1
use contact_33  contact_33_4370
timestamp 1624857261
transform 1 0 23528 0 1 70317
box 0 0 1 1
use contact_33  contact_33_4371
timestamp 1624857261
transform 1 0 23528 0 1 70045
box 0 0 1 1
use contact_33  contact_33_4460
timestamp 1624857261
transform 1 0 23392 0 1 69909
box 0 0 1 1
use contact_33  contact_33_4482
timestamp 1624857261
transform 1 0 23392 0 1 70453
box 0 0 1 1
use contact_33  contact_33_4483
timestamp 1624857261
transform 1 0 23392 0 1 70725
box 0 0 1 1
use contact_33  contact_33_4485
timestamp 1624857261
transform 1 0 23528 0 1 70861
box 0 0 1 1
use contact_13  contact_13_565
timestamp 1624857261
transform 1 0 1801 0 1 71235
box 0 0 1 1
use contact_19  contact_19_565
timestamp 1624857261
transform 1 0 1794 0 1 71244
box 0 0 1 1
use contact_14  contact_14_565
timestamp 1624857261
transform 1 0 1797 0 1 71243
box 0 0 1 1
use contact_13  contact_13_564
timestamp 1624857261
transform 1 0 1801 0 1 71571
box 0 0 1 1
use contact_19  contact_19_564
timestamp 1624857261
transform 1 0 1794 0 1 71580
box 0 0 1 1
use contact_14  contact_14_564
timestamp 1624857261
transform 1 0 1797 0 1 71579
box 0 0 1 1
use contact_13  contact_13_563
timestamp 1624857261
transform 1 0 1801 0 1 71907
box 0 0 1 1
use contact_19  contact_19_563
timestamp 1624857261
transform 1 0 1794 0 1 71916
box 0 0 1 1
use contact_14  contact_14_563
timestamp 1624857261
transform 1 0 1797 0 1 71915
box 0 0 1 1
use contact_13  contact_13_562
timestamp 1624857261
transform 1 0 1801 0 1 72243
box 0 0 1 1
use contact_19  contact_19_562
timestamp 1624857261
transform 1 0 1794 0 1 72252
box 0 0 1 1
use contact_14  contact_14_562
timestamp 1624857261
transform 1 0 1797 0 1 72251
box 0 0 1 1
use contact_33  contact_33_1973
timestamp 1624857261
transform 1 0 21896 0 1 71949
box 0 0 1 1
use contact_33  contact_33_1974
timestamp 1624857261
transform 1 0 21896 0 1 71677
box 0 0 1 1
use contact_33  contact_33_1975
timestamp 1624857261
transform 1 0 21896 0 1 71269
box 0 0 1 1
use contact_33  contact_33_1976
timestamp 1624857261
transform 1 0 21896 0 1 71541
box 0 0 1 1
use contact_33  contact_33_2121
timestamp 1624857261
transform 1 0 21760 0 1 72085
box 0 0 1 1
use contact_33  contact_33_2122
timestamp 1624857261
transform 1 0 21760 0 1 72357
box 0 0 1 1
use contact_33  contact_33_2221
timestamp 1624857261
transform 1 0 21760 0 1 71133
box 0 0 1 1
use contact_33  contact_33_5055
timestamp 1624857261
transform 1 0 22168 0 1 71133
box 0 0 1 1
use contact_33  contact_33_5053
timestamp 1624857261
transform 1 0 22440 0 1 71269
box 0 0 1 1
use contact_33  contact_33_4810
timestamp 1624857261
transform 1 0 22576 0 1 71133
box 0 0 1 1
use contact_33  contact_33_4726
timestamp 1624857261
transform 1 0 22712 0 1 71269
box 0 0 1 1
use contact_33  contact_33_1874
timestamp 1624857261
transform 1 0 22984 0 1 71269
box 0 0 1 1
use contact_33  contact_33_1872
timestamp 1624857261
transform 1 0 22984 0 1 71133
box 0 0 1 1
use contact_33  contact_33_5052
timestamp 1624857261
transform 1 0 22440 0 1 71541
box 0 0 1 1
use contact_33  contact_33_4727
timestamp 1624857261
transform 1 0 22712 0 1 71541
box 0 0 1 1
use contact_33  contact_33_1873
timestamp 1624857261
transform 1 0 22984 0 1 71541
box 0 0 1 1
use contact_33  contact_33_5011
timestamp 1624857261
transform 1 0 22168 0 1 72085
box 0 0 1 1
use contact_33  contact_33_4825
timestamp 1624857261
transform 1 0 22576 0 1 72085
box 0 0 1 1
use contact_33  contact_33_5010
timestamp 1624857261
transform 1 0 22168 0 1 72357
box 0 0 1 1
use contact_33  contact_33_4824
timestamp 1624857261
transform 1 0 22576 0 1 72357
box 0 0 1 1
use contact_33  contact_33_4406
timestamp 1624857261
transform 1 0 23528 0 1 71541
box 0 0 1 1
use contact_33  contact_33_4407
timestamp 1624857261
transform 1 0 23528 0 1 71269
box 0 0 1 1
use contact_33  contact_33_4484
timestamp 1624857261
transform 1 0 23528 0 1 71133
box 0 0 1 1
use contact_33  contact_33_1467
timestamp 1624857261
transform 1 0 28288 0 1 71813
box 0 0 1 1
use contact_33  contact_33_1468
timestamp 1624857261
transform 1 0 28288 0 1 72085
box 0 0 1 1
use contact_33  contact_33_1517
timestamp 1624857261
transform 1 0 28424 0 1 72221
box 0 0 1 1
use contact_33  contact_33_5355
timestamp 1624857261
transform 1 0 1224 0 1 72629
box 0 0 1 1
use contact_13  contact_13_561
timestamp 1624857261
transform 1 0 1801 0 1 72579
box 0 0 1 1
use contact_19  contact_19_561
timestamp 1624857261
transform 1 0 1794 0 1 72588
box 0 0 1 1
use contact_14  contact_14_561
timestamp 1624857261
transform 1 0 1797 0 1 72587
box 0 0 1 1
use contact_7  contact_7_113
timestamp 1624857261
transform 1 0 1793 0 1 72583
box 0 0 1 1
use contact_13  contact_13_560
timestamp 1624857261
transform 1 0 1801 0 1 72915
box 0 0 1 1
use contact_19  contact_19_560
timestamp 1624857261
transform 1 0 1794 0 1 72924
box 0 0 1 1
use contact_14  contact_14_560
timestamp 1624857261
transform 1 0 1797 0 1 72923
box 0 0 1 1
use contact_13  contact_13_559
timestamp 1624857261
transform 1 0 1801 0 1 73251
box 0 0 1 1
use contact_19  contact_19_559
timestamp 1624857261
transform 1 0 1794 0 1 73260
box 0 0 1 1
use contact_14  contact_14_559
timestamp 1624857261
transform 1 0 1797 0 1 73259
box 0 0 1 1
use contact_13  contact_13_558
timestamp 1624857261
transform 1 0 1801 0 1 73587
box 0 0 1 1
use contact_19  contact_19_558
timestamp 1624857261
transform 1 0 1794 0 1 73596
box 0 0 1 1
use contact_14  contact_14_558
timestamp 1624857261
transform 1 0 1797 0 1 73595
box 0 0 1 1
use contact_33  contact_33_2123
timestamp 1624857261
transform 1 0 21896 0 1 72765
box 0 0 1 1
use contact_33  contact_33_2124
timestamp 1624857261
transform 1 0 21896 0 1 72493
box 0 0 1 1
use contact_33  contact_33_2179
timestamp 1624857261
transform 1 0 21896 0 1 73173
box 0 0 1 1
use contact_33  contact_33_2180
timestamp 1624857261
transform 1 0 21896 0 1 73445
box 0 0 1 1
use contact_33  contact_33_4961
timestamp 1624857261
transform 1 0 22440 0 1 72765
box 0 0 1 1
use contact_33  contact_33_1698
timestamp 1624857261
transform 1 0 22984 0 1 72765
box 0 0 1 1
use contact_33  contact_33_5035
timestamp 1624857261
transform 1 0 22168 0 1 73173
box 0 0 1 1
use contact_33  contact_33_4960
timestamp 1624857261
transform 1 0 22440 0 1 73037
box 0 0 1 1
use contact_33  contact_33_1697
timestamp 1624857261
transform 1 0 22984 0 1 73037
box 0 0 1 1
use contact_33  contact_33_1627
timestamp 1624857261
transform 1 0 22984 0 1 73173
box 0 0 1 1
use contact_33  contact_33_5034
timestamp 1624857261
transform 1 0 22168 0 1 73445
box 0 0 1 1
use contact_33  contact_33_4851
timestamp 1624857261
transform 1 0 22712 0 1 73581
box 0 0 1 1
use contact_33  contact_33_1657
timestamp 1624857261
transform 1 0 22984 0 1 73581
box 0 0 1 1
use contact_33  contact_33_1628
timestamp 1624857261
transform 1 0 22984 0 1 73445
box 0 0 1 1
use contact_33  contact_33_4528
timestamp 1624857261
transform 1 0 23528 0 1 73173
box 0 0 1 1
use contact_33  contact_33_4529
timestamp 1624857261
transform 1 0 23528 0 1 73445
box 0 0 1 1
use contact_33  contact_33_4554
timestamp 1624857261
transform 1 0 23392 0 1 73037
box 0 0 1 1
use contact_33  contact_33_4555
timestamp 1624857261
transform 1 0 23392 0 1 72765
box 0 0 1 1
use contact_33  contact_33_4564
timestamp 1624857261
transform 1 0 23392 0 1 73581
box 0 0 1 1
use contact_33  contact_33_1515
timestamp 1624857261
transform 1 0 28424 0 1 72901
box 0 0 1 1
use contact_33  contact_33_1516
timestamp 1624857261
transform 1 0 28424 0 1 72629
box 0 0 1 1
use contact_33  contact_33_1518
timestamp 1624857261
transform 1 0 28424 0 1 72493
box 0 0 1 1
use contact_33  contact_33_5343
timestamp 1624857261
transform 1 0 1224 0 1 74125
box 0 0 1 1
use contact_13  contact_13_557
timestamp 1624857261
transform 1 0 1801 0 1 73923
box 0 0 1 1
use contact_19  contact_19_557
timestamp 1624857261
transform 1 0 1794 0 1 73932
box 0 0 1 1
use contact_14  contact_14_557
timestamp 1624857261
transform 1 0 1797 0 1 73931
box 0 0 1 1
use contact_13  contact_13_556
timestamp 1624857261
transform 1 0 1801 0 1 74259
box 0 0 1 1
use contact_19  contact_19_556
timestamp 1624857261
transform 1 0 1794 0 1 74268
box 0 0 1 1
use contact_14  contact_14_556
timestamp 1624857261
transform 1 0 1797 0 1 74267
box 0 0 1 1
use contact_7  contact_7_112
timestamp 1624857261
transform 1 0 1793 0 1 74263
box 0 0 1 1
use contact_13  contact_13_555
timestamp 1624857261
transform 1 0 1801 0 1 74595
box 0 0 1 1
use contact_19  contact_19_555
timestamp 1624857261
transform 1 0 1794 0 1 74604
box 0 0 1 1
use contact_14  contact_14_555
timestamp 1624857261
transform 1 0 1797 0 1 74603
box 0 0 1 1
use contact_13  contact_13_554
timestamp 1624857261
transform 1 0 1801 0 1 74931
box 0 0 1 1
use contact_19  contact_19_554
timestamp 1624857261
transform 1 0 1794 0 1 74940
box 0 0 1 1
use contact_14  contact_14_554
timestamp 1624857261
transform 1 0 1797 0 1 74939
box 0 0 1 1
use contact_33  contact_33_2033
timestamp 1624857261
transform 1 0 21896 0 1 74805
box 0 0 1 1
use contact_33  contact_33_2034
timestamp 1624857261
transform 1 0 21896 0 1 75077
box 0 0 1 1
use contact_33  contact_33_2259
timestamp 1624857261
transform 1 0 21760 0 1 74669
box 0 0 1 1
use contact_33  contact_33_2260
timestamp 1624857261
transform 1 0 21760 0 1 74397
box 0 0 1 1
use contact_33  contact_33_2261
timestamp 1624857261
transform 1 0 21760 0 1 73989
box 0 0 1 1
use contact_33  contact_33_2262
timestamp 1624857261
transform 1 0 21760 0 1 74261
box 0 0 1 1
use contact_33  contact_33_4836
timestamp 1624857261
transform 1 0 22576 0 1 73989
box 0 0 1 1
use contact_33  contact_33_4850
timestamp 1624857261
transform 1 0 22712 0 1 73853
box 0 0 1 1
use contact_33  contact_33_1658
timestamp 1624857261
transform 1 0 22984 0 1 73853
box 0 0 1 1
use contact_33  contact_33_1656
timestamp 1624857261
transform 1 0 22984 0 1 73989
box 0 0 1 1
use contact_33  contact_33_5101
timestamp 1624857261
transform 1 0 22168 0 1 74397
box 0 0 1 1
use contact_33  contact_33_5042
timestamp 1624857261
transform 1 0 22440 0 1 74397
box 0 0 1 1
use contact_33  contact_33_4837
timestamp 1624857261
transform 1 0 22576 0 1 74261
box 0 0 1 1
use contact_33  contact_33_1655
timestamp 1624857261
transform 1 0 22984 0 1 74261
box 0 0 1 1
use contact_33  contact_33_1612
timestamp 1624857261
transform 1 0 23120 0 1 74397
box 0 0 1 1
use contact_33  contact_33_5100
timestamp 1624857261
transform 1 0 22168 0 1 74669
box 0 0 1 1
use contact_33  contact_33_5043
timestamp 1624857261
transform 1 0 22440 0 1 74669
box 0 0 1 1
use contact_33  contact_33_1611
timestamp 1624857261
transform 1 0 23120 0 1 74669
box 0 0 1 1
use contact_33  contact_33_4783
timestamp 1624857261
transform 1 0 22712 0 1 74805
box 0 0 1 1
use contact_33  contact_33_4782
timestamp 1624857261
transform 1 0 22712 0 1 75077
box 0 0 1 1
use contact_33  contact_33_1594
timestamp 1624857261
transform 1 0 23120 0 1 74805
box 0 0 1 1
use contact_33  contact_33_1593
timestamp 1624857261
transform 1 0 23120 0 1 75077
box 0 0 1 1
use contact_33  contact_33_4548
timestamp 1624857261
transform 1 0 23392 0 1 74397
box 0 0 1 1
use contact_33  contact_33_4549
timestamp 1624857261
transform 1 0 23392 0 1 74669
box 0 0 1 1
use contact_33  contact_33_4550
timestamp 1624857261
transform 1 0 23392 0 1 75077
box 0 0 1 1
use contact_33  contact_33_4551
timestamp 1624857261
transform 1 0 23392 0 1 74805
box 0 0 1 1
use contact_33  contact_33_4562
timestamp 1624857261
transform 1 0 23392 0 1 74261
box 0 0 1 1
use contact_33  contact_33_4563
timestamp 1624857261
transform 1 0 23392 0 1 73989
box 0 0 1 1
use contact_33  contact_33_4565
timestamp 1624857261
transform 1 0 23392 0 1 73853
box 0 0 1 1
use contact_33  contact_33_1464
timestamp 1624857261
transform 1 0 28424 0 1 74941
box 0 0 1 1
use contact_33  contact_33_5301
timestamp 1624857261
transform 1 0 1224 0 1 75893
box 0 0 1 1
use contact_13  contact_13_553
timestamp 1624857261
transform 1 0 1801 0 1 75267
box 0 0 1 1
use contact_19  contact_19_553
timestamp 1624857261
transform 1 0 1794 0 1 75276
box 0 0 1 1
use contact_14  contact_14_553
timestamp 1624857261
transform 1 0 1797 0 1 75275
box 0 0 1 1
use contact_13  contact_13_552
timestamp 1624857261
transform 1 0 1801 0 1 75603
box 0 0 1 1
use contact_19  contact_19_552
timestamp 1624857261
transform 1 0 1794 0 1 75612
box 0 0 1 1
use contact_14  contact_14_552
timestamp 1624857261
transform 1 0 1797 0 1 75611
box 0 0 1 1
use contact_13  contact_13_551
timestamp 1624857261
transform 1 0 1801 0 1 75939
box 0 0 1 1
use contact_19  contact_19_551
timestamp 1624857261
transform 1 0 1794 0 1 75948
box 0 0 1 1
use contact_14  contact_14_551
timestamp 1624857261
transform 1 0 1797 0 1 75947
box 0 0 1 1
use contact_7  contact_7_111
timestamp 1624857261
transform 1 0 1793 0 1 75943
box 0 0 1 1
use contact_13  contact_13_550
timestamp 1624857261
transform 1 0 1801 0 1 76275
box 0 0 1 1
use contact_19  contact_19_550
timestamp 1624857261
transform 1 0 1794 0 1 76284
box 0 0 1 1
use contact_14  contact_14_550
timestamp 1624857261
transform 1 0 1797 0 1 76283
box 0 0 1 1
use contact_33  contact_33_2054
timestamp 1624857261
transform 1 0 21760 0 1 76437
box 0 0 1 1
use contact_33  contact_33_2061
timestamp 1624857261
transform 1 0 21896 0 1 76301
box 0 0 1 1
use contact_33  contact_33_2062
timestamp 1624857261
transform 1 0 21896 0 1 76029
box 0 0 1 1
use contact_33  contact_33_2063
timestamp 1624857261
transform 1 0 21760 0 1 75213
box 0 0 1 1
use contact_33  contact_33_2064
timestamp 1624857261
transform 1 0 21760 0 1 75485
box 0 0 1 1
use contact_33  contact_33_2065
timestamp 1624857261
transform 1 0 21760 0 1 75893
box 0 0 1 1
use contact_33  contact_33_2066
timestamp 1624857261
transform 1 0 21760 0 1 75621
box 0 0 1 1
use contact_33  contact_33_1745
timestamp 1624857261
transform 1 0 22984 0 1 75213
box 0 0 1 1
use contact_33  contact_33_1746
timestamp 1624857261
transform 1 0 22984 0 1 75485
box 0 0 1 1
use contact_33  contact_33_4764
timestamp 1624857261
transform 1 0 22576 0 1 76029
box 0 0 1 1
use contact_33  contact_33_4765
timestamp 1624857261
transform 1 0 22576 0 1 76301
box 0 0 1 1
use contact_33  contact_33_4992
timestamp 1624857261
transform 1 0 22440 0 1 75485
box 0 0 1 1
use contact_33  contact_33_4993
timestamp 1624857261
transform 1 0 22440 0 1 75213
box 0 0 1 1
use contact_33  contact_33_4510
timestamp 1624857261
transform 1 0 23528 0 1 75485
box 0 0 1 1
use contact_33  contact_33_4511
timestamp 1624857261
transform 1 0 23528 0 1 75213
box 0 0 1 1
use contact_33  contact_33_1411
timestamp 1624857261
transform 1 0 28560 0 1 75757
box 0 0 1 1
use contact_33  contact_33_1412
timestamp 1624857261
transform 1 0 28560 0 1 76029
box 0 0 1 1
use contact_33  contact_33_1413
timestamp 1624857261
transform 1 0 28288 0 1 76437
box 0 0 1 1
use contact_33  contact_33_1414
timestamp 1624857261
transform 1 0 28288 0 1 76165
box 0 0 1 1
use contact_33  contact_33_1463
timestamp 1624857261
transform 1 0 28424 0 1 75213
box 0 0 1 1
use contact_33  contact_33_5360
timestamp 1624857261
transform 1 0 1224 0 1 77661
box 0 0 1 1
use contact_13  contact_13_549
timestamp 1624857261
transform 1 0 1801 0 1 76611
box 0 0 1 1
use contact_19  contact_19_549
timestamp 1624857261
transform 1 0 1794 0 1 76620
box 0 0 1 1
use contact_14  contact_14_549
timestamp 1624857261
transform 1 0 1797 0 1 76619
box 0 0 1 1
use contact_13  contact_13_548
timestamp 1624857261
transform 1 0 1801 0 1 76947
box 0 0 1 1
use contact_19  contact_19_548
timestamp 1624857261
transform 1 0 1794 0 1 76956
box 0 0 1 1
use contact_14  contact_14_548
timestamp 1624857261
transform 1 0 1797 0 1 76955
box 0 0 1 1
use contact_13  contact_13_547
timestamp 1624857261
transform 1 0 1801 0 1 77283
box 0 0 1 1
use contact_19  contact_19_547
timestamp 1624857261
transform 1 0 1794 0 1 77292
box 0 0 1 1
use contact_14  contact_14_547
timestamp 1624857261
transform 1 0 1797 0 1 77291
box 0 0 1 1
use contact_13  contact_13_546
timestamp 1624857261
transform 1 0 1801 0 1 77619
box 0 0 1 1
use contact_19  contact_19_546
timestamp 1624857261
transform 1 0 1794 0 1 77628
box 0 0 1 1
use contact_14  contact_14_546
timestamp 1624857261
transform 1 0 1797 0 1 77627
box 0 0 1 1
use contact_7  contact_7_110
timestamp 1624857261
transform 1 0 1793 0 1 77623
box 0 0 1 1
use contact_33  contact_33_2053
timestamp 1624857261
transform 1 0 21760 0 1 76709
box 0 0 1 1
use contact_33  contact_33_4839
timestamp 1624857261
transform 1 0 22576 0 1 76709
box 0 0 1 1
use contact_33  contact_33_1862
timestamp 1624857261
transform 1 0 22984 0 1 76709
box 0 0 1 1
use contact_33  contact_33_4838
timestamp 1624857261
transform 1 0 22576 0 1 76981
box 0 0 1 1
use contact_33  contact_33_1861
timestamp 1624857261
transform 1 0 22984 0 1 76981
box 0 0 1 1
use contact_33  contact_33_1822
timestamp 1624857261
transform 1 0 22984 0 1 77117
box 0 0 1 1
use contact_33  contact_33_5048
timestamp 1624857261
transform 1 0 22440 0 1 77525
box 0 0 1 1
use contact_33  contact_33_1821
timestamp 1624857261
transform 1 0 22984 0 1 77389
box 0 0 1 1
use contact_33  contact_33_1654
timestamp 1624857261
transform 1 0 23120 0 1 77525
box 0 0 1 1
use contact_33  contact_33_5049
timestamp 1624857261
transform 1 0 22440 0 1 77797
box 0 0 1 1
use contact_33  contact_33_1653
timestamp 1624857261
transform 1 0 23120 0 1 77797
box 0 0 1 1
use contact_33  contact_33_4418
timestamp 1624857261
transform 1 0 23528 0 1 77797
box 0 0 1 1
use contact_33  contact_33_4419
timestamp 1624857261
transform 1 0 23528 0 1 77525
box 0 0 1 1
use contact_33  contact_33_4436
timestamp 1624857261
transform 1 0 23392 0 1 77389
box 0 0 1 1
use contact_33  contact_33_4437
timestamp 1624857261
transform 1 0 23392 0 1 77117
box 0 0 1 1
use contact_33  contact_33_4448
timestamp 1624857261
transform 1 0 23528 0 1 76981
box 0 0 1 1
use contact_33  contact_33_4449
timestamp 1624857261
transform 1 0 23528 0 1 76709
box 0 0 1 1
use contact_33  contact_33_1507
timestamp 1624857261
transform 1 0 28288 0 1 77661
box 0 0 1 1
use contact_33  contact_33_1508
timestamp 1624857261
transform 1 0 28288 0 1 77389
box 0 0 1 1
use contact_13  contact_13_545
timestamp 1624857261
transform 1 0 1801 0 1 77955
box 0 0 1 1
use contact_19  contact_19_545
timestamp 1624857261
transform 1 0 1794 0 1 77964
box 0 0 1 1
use contact_14  contact_14_545
timestamp 1624857261
transform 1 0 1797 0 1 77963
box 0 0 1 1
use contact_13  contact_13_544
timestamp 1624857261
transform 1 0 1801 0 1 78291
box 0 0 1 1
use contact_19  contact_19_544
timestamp 1624857261
transform 1 0 1794 0 1 78300
box 0 0 1 1
use contact_14  contact_14_544
timestamp 1624857261
transform 1 0 1797 0 1 78299
box 0 0 1 1
use contact_13  contact_13_543
timestamp 1624857261
transform 1 0 1801 0 1 78627
box 0 0 1 1
use contact_13  contact_13_542
timestamp 1624857261
transform 1 0 1801 0 1 78963
box 0 0 1 1
use contact_19  contact_19_543
timestamp 1624857261
transform 1 0 1794 0 1 78636
box 0 0 1 1
use contact_19  contact_19_542
timestamp 1624857261
transform 1 0 1794 0 1 78972
box 0 0 1 1
use contact_14  contact_14_543
timestamp 1624857261
transform 1 0 1797 0 1 78635
box 0 0 1 1
use contact_14  contact_14_542
timestamp 1624857261
transform 1 0 1797 0 1 78971
box 0 0 1 1
use contact_33  contact_33_2025
timestamp 1624857261
transform 1 0 21760 0 1 79021
box 0 0 1 1
use contact_33  contact_33_2026
timestamp 1624857261
transform 1 0 21760 0 1 78749
box 0 0 1 1
use contact_33  contact_33_2233
timestamp 1624857261
transform 1 0 21896 0 1 79157
box 0 0 1 1
use contact_33  contact_33_2239
timestamp 1624857261
transform 1 0 21896 0 1 78613
box 0 0 1 1
use contact_33  contact_33_2240
timestamp 1624857261
transform 1 0 21896 0 1 78341
box 0 0 1 1
use contact_33  contact_33_2241
timestamp 1624857261
transform 1 0 21896 0 1 77933
box 0 0 1 1
use contact_33  contact_33_2242
timestamp 1624857261
transform 1 0 21896 0 1 78205
box 0 0 1 1
use contact_33  contact_33_5084
timestamp 1624857261
transform 1 0 22304 0 1 77933
box 0 0 1 1
use contact_33  contact_33_1663
timestamp 1624857261
transform 1 0 22984 0 1 77933
box 0 0 1 1
use contact_33  contact_33_5085
timestamp 1624857261
transform 1 0 22304 0 1 78205
box 0 0 1 1
use contact_33  contact_33_5083
timestamp 1624857261
transform 1 0 22304 0 1 78341
box 0 0 1 1
use contact_33  contact_33_4774
timestamp 1624857261
transform 1 0 22576 0 1 78341
box 0 0 1 1
use contact_33  contact_33_1664
timestamp 1624857261
transform 1 0 22984 0 1 78205
box 0 0 1 1
use contact_33  contact_33_1662
timestamp 1624857261
transform 1 0 22984 0 1 78341
box 0 0 1 1
use contact_33  contact_33_5082
timestamp 1624857261
transform 1 0 22304 0 1 78613
box 0 0 1 1
use contact_33  contact_33_4775
timestamp 1624857261
transform 1 0 22576 0 1 78613
box 0 0 1 1
use contact_33  contact_33_1889
timestamp 1624857261
transform 1 0 23120 0 1 78749
box 0 0 1 1
use contact_33  contact_33_1661
timestamp 1624857261
transform 1 0 22984 0 1 78613
box 0 0 1 1
use contact_33  contact_33_4897
timestamp 1624857261
transform 1 0 22712 0 1 79157
box 0 0 1 1
use contact_33  contact_33_1892
timestamp 1624857261
transform 1 0 23120 0 1 79157
box 0 0 1 1
use contact_33  contact_33_1890
timestamp 1624857261
transform 1 0 23120 0 1 79021
box 0 0 1 1
use contact_33  contact_33_4632
timestamp 1624857261
transform 1 0 23392 0 1 78749
box 0 0 1 1
use contact_33  contact_33_4633
timestamp 1624857261
transform 1 0 23392 0 1 79021
box 0 0 1 1
use contact_33  contact_33_4635
timestamp 1624857261
transform 1 0 23392 0 1 79157
box 0 0 1 1
use contact_33  contact_33_4690
timestamp 1624857261
transform 1 0 23392 0 1 77933
box 0 0 1 1
use contact_33  contact_33_4691
timestamp 1624857261
transform 1 0 23392 0 1 78205
box 0 0 1 1
use contact_33  contact_33_4692
timestamp 1624857261
transform 1 0 23392 0 1 78613
box 0 0 1 1
use contact_33  contact_33_4693
timestamp 1624857261
transform 1 0 23392 0 1 78341
box 0 0 1 1
use contact_33  contact_33_1433
timestamp 1624857261
transform 1 0 28288 0 1 79157
box 0 0 1 1
use contact_33  contact_33_1434
timestamp 1624857261
transform 1 0 28288 0 1 78885
box 0 0 1 1
use contact_33  contact_33_5300
timestamp 1624857261
transform 1 0 1224 0 1 79429
box 0 0 1 1
use contact_13  contact_13_541
timestamp 1624857261
transform 1 0 1801 0 1 79299
box 0 0 1 1
use contact_19  contact_19_541
timestamp 1624857261
transform 1 0 1794 0 1 79308
box 0 0 1 1
use contact_14  contact_14_541
timestamp 1624857261
transform 1 0 1797 0 1 79307
box 0 0 1 1
use contact_7  contact_7_109
timestamp 1624857261
transform 1 0 1793 0 1 79303
box 0 0 1 1
use contact_13  contact_13_540
timestamp 1624857261
transform 1 0 1801 0 1 79635
box 0 0 1 1
use contact_19  contact_19_540
timestamp 1624857261
transform 1 0 1794 0 1 79644
box 0 0 1 1
use contact_14  contact_14_540
timestamp 1624857261
transform 1 0 1797 0 1 79643
box 0 0 1 1
use contact_13  contact_13_539
timestamp 1624857261
transform 1 0 1801 0 1 79971
box 0 0 1 1
use contact_13  contact_13_538
timestamp 1624857261
transform 1 0 1801 0 1 80307
box 0 0 1 1
use contact_19  contact_19_539
timestamp 1624857261
transform 1 0 1794 0 1 79980
box 0 0 1 1
use contact_19  contact_19_538
timestamp 1624857261
transform 1 0 1794 0 1 80316
box 0 0 1 1
use contact_14  contact_14_539
timestamp 1624857261
transform 1 0 1797 0 1 79979
box 0 0 1 1
use contact_14  contact_14_538
timestamp 1624857261
transform 1 0 1797 0 1 80315
box 0 0 1 1
use contact_33  contact_33_2183
timestamp 1624857261
transform 1 0 21896 0 1 79973
box 0 0 1 1
use contact_33  contact_33_2184
timestamp 1624857261
transform 1 0 21896 0 1 80245
box 0 0 1 1
use contact_33  contact_33_2186
timestamp 1624857261
transform 1 0 21896 0 1 80381
box 0 0 1 1
use contact_33  contact_33_2231
timestamp 1624857261
transform 1 0 21760 0 1 79837
box 0 0 1 1
use contact_33  contact_33_2232
timestamp 1624857261
transform 1 0 21760 0 1 79565
box 0 0 1 1
use contact_33  contact_33_2234
timestamp 1624857261
transform 1 0 21896 0 1 79429
box 0 0 1 1
use contact_33  contact_33_1787
timestamp 1624857261
transform 1 0 22984 0 1 79565
box 0 0 1 1
use contact_33  contact_33_1788
timestamp 1624857261
transform 1 0 22984 0 1 79837
box 0 0 1 1
use contact_33  contact_33_1891
timestamp 1624857261
transform 1 0 23120 0 1 79429
box 0 0 1 1
use contact_33  contact_33_4714
timestamp 1624857261
transform 1 0 22712 0 1 79973
box 0 0 1 1
use contact_33  contact_33_4715
timestamp 1624857261
transform 1 0 22712 0 1 80245
box 0 0 1 1
use contact_33  contact_33_4896
timestamp 1624857261
transform 1 0 22712 0 1 79429
box 0 0 1 1
use contact_33  contact_33_4976
timestamp 1624857261
transform 1 0 22440 0 1 80517
box 0 0 1 1
use contact_33  contact_33_4977
timestamp 1624857261
transform 1 0 22440 0 1 80245
box 0 0 1 1
use contact_33  contact_33_4466
timestamp 1624857261
transform 1 0 23528 0 1 79837
box 0 0 1 1
use contact_33  contact_33_4467
timestamp 1624857261
transform 1 0 23528 0 1 79565
box 0 0 1 1
use contact_33  contact_33_4634
timestamp 1624857261
transform 1 0 23392 0 1 79429
box 0 0 1 1
use contact_33  contact_33_1377
timestamp 1624857261
transform 1 0 28560 0 1 80517
box 0 0 1 1
use contact_33  contact_33_1429
timestamp 1624857261
transform 1 0 28288 0 1 80381
box 0 0 1 1
use contact_33  contact_33_1430
timestamp 1624857261
transform 1 0 28288 0 1 80109
box 0 0 1 1
use contact_33  contact_33_5297
timestamp 1624857261
transform 1 0 1224 0 1 81061
box 0 0 1 1
use contact_13  contact_13_537
timestamp 1624857261
transform 1 0 1801 0 1 80643
box 0 0 1 1
use contact_19  contact_19_537
timestamp 1624857261
transform 1 0 1794 0 1 80652
box 0 0 1 1
use contact_14  contact_14_537
timestamp 1624857261
transform 1 0 1797 0 1 80651
box 0 0 1 1
use contact_13  contact_13_536
timestamp 1624857261
transform 1 0 1801 0 1 80979
box 0 0 1 1
use contact_19  contact_19_536
timestamp 1624857261
transform 1 0 1794 0 1 80988
box 0 0 1 1
use contact_14  contact_14_536
timestamp 1624857261
transform 1 0 1797 0 1 80987
box 0 0 1 1
use contact_7  contact_7_108
timestamp 1624857261
transform 1 0 1793 0 1 80983
box 0 0 1 1
use contact_13  contact_13_535
timestamp 1624857261
transform 1 0 1801 0 1 81315
box 0 0 1 1
use contact_13  contact_13_534
timestamp 1624857261
transform 1 0 1801 0 1 81651
box 0 0 1 1
use contact_19  contact_19_535
timestamp 1624857261
transform 1 0 1794 0 1 81324
box 0 0 1 1
use contact_19  contact_19_534
timestamp 1624857261
transform 1 0 1794 0 1 81660
box 0 0 1 1
use contact_14  contact_14_535
timestamp 1624857261
transform 1 0 1797 0 1 81323
box 0 0 1 1
use contact_14  contact_14_534
timestamp 1624857261
transform 1 0 1797 0 1 81659
box 0 0 1 1
use contact_33  contact_33_2185
timestamp 1624857261
transform 1 0 21896 0 1 80653
box 0 0 1 1
use contact_33  contact_33_2227
timestamp 1624857261
transform 1 0 21760 0 1 81877
box 0 0 1 1
use contact_33  contact_33_5099
timestamp 1624857261
transform 1 0 22168 0 1 80653
box 0 0 1 1
use contact_33  contact_33_5098
timestamp 1624857261
transform 1 0 22168 0 1 80925
box 0 0 1 1
use contact_33  contact_33_1838
timestamp 1624857261
transform 1 0 22984 0 1 81061
box 0 0 1 1
use contact_33  contact_33_5105
timestamp 1624857261
transform 1 0 22304 0 1 81469
box 0 0 1 1
use contact_33  contact_33_4788
timestamp 1624857261
transform 1 0 22576 0 1 81469
box 0 0 1 1
use contact_33  contact_33_1837
timestamp 1624857261
transform 1 0 22984 0 1 81333
box 0 0 1 1
use contact_33  contact_33_1833
timestamp 1624857261
transform 1 0 23120 0 1 81469
box 0 0 1 1
use contact_33  contact_33_5104
timestamp 1624857261
transform 1 0 22304 0 1 81741
box 0 0 1 1
use contact_33  contact_33_4789
timestamp 1624857261
transform 1 0 22576 0 1 81741
box 0 0 1 1
use contact_33  contact_33_4787
timestamp 1624857261
transform 1 0 22576 0 1 81877
box 0 0 1 1
use contact_33  contact_33_1836
timestamp 1624857261
transform 1 0 23120 0 1 81877
box 0 0 1 1
use contact_33  contact_33_1834
timestamp 1624857261
transform 1 0 23120 0 1 81741
box 0 0 1 1
use contact_33  contact_33_4402
timestamp 1624857261
transform 1 0 23528 0 1 81333
box 0 0 1 1
use contact_33  contact_33_4403
timestamp 1624857261
transform 1 0 23528 0 1 81061
box 0 0 1 1
use contact_33  contact_33_4473
timestamp 1624857261
transform 1 0 23528 0 1 81877
box 0 0 1 1
use contact_33  contact_33_4474
timestamp 1624857261
transform 1 0 23528 0 1 81469
box 0 0 1 1
use contact_33  contact_33_4475
timestamp 1624857261
transform 1 0 23528 0 1 81741
box 0 0 1 1
use contact_33  contact_33_1378
timestamp 1624857261
transform 1 0 28560 0 1 80789
box 0 0 1 1
use contact_33  contact_33_1453
timestamp 1624857261
transform 1 0 28288 0 1 81061
box 0 0 1 1
use contact_33  contact_33_1454
timestamp 1624857261
transform 1 0 28288 0 1 80789
box 0 0 1 1
use contact_33  contact_33_5304
timestamp 1624857261
transform 1 0 1224 0 1 82693
box 0 0 1 1
use contact_13  contact_13_533
timestamp 1624857261
transform 1 0 1801 0 1 81987
box 0 0 1 1
use contact_19  contact_19_533
timestamp 1624857261
transform 1 0 1794 0 1 81996
box 0 0 1 1
use contact_14  contact_14_533
timestamp 1624857261
transform 1 0 1797 0 1 81995
box 0 0 1 1
use contact_13  contact_13_532
timestamp 1624857261
transform 1 0 1801 0 1 82323
box 0 0 1 1
use contact_13  contact_13_531
timestamp 1624857261
transform 1 0 1801 0 1 82659
box 0 0 1 1
use contact_19  contact_19_532
timestamp 1624857261
transform 1 0 1794 0 1 82332
box 0 0 1 1
use contact_14  contact_14_532
timestamp 1624857261
transform 1 0 1797 0 1 82331
box 0 0 1 1
use contact_13  contact_13_530
timestamp 1624857261
transform 1 0 1801 0 1 82995
box 0 0 1 1
use contact_19  contact_19_531
timestamp 1624857261
transform 1 0 1794 0 1 82668
box 0 0 1 1
use contact_19  contact_19_530
timestamp 1624857261
transform 1 0 1794 0 1 83004
box 0 0 1 1
use contact_14  contact_14_531
timestamp 1624857261
transform 1 0 1797 0 1 82667
box 0 0 1 1
use contact_14  contact_14_530
timestamp 1624857261
transform 1 0 1797 0 1 83003
box 0 0 1 1
use contact_7  contact_7_107
timestamp 1624857261
transform 1 0 1793 0 1 82663
box 0 0 1 1
use contact_33  contact_33_2110
timestamp 1624857261
transform 1 0 21760 0 1 83101
box 0 0 1 1
use contact_33  contact_33_2111
timestamp 1624857261
transform 1 0 21760 0 1 82693
box 0 0 1 1
use contact_33  contact_33_2112
timestamp 1624857261
transform 1 0 21760 0 1 82965
box 0 0 1 1
use contact_33  contact_33_2228
timestamp 1624857261
transform 1 0 21760 0 1 82149
box 0 0 1 1
use contact_33  contact_33_2229
timestamp 1624857261
transform 1 0 21896 0 1 82557
box 0 0 1 1
use contact_33  contact_33_2230
timestamp 1624857261
transform 1 0 21896 0 1 82285
box 0 0 1 1
use contact_33  contact_33_4786
timestamp 1624857261
transform 1 0 22576 0 1 82149
box 0 0 1 1
use contact_33  contact_33_1835
timestamp 1624857261
transform 1 0 23120 0 1 82149
box 0 0 1 1
use contact_33  contact_33_4945
timestamp 1624857261
transform 1 0 22440 0 1 82285
box 0 0 1 1
use contact_33  contact_33_4944
timestamp 1624857261
transform 1 0 22440 0 1 82557
box 0 0 1 1
use contact_33  contact_33_1774
timestamp 1624857261
transform 1 0 23120 0 1 82285
box 0 0 1 1
use contact_33  contact_33_1773
timestamp 1624857261
transform 1 0 23120 0 1 82557
box 0 0 1 1
use contact_33  contact_33_5031
timestamp 1624857261
transform 1 0 22168 0 1 82965
box 0 0 1 1
use contact_33  contact_33_5030
timestamp 1624857261
transform 1 0 22168 0 1 82693
box 0 0 1 1
use contact_33  contact_33_4881
timestamp 1624857261
transform 1 0 22576 0 1 82965
box 0 0 1 1
use contact_33  contact_33_4880
timestamp 1624857261
transform 1 0 22576 0 1 82693
box 0 0 1 1
use contact_33  contact_33_1760
timestamp 1624857261
transform 1 0 22984 0 1 82693
box 0 0 1 1
use contact_33  contact_33_1759
timestamp 1624857261
transform 1 0 22984 0 1 82965
box 0 0 1 1
use contact_33  contact_33_5056
timestamp 1624857261
transform 1 0 22304 0 1 83101
box 0 0 1 1
use contact_33  contact_33_1722
timestamp 1624857261
transform 1 0 22984 0 1 83101
box 0 0 1 1
use contact_33  contact_33_4342
timestamp 1624857261
transform 1 0 23392 0 1 83101
box 0 0 1 1
use contact_33  contact_33_4362
timestamp 1624857261
transform 1 0 23392 0 1 82285
box 0 0 1 1
use contact_33  contact_33_4363
timestamp 1624857261
transform 1 0 23392 0 1 82557
box 0 0 1 1
use contact_33  contact_33_4364
timestamp 1624857261
transform 1 0 23392 0 1 82965
box 0 0 1 1
use contact_33  contact_33_4365
timestamp 1624857261
transform 1 0 23392 0 1 82693
box 0 0 1 1
use contact_33  contact_33_4472
timestamp 1624857261
transform 1 0 23528 0 1 82149
box 0 0 1 1
use contact_33  contact_33_5308
timestamp 1624857261
transform 1 0 1224 0 1 84325
box 0 0 1 1
use contact_13  contact_13_529
timestamp 1624857261
transform 1 0 1801 0 1 83331
box 0 0 1 1
use contact_19  contact_19_529
timestamp 1624857261
transform 1 0 1794 0 1 83340
box 0 0 1 1
use contact_14  contact_14_529
timestamp 1624857261
transform 1 0 1797 0 1 83339
box 0 0 1 1
use contact_13  contact_13_528
timestamp 1624857261
transform 1 0 1801 0 1 83667
box 0 0 1 1
use contact_13  contact_13_527
timestamp 1624857261
transform 1 0 1801 0 1 84003
box 0 0 1 1
use contact_19  contact_19_528
timestamp 1624857261
transform 1 0 1794 0 1 83676
box 0 0 1 1
use contact_19  contact_19_527
timestamp 1624857261
transform 1 0 1794 0 1 84012
box 0 0 1 1
use contact_14  contact_14_528
timestamp 1624857261
transform 1 0 1797 0 1 83675
box 0 0 1 1
use contact_14  contact_14_527
timestamp 1624857261
transform 1 0 1797 0 1 84011
box 0 0 1 1
use contact_13  contact_13_526
timestamp 1624857261
transform 1 0 1801 0 1 84339
box 0 0 1 1
use contact_19  contact_19_526
timestamp 1624857261
transform 1 0 1794 0 1 84348
box 0 0 1 1
use contact_14  contact_14_526
timestamp 1624857261
transform 1 0 1797 0 1 84347
box 0 0 1 1
use contact_7  contact_7_106
timestamp 1624857261
transform 1 0 1793 0 1 84343
box 0 0 1 1
use contact_33  contact_33_1999
timestamp 1624857261
transform 1 0 21896 0 1 83509
box 0 0 1 1
use contact_33  contact_33_2000
timestamp 1624857261
transform 1 0 21896 0 1 83781
box 0 0 1 1
use contact_33  contact_33_2001
timestamp 1624857261
transform 1 0 21760 0 1 84189
box 0 0 1 1
use contact_33  contact_33_2002
timestamp 1624857261
transform 1 0 21760 0 1 83917
box 0 0 1 1
use contact_33  contact_33_2055
timestamp 1624857261
transform 1 0 21896 0 1 84325
box 0 0 1 1
use contact_33  contact_33_2056
timestamp 1624857261
transform 1 0 21896 0 1 84597
box 0 0 1 1
use contact_33  contact_33_2109
timestamp 1624857261
transform 1 0 21760 0 1 83373
box 0 0 1 1
use contact_33  contact_33_1545
timestamp 1624857261
transform 1 0 23120 0 1 83781
box 0 0 1 1
use contact_33  contact_33_1546
timestamp 1624857261
transform 1 0 23120 0 1 83509
box 0 0 1 1
use contact_33  contact_33_1721
timestamp 1624857261
transform 1 0 22984 0 1 83373
box 0 0 1 1
use contact_33  contact_33_4741
timestamp 1624857261
transform 1 0 22712 0 1 84597
box 0 0 1 1
use contact_33  contact_33_4760
timestamp 1624857261
transform 1 0 22576 0 1 84189
box 0 0 1 1
use contact_33  contact_33_4761
timestamp 1624857261
transform 1 0 22576 0 1 83917
box 0 0 1 1
use contact_33  contact_33_5057
timestamp 1624857261
transform 1 0 22304 0 1 83373
box 0 0 1 1
use contact_33  contact_33_4343
timestamp 1624857261
transform 1 0 23392 0 1 83373
box 0 0 1 1
use contact_33  contact_33_4426
timestamp 1624857261
transform 1 0 23392 0 1 83509
box 0 0 1 1
use contact_33  contact_33_4427
timestamp 1624857261
transform 1 0 23392 0 1 83781
box 0 0 1 1
use contact_33  contact_33_1371
timestamp 1624857261
transform 1 0 28424 0 1 83917
box 0 0 1 1
use contact_33  contact_33_1372
timestamp 1624857261
transform 1 0 28424 0 1 83645
box 0 0 1 1
use contact_33  contact_33_1401
timestamp 1624857261
transform 1 0 28424 0 1 84053
box 0 0 1 1
use contact_33  contact_33_1402
timestamp 1624857261
transform 1 0 28424 0 1 84325
box 0 0 1 1
use contact_33  contact_33_1439
timestamp 1624857261
transform 1 0 28560 0 1 84461
box 0 0 1 1
use contact_13  contact_13_525
timestamp 1624857261
transform 1 0 1801 0 1 84675
box 0 0 1 1
use contact_13  contact_13_524
timestamp 1624857261
transform 1 0 1801 0 1 85011
box 0 0 1 1
use contact_19  contact_19_525
timestamp 1624857261
transform 1 0 1794 0 1 84684
box 0 0 1 1
use contact_14  contact_14_525
timestamp 1624857261
transform 1 0 1797 0 1 84683
box 0 0 1 1
use contact_13  contact_13_523
timestamp 1624857261
transform 1 0 1801 0 1 85347
box 0 0 1 1
use contact_19  contact_19_524
timestamp 1624857261
transform 1 0 1794 0 1 85020
box 0 0 1 1
use contact_19  contact_19_523
timestamp 1624857261
transform 1 0 1794 0 1 85356
box 0 0 1 1
use contact_14  contact_14_524
timestamp 1624857261
transform 1 0 1797 0 1 85019
box 0 0 1 1
use contact_14  contact_14_523
timestamp 1624857261
transform 1 0 1797 0 1 85355
box 0 0 1 1
use contact_13  contact_13_522
timestamp 1624857261
transform 1 0 1801 0 1 85683
box 0 0 1 1
use contact_19  contact_19_522
timestamp 1624857261
transform 1 0 1794 0 1 85692
box 0 0 1 1
use contact_14  contact_14_522
timestamp 1624857261
transform 1 0 1797 0 1 85691
box 0 0 1 1
use contact_33  contact_33_1955
timestamp 1624857261
transform 1 0 21760 0 1 85141
box 0 0 1 1
use contact_33  contact_33_1956
timestamp 1624857261
transform 1 0 21760 0 1 85413
box 0 0 1 1
use contact_33  contact_33_2277
timestamp 1624857261
transform 1 0 21760 0 1 85821
box 0 0 1 1
use contact_33  contact_33_4740
timestamp 1624857261
transform 1 0 22712 0 1 84869
box 0 0 1 1
use contact_33  contact_33_1783
timestamp 1624857261
transform 1 0 22984 0 1 85005
box 0 0 1 1
use contact_33  contact_33_5069
timestamp 1624857261
transform 1 0 22440 0 1 85413
box 0 0 1 1
use contact_33  contact_33_4874
timestamp 1624857261
transform 1 0 22712 0 1 85413
box 0 0 1 1
use contact_33  contact_33_1784
timestamp 1624857261
transform 1 0 22984 0 1 85277
box 0 0 1 1
use contact_33  contact_33_1782
timestamp 1624857261
transform 1 0 22984 0 1 85413
box 0 0 1 1
use contact_33  contact_33_5093
timestamp 1624857261
transform 1 0 22304 0 1 85821
box 0 0 1 1
use contact_33  contact_33_5068
timestamp 1624857261
transform 1 0 22440 0 1 85685
box 0 0 1 1
use contact_33  contact_33_4875
timestamp 1624857261
transform 1 0 22712 0 1 85685
box 0 0 1 1
use contact_33  contact_33_1781
timestamp 1624857261
transform 1 0 22984 0 1 85685
box 0 0 1 1
use contact_33  contact_33_1636
timestamp 1624857261
transform 1 0 22984 0 1 85821
box 0 0 1 1
use contact_33  contact_33_4400
timestamp 1624857261
transform 1 0 23528 0 1 85685
box 0 0 1 1
use contact_33  contact_33_4401
timestamp 1624857261
transform 1 0 23528 0 1 85413
box 0 0 1 1
use contact_33  contact_33_4556
timestamp 1624857261
transform 1 0 23528 0 1 85821
box 0 0 1 1
use contact_33  contact_33_4708
timestamp 1624857261
transform 1 0 23528 0 1 85277
box 0 0 1 1
use contact_33  contact_33_4709
timestamp 1624857261
transform 1 0 23528 0 1 85005
box 0 0 1 1
use contact_33  contact_33_1440
timestamp 1624857261
transform 1 0 28560 0 1 84733
box 0 0 1 1
use contact_33  contact_33_5331
timestamp 1624857261
transform 1 0 1224 0 1 86093
box 0 0 1 1
use contact_13  contact_13_521
timestamp 1624857261
transform 1 0 1801 0 1 86019
box 0 0 1 1
use contact_13  contact_13_520
timestamp 1624857261
transform 1 0 1801 0 1 86355
box 0 0 1 1
use contact_19  contact_19_521
timestamp 1624857261
transform 1 0 1794 0 1 86028
box 0 0 1 1
use contact_14  contact_14_521
timestamp 1624857261
transform 1 0 1797 0 1 86027
box 0 0 1 1
use contact_7  contact_7_105
timestamp 1624857261
transform 1 0 1793 0 1 86023
box 0 0 1 1
use contact_13  contact_13_519
timestamp 1624857261
transform 1 0 1801 0 1 86691
box 0 0 1 1
use contact_19  contact_19_520
timestamp 1624857261
transform 1 0 1794 0 1 86364
box 0 0 1 1
use contact_19  contact_19_519
timestamp 1624857261
transform 1 0 1794 0 1 86700
box 0 0 1 1
use contact_14  contact_14_520
timestamp 1624857261
transform 1 0 1797 0 1 86363
box 0 0 1 1
use contact_14  contact_14_519
timestamp 1624857261
transform 1 0 1797 0 1 86699
box 0 0 1 1
use contact_13  contact_13_518
timestamp 1624857261
transform 1 0 1801 0 1 87027
box 0 0 1 1
use contact_19  contact_19_518
timestamp 1624857261
transform 1 0 1794 0 1 87036
box 0 0 1 1
use contact_14  contact_14_518
timestamp 1624857261
transform 1 0 1797 0 1 87035
box 0 0 1 1
use contact_33  contact_33_2225
timestamp 1624857261
transform 1 0 21896 0 1 86637
box 0 0 1 1
use contact_33  contact_33_2226
timestamp 1624857261
transform 1 0 21896 0 1 86909
box 0 0 1 1
use contact_33  contact_33_2247
timestamp 1624857261
transform 1 0 21760 0 1 87045
box 0 0 1 1
use contact_33  contact_33_2248
timestamp 1624857261
transform 1 0 21760 0 1 87317
box 0 0 1 1
use contact_33  contact_33_2278
timestamp 1624857261
transform 1 0 21760 0 1 86093
box 0 0 1 1
use contact_33  contact_33_2279
timestamp 1624857261
transform 1 0 21760 0 1 86501
box 0 0 1 1
use contact_33  contact_33_2280
timestamp 1624857261
transform 1 0 21760 0 1 86229
box 0 0 1 1
use contact_33  contact_33_5092
timestamp 1624857261
transform 1 0 22304 0 1 86093
box 0 0 1 1
use contact_33  contact_33_5000
timestamp 1624857261
transform 1 0 22440 0 1 86229
box 0 0 1 1
use contact_33  contact_33_1741
timestamp 1624857261
transform 1 0 22984 0 1 86229
box 0 0 1 1
use contact_33  contact_33_1635
timestamp 1624857261
transform 1 0 22984 0 1 86093
box 0 0 1 1
use contact_33  contact_33_5001
timestamp 1624857261
transform 1 0 22440 0 1 86501
box 0 0 1 1
use contact_33  contact_33_1744
timestamp 1624857261
transform 1 0 23120 0 1 86637
box 0 0 1 1
use contact_33  contact_33_1742
timestamp 1624857261
transform 1 0 22984 0 1 86501
box 0 0 1 1
use contact_33  contact_33_5006
timestamp 1624857261
transform 1 0 22168 0 1 87045
box 0 0 1 1
use contact_33  contact_33_4790
timestamp 1624857261
transform 1 0 22576 0 1 87045
box 0 0 1 1
use contact_33  contact_33_1743
timestamp 1624857261
transform 1 0 23120 0 1 86909
box 0 0 1 1
use contact_33  contact_33_1690
timestamp 1624857261
transform 1 0 22984 0 1 87045
box 0 0 1 1
use contact_33  contact_33_5007
timestamp 1624857261
transform 1 0 22168 0 1 87317
box 0 0 1 1
use contact_33  contact_33_4791
timestamp 1624857261
transform 1 0 22576 0 1 87317
box 0 0 1 1
use contact_33  contact_33_1689
timestamp 1624857261
transform 1 0 22984 0 1 87317
box 0 0 1 1
use contact_33  contact_33_4408
timestamp 1624857261
transform 1 0 23392 0 1 86909
box 0 0 1 1
use contact_33  contact_33_4409
timestamp 1624857261
transform 1 0 23392 0 1 86637
box 0 0 1 1
use contact_33  contact_33_4557
timestamp 1624857261
transform 1 0 23528 0 1 86093
box 0 0 1 1
use contact_33  contact_33_4558
timestamp 1624857261
transform 1 0 23528 0 1 86501
box 0 0 1 1
use contact_33  contact_33_4559
timestamp 1624857261
transform 1 0 23528 0 1 86229
box 0 0 1 1
use contact_33  contact_33_4660
timestamp 1624857261
transform 1 0 23528 0 1 87045
box 0 0 1 1
use contact_33  contact_33_4661
timestamp 1624857261
transform 1 0 23528 0 1 87317
box 0 0 1 1
use contact_33  contact_33_5326
timestamp 1624857261
transform 1 0 1224 0 1 87589
box 0 0 1 1
use contact_13  contact_13_517
timestamp 1624857261
transform 1 0 1801 0 1 87363
box 0 0 1 1
use contact_13  contact_13_516
timestamp 1624857261
transform 1 0 1801 0 1 87699
box 0 0 1 1
use contact_19  contact_19_517
timestamp 1624857261
transform 1 0 1794 0 1 87372
box 0 0 1 1
use contact_19  contact_19_516
timestamp 1624857261
transform 1 0 1794 0 1 87708
box 0 0 1 1
use contact_14  contact_14_517
timestamp 1624857261
transform 1 0 1797 0 1 87371
box 0 0 1 1
use contact_14  contact_14_516
timestamp 1624857261
transform 1 0 1797 0 1 87707
box 0 0 1 1
use contact_7  contact_7_104
timestamp 1624857261
transform 1 0 1793 0 1 87703
box 0 0 1 1
use contact_13  contact_13_515
timestamp 1624857261
transform 1 0 1801 0 1 88035
box 0 0 1 1
use contact_19  contact_19_515
timestamp 1624857261
transform 1 0 1794 0 1 88044
box 0 0 1 1
use contact_14  contact_14_515
timestamp 1624857261
transform 1 0 1797 0 1 88043
box 0 0 1 1
use contact_13  contact_13_514
timestamp 1624857261
transform 1 0 1801 0 1 88371
box 0 0 1 1
use contact_19  contact_19_514
timestamp 1624857261
transform 1 0 1794 0 1 88380
box 0 0 1 1
use contact_14  contact_14_514
timestamp 1624857261
transform 1 0 1797 0 1 88379
box 0 0 1 1
use contact_33  contact_33_1903
timestamp 1624857261
transform 1 0 21760 0 1 88541
box 0 0 1 1
use contact_33  contact_33_1904
timestamp 1624857261
transform 1 0 21760 0 1 88269
box 0 0 1 1
use contact_33  contact_33_1919
timestamp 1624857261
transform 1 0 21896 0 1 88677
box 0 0 1 1
use contact_33  contact_33_1949
timestamp 1624857261
transform 1 0 21896 0 1 88133
box 0 0 1 1
use contact_33  contact_33_1950
timestamp 1624857261
transform 1 0 21896 0 1 87861
box 0 0 1 1
use contact_33  contact_33_2245
timestamp 1624857261
transform 1 0 21760 0 1 87725
box 0 0 1 1
use contact_33  contact_33_2246
timestamp 1624857261
transform 1 0 21760 0 1 87453
box 0 0 1 1
use contact_33  contact_33_1829
timestamp 1624857261
transform 1 0 23120 0 1 88133
box 0 0 1 1
use contact_33  contact_33_1830
timestamp 1624857261
transform 1 0 23120 0 1 87861
box 0 0 1 1
use contact_33  contact_33_1831
timestamp 1624857261
transform 1 0 23120 0 1 87453
box 0 0 1 1
use contact_33  contact_33_1832
timestamp 1624857261
transform 1 0 23120 0 1 87725
box 0 0 1 1
use contact_33  contact_33_4856
timestamp 1624857261
transform 1 0 22712 0 1 88133
box 0 0 1 1
use contact_33  contact_33_4857
timestamp 1624857261
transform 1 0 22712 0 1 87861
box 0 0 1 1
use contact_33  contact_33_5147
timestamp 1624857261
transform 1 0 22168 0 1 88541
box 0 0 1 1
use contact_33  contact_33_4422
timestamp 1624857261
transform 1 0 23392 0 1 88133
box 0 0 1 1
use contact_33  contact_33_4423
timestamp 1624857261
transform 1 0 23392 0 1 87861
box 0 0 1 1
use contact_33  contact_33_4662
timestamp 1624857261
transform 1 0 23528 0 1 87725
box 0 0 1 1
use contact_33  contact_33_4663
timestamp 1624857261
transform 1 0 23528 0 1 87453
box 0 0 1 1
use contact_33  contact_33_1475
timestamp 1624857261
transform 1 0 28288 0 1 87861
box 0 0 1 1
use contact_33  contact_33_1476
timestamp 1624857261
transform 1 0 28288 0 1 87589
box 0 0 1 1
use contact_33  contact_33_5337
timestamp 1624857261
transform 1 0 1224 0 1 89493
box 0 0 1 1
use contact_13  contact_13_513
timestamp 1624857261
transform 1 0 1801 0 1 88707
box 0 0 1 1
use contact_13  contact_13_512
timestamp 1624857261
transform 1 0 1801 0 1 89043
box 0 0 1 1
use contact_19  contact_19_513
timestamp 1624857261
transform 1 0 1794 0 1 88716
box 0 0 1 1
use contact_14  contact_14_513
timestamp 1624857261
transform 1 0 1797 0 1 88715
box 0 0 1 1
use contact_13  contact_13_511
timestamp 1624857261
transform 1 0 1801 0 1 89379
box 0 0 1 1
use contact_19  contact_19_512
timestamp 1624857261
transform 1 0 1794 0 1 89052
box 0 0 1 1
use contact_14  contact_14_512
timestamp 1624857261
transform 1 0 1797 0 1 89051
box 0 0 1 1
use contact_7  contact_7_103
timestamp 1624857261
transform 1 0 1793 0 1 89383
box 0 0 1 1
use contact_13  contact_13_510
timestamp 1624857261
transform 1 0 1801 0 1 89715
box 0 0 1 1
use contact_19  contact_19_511
timestamp 1624857261
transform 1 0 1794 0 1 89388
box 0 0 1 1
use contact_19  contact_19_510
timestamp 1624857261
transform 1 0 1794 0 1 89724
box 0 0 1 1
use contact_14  contact_14_511
timestamp 1624857261
transform 1 0 1797 0 1 89387
box 0 0 1 1
use contact_14  contact_14_510
timestamp 1624857261
transform 1 0 1797 0 1 89723
box 0 0 1 1
use contact_13  contact_13_509
timestamp 1624857261
transform 1 0 1801 0 1 90051
box 0 0 1 1
use contact_19  contact_19_509
timestamp 1624857261
transform 1 0 1794 0 1 90060
box 0 0 1 1
use contact_14  contact_14_509
timestamp 1624857261
transform 1 0 1797 0 1 90059
box 0 0 1 1
use contact_33  contact_33_1920
timestamp 1624857261
transform 1 0 21896 0 1 88949
box 0 0 1 1
use contact_33  contact_33_2007
timestamp 1624857261
transform 1 0 21760 0 1 89765
box 0 0 1 1
use contact_33  contact_33_2008
timestamp 1624857261
transform 1 0 21760 0 1 90037
box 0 0 1 1
use contact_33  contact_33_2243
timestamp 1624857261
transform 1 0 21760 0 1 89085
box 0 0 1 1
use contact_33  contact_33_2244
timestamp 1624857261
transform 1 0 21760 0 1 89357
box 0 0 1 1
use contact_33  contact_33_5146
timestamp 1624857261
transform 1 0 22168 0 1 88949
box 0 0 1 1
use contact_33  contact_33_5033
timestamp 1624857261
transform 1 0 22440 0 1 88949
box 0 0 1 1
use contact_33  contact_33_5032
timestamp 1624857261
transform 1 0 22440 0 1 89221
box 0 0 1 1
use contact_33  contact_33_4826
timestamp 1624857261
transform 1 0 22576 0 1 89357
box 0 0 1 1
use contact_33  contact_33_1885
timestamp 1624857261
transform 1 0 22984 0 1 89357
box 0 0 1 1
use contact_33  contact_33_4973
timestamp 1624857261
transform 1 0 22168 0 1 89765
box 0 0 1 1
use contact_33  contact_33_4827
timestamp 1624857261
transform 1 0 22576 0 1 89629
box 0 0 1 1
use contact_33  contact_33_1886
timestamp 1624857261
transform 1 0 22984 0 1 89629
box 0 0 1 1
use contact_33  contact_33_1884
timestamp 1624857261
transform 1 0 22984 0 1 89765
box 0 0 1 1
use contact_33  contact_33_4972
timestamp 1624857261
transform 1 0 22168 0 1 90037
box 0 0 1 1
use contact_33  contact_33_1883
timestamp 1624857261
transform 1 0 22984 0 1 90037
box 0 0 1 1
use contact_33  contact_33_4666
timestamp 1624857261
transform 1 0 23528 0 1 90037
box 0 0 1 1
use contact_33  contact_33_4667
timestamp 1624857261
transform 1 0 23528 0 1 89765
box 0 0 1 1
use contact_33  contact_33_4668
timestamp 1624857261
transform 1 0 23528 0 1 89357
box 0 0 1 1
use contact_33  contact_33_4669
timestamp 1624857261
transform 1 0 23528 0 1 89629
box 0 0 1 1
use contact_33  contact_33_1437
timestamp 1624857261
transform 1 0 28288 0 1 89493
box 0 0 1 1
use contact_33  contact_33_1438
timestamp 1624857261
transform 1 0 28288 0 1 89221
box 0 0 1 1
use contact_33  contact_33_5361
timestamp 1624857261
transform 1 0 1224 0 1 91125
box 0 0 1 1
use contact_13  contact_13_508
timestamp 1624857261
transform 1 0 1801 0 1 90387
box 0 0 1 1
use contact_19  contact_19_508
timestamp 1624857261
transform 1 0 1794 0 1 90396
box 0 0 1 1
use contact_14  contact_14_508
timestamp 1624857261
transform 1 0 1797 0 1 90395
box 0 0 1 1
use contact_13  contact_13_507
timestamp 1624857261
transform 1 0 1801 0 1 90723
box 0 0 1 1
use contact_19  contact_19_507
timestamp 1624857261
transform 1 0 1794 0 1 90732
box 0 0 1 1
use contact_14  contact_14_507
timestamp 1624857261
transform 1 0 1797 0 1 90731
box 0 0 1 1
use contact_13  contact_13_506
timestamp 1624857261
transform 1 0 1801 0 1 91059
box 0 0 1 1
use contact_19  contact_19_506
timestamp 1624857261
transform 1 0 1794 0 1 91068
box 0 0 1 1
use contact_14  contact_14_506
timestamp 1624857261
transform 1 0 1797 0 1 91067
box 0 0 1 1
use contact_7  contact_7_102
timestamp 1624857261
transform 1 0 1793 0 1 91063
box 0 0 1 1
use contact_13  contact_13_505
timestamp 1624857261
transform 1 0 1801 0 1 91395
box 0 0 1 1
use contact_19  contact_19_505
timestamp 1624857261
transform 1 0 1794 0 1 91404
box 0 0 1 1
use contact_14  contact_14_505
timestamp 1624857261
transform 1 0 1797 0 1 91403
box 0 0 1 1
use contact_33  contact_33_2105
timestamp 1624857261
transform 1 0 21760 0 1 90581
box 0 0 1 1
use contact_33  contact_33_2106
timestamp 1624857261
transform 1 0 21760 0 1 90853
box 0 0 1 1
use contact_33  contact_33_2107
timestamp 1624857261
transform 1 0 21896 0 1 91261
box 0 0 1 1
use contact_33  contact_33_2108
timestamp 1624857261
transform 1 0 21896 0 1 90989
box 0 0 1 1
use contact_33  contact_33_2147
timestamp 1624857261
transform 1 0 21760 0 1 91397
box 0 0 1 1
use contact_33  contact_33_4917
timestamp 1624857261
transform 1 0 22440 0 1 90173
box 0 0 1 1
use contact_33  contact_33_1597
timestamp 1624857261
transform 1 0 23120 0 1 90173
box 0 0 1 1
use contact_33  contact_33_5178
timestamp 1624857261
transform 1 0 22168 0 1 90581
box 0 0 1 1
use contact_33  contact_33_4916
timestamp 1624857261
transform 1 0 22440 0 1 90445
box 0 0 1 1
use contact_33  contact_33_4872
timestamp 1624857261
transform 1 0 22576 0 1 90581
box 0 0 1 1
use contact_33  contact_33_1619
timestamp 1624857261
transform 1 0 22984 0 1 90581
box 0 0 1 1
use contact_33  contact_33_1598
timestamp 1624857261
transform 1 0 23120 0 1 90445
box 0 0 1 1
use contact_33  contact_33_5181
timestamp 1624857261
transform 1 0 22168 0 1 90989
box 0 0 1 1
use contact_33  contact_33_5179
timestamp 1624857261
transform 1 0 22168 0 1 90853
box 0 0 1 1
use contact_33  contact_33_4873
timestamp 1624857261
transform 1 0 22576 0 1 90853
box 0 0 1 1
use contact_33  contact_33_4871
timestamp 1624857261
transform 1 0 22712 0 1 90989
box 0 0 1 1
use contact_33  contact_33_1735
timestamp 1624857261
transform 1 0 22984 0 1 90989
box 0 0 1 1
use contact_33  contact_33_1620
timestamp 1624857261
transform 1 0 22984 0 1 90853
box 0 0 1 1
use contact_33  contact_33_5180
timestamp 1624857261
transform 1 0 22168 0 1 91261
box 0 0 1 1
use contact_33  contact_33_4870
timestamp 1624857261
transform 1 0 22712 0 1 91261
box 0 0 1 1
use contact_33  contact_33_1736
timestamp 1624857261
transform 1 0 22984 0 1 91261
box 0 0 1 1
use contact_33  contact_33_5173
timestamp 1624857261
transform 1 0 22304 0 1 91397
box 0 0 1 1
use contact_33  contact_33_4799
timestamp 1624857261
transform 1 0 22712 0 1 91397
box 0 0 1 1
use contact_33  contact_33_1738
timestamp 1624857261
transform 1 0 22984 0 1 91397
box 0 0 1 1
use contact_33  contact_33_4344
timestamp 1624857261
transform 1 0 23392 0 1 90989
box 0 0 1 1
use contact_33  contact_33_4345
timestamp 1624857261
transform 1 0 23392 0 1 91261
box 0 0 1 1
use contact_33  contact_33_4506
timestamp 1624857261
transform 1 0 23528 0 1 91397
box 0 0 1 1
use contact_33  contact_33_4614
timestamp 1624857261
transform 1 0 23528 0 1 90853
box 0 0 1 1
use contact_33  contact_33_4615
timestamp 1624857261
transform 1 0 23528 0 1 90581
box 0 0 1 1
use contact_33  contact_33_4616
timestamp 1624857261
transform 1 0 23528 0 1 90173
box 0 0 1 1
use contact_33  contact_33_4617
timestamp 1624857261
transform 1 0 23528 0 1 90445
box 0 0 1 1
use contact_13  contact_13_504
timestamp 1624857261
transform 1 0 1801 0 1 91731
box 0 0 1 1
use contact_19  contact_19_504
timestamp 1624857261
transform 1 0 1794 0 1 91740
box 0 0 1 1
use contact_14  contact_14_504
timestamp 1624857261
transform 1 0 1797 0 1 91739
box 0 0 1 1
use contact_13  contact_13_503
timestamp 1624857261
transform 1 0 1801 0 1 92067
box 0 0 1 1
use contact_19  contact_19_503
timestamp 1624857261
transform 1 0 1794 0 1 92076
box 0 0 1 1
use contact_14  contact_14_503
timestamp 1624857261
transform 1 0 1797 0 1 92075
box 0 0 1 1
use contact_13  contact_13_502
timestamp 1624857261
transform 1 0 1801 0 1 92403
box 0 0 1 1
use contact_19  contact_19_502
timestamp 1624857261
transform 1 0 1794 0 1 92412
box 0 0 1 1
use contact_14  contact_14_502
timestamp 1624857261
transform 1 0 1797 0 1 92411
box 0 0 1 1
use contact_13  contact_13_501
timestamp 1624857261
transform 1 0 1801 0 1 92739
box 0 0 1 1
use contact_19  contact_19_501
timestamp 1624857261
transform 1 0 1794 0 1 92748
box 0 0 1 1
use contact_14  contact_14_501
timestamp 1624857261
transform 1 0 1797 0 1 92747
box 0 0 1 1
use contact_7  contact_7_101
timestamp 1624857261
transform 1 0 1793 0 1 92743
box 0 0 1 1
use contact_33  contact_33_2145
timestamp 1624857261
transform 1 0 21760 0 1 92077
box 0 0 1 1
use contact_33  contact_33_2146
timestamp 1624857261
transform 1 0 21760 0 1 91805
box 0 0 1 1
use contact_33  contact_33_2148
timestamp 1624857261
transform 1 0 21760 0 1 91669
box 0 0 1 1
use contact_33  contact_33_2198
timestamp 1624857261
transform 1 0 21760 0 1 92621
box 0 0 1 1
use contact_33  contact_33_2199
timestamp 1624857261
transform 1 0 21896 0 1 92213
box 0 0 1 1
use contact_33  contact_33_2200
timestamp 1624857261
transform 1 0 21896 0 1 92485
box 0 0 1 1
use contact_33  contact_33_1675
timestamp 1624857261
transform 1 0 23120 0 1 91805
box 0 0 1 1
use contact_33  contact_33_1676
timestamp 1624857261
transform 1 0 23120 0 1 92077
box 0 0 1 1
use contact_33  contact_33_1737
timestamp 1624857261
transform 1 0 22984 0 1 91669
box 0 0 1 1
use contact_33  contact_33_4792
timestamp 1624857261
transform 1 0 22576 0 1 92621
box 0 0 1 1
use contact_33  contact_33_4798
timestamp 1624857261
transform 1 0 22712 0 1 91669
box 0 0 1 1
use contact_33  contact_33_4928
timestamp 1624857261
transform 1 0 22440 0 1 91805
box 0 0 1 1
use contact_33  contact_33_4929
timestamp 1624857261
transform 1 0 22440 0 1 92077
box 0 0 1 1
use contact_33  contact_33_5172
timestamp 1624857261
transform 1 0 22304 0 1 91669
box 0 0 1 1
use contact_33  contact_33_4507
timestamp 1624857261
transform 1 0 23528 0 1 91669
box 0 0 1 1
use contact_33  contact_33_4508
timestamp 1624857261
transform 1 0 23528 0 1 92077
box 0 0 1 1
use contact_33  contact_33_4509
timestamp 1624857261
transform 1 0 23528 0 1 91805
box 0 0 1 1
use contact_33  contact_33_1389
timestamp 1624857261
transform 1 0 28424 0 1 92077
box 0 0 1 1
use contact_33  contact_33_1390
timestamp 1624857261
transform 1 0 28424 0 1 92349
box 0 0 1 1
use contact_33  contact_33_1479
timestamp 1624857261
transform 1 0 28560 0 1 92349
box 0 0 1 1
use contact_33  contact_33_1480
timestamp 1624857261
transform 1 0 28560 0 1 92621
box 0 0 1 1
use contact_33  contact_33_1482
timestamp 1624857261
transform 1 0 28288 0 1 92757
box 0 0 1 1
use contact_33  contact_33_5314
timestamp 1624857261
transform 1 0 1224 0 1 92893
box 0 0 1 1
use contact_13  contact_13_500
timestamp 1624857261
transform 1 0 1801 0 1 93075
box 0 0 1 1
use contact_19  contact_19_500
timestamp 1624857261
transform 1 0 1794 0 1 93084
box 0 0 1 1
use contact_14  contact_14_500
timestamp 1624857261
transform 1 0 1797 0 1 93083
box 0 0 1 1
use contact_13  contact_13_499
timestamp 1624857261
transform 1 0 1801 0 1 93411
box 0 0 1 1
use contact_19  contact_19_499
timestamp 1624857261
transform 1 0 1794 0 1 93420
box 0 0 1 1
use contact_14  contact_14_499
timestamp 1624857261
transform 1 0 1797 0 1 93419
box 0 0 1 1
use contact_13  contact_13_498
timestamp 1624857261
transform 1 0 1801 0 1 93747
box 0 0 1 1
use contact_19  contact_19_498
timestamp 1624857261
transform 1 0 1794 0 1 93756
box 0 0 1 1
use contact_14  contact_14_498
timestamp 1624857261
transform 1 0 1797 0 1 93755
box 0 0 1 1
use contact_13  contact_13_497
timestamp 1624857261
transform 1 0 1801 0 1 94083
box 0 0 1 1
use contact_19  contact_19_497
timestamp 1624857261
transform 1 0 1794 0 1 94092
box 0 0 1 1
use contact_14  contact_14_497
timestamp 1624857261
transform 1 0 1797 0 1 94091
box 0 0 1 1
use contact_33  contact_33_1953
timestamp 1624857261
transform 1 0 21896 0 1 93029
box 0 0 1 1
use contact_33  contact_33_1954
timestamp 1624857261
transform 1 0 21896 0 1 93301
box 0 0 1 1
use contact_33  contact_33_2197
timestamp 1624857261
transform 1 0 21760 0 1 92893
box 0 0 1 1
use contact_33  contact_33_1717
timestamp 1624857261
transform 1 0 23120 0 1 93981
box 0 0 1 1
use contact_33  contact_33_1718
timestamp 1624857261
transform 1 0 23120 0 1 93709
box 0 0 1 1
use contact_33  contact_33_1719
timestamp 1624857261
transform 1 0 22984 0 1 93301
box 0 0 1 1
use contact_33  contact_33_1720
timestamp 1624857261
transform 1 0 22984 0 1 93573
box 0 0 1 1
use contact_33  contact_33_1801
timestamp 1624857261
transform 1 0 23120 0 1 94117
box 0 0 1 1
use contact_33  contact_33_4793
timestamp 1624857261
transform 1 0 22576 0 1 92893
box 0 0 1 1
use contact_33  contact_33_4861
timestamp 1624857261
transform 1 0 22576 0 1 94117
box 0 0 1 1
use contact_33  contact_33_4966
timestamp 1624857261
transform 1 0 22440 0 1 93573
box 0 0 1 1
use contact_33  contact_33_4967
timestamp 1624857261
transform 1 0 22440 0 1 93301
box 0 0 1 1
use contact_33  contact_33_4384
timestamp 1624857261
transform 1 0 23392 0 1 94117
box 0 0 1 1
use contact_33  contact_33_4394
timestamp 1624857261
transform 1 0 23392 0 1 93301
box 0 0 1 1
use contact_33  contact_33_4395
timestamp 1624857261
transform 1 0 23392 0 1 93573
box 0 0 1 1
use contact_33  contact_33_4396
timestamp 1624857261
transform 1 0 23528 0 1 93981
box 0 0 1 1
use contact_33  contact_33_4397
timestamp 1624857261
transform 1 0 23528 0 1 93709
box 0 0 1 1
use contact_33  contact_33_1427
timestamp 1624857261
transform 1 0 28560 0 1 93165
box 0 0 1 1
use contact_33  contact_33_1428
timestamp 1624857261
transform 1 0 28560 0 1 93437
box 0 0 1 1
use contact_33  contact_33_1481
timestamp 1624857261
transform 1 0 28288 0 1 93029
box 0 0 1 1
use contact_33  contact_33_5296
timestamp 1624857261
transform 1 0 1224 0 1 94525
box 0 0 1 1
use contact_13  contact_13_496
timestamp 1624857261
transform 1 0 1801 0 1 94419
box 0 0 1 1
use contact_19  contact_19_496
timestamp 1624857261
transform 1 0 1794 0 1 94428
box 0 0 1 1
use contact_14  contact_14_496
timestamp 1624857261
transform 1 0 1797 0 1 94427
box 0 0 1 1
use contact_7  contact_7_100
timestamp 1624857261
transform 1 0 1793 0 1 94423
box 0 0 1 1
use contact_13  contact_13_495
timestamp 1624857261
transform 1 0 1801 0 1 94755
box 0 0 1 1
use contact_19  contact_19_495
timestamp 1624857261
transform 1 0 1794 0 1 94764
box 0 0 1 1
use contact_14  contact_14_495
timestamp 1624857261
transform 1 0 1797 0 1 94763
box 0 0 1 1
use contact_13  contact_13_494
timestamp 1624857261
transform 1 0 1801 0 1 95091
box 0 0 1 1
use contact_19  contact_19_494
timestamp 1624857261
transform 1 0 1794 0 1 95100
box 0 0 1 1
use contact_14  contact_14_494
timestamp 1624857261
transform 1 0 1797 0 1 95099
box 0 0 1 1
use contact_13  contact_13_493
timestamp 1624857261
transform 1 0 1801 0 1 95427
box 0 0 1 1
use contact_19  contact_19_493
timestamp 1624857261
transform 1 0 1794 0 1 95436
box 0 0 1 1
use contact_14  contact_14_493
timestamp 1624857261
transform 1 0 1797 0 1 95435
box 0 0 1 1
use contact_33  contact_33_1935
timestamp 1624857261
transform 1 0 21896 0 1 94797
box 0 0 1 1
use contact_33  contact_33_1936
timestamp 1624857261
transform 1 0 21896 0 1 94525
box 0 0 1 1
use contact_33  contact_33_2213
timestamp 1624857261
transform 1 0 21760 0 1 94933
box 0 0 1 1
use contact_33  contact_33_2214
timestamp 1624857261
transform 1 0 21760 0 1 95205
box 0 0 1 1
use contact_33  contact_33_2216
timestamp 1624857261
transform 1 0 21896 0 1 95341
box 0 0 1 1
use contact_33  contact_33_4860
timestamp 1624857261
transform 1 0 22576 0 1 94389
box 0 0 1 1
use contact_33  contact_33_1802
timestamp 1624857261
transform 1 0 23120 0 1 94389
box 0 0 1 1
use contact_33  contact_33_5167
timestamp 1624857261
transform 1 0 22304 0 1 94525
box 0 0 1 1
use contact_33  contact_33_5166
timestamp 1624857261
transform 1 0 22304 0 1 94797
box 0 0 1 1
use contact_33  contact_33_1804
timestamp 1624857261
transform 1 0 23120 0 1 94525
box 0 0 1 1
use contact_33  contact_33_1803
timestamp 1624857261
transform 1 0 23120 0 1 94797
box 0 0 1 1
use contact_33  contact_33_5141
timestamp 1624857261
transform 1 0 22168 0 1 94933
box 0 0 1 1
use contact_33  contact_33_5140
timestamp 1624857261
transform 1 0 22168 0 1 95205
box 0 0 1 1
use contact_33  contact_33_4747
timestamp 1624857261
transform 1 0 22576 0 1 95205
box 0 0 1 1
use contact_33  contact_33_4746
timestamp 1624857261
transform 1 0 22576 0 1 94933
box 0 0 1 1
use contact_33  contact_33_1786
timestamp 1624857261
transform 1 0 23120 0 1 94933
box 0 0 1 1
use contact_33  contact_33_1785
timestamp 1624857261
transform 1 0 23120 0 1 95205
box 0 0 1 1
use contact_33  contact_33_1695
timestamp 1624857261
transform 1 0 22984 0 1 95341
box 0 0 1 1
use contact_33  contact_33_4385
timestamp 1624857261
transform 1 0 23392 0 1 94389
box 0 0 1 1
use contact_33  contact_33_4390
timestamp 1624857261
transform 1 0 23528 0 1 95205
box 0 0 1 1
use contact_33  contact_33_4391
timestamp 1624857261
transform 1 0 23528 0 1 94933
box 0 0 1 1
use contact_33  contact_33_4392
timestamp 1624857261
transform 1 0 23528 0 1 94525
box 0 0 1 1
use contact_33  contact_33_4393
timestamp 1624857261
transform 1 0 23528 0 1 94797
box 0 0 1 1
use contact_33  contact_33_4704
timestamp 1624857261
transform 1 0 23392 0 1 95341
box 0 0 1 1
use contact_33  contact_33_1505
timestamp 1624857261
transform 1 0 28424 0 1 95477
box 0 0 1 1
use contact_33  contact_33_5322
timestamp 1624857261
transform 1 0 1224 0 1 96157
box 0 0 1 1
use contact_13  contact_13_492
timestamp 1624857261
transform 1 0 1801 0 1 95763
box 0 0 1 1
use contact_19  contact_19_492
timestamp 1624857261
transform 1 0 1794 0 1 95772
box 0 0 1 1
use contact_14  contact_14_492
timestamp 1624857261
transform 1 0 1797 0 1 95771
box 0 0 1 1
use contact_13  contact_13_491
timestamp 1624857261
transform 1 0 1801 0 1 96099
box 0 0 1 1
use contact_19  contact_19_491
timestamp 1624857261
transform 1 0 1794 0 1 96108
box 0 0 1 1
use contact_14  contact_14_491
timestamp 1624857261
transform 1 0 1797 0 1 96107
box 0 0 1 1
use contact_7  contact_7_99
timestamp 1624857261
transform 1 0 1793 0 1 96103
box 0 0 1 1
use contact_13  contact_13_490
timestamp 1624857261
transform 1 0 1801 0 1 96435
box 0 0 1 1
use contact_19  contact_19_490
timestamp 1624857261
transform 1 0 1794 0 1 96444
box 0 0 1 1
use contact_14  contact_14_490
timestamp 1624857261
transform 1 0 1797 0 1 96443
box 0 0 1 1
use contact_13  contact_13_489
timestamp 1624857261
transform 1 0 1801 0 1 96771
box 0 0 1 1
use contact_19  contact_19_489
timestamp 1624857261
transform 1 0 1794 0 1 96780
box 0 0 1 1
use contact_14  contact_14_489
timestamp 1624857261
transform 1 0 1797 0 1 96779
box 0 0 1 1
use contact_33  contact_33_1993
timestamp 1624857261
transform 1 0 21760 0 1 96429
box 0 0 1 1
use contact_33  contact_33_1994
timestamp 1624857261
transform 1 0 21760 0 1 96157
box 0 0 1 1
use contact_33  contact_33_2149
timestamp 1624857261
transform 1 0 21896 0 1 96565
box 0 0 1 1
use contact_33  contact_33_2150
timestamp 1624857261
transform 1 0 21896 0 1 96837
box 0 0 1 1
use contact_33  contact_33_2211
timestamp 1624857261
transform 1 0 21896 0 1 96021
box 0 0 1 1
use contact_33  contact_33_2212
timestamp 1624857261
transform 1 0 21896 0 1 95749
box 0 0 1 1
use contact_33  contact_33_2215
timestamp 1624857261
transform 1 0 21896 0 1 95613
box 0 0 1 1
use contact_33  contact_33_5028
timestamp 1624857261
transform 1 0 22168 0 1 95749
box 0 0 1 1
use contact_33  contact_33_4819
timestamp 1624857261
transform 1 0 22712 0 1 95749
box 0 0 1 1
use contact_33  contact_33_1869
timestamp 1624857261
transform 1 0 22984 0 1 95749
box 0 0 1 1
use contact_33  contact_33_1696
timestamp 1624857261
transform 1 0 22984 0 1 95613
box 0 0 1 1
use contact_33  contact_33_5029
timestamp 1624857261
transform 1 0 22168 0 1 96021
box 0 0 1 1
use contact_33  contact_33_4818
timestamp 1624857261
transform 1 0 22712 0 1 96021
box 0 0 1 1
use contact_33  contact_33_1870
timestamp 1624857261
transform 1 0 22984 0 1 96021
box 0 0 1 1
use contact_33  contact_33_1868
timestamp 1624857261
transform 1 0 22984 0 1 96157
box 0 0 1 1
use contact_33  contact_33_4892
timestamp 1624857261
transform 1 0 22712 0 1 96565
box 0 0 1 1
use contact_33  contact_33_1867
timestamp 1624857261
transform 1 0 22984 0 1 96429
box 0 0 1 1
use contact_33  contact_33_4893
timestamp 1624857261
transform 1 0 22712 0 1 96837
box 0 0 1 1
use contact_33  contact_33_4546
timestamp 1624857261
transform 1 0 23528 0 1 96429
box 0 0 1 1
use contact_33  contact_33_4547
timestamp 1624857261
transform 1 0 23528 0 1 96157
box 0 0 1 1
use contact_33  contact_33_4705
timestamp 1624857261
transform 1 0 23392 0 1 95613
box 0 0 1 1
use contact_33  contact_33_4706
timestamp 1624857261
transform 1 0 23392 0 1 96021
box 0 0 1 1
use contact_33  contact_33_4707
timestamp 1624857261
transform 1 0 23392 0 1 95749
box 0 0 1 1
use contact_33  contact_33_1446
timestamp 1624857261
transform 1 0 28424 0 1 96701
box 0 0 1 1
use contact_33  contact_33_1506
timestamp 1624857261
transform 1 0 28424 0 1 95749
box 0 0 1 1
use contact_33  contact_33_5299
timestamp 1624857261
transform 1 0 1224 0 1 97789
box 0 0 1 1
use contact_13  contact_13_488
timestamp 1624857261
transform 1 0 1801 0 1 97107
box 0 0 1 1
use contact_19  contact_19_488
timestamp 1624857261
transform 1 0 1794 0 1 97116
box 0 0 1 1
use contact_14  contact_14_488
timestamp 1624857261
transform 1 0 1797 0 1 97115
box 0 0 1 1
use contact_13  contact_13_487
timestamp 1624857261
transform 1 0 1801 0 1 97443
box 0 0 1 1
use contact_19  contact_19_487
timestamp 1624857261
transform 1 0 1794 0 1 97452
box 0 0 1 1
use contact_14  contact_14_487
timestamp 1624857261
transform 1 0 1797 0 1 97451
box 0 0 1 1
use contact_13  contact_13_486
timestamp 1624857261
transform 1 0 1801 0 1 97779
box 0 0 1 1
use contact_19  contact_19_486
timestamp 1624857261
transform 1 0 1794 0 1 97788
box 0 0 1 1
use contact_14  contact_14_486
timestamp 1624857261
transform 1 0 1797 0 1 97787
box 0 0 1 1
use contact_7  contact_7_98
timestamp 1624857261
transform 1 0 1793 0 1 97783
box 0 0 1 1
use contact_13  contact_13_485
timestamp 1624857261
transform 1 0 1801 0 1 98115
box 0 0 1 1
use contact_19  contact_19_485
timestamp 1624857261
transform 1 0 1794 0 1 98124
box 0 0 1 1
use contact_14  contact_14_485
timestamp 1624857261
transform 1 0 1797 0 1 98123
box 0 0 1 1
use contact_33  contact_33_2151
timestamp 1624857261
transform 1 0 21760 0 1 97245
box 0 0 1 1
use contact_33  contact_33_2152
timestamp 1624857261
transform 1 0 21760 0 1 96973
box 0 0 1 1
use contact_33  contact_33_1535
timestamp 1624857261
transform 1 0 22984 0 1 98061
box 0 0 1 1
use contact_33  contact_33_1793
timestamp 1624857261
transform 1 0 23120 0 1 97925
box 0 0 1 1
use contact_33  contact_33_1794
timestamp 1624857261
transform 1 0 23120 0 1 97653
box 0 0 1 1
use contact_33  contact_33_1795
timestamp 1624857261
transform 1 0 23120 0 1 97245
box 0 0 1 1
use contact_33  contact_33_1796
timestamp 1624857261
transform 1 0 23120 0 1 97517
box 0 0 1 1
use contact_33  contact_33_4808
timestamp 1624857261
transform 1 0 22576 0 1 97517
box 0 0 1 1
use contact_33  contact_33_4809
timestamp 1624857261
transform 1 0 22576 0 1 97245
box 0 0 1 1
use contact_33  contact_33_4816
timestamp 1624857261
transform 1 0 22576 0 1 98061
box 0 0 1 1
use contact_33  contact_33_5074
timestamp 1624857261
transform 1 0 22168 0 1 98061
box 0 0 1 1
use contact_33  contact_33_4496
timestamp 1624857261
transform 1 0 23392 0 1 97245
box 0 0 1 1
use contact_33  contact_33_4497
timestamp 1624857261
transform 1 0 23392 0 1 97517
box 0 0 1 1
use contact_33  contact_33_4498
timestamp 1624857261
transform 1 0 23392 0 1 97925
box 0 0 1 1
use contact_33  contact_33_4499
timestamp 1624857261
transform 1 0 23392 0 1 97653
box 0 0 1 1
use contact_33  contact_33_4618
timestamp 1624857261
transform 1 0 23528 0 1 98061
box 0 0 1 1
use contact_33  contact_33_1445
timestamp 1624857261
transform 1 0 28424 0 1 96973
box 0 0 1 1
use contact_33  contact_33_1491
timestamp 1624857261
transform 1 0 28288 0 1 97517
box 0 0 1 1
use contact_33  contact_33_1492
timestamp 1624857261
transform 1 0 28288 0 1 97925
box 0 0 1 1
use contact_33  contact_33_5349
timestamp 1624857261
transform 1 0 1224 0 1 99557
box 0 0 1 1
use contact_13  contact_13_484
timestamp 1624857261
transform 1 0 1801 0 1 98451
box 0 0 1 1
use contact_19  contact_19_484
timestamp 1624857261
transform 1 0 1794 0 1 98460
box 0 0 1 1
use contact_14  contact_14_484
timestamp 1624857261
transform 1 0 1797 0 1 98459
box 0 0 1 1
use contact_13  contact_13_483
timestamp 1624857261
transform 1 0 1801 0 1 98787
box 0 0 1 1
use contact_19  contact_19_483
timestamp 1624857261
transform 1 0 1794 0 1 98796
box 0 0 1 1
use contact_14  contact_14_483
timestamp 1624857261
transform 1 0 1797 0 1 98795
box 0 0 1 1
use contact_13  contact_13_482
timestamp 1624857261
transform 1 0 1801 0 1 99123
box 0 0 1 1
use contact_19  contact_19_482
timestamp 1624857261
transform 1 0 1794 0 1 99132
box 0 0 1 1
use contact_14  contact_14_482
timestamp 1624857261
transform 1 0 1797 0 1 99131
box 0 0 1 1
use contact_13  contact_13_481
timestamp 1624857261
transform 1 0 1801 0 1 99459
box 0 0 1 1
use contact_19  contact_19_481
timestamp 1624857261
transform 1 0 1794 0 1 99468
box 0 0 1 1
use contact_14  contact_14_481
timestamp 1624857261
transform 1 0 1797 0 1 99467
box 0 0 1 1
use contact_7  contact_7_97
timestamp 1624857261
transform 1 0 1793 0 1 99463
box 0 0 1 1
use contact_33  contact_33_1907
timestamp 1624857261
transform 1 0 21760 0 1 99557
box 0 0 1 1
use contact_33  contact_33_1908
timestamp 1624857261
transform 1 0 21760 0 1 99285
box 0 0 1 1
use contact_33  contact_33_2057
timestamp 1624857261
transform 1 0 21896 0 1 99149
box 0 0 1 1
use contact_33  contact_33_2058
timestamp 1624857261
transform 1 0 21896 0 1 98877
box 0 0 1 1
use contact_33  contact_33_2059
timestamp 1624857261
transform 1 0 21896 0 1 98469
box 0 0 1 1
use contact_33  contact_33_2060
timestamp 1624857261
transform 1 0 21896 0 1 98741
box 0 0 1 1
use contact_33  contact_33_5075
timestamp 1624857261
transform 1 0 22168 0 1 98333
box 0 0 1 1
use contact_33  contact_33_5073
timestamp 1624857261
transform 1 0 22168 0 1 98469
box 0 0 1 1
use contact_33  contact_33_4817
timestamp 1624857261
transform 1 0 22576 0 1 98333
box 0 0 1 1
use contact_33  contact_33_1536
timestamp 1624857261
transform 1 0 22984 0 1 98333
box 0 0 1 1
use contact_33  contact_33_1813
timestamp 1624857261
transform 1 0 23120 0 1 98469
box 0 0 1 1
use contact_33  contact_33_5072
timestamp 1624857261
transform 1 0 22168 0 1 98741
box 0 0 1 1
use contact_33  contact_33_4756
timestamp 1624857261
transform 1 0 22576 0 1 98877
box 0 0 1 1
use contact_33  contact_33_1816
timestamp 1624857261
transform 1 0 22984 0 1 98877
box 0 0 1 1
use contact_33  contact_33_1814
timestamp 1624857261
transform 1 0 23120 0 1 98741
box 0 0 1 1
use contact_33  contact_33_4757
timestamp 1624857261
transform 1 0 22576 0 1 99149
box 0 0 1 1
use contact_33  contact_33_1815
timestamp 1624857261
transform 1 0 22984 0 1 99149
box 0 0 1 1
use contact_33  contact_33_4986
timestamp 1624857261
transform 1 0 22168 0 1 99285
box 0 0 1 1
use contact_33  contact_33_4982
timestamp 1624857261
transform 1 0 22440 0 1 99285
box 0 0 1 1
use contact_33  contact_33_1779
timestamp 1624857261
transform 1 0 22984 0 1 99285
box 0 0 1 1
use contact_33  contact_33_4987
timestamp 1624857261
transform 1 0 22168 0 1 99557
box 0 0 1 1
use contact_33  contact_33_4983
timestamp 1624857261
transform 1 0 22440 0 1 99557
box 0 0 1 1
use contact_33  contact_33_1780
timestamp 1624857261
transform 1 0 22984 0 1 99557
box 0 0 1 1
use contact_33  contact_33_4500
timestamp 1624857261
transform 1 0 23528 0 1 99557
box 0 0 1 1
use contact_33  contact_33_4501
timestamp 1624857261
transform 1 0 23528 0 1 99285
box 0 0 1 1
use contact_33  contact_33_4619
timestamp 1624857261
transform 1 0 23528 0 1 98333
box 0 0 1 1
use contact_33  contact_33_4620
timestamp 1624857261
transform 1 0 23392 0 1 99149
box 0 0 1 1
use contact_33  contact_33_4621
timestamp 1624857261
transform 1 0 23392 0 1 98877
box 0 0 1 1
use contact_33  contact_33_4622
timestamp 1624857261
transform 1 0 23392 0 1 98469
box 0 0 1 1
use contact_33  contact_33_4623
timestamp 1624857261
transform 1 0 23392 0 1 98741
box 0 0 1 1
use contact_33  contact_33_1393
timestamp 1624857261
transform 1 0 28560 0 1 99421
box 0 0 1 1
use contact_13  contact_13_480
timestamp 1624857261
transform 1 0 1801 0 1 99795
box 0 0 1 1
use contact_19  contact_19_480
timestamp 1624857261
transform 1 0 1794 0 1 99804
box 0 0 1 1
use contact_14  contact_14_480
timestamp 1624857261
transform 1 0 1797 0 1 99803
box 0 0 1 1
use contact_13  contact_13_479
timestamp 1624857261
transform 1 0 1801 0 1 100131
box 0 0 1 1
use contact_19  contact_19_479
timestamp 1624857261
transform 1 0 1794 0 1 100140
box 0 0 1 1
use contact_14  contact_14_479
timestamp 1624857261
transform 1 0 1797 0 1 100139
box 0 0 1 1
use contact_13  contact_13_478
timestamp 1624857261
transform 1 0 1801 0 1 100467
box 0 0 1 1
use contact_19  contact_19_478
timestamp 1624857261
transform 1 0 1794 0 1 100476
box 0 0 1 1
use contact_14  contact_14_478
timestamp 1624857261
transform 1 0 1797 0 1 100475
box 0 0 1 1
use contact_13  contact_13_477
timestamp 1624857261
transform 1 0 1801 0 1 100803
box 0 0 1 1
use contact_19  contact_19_477
timestamp 1624857261
transform 1 0 1794 0 1 100812
box 0 0 1 1
use contact_14  contact_14_477
timestamp 1624857261
transform 1 0 1797 0 1 100811
box 0 0 1 1
use contact_33  contact_33_1917
timestamp 1624857261
transform 1 0 21896 0 1 99693
box 0 0 1 1
use contact_33  contact_33_1918
timestamp 1624857261
transform 1 0 21896 0 1 99965
box 0 0 1 1
use contact_33  contact_33_1969
timestamp 1624857261
transform 1 0 21760 0 1 100101
box 0 0 1 1
use contact_33  contact_33_1970
timestamp 1624857261
transform 1 0 21760 0 1 100373
box 0 0 1 1
use contact_33  contact_33_1971
timestamp 1624857261
transform 1 0 21760 0 1 100781
box 0 0 1 1
use contact_33  contact_33_1972
timestamp 1624857261
transform 1 0 21760 0 1 100509
box 0 0 1 1
use contact_33  contact_33_2119
timestamp 1624857261
transform 1 0 21896 0 1 100917
box 0 0 1 1
use contact_33  contact_33_1797
timestamp 1624857261
transform 1 0 22984 0 1 100373
box 0 0 1 1
use contact_33  contact_33_1798
timestamp 1624857261
transform 1 0 22984 0 1 100101
box 0 0 1 1
use contact_33  contact_33_1799
timestamp 1624857261
transform 1 0 22984 0 1 99693
box 0 0 1 1
use contact_33  contact_33_1800
timestamp 1624857261
transform 1 0 22984 0 1 99965
box 0 0 1 1
use contact_33  contact_33_4974
timestamp 1624857261
transform 1 0 22440 0 1 100509
box 0 0 1 1
use contact_33  contact_33_4975
timestamp 1624857261
transform 1 0 22440 0 1 100781
box 0 0 1 1
use contact_33  contact_33_4984
timestamp 1624857261
transform 1 0 22168 0 1 99965
box 0 0 1 1
use contact_33  contact_33_4985
timestamp 1624857261
transform 1 0 22168 0 1 99693
box 0 0 1 1
use contact_33  contact_33_4648
timestamp 1624857261
transform 1 0 23392 0 1 99693
box 0 0 1 1
use contact_33  contact_33_4649
timestamp 1624857261
transform 1 0 23392 0 1 99965
box 0 0 1 1
use contact_33  contact_33_4650
timestamp 1624857261
transform 1 0 23392 0 1 100373
box 0 0 1 1
use contact_33  contact_33_4651
timestamp 1624857261
transform 1 0 23392 0 1 100101
box 0 0 1 1
use contact_33  contact_33_1387
timestamp 1624857261
transform 1 0 28288 0 1 100917
box 0 0 1 1
use contact_33  contact_33_1388
timestamp 1624857261
transform 1 0 28288 0 1 100645
box 0 0 1 1
use contact_33  contact_33_1394
timestamp 1624857261
transform 1 0 28560 0 1 99693
box 0 0 1 1
use contact_33  contact_33_1417
timestamp 1624857261
transform 1 0 28424 0 1 99965
box 0 0 1 1
use contact_33  contact_33_1418
timestamp 1624857261
transform 1 0 28424 0 1 100373
box 0 0 1 1
use contact_33  contact_33_5325
timestamp 1624857261
transform 1 0 1224 0 1 101189
box 0 0 1 1
use contact_13  contact_13_476
timestamp 1624857261
transform 1 0 1801 0 1 101139
box 0 0 1 1
use contact_19  contact_19_476
timestamp 1624857261
transform 1 0 1794 0 1 101148
box 0 0 1 1
use contact_14  contact_14_476
timestamp 1624857261
transform 1 0 1797 0 1 101147
box 0 0 1 1
use contact_7  contact_7_96
timestamp 1624857261
transform 1 0 1793 0 1 101143
box 0 0 1 1
use contact_13  contact_13_475
timestamp 1624857261
transform 1 0 1801 0 1 101475
box 0 0 1 1
use contact_19  contact_19_475
timestamp 1624857261
transform 1 0 1794 0 1 101484
box 0 0 1 1
use contact_14  contact_14_475
timestamp 1624857261
transform 1 0 1797 0 1 101483
box 0 0 1 1
use contact_13  contact_13_474
timestamp 1624857261
transform 1 0 1801 0 1 101811
box 0 0 1 1
use contact_19  contact_19_474
timestamp 1624857261
transform 1 0 1794 0 1 101820
box 0 0 1 1
use contact_14  contact_14_474
timestamp 1624857261
transform 1 0 1797 0 1 101819
box 0 0 1 1
use contact_13  contact_13_473
timestamp 1624857261
transform 1 0 1801 0 1 102147
box 0 0 1 1
use contact_19  contact_19_473
timestamp 1624857261
transform 1 0 1794 0 1 102156
box 0 0 1 1
use contact_14  contact_14_473
timestamp 1624857261
transform 1 0 1797 0 1 102155
box 0 0 1 1
use contact_33  contact_33_2120
timestamp 1624857261
transform 1 0 21896 0 1 101189
box 0 0 1 1
use contact_33  contact_33_2195
timestamp 1624857261
transform 1 0 21760 0 1 102005
box 0 0 1 1
use contact_33  contact_33_2196
timestamp 1624857261
transform 1 0 21760 0 1 101733
box 0 0 1 1
use contact_33  contact_33_4753
timestamp 1624857261
transform 1 0 22712 0 1 101189
box 0 0 1 1
use contact_33  contact_33_4752
timestamp 1624857261
transform 1 0 22712 0 1 101461
box 0 0 1 1
use contact_33  contact_33_1665
timestamp 1624857261
transform 1 0 23120 0 1 101597
box 0 0 1 1
use contact_33  contact_33_5122
timestamp 1624857261
transform 1 0 22304 0 1 102005
box 0 0 1 1
use contact_33  contact_33_4989
timestamp 1624857261
transform 1 0 22440 0 1 102005
box 0 0 1 1
use contact_33  contact_33_4988
timestamp 1624857261
transform 1 0 22440 0 1 101733
box 0 0 1 1
use contact_33  contact_33_4797
timestamp 1624857261
transform 1 0 22712 0 1 102005
box 0 0 1 1
use contact_33  contact_33_1669
timestamp 1624857261
transform 1 0 22984 0 1 102005
box 0 0 1 1
use contact_33  contact_33_1666
timestamp 1624857261
transform 1 0 23120 0 1 101869
box 0 0 1 1
use contact_33  contact_33_5123
timestamp 1624857261
transform 1 0 22304 0 1 102277
box 0 0 1 1
use contact_33  contact_33_4796
timestamp 1624857261
transform 1 0 22712 0 1 102277
box 0 0 1 1
use contact_33  contact_33_1670
timestamp 1624857261
transform 1 0 22984 0 1 102277
box 0 0 1 1
use contact_33  contact_33_4348
timestamp 1624857261
transform 1 0 23392 0 1 102005
box 0 0 1 1
use contact_33  contact_33_4349
timestamp 1624857261
transform 1 0 23392 0 1 102277
box 0 0 1 1
use contact_33  contact_33_4682
timestamp 1624857261
transform 1 0 23528 0 1 101869
box 0 0 1 1
use contact_33  contact_33_4683
timestamp 1624857261
transform 1 0 23528 0 1 101597
box 0 0 1 1
use contact_33  contact_33_1441
timestamp 1624857261
transform 1 0 28560 0 1 101053
box 0 0 1 1
use contact_33  contact_33_1442
timestamp 1624857261
transform 1 0 28560 0 1 101325
box 0 0 1 1
use contact_33  contact_33_1469
timestamp 1624857261
transform 1 0 28288 0 1 101325
box 0 0 1 1
use contact_33  contact_33_1470
timestamp 1624857261
transform 1 0 28288 0 1 101597
box 0 0 1 1
use contact_33  contact_33_5357
timestamp 1624857261
transform 1 0 1224 0 1 102685
box 0 0 1 1
use contact_13  contact_13_472
timestamp 1624857261
transform 1 0 1801 0 1 102483
box 0 0 1 1
use contact_19  contact_19_472
timestamp 1624857261
transform 1 0 1794 0 1 102492
box 0 0 1 1
use contact_14  contact_14_472
timestamp 1624857261
transform 1 0 1797 0 1 102491
box 0 0 1 1
use contact_13  contact_13_471
timestamp 1624857261
transform 1 0 1801 0 1 102819
box 0 0 1 1
use contact_19  contact_19_471
timestamp 1624857261
transform 1 0 1794 0 1 102828
box 0 0 1 1
use contact_14  contact_14_471
timestamp 1624857261
transform 1 0 1797 0 1 102827
box 0 0 1 1
use contact_7  contact_7_95
timestamp 1624857261
transform 1 0 1793 0 1 102823
box 0 0 1 1
use contact_13  contact_13_470
timestamp 1624857261
transform 1 0 1801 0 1 103155
box 0 0 1 1
use contact_19  contact_19_470
timestamp 1624857261
transform 1 0 1794 0 1 103164
box 0 0 1 1
use contact_14  contact_14_470
timestamp 1624857261
transform 1 0 1797 0 1 103163
box 0 0 1 1
use contact_13  contact_13_469
timestamp 1624857261
transform 1 0 1801 0 1 103491
box 0 0 1 1
use contact_19  contact_19_469
timestamp 1624857261
transform 1 0 1794 0 1 103500
box 0 0 1 1
use contact_14  contact_14_469
timestamp 1624857261
transform 1 0 1797 0 1 103499
box 0 0 1 1
use contact_33  contact_33_2087
timestamp 1624857261
transform 1 0 21896 0 1 102821
box 0 0 1 1
use contact_33  contact_33_2088
timestamp 1624857261
transform 1 0 21896 0 1 103093
box 0 0 1 1
use contact_33  contact_33_2163
timestamp 1624857261
transform 1 0 21760 0 1 102685
box 0 0 1 1
use contact_33  contact_33_2164
timestamp 1624857261
transform 1 0 21760 0 1 102413
box 0 0 1 1
use contact_33  contact_33_2191
timestamp 1624857261
transform 1 0 21760 0 1 103229
box 0 0 1 1
use contact_33  contact_33_2192
timestamp 1624857261
transform 1 0 21760 0 1 103501
box 0 0 1 1
use contact_33  contact_33_2194
timestamp 1624857261
transform 1 0 21760 0 1 103637
box 0 0 1 1
use contact_33  contact_33_4876
timestamp 1624857261
transform 1 0 22576 0 1 102413
box 0 0 1 1
use contact_33  contact_33_1668
timestamp 1624857261
transform 1 0 23120 0 1 102413
box 0 0 1 1
use contact_33  contact_33_5155
timestamp 1624857261
transform 1 0 22168 0 1 102821
box 0 0 1 1
use contact_33  contact_33_4996
timestamp 1624857261
transform 1 0 22440 0 1 102821
box 0 0 1 1
use contact_33  contact_33_4877
timestamp 1624857261
transform 1 0 22576 0 1 102685
box 0 0 1 1
use contact_33  contact_33_1529
timestamp 1624857261
transform 1 0 22984 0 1 102821
box 0 0 1 1
use contact_33  contact_33_1667
timestamp 1624857261
transform 1 0 23120 0 1 102685
box 0 0 1 1
use contact_33  contact_33_5154
timestamp 1624857261
transform 1 0 22168 0 1 103093
box 0 0 1 1
use contact_33  contact_33_4999
timestamp 1624857261
transform 1 0 22304 0 1 103229
box 0 0 1 1
use contact_33  contact_33_4997
timestamp 1624857261
transform 1 0 22440 0 1 103093
box 0 0 1 1
use contact_33  contact_33_1530
timestamp 1624857261
transform 1 0 22984 0 1 103093
box 0 0 1 1
use contact_33  contact_33_1751
timestamp 1624857261
transform 1 0 23120 0 1 103229
box 0 0 1 1
use contact_33  contact_33_5124
timestamp 1624857261
transform 1 0 22168 0 1 103637
box 0 0 1 1
use contact_33  contact_33_4998
timestamp 1624857261
transform 1 0 22304 0 1 103501
box 0 0 1 1
use contact_33  contact_33_1754
timestamp 1624857261
transform 1 0 23120 0 1 103637
box 0 0 1 1
use contact_33  contact_33_1752
timestamp 1624857261
transform 1 0 23120 0 1 103501
box 0 0 1 1
use contact_33  contact_33_4346
timestamp 1624857261
transform 1 0 23528 0 1 102685
box 0 0 1 1
use contact_33  contact_33_4347
timestamp 1624857261
transform 1 0 23528 0 1 102413
box 0 0 1 1
use contact_33  contact_33_4439
timestamp 1624857261
transform 1 0 23528 0 1 103637
box 0 0 1 1
use contact_33  contact_33_4652
timestamp 1624857261
transform 1 0 23392 0 1 102821
box 0 0 1 1
use contact_33  contact_33_4653
timestamp 1624857261
transform 1 0 23392 0 1 103093
box 0 0 1 1
use contact_33  contact_33_4654
timestamp 1624857261
transform 1 0 23392 0 1 103501
box 0 0 1 1
use contact_33  contact_33_4655
timestamp 1624857261
transform 1 0 23392 0 1 103229
box 0 0 1 1
use contact_33  contact_33_5372
timestamp 1624857261
transform 1 0 1224 0 1 104589
box 0 0 1 1
use contact_13  contact_13_468
timestamp 1624857261
transform 1 0 1801 0 1 103827
box 0 0 1 1
use contact_19  contact_19_468
timestamp 1624857261
transform 1 0 1794 0 1 103836
box 0 0 1 1
use contact_14  contact_14_468
timestamp 1624857261
transform 1 0 1797 0 1 103835
box 0 0 1 1
use contact_13  contact_13_467
timestamp 1624857261
transform 1 0 1801 0 1 104163
box 0 0 1 1
use contact_19  contact_19_467
timestamp 1624857261
transform 1 0 1794 0 1 104172
box 0 0 1 1
use contact_14  contact_14_467
timestamp 1624857261
transform 1 0 1797 0 1 104171
box 0 0 1 1
use contact_13  contact_13_466
timestamp 1624857261
transform 1 0 1801 0 1 104499
box 0 0 1 1
use contact_19  contact_19_466
timestamp 1624857261
transform 1 0 1794 0 1 104508
box 0 0 1 1
use contact_14  contact_14_466
timestamp 1624857261
transform 1 0 1797 0 1 104507
box 0 0 1 1
use contact_7  contact_7_94
timestamp 1624857261
transform 1 0 1793 0 1 104503
box 0 0 1 1
use contact_13  contact_13_465
timestamp 1624857261
transform 1 0 1801 0 1 104835
box 0 0 1 1
use contact_19  contact_19_465
timestamp 1624857261
transform 1 0 1794 0 1 104844
box 0 0 1 1
use contact_14  contact_14_465
timestamp 1624857261
transform 1 0 1797 0 1 104843
box 0 0 1 1
use contact_33  contact_33_1939
timestamp 1624857261
transform 1 0 21896 0 1 104861
box 0 0 1 1
use contact_33  contact_33_1983
timestamp 1624857261
transform 1 0 21896 0 1 104725
box 0 0 1 1
use contact_33  contact_33_1984
timestamp 1624857261
transform 1 0 21896 0 1 104453
box 0 0 1 1
use contact_33  contact_33_2181
timestamp 1624857261
transform 1 0 21896 0 1 104317
box 0 0 1 1
use contact_33  contact_33_2182
timestamp 1624857261
transform 1 0 21896 0 1 104045
box 0 0 1 1
use contact_33  contact_33_2193
timestamp 1624857261
transform 1 0 21760 0 1 103909
box 0 0 1 1
use contact_33  contact_33_1753
timestamp 1624857261
transform 1 0 23120 0 1 103909
box 0 0 1 1
use contact_33  contact_33_1817
timestamp 1624857261
transform 1 0 22984 0 1 104725
box 0 0 1 1
use contact_33  contact_33_1818
timestamp 1624857261
transform 1 0 22984 0 1 104453
box 0 0 1 1
use contact_33  contact_33_1819
timestamp 1624857261
transform 1 0 22984 0 1 104045
box 0 0 1 1
use contact_33  contact_33_1820
timestamp 1624857261
transform 1 0 22984 0 1 104317
box 0 0 1 1
use contact_33  contact_33_4772
timestamp 1624857261
transform 1 0 22576 0 1 104453
box 0 0 1 1
use contact_33  contact_33_4773
timestamp 1624857261
transform 1 0 22576 0 1 104725
box 0 0 1 1
use contact_33  contact_33_5125
timestamp 1624857261
transform 1 0 22168 0 1 103909
box 0 0 1 1
use contact_33  contact_33_4438
timestamp 1624857261
transform 1 0 23528 0 1 103909
box 0 0 1 1
use contact_33  contact_33_4492
timestamp 1624857261
transform 1 0 23392 0 1 104045
box 0 0 1 1
use contact_33  contact_33_4493
timestamp 1624857261
transform 1 0 23392 0 1 104317
box 0 0 1 1
use contact_33  contact_33_4612
timestamp 1624857261
transform 1 0 23528 0 1 104453
box 0 0 1 1
use contact_33  contact_33_4613
timestamp 1624857261
transform 1 0 23528 0 1 104725
box 0 0 1 1
use contact_33  contact_33_1403
timestamp 1624857261
transform 1 0 28560 0 1 104861
box 0 0 1 1
use contact_33  contact_33_1404
timestamp 1624857261
transform 1 0 28560 0 1 104453
box 0 0 1 1
use contact_33  contact_33_1421
timestamp 1624857261
transform 1 0 28424 0 1 104181
box 0 0 1 1
use contact_33  contact_33_1422
timestamp 1624857261
transform 1 0 28424 0 1 104453
box 0 0 1 1
use contact_33  contact_33_1465
timestamp 1624857261
transform 1 0 28288 0 1 104725
box 0 0 1 1
use contact_33  contact_33_1466
timestamp 1624857261
transform 1 0 28288 0 1 104997
box 0 0 1 1
use contact_33  contact_33_5376
timestamp 1624857261
transform 1 0 1224 0 1 106085
box 0 0 1 1
use contact_13  contact_13_464
timestamp 1624857261
transform 1 0 1801 0 1 105171
box 0 0 1 1
use contact_19  contact_19_464
timestamp 1624857261
transform 1 0 1794 0 1 105180
box 0 0 1 1
use contact_14  contact_14_464
timestamp 1624857261
transform 1 0 1797 0 1 105179
box 0 0 1 1
use contact_13  contact_13_463
timestamp 1624857261
transform 1 0 1801 0 1 105507
box 0 0 1 1
use contact_19  contact_19_463
timestamp 1624857261
transform 1 0 1794 0 1 105516
box 0 0 1 1
use contact_14  contact_14_463
timestamp 1624857261
transform 1 0 1797 0 1 105515
box 0 0 1 1
use contact_13  contact_13_462
timestamp 1624857261
transform 1 0 1801 0 1 105843
box 0 0 1 1
use contact_19  contact_19_462
timestamp 1624857261
transform 1 0 1794 0 1 105852
box 0 0 1 1
use contact_14  contact_14_462
timestamp 1624857261
transform 1 0 1797 0 1 105851
box 0 0 1 1
use contact_13  contact_13_461
timestamp 1624857261
transform 1 0 1801 0 1 106179
box 0 0 1 1
use contact_19  contact_19_461
timestamp 1624857261
transform 1 0 1794 0 1 106188
box 0 0 1 1
use contact_14  contact_14_461
timestamp 1624857261
transform 1 0 1797 0 1 106187
box 0 0 1 1
use contact_7  contact_7_93
timestamp 1624857261
transform 1 0 1793 0 1 106183
box 0 0 1 1
use contact_33  contact_33_1940
timestamp 1624857261
transform 1 0 21896 0 1 105133
box 0 0 1 1
use contact_33  contact_33_2027
timestamp 1624857261
transform 1 0 21760 0 1 105949
box 0 0 1 1
use contact_33  contact_33_2028
timestamp 1624857261
transform 1 0 21760 0 1 105677
box 0 0 1 1
use contact_33  contact_33_2047
timestamp 1624857261
transform 1 0 21896 0 1 106357
box 0 0 1 1
use contact_33  contact_33_4971
timestamp 1624857261
transform 1 0 22304 0 1 105405
box 0 0 1 1
use contact_33  contact_33_4970
timestamp 1624857261
transform 1 0 22304 0 1 105133
box 0 0 1 1
use contact_33  contact_33_4969
timestamp 1624857261
transform 1 0 22440 0 1 105405
box 0 0 1 1
use contact_33  contact_33_4968
timestamp 1624857261
transform 1 0 22440 0 1 105133
box 0 0 1 1
use contact_33  contact_33_1894
timestamp 1624857261
transform 1 0 22984 0 1 105541
box 0 0 1 1
use contact_33  contact_33_5134
timestamp 1624857261
transform 1 0 22440 0 1 105949
box 0 0 1 1
use contact_33  contact_33_1893
timestamp 1624857261
transform 1 0 22984 0 1 105813
box 0 0 1 1
use contact_33  contact_33_1789
timestamp 1624857261
transform 1 0 23120 0 1 105949
box 0 0 1 1
use contact_33  contact_33_5135
timestamp 1624857261
transform 1 0 22440 0 1 106221
box 0 0 1 1
use contact_33  contact_33_4751
timestamp 1624857261
transform 1 0 22712 0 1 106357
box 0 0 1 1
use contact_33  contact_33_1792
timestamp 1624857261
transform 1 0 23120 0 1 106357
box 0 0 1 1
use contact_33  contact_33_1790
timestamp 1624857261
transform 1 0 23120 0 1 106221
box 0 0 1 1
use contact_33  contact_33_4566
timestamp 1624857261
transform 1 0 23528 0 1 105541
box 0 0 1 1
use contact_33  contact_33_4567
timestamp 1624857261
transform 1 0 23528 0 1 105813
box 0 0 1 1
use contact_33  contact_33_4568
timestamp 1624857261
transform 1 0 23528 0 1 106221
box 0 0 1 1
use contact_33  contact_33_4569
timestamp 1624857261
transform 1 0 23528 0 1 105949
box 0 0 1 1
use contact_33  contact_33_4602
timestamp 1624857261
transform 1 0 23392 0 1 106357
box 0 0 1 1
use contact_13  contact_13_460
timestamp 1624857261
transform 1 0 1801 0 1 106515
box 0 0 1 1
use contact_19  contact_19_460
timestamp 1624857261
transform 1 0 1794 0 1 106524
box 0 0 1 1
use contact_14  contact_14_460
timestamp 1624857261
transform 1 0 1797 0 1 106523
box 0 0 1 1
use contact_13  contact_13_459
timestamp 1624857261
transform 1 0 1801 0 1 106851
box 0 0 1 1
use contact_19  contact_19_459
timestamp 1624857261
transform 1 0 1794 0 1 106860
box 0 0 1 1
use contact_14  contact_14_459
timestamp 1624857261
transform 1 0 1797 0 1 106859
box 0 0 1 1
use contact_13  contact_13_458
timestamp 1624857261
transform 1 0 1801 0 1 107187
box 0 0 1 1
use contact_13  contact_13_457
timestamp 1624857261
transform 1 0 1801 0 1 107523
box 0 0 1 1
use contact_19  contact_19_458
timestamp 1624857261
transform 1 0 1794 0 1 107196
box 0 0 1 1
use contact_19  contact_19_457
timestamp 1624857261
transform 1 0 1794 0 1 107532
box 0 0 1 1
use contact_14  contact_14_458
timestamp 1624857261
transform 1 0 1797 0 1 107195
box 0 0 1 1
use contact_14  contact_14_457
timestamp 1624857261
transform 1 0 1797 0 1 107531
box 0 0 1 1
use contact_33  contact_33_2048
timestamp 1624857261
transform 1 0 21896 0 1 106629
box 0 0 1 1
use contact_33  contact_33_2073
timestamp 1624857261
transform 1 0 21896 0 1 107173
box 0 0 1 1
use contact_33  contact_33_2074
timestamp 1624857261
transform 1 0 21896 0 1 107445
box 0 0 1 1
use contact_33  contact_33_2076
timestamp 1624857261
transform 1 0 21896 0 1 107581
box 0 0 1 1
use contact_33  contact_33_4750
timestamp 1624857261
transform 1 0 22712 0 1 106629
box 0 0 1 1
use contact_33  contact_33_1791
timestamp 1624857261
transform 1 0 23120 0 1 106629
box 0 0 1 1
use contact_33  contact_33_4965
timestamp 1624857261
transform 1 0 22168 0 1 107037
box 0 0 1 1
use contact_33  contact_33_4964
timestamp 1624857261
transform 1 0 22168 0 1 106765
box 0 0 1 1
use contact_33  contact_33_4739
timestamp 1624857261
transform 1 0 22576 0 1 107037
box 0 0 1 1
use contact_33  contact_33_4738
timestamp 1624857261
transform 1 0 22576 0 1 106765
box 0 0 1 1
use contact_33  contact_33_1624
timestamp 1624857261
transform 1 0 23120 0 1 106765
box 0 0 1 1
use contact_33  contact_33_1623
timestamp 1624857261
transform 1 0 23120 0 1 107037
box 0 0 1 1
use contact_33  contact_33_4963
timestamp 1624857261
transform 1 0 22440 0 1 107173
box 0 0 1 1
use contact_33  contact_33_4737
timestamp 1624857261
transform 1 0 22576 0 1 107173
box 0 0 1 1
use contact_33  contact_33_1618
timestamp 1624857261
transform 1 0 22984 0 1 107173
box 0 0 1 1
use contact_33  contact_33_5145
timestamp 1624857261
transform 1 0 22304 0 1 107581
box 0 0 1 1
use contact_33  contact_33_4962
timestamp 1624857261
transform 1 0 22440 0 1 107445
box 0 0 1 1
use contact_33  contact_33_4754
timestamp 1624857261
transform 1 0 22576 0 1 107581
box 0 0 1 1
use contact_33  contact_33_4736
timestamp 1624857261
transform 1 0 22576 0 1 107445
box 0 0 1 1
use contact_33  contact_33_1617
timestamp 1624857261
transform 1 0 22984 0 1 107445
box 0 0 1 1
use contact_33  contact_33_1615
timestamp 1624857261
transform 1 0 23120 0 1 107581
box 0 0 1 1
use contact_33  contact_33_4465
timestamp 1624857261
transform 1 0 23392 0 1 107581
box 0 0 1 1
use contact_33  contact_33_4544
timestamp 1624857261
transform 1 0 23528 0 1 107445
box 0 0 1 1
use contact_33  contact_33_4545
timestamp 1624857261
transform 1 0 23528 0 1 107173
box 0 0 1 1
use contact_33  contact_33_4600
timestamp 1624857261
transform 1 0 23528 0 1 107037
box 0 0 1 1
use contact_33  contact_33_4601
timestamp 1624857261
transform 1 0 23528 0 1 106765
box 0 0 1 1
use contact_33  contact_33_4603
timestamp 1624857261
transform 1 0 23392 0 1 106629
box 0 0 1 1
use contact_33  contact_33_5362
timestamp 1624857261
transform 1 0 1224 0 1 107989
box 0 0 1 1
use contact_13  contact_13_456
timestamp 1624857261
transform 1 0 1801 0 1 107859
box 0 0 1 1
use contact_19  contact_19_456
timestamp 1624857261
transform 1 0 1794 0 1 107868
box 0 0 1 1
use contact_14  contact_14_456
timestamp 1624857261
transform 1 0 1797 0 1 107867
box 0 0 1 1
use contact_7  contact_7_92
timestamp 1624857261
transform 1 0 1793 0 1 107863
box 0 0 1 1
use contact_13  contact_13_455
timestamp 1624857261
transform 1 0 1801 0 1 108195
box 0 0 1 1
use contact_19  contact_19_455
timestamp 1624857261
transform 1 0 1794 0 1 108204
box 0 0 1 1
use contact_14  contact_14_455
timestamp 1624857261
transform 1 0 1797 0 1 108203
box 0 0 1 1
use contact_13  contact_13_454
timestamp 1624857261
transform 1 0 1801 0 1 108531
box 0 0 1 1
use contact_13  contact_13_453
timestamp 1624857261
transform 1 0 1801 0 1 108867
box 0 0 1 1
use contact_19  contact_19_454
timestamp 1624857261
transform 1 0 1794 0 1 108540
box 0 0 1 1
use contact_19  contact_19_453
timestamp 1624857261
transform 1 0 1794 0 1 108876
box 0 0 1 1
use contact_14  contact_14_454
timestamp 1624857261
transform 1 0 1797 0 1 108539
box 0 0 1 1
use contact_14  contact_14_453
timestamp 1624857261
transform 1 0 1797 0 1 108875
box 0 0 1 1
use contact_33  contact_33_1931
timestamp 1624857261
transform 1 0 21760 0 1 108261
box 0 0 1 1
use contact_33  contact_33_1932
timestamp 1624857261
transform 1 0 21760 0 1 107989
box 0 0 1 1
use contact_33  contact_33_2075
timestamp 1624857261
transform 1 0 21896 0 1 107853
box 0 0 1 1
use contact_33  contact_33_2093
timestamp 1624857261
transform 1 0 21896 0 1 108397
box 0 0 1 1
use contact_33  contact_33_2094
timestamp 1624857261
transform 1 0 21896 0 1 108669
box 0 0 1 1
use contact_33  contact_33_2095
timestamp 1624857261
transform 1 0 21896 0 1 109077
box 0 0 1 1
use contact_33  contact_33_2096
timestamp 1624857261
transform 1 0 21896 0 1 108805
box 0 0 1 1
use contact_33  contact_33_5144
timestamp 1624857261
transform 1 0 22304 0 1 107853
box 0 0 1 1
use contact_33  contact_33_5090
timestamp 1624857261
transform 1 0 22168 0 1 107989
box 0 0 1 1
use contact_33  contact_33_4755
timestamp 1624857261
transform 1 0 22576 0 1 107853
box 0 0 1 1
use contact_33  contact_33_1769
timestamp 1624857261
transform 1 0 22984 0 1 107989
box 0 0 1 1
use contact_33  contact_33_1616
timestamp 1624857261
transform 1 0 23120 0 1 107853
box 0 0 1 1
use contact_33  contact_33_5106
timestamp 1624857261
transform 1 0 22304 0 1 108397
box 0 0 1 1
use contact_33  contact_33_5091
timestamp 1624857261
transform 1 0 22168 0 1 108261
box 0 0 1 1
use contact_33  contact_33_1772
timestamp 1624857261
transform 1 0 23120 0 1 108397
box 0 0 1 1
use contact_33  contact_33_1770
timestamp 1624857261
transform 1 0 22984 0 1 108261
box 0 0 1 1
use contact_33  contact_33_5107
timestamp 1624857261
transform 1 0 22304 0 1 108669
box 0 0 1 1
use contact_33  contact_33_1771
timestamp 1624857261
transform 1 0 23120 0 1 108669
box 0 0 1 1
use contact_33  contact_33_4328
timestamp 1624857261
transform 1 0 23528 0 1 107989
box 0 0 1 1
use contact_33  contact_33_4329
timestamp 1624857261
transform 1 0 23528 0 1 108261
box 0 0 1 1
use contact_33  contact_33_4414
timestamp 1624857261
transform 1 0 23392 0 1 108397
box 0 0 1 1
use contact_33  contact_33_4415
timestamp 1624857261
transform 1 0 23392 0 1 108669
box 0 0 1 1
use contact_33  contact_33_4464
timestamp 1624857261
transform 1 0 23392 0 1 107853
box 0 0 1 1
use contact_33  contact_33_1363
timestamp 1624857261
transform 1 0 28424 0 1 108397
box 0 0 1 1
use contact_33  contact_33_1364
timestamp 1624857261
transform 1 0 28424 0 1 108805
box 0 0 1 1
use contact_33  contact_33_1447
timestamp 1624857261
transform 1 0 28288 0 1 108941
box 0 0 1 1
use contact_33  contact_33_1503
timestamp 1624857261
transform 1 0 28560 0 1 108397
box 0 0 1 1
use contact_33  contact_33_1504
timestamp 1624857261
transform 1 0 28560 0 1 108125
box 0 0 1 1
use contact_33  contact_33_5316
timestamp 1624857261
transform 1 0 1224 0 1 109621
box 0 0 1 1
use contact_13  contact_13_452
timestamp 1624857261
transform 1 0 1801 0 1 109203
box 0 0 1 1
use contact_19  contact_19_452
timestamp 1624857261
transform 1 0 1794 0 1 109212
box 0 0 1 1
use contact_14  contact_14_452
timestamp 1624857261
transform 1 0 1797 0 1 109211
box 0 0 1 1
use contact_13  contact_13_451
timestamp 1624857261
transform 1 0 1801 0 1 109539
box 0 0 1 1
use contact_19  contact_19_451
timestamp 1624857261
transform 1 0 1794 0 1 109548
box 0 0 1 1
use contact_14  contact_14_451
timestamp 1624857261
transform 1 0 1797 0 1 109547
box 0 0 1 1
use contact_7  contact_7_91
timestamp 1624857261
transform 1 0 1793 0 1 109543
box 0 0 1 1
use contact_13  contact_13_450
timestamp 1624857261
transform 1 0 1801 0 1 109875
box 0 0 1 1
use contact_13  contact_13_449
timestamp 1624857261
transform 1 0 1801 0 1 110211
box 0 0 1 1
use contact_19  contact_19_450
timestamp 1624857261
transform 1 0 1794 0 1 109884
box 0 0 1 1
use contact_19  contact_19_449
timestamp 1624857261
transform 1 0 1794 0 1 110220
box 0 0 1 1
use contact_14  contact_14_450
timestamp 1624857261
transform 1 0 1797 0 1 109883
box 0 0 1 1
use contact_14  contact_14_449
timestamp 1624857261
transform 1 0 1797 0 1 110219
box 0 0 1 1
use contact_33  contact_33_1957
timestamp 1624857261
transform 1 0 21896 0 1 109621
box 0 0 1 1
use contact_33  contact_33_1958
timestamp 1624857261
transform 1 0 21896 0 1 109893
box 0 0 1 1
use contact_33  contact_33_1967
timestamp 1624857261
transform 1 0 21760 0 1 109485
box 0 0 1 1
use contact_33  contact_33_1968
timestamp 1624857261
transform 1 0 21760 0 1 109213
box 0 0 1 1
use contact_33  contact_33_1525
timestamp 1624857261
transform 1 0 22984 0 1 110165
box 0 0 1 1
use contact_33  contact_33_1526
timestamp 1624857261
transform 1 0 22984 0 1 109893
box 0 0 1 1
use contact_33  contact_33_1573
timestamp 1624857261
transform 1 0 23120 0 1 110301
box 0 0 1 1
use contact_33  contact_33_4920
timestamp 1624857261
transform 1 0 22440 0 1 109213
box 0 0 1 1
use contact_33  contact_33_4921
timestamp 1624857261
transform 1 0 22440 0 1 109485
box 0 0 1 1
use contact_33  contact_33_4956
timestamp 1624857261
transform 1 0 22440 0 1 109621
box 0 0 1 1
use contact_33  contact_33_4957
timestamp 1624857261
transform 1 0 22304 0 1 109757
box 0 0 1 1
use contact_33  contact_33_4958
timestamp 1624857261
transform 1 0 22440 0 1 110165
box 0 0 1 1
use contact_33  contact_33_4959
timestamp 1624857261
transform 1 0 22440 0 1 109893
box 0 0 1 1
use contact_33  contact_33_4354
timestamp 1624857261
transform 1 0 23528 0 1 109893
box 0 0 1 1
use contact_33  contact_33_4355
timestamp 1624857261
transform 1 0 23528 0 1 110165
box 0 0 1 1
use contact_33  contact_33_4386
timestamp 1624857261
transform 1 0 23392 0 1 110301
box 0 0 1 1
use contact_33  contact_33_1448
timestamp 1624857261
transform 1 0 28288 0 1 109213
box 0 0 1 1
use contact_33  contact_33_1449
timestamp 1624857261
transform 1 0 28288 0 1 109621
box 0 0 1 1
use contact_33  contact_33_1450
timestamp 1624857261
transform 1 0 28288 0 1 109349
box 0 0 1 1
use contact_33  contact_33_1461
timestamp 1624857261
transform 1 0 28560 0 1 109757
box 0 0 1 1
use contact_33  contact_33_1462
timestamp 1624857261
transform 1 0 28560 0 1 110029
box 0 0 1 1
use contact_33  contact_33_5341
timestamp 1624857261
transform 1 0 1224 0 1 111253
box 0 0 1 1
use contact_13  contact_13_448
timestamp 1624857261
transform 1 0 1801 0 1 110547
box 0 0 1 1
use contact_19  contact_19_448
timestamp 1624857261
transform 1 0 1794 0 1 110556
box 0 0 1 1
use contact_14  contact_14_448
timestamp 1624857261
transform 1 0 1797 0 1 110555
box 0 0 1 1
use contact_13  contact_13_447
timestamp 1624857261
transform 1 0 1801 0 1 110883
box 0 0 1 1
use contact_13  contact_13_446
timestamp 1624857261
transform 1 0 1801 0 1 111219
box 0 0 1 1
use contact_19  contact_19_447
timestamp 1624857261
transform 1 0 1794 0 1 110892
box 0 0 1 1
use contact_14  contact_14_447
timestamp 1624857261
transform 1 0 1797 0 1 110891
box 0 0 1 1
use contact_13  contact_13_445
timestamp 1624857261
transform 1 0 1801 0 1 111555
box 0 0 1 1
use contact_19  contact_19_446
timestamp 1624857261
transform 1 0 1794 0 1 111228
box 0 0 1 1
use contact_19  contact_19_445
timestamp 1624857261
transform 1 0 1794 0 1 111564
box 0 0 1 1
use contact_14  contact_14_446
timestamp 1624857261
transform 1 0 1797 0 1 111227
box 0 0 1 1
use contact_14  contact_14_445
timestamp 1624857261
transform 1 0 1797 0 1 111563
box 0 0 1 1
use contact_7  contact_7_90
timestamp 1624857261
transform 1 0 1793 0 1 111223
box 0 0 1 1
use contact_33  contact_33_2153
timestamp 1624857261
transform 1 0 21896 0 1 111525
box 0 0 1 1
use contact_33  contact_33_2154
timestamp 1624857261
transform 1 0 21896 0 1 111797
box 0 0 1 1
use contact_33  contact_33_2161
timestamp 1624857261
transform 1 0 21760 0 1 111389
box 0 0 1 1
use contact_33  contact_33_2162
timestamp 1624857261
transform 1 0 21760 0 1 111117
box 0 0 1 1
use contact_33  contact_33_5040
timestamp 1624857261
transform 1 0 22304 0 1 110709
box 0 0 1 1
use contact_33  contact_33_5038
timestamp 1624857261
transform 1 0 22440 0 1 110709
box 0 0 1 1
use contact_33  contact_33_1576
timestamp 1624857261
transform 1 0 23120 0 1 110709
box 0 0 1 1
use contact_33  contact_33_1574
timestamp 1624857261
transform 1 0 23120 0 1 110573
box 0 0 1 1
use contact_33  contact_33_5041
timestamp 1624857261
transform 1 0 22304 0 1 110981
box 0 0 1 1
use contact_33  contact_33_5039
timestamp 1624857261
transform 1 0 22440 0 1 110981
box 0 0 1 1
use contact_33  contact_33_4821
timestamp 1624857261
transform 1 0 22576 0 1 111117
box 0 0 1 1
use contact_33  contact_33_1575
timestamp 1624857261
transform 1 0 23120 0 1 110981
box 0 0 1 1
use contact_33  contact_33_1558
timestamp 1624857261
transform 1 0 23120 0 1 111117
box 0 0 1 1
use contact_33  contact_33_4820
timestamp 1624857261
transform 1 0 22576 0 1 111389
box 0 0 1 1
use contact_33  contact_33_1557
timestamp 1624857261
transform 1 0 23120 0 1 111389
box 0 0 1 1
use contact_33  contact_33_5067
timestamp 1624857261
transform 1 0 22168 0 1 111525
box 0 0 1 1
use contact_33  contact_33_4858
timestamp 1624857261
transform 1 0 22712 0 1 111525
box 0 0 1 1
use contact_33  contact_33_1537
timestamp 1624857261
transform 1 0 22984 0 1 111525
box 0 0 1 1
use contact_33  contact_33_5066
timestamp 1624857261
transform 1 0 22168 0 1 111797
box 0 0 1 1
use contact_33  contact_33_4859
timestamp 1624857261
transform 1 0 22712 0 1 111797
box 0 0 1 1
use contact_33  contact_33_1538
timestamp 1624857261
transform 1 0 22984 0 1 111797
box 0 0 1 1
use contact_33  contact_33_4387
timestamp 1624857261
transform 1 0 23392 0 1 110573
box 0 0 1 1
use contact_33  contact_33_4388
timestamp 1624857261
transform 1 0 23392 0 1 110981
box 0 0 1 1
use contact_33  contact_33_4389
timestamp 1624857261
transform 1 0 23392 0 1 110709
box 0 0 1 1
use contact_33  contact_33_4456
timestamp 1624857261
transform 1 0 23528 0 1 111117
box 0 0 1 1
use contact_33  contact_33_4457
timestamp 1624857261
transform 1 0 23528 0 1 111389
box 0 0 1 1
use contact_33  contact_33_4586
timestamp 1624857261
transform 1 0 23392 0 1 111525
box 0 0 1 1
use contact_33  contact_33_4587
timestamp 1624857261
transform 1 0 23392 0 1 111797
box 0 0 1 1
use contact_33  contact_33_1365
timestamp 1624857261
transform 1 0 28288 0 1 110845
box 0 0 1 1
use contact_33  contact_33_1366
timestamp 1624857261
transform 1 0 28288 0 1 110573
box 0 0 1 1
use contact_33  contact_33_5351
timestamp 1624857261
transform 1 0 1224 0 1 113021
box 0 0 1 1
use contact_13  contact_13_444
timestamp 1624857261
transform 1 0 1801 0 1 111891
box 0 0 1 1
use contact_19  contact_19_444
timestamp 1624857261
transform 1 0 1794 0 1 111900
box 0 0 1 1
use contact_14  contact_14_444
timestamp 1624857261
transform 1 0 1797 0 1 111899
box 0 0 1 1
use contact_13  contact_13_443
timestamp 1624857261
transform 1 0 1801 0 1 112227
box 0 0 1 1
use contact_13  contact_13_442
timestamp 1624857261
transform 1 0 1801 0 1 112563
box 0 0 1 1
use contact_19  contact_19_443
timestamp 1624857261
transform 1 0 1794 0 1 112236
box 0 0 1 1
use contact_19  contact_19_442
timestamp 1624857261
transform 1 0 1794 0 1 112572
box 0 0 1 1
use contact_14  contact_14_443
timestamp 1624857261
transform 1 0 1797 0 1 112235
box 0 0 1 1
use contact_14  contact_14_442
timestamp 1624857261
transform 1 0 1797 0 1 112571
box 0 0 1 1
use contact_13  contact_13_441
timestamp 1624857261
transform 1 0 1801 0 1 112899
box 0 0 1 1
use contact_19  contact_19_441
timestamp 1624857261
transform 1 0 1794 0 1 112908
box 0 0 1 1
use contact_14  contact_14_441
timestamp 1624857261
transform 1 0 1797 0 1 112907
box 0 0 1 1
use contact_7  contact_7_89
timestamp 1624857261
transform 1 0 1793 0 1 112903
box 0 0 1 1
use contact_33  contact_33_1923
timestamp 1624857261
transform 1 0 21760 0 1 112613
box 0 0 1 1
use contact_33  contact_33_1924
timestamp 1624857261
transform 1 0 21760 0 1 112341
box 0 0 1 1
use contact_33  contact_33_2017
timestamp 1624857261
transform 1 0 21896 0 1 112749
box 0 0 1 1
use contact_33  contact_33_2018
timestamp 1624857261
transform 1 0 21896 0 1 113021
box 0 0 1 1
use contact_33  contact_33_2020
timestamp 1624857261
transform 1 0 21896 0 1 113157
box 0 0 1 1
use contact_33  contact_33_2155
timestamp 1624857261
transform 1 0 21896 0 1 112205
box 0 0 1 1
use contact_33  contact_33_2156
timestamp 1624857261
transform 1 0 21896 0 1 111933
box 0 0 1 1
use contact_33  contact_33_4991
timestamp 1624857261
transform 1 0 22304 0 1 111933
box 0 0 1 1
use contact_33  contact_33_4990
timestamp 1624857261
transform 1 0 22304 0 1 112205
box 0 0 1 1
use contact_33  contact_33_1590
timestamp 1624857261
transform 1 0 23120 0 1 112205
box 0 0 1 1
use contact_33  contact_33_1589
timestamp 1624857261
transform 1 0 23120 0 1 111933
box 0 0 1 1
use contact_33  contact_33_4942
timestamp 1624857261
transform 1 0 22168 0 1 112341
box 0 0 1 1
use contact_33  contact_33_1588
timestamp 1624857261
transform 1 0 23120 0 1 112341
box 0 0 1 1
use contact_33  contact_33_4943
timestamp 1624857261
transform 1 0 22168 0 1 112613
box 0 0 1 1
use contact_33  contact_33_1587
timestamp 1624857261
transform 1 0 23120 0 1 112613
box 0 0 1 1
use contact_33  contact_33_1533
timestamp 1624857261
transform 1 0 22984 0 1 112749
box 0 0 1 1
use contact_33  contact_33_5148
timestamp 1624857261
transform 1 0 22168 0 1 113157
box 0 0 1 1
use contact_33  contact_33_4931
timestamp 1624857261
transform 1 0 22440 0 1 113157
box 0 0 1 1
use contact_33  contact_33_1534
timestamp 1624857261
transform 1 0 22984 0 1 113021
box 0 0 1 1
use contact_33  contact_33_4584
timestamp 1624857261
transform 1 0 23392 0 1 112205
box 0 0 1 1
use contact_33  contact_33_4585
timestamp 1624857261
transform 1 0 23392 0 1 111933
box 0 0 1 1
use contact_33  contact_33_4684
timestamp 1624857261
transform 1 0 23392 0 1 113021
box 0 0 1 1
use contact_33  contact_33_4685
timestamp 1624857261
transform 1 0 23392 0 1 112749
box 0 0 1 1
use contact_33  contact_33_4686
timestamp 1624857261
transform 1 0 23528 0 1 112341
box 0 0 1 1
use contact_33  contact_33_4687
timestamp 1624857261
transform 1 0 23528 0 1 112613
box 0 0 1 1
use contact_33  contact_33_1457
timestamp 1624857261
transform 1 0 28424 0 1 112069
box 0 0 1 1
use contact_33  contact_33_1458
timestamp 1624857261
transform 1 0 28424 0 1 112341
box 0 0 1 1
use contact_33  contact_33_1471
timestamp 1624857261
transform 1 0 28288 0 1 113157
box 0 0 1 1
use contact_33  contact_33_1472
timestamp 1624857261
transform 1 0 28288 0 1 112885
box 0 0 1 1
use contact_13  contact_13_440
timestamp 1624857261
transform 1 0 1801 0 1 113235
box 0 0 1 1
use contact_13  contact_13_439
timestamp 1624857261
transform 1 0 1801 0 1 113571
box 0 0 1 1
use contact_19  contact_19_440
timestamp 1624857261
transform 1 0 1794 0 1 113244
box 0 0 1 1
use contact_14  contact_14_440
timestamp 1624857261
transform 1 0 1797 0 1 113243
box 0 0 1 1
use contact_13  contact_13_438
timestamp 1624857261
transform 1 0 1801 0 1 113907
box 0 0 1 1
use contact_19  contact_19_439
timestamp 1624857261
transform 1 0 1794 0 1 113580
box 0 0 1 1
use contact_19  contact_19_438
timestamp 1624857261
transform 1 0 1794 0 1 113916
box 0 0 1 1
use contact_14  contact_14_439
timestamp 1624857261
transform 1 0 1797 0 1 113579
box 0 0 1 1
use contact_14  contact_14_438
timestamp 1624857261
transform 1 0 1797 0 1 113915
box 0 0 1 1
use contact_13  contact_13_437
timestamp 1624857261
transform 1 0 1801 0 1 114243
box 0 0 1 1
use contact_19  contact_19_437
timestamp 1624857261
transform 1 0 1794 0 1 114252
box 0 0 1 1
use contact_14  contact_14_437
timestamp 1624857261
transform 1 0 1797 0 1 114251
box 0 0 1 1
use contact_33  contact_33_1951
timestamp 1624857261
transform 1 0 21760 0 1 113837
box 0 0 1 1
use contact_33  contact_33_1952
timestamp 1624857261
transform 1 0 21760 0 1 113565
box 0 0 1 1
use contact_33  contact_33_2019
timestamp 1624857261
transform 1 0 21896 0 1 113429
box 0 0 1 1
use contact_33  contact_33_1807
timestamp 1624857261
transform 1 0 22984 0 1 114517
box 0 0 1 1
use contact_33  contact_33_1808
timestamp 1624857261
transform 1 0 22984 0 1 114245
box 0 0 1 1
use contact_33  contact_33_1899
timestamp 1624857261
transform 1 0 23120 0 1 114109
box 0 0 1 1
use contact_33  contact_33_1900
timestamp 1624857261
transform 1 0 23120 0 1 113837
box 0 0 1 1
use contact_33  contact_33_4926
timestamp 1624857261
transform 1 0 22440 0 1 113837
box 0 0 1 1
use contact_33  contact_33_4927
timestamp 1624857261
transform 1 0 22440 0 1 114109
box 0 0 1 1
use contact_33  contact_33_4930
timestamp 1624857261
transform 1 0 22440 0 1 113429
box 0 0 1 1
use contact_33  contact_33_5149
timestamp 1624857261
transform 1 0 22168 0 1 113429
box 0 0 1 1
use contact_33  contact_33_4428
timestamp 1624857261
transform 1 0 23392 0 1 114517
box 0 0 1 1
use contact_33  contact_33_4429
timestamp 1624857261
transform 1 0 23392 0 1 114245
box 0 0 1 1
use contact_33  contact_33_4514
timestamp 1624857261
transform 1 0 23392 0 1 114109
box 0 0 1 1
use contact_33  contact_33_4515
timestamp 1624857261
transform 1 0 23392 0 1 113837
box 0 0 1 1
use contact_33  contact_33_1455
timestamp 1624857261
transform 1 0 28560 0 1 113973
box 0 0 1 1
use contact_33  contact_33_1456
timestamp 1624857261
transform 1 0 28560 0 1 113701
box 0 0 1 1
use contact_33  contact_33_1459
timestamp 1624857261
transform 1 0 28288 0 1 113293
box 0 0 1 1
use contact_33  contact_33_1460
timestamp 1624857261
transform 1 0 28288 0 1 113701
box 0 0 1 1
use contact_33  contact_33_5352
timestamp 1624857261
transform 1 0 1224 0 1 114653
box 0 0 1 1
use contact_13  contact_13_436
timestamp 1624857261
transform 1 0 1801 0 1 114579
box 0 0 1 1
use contact_13  contact_13_435
timestamp 1624857261
transform 1 0 1801 0 1 114915
box 0 0 1 1
use contact_19  contact_19_436
timestamp 1624857261
transform 1 0 1794 0 1 114588
box 0 0 1 1
use contact_14  contact_14_436
timestamp 1624857261
transform 1 0 1797 0 1 114587
box 0 0 1 1
use contact_7  contact_7_88
timestamp 1624857261
transform 1 0 1793 0 1 114583
box 0 0 1 1
use contact_13  contact_13_434
timestamp 1624857261
transform 1 0 1801 0 1 115251
box 0 0 1 1
use contact_19  contact_19_435
timestamp 1624857261
transform 1 0 1794 0 1 114924
box 0 0 1 1
use contact_19  contact_19_434
timestamp 1624857261
transform 1 0 1794 0 1 115260
box 0 0 1 1
use contact_14  contact_14_435
timestamp 1624857261
transform 1 0 1797 0 1 114923
box 0 0 1 1
use contact_14  contact_14_434
timestamp 1624857261
transform 1 0 1797 0 1 115259
box 0 0 1 1
use contact_13  contact_13_433
timestamp 1624857261
transform 1 0 1801 0 1 115587
box 0 0 1 1
use contact_19  contact_19_433
timestamp 1624857261
transform 1 0 1794 0 1 115596
box 0 0 1 1
use contact_14  contact_14_433
timestamp 1624857261
transform 1 0 1797 0 1 115595
box 0 0 1 1
use contact_33  contact_33_2113
timestamp 1624857261
transform 1 0 21760 0 1 115741
box 0 0 1 1
use contact_33  contact_33_2114
timestamp 1624857261
transform 1 0 21760 0 1 115469
box 0 0 1 1
use contact_33  contact_33_2125
timestamp 1624857261
transform 1 0 21896 0 1 115877
box 0 0 1 1
use contact_33  contact_33_2171
timestamp 1624857261
transform 1 0 21896 0 1 115333
box 0 0 1 1
use contact_33  contact_33_2172
timestamp 1624857261
transform 1 0 21896 0 1 115061
box 0 0 1 1
use contact_33  contact_33_1895
timestamp 1624857261
transform 1 0 23120 0 1 114653
box 0 0 1 1
use contact_33  contact_33_4835
timestamp 1624857261
transform 1 0 22712 0 1 115061
box 0 0 1 1
use contact_33  contact_33_1898
timestamp 1624857261
transform 1 0 23120 0 1 115061
box 0 0 1 1
use contact_33  contact_33_1896
timestamp 1624857261
transform 1 0 23120 0 1 114925
box 0 0 1 1
use contact_33  contact_33_5169
timestamp 1624857261
transform 1 0 22168 0 1 115469
box 0 0 1 1
use contact_33  contact_33_4834
timestamp 1624857261
transform 1 0 22712 0 1 115333
box 0 0 1 1
use contact_33  contact_33_4807
timestamp 1624857261
transform 1 0 22576 0 1 115469
box 0 0 1 1
use contact_33  contact_33_1897
timestamp 1624857261
transform 1 0 23120 0 1 115333
box 0 0 1 1
use contact_33  contact_33_1704
timestamp 1624857261
transform 1 0 23120 0 1 115469
box 0 0 1 1
use contact_33  contact_33_5168
timestamp 1624857261
transform 1 0 22168 0 1 115741
box 0 0 1 1
use contact_33  contact_33_4923
timestamp 1624857261
transform 1 0 22440 0 1 115877
box 0 0 1 1
use contact_33  contact_33_4806
timestamp 1624857261
transform 1 0 22576 0 1 115741
box 0 0 1 1
use contact_33  contact_33_1703
timestamp 1624857261
transform 1 0 23120 0 1 115741
box 0 0 1 1
use contact_33  contact_33_1581
timestamp 1624857261
transform 1 0 22984 0 1 115877
box 0 0 1 1
use contact_33  contact_33_4350
timestamp 1624857261
transform 1 0 23528 0 1 115469
box 0 0 1 1
use contact_33  contact_33_4351
timestamp 1624857261
transform 1 0 23528 0 1 115741
box 0 0 1 1
use contact_33  contact_33_4360
timestamp 1624857261
transform 1 0 23392 0 1 115333
box 0 0 1 1
use contact_33  contact_33_4361
timestamp 1624857261
transform 1 0 23392 0 1 115061
box 0 0 1 1
use contact_33  contact_33_4380
timestamp 1624857261
transform 1 0 23528 0 1 114925
box 0 0 1 1
use contact_33  contact_33_4381
timestamp 1624857261
transform 1 0 23528 0 1 114653
box 0 0 1 1
use contact_33  contact_33_4530
timestamp 1624857261
transform 1 0 23392 0 1 115877
box 0 0 1 1
use contact_33  contact_33_5303
timestamp 1624857261
transform 1 0 1224 0 1 116285
box 0 0 1 1
use contact_13  contact_13_432
timestamp 1624857261
transform 1 0 1801 0 1 115923
box 0 0 1 1
use contact_13  contact_13_431
timestamp 1624857261
transform 1 0 1801 0 1 116259
box 0 0 1 1
use contact_19  contact_19_432
timestamp 1624857261
transform 1 0 1794 0 1 115932
box 0 0 1 1
use contact_19  contact_19_431
timestamp 1624857261
transform 1 0 1794 0 1 116268
box 0 0 1 1
use contact_14  contact_14_432
timestamp 1624857261
transform 1 0 1797 0 1 115931
box 0 0 1 1
use contact_14  contact_14_431
timestamp 1624857261
transform 1 0 1797 0 1 116267
box 0 0 1 1
use contact_7  contact_7_87
timestamp 1624857261
transform 1 0 1793 0 1 116263
box 0 0 1 1
use contact_13  contact_13_430
timestamp 1624857261
transform 1 0 1801 0 1 116595
box 0 0 1 1
use contact_19  contact_19_430
timestamp 1624857261
transform 1 0 1794 0 1 116604
box 0 0 1 1
use contact_14  contact_14_430
timestamp 1624857261
transform 1 0 1797 0 1 116603
box 0 0 1 1
use contact_13  contact_13_429
timestamp 1624857261
transform 1 0 1801 0 1 116931
box 0 0 1 1
use contact_19  contact_19_429
timestamp 1624857261
transform 1 0 1794 0 1 116940
box 0 0 1 1
use contact_14  contact_14_429
timestamp 1624857261
transform 1 0 1797 0 1 116939
box 0 0 1 1
use contact_33  contact_33_1930
timestamp 1624857261
transform 1 0 21896 0 1 117101
box 0 0 1 1
use contact_33  contact_33_2049
timestamp 1624857261
transform 1 0 21760 0 1 116965
box 0 0 1 1
use contact_33  contact_33_2050
timestamp 1624857261
transform 1 0 21760 0 1 116693
box 0 0 1 1
use contact_33  contact_33_2126
timestamp 1624857261
transform 1 0 21896 0 1 116149
box 0 0 1 1
use contact_33  contact_33_2127
timestamp 1624857261
transform 1 0 21896 0 1 116557
box 0 0 1 1
use contact_33  contact_33_2128
timestamp 1624857261
transform 1 0 21896 0 1 116285
box 0 0 1 1
use contact_33  contact_33_1582
timestamp 1624857261
transform 1 0 22984 0 1 116149
box 0 0 1 1
use contact_33  contact_33_1755
timestamp 1624857261
transform 1 0 23120 0 1 116285
box 0 0 1 1
use contact_33  contact_33_1756
timestamp 1624857261
transform 1 0 23120 0 1 116557
box 0 0 1 1
use contact_33  contact_33_1805
timestamp 1624857261
transform 1 0 22984 0 1 116693
box 0 0 1 1
use contact_33  contact_33_1806
timestamp 1624857261
transform 1 0 22984 0 1 116965
box 0 0 1 1
use contact_33  contact_33_4922
timestamp 1624857261
transform 1 0 22440 0 1 116149
box 0 0 1 1
use contact_33  contact_33_5064
timestamp 1624857261
transform 1 0 22440 0 1 117101
box 0 0 1 1
use contact_33  contact_33_4356
timestamp 1624857261
transform 1 0 23528 0 1 116965
box 0 0 1 1
use contact_33  contact_33_4357
timestamp 1624857261
transform 1 0 23528 0 1 116693
box 0 0 1 1
use contact_33  contact_33_4531
timestamp 1624857261
transform 1 0 23392 0 1 116149
box 0 0 1 1
use contact_33  contact_33_4532
timestamp 1624857261
transform 1 0 23392 0 1 116557
box 0 0 1 1
use contact_33  contact_33_4533
timestamp 1624857261
transform 1 0 23392 0 1 116285
box 0 0 1 1
use contact_33  contact_33_1407
timestamp 1624857261
transform 1 0 28560 0 1 116693
box 0 0 1 1
use contact_33  contact_33_1408
timestamp 1624857261
transform 1 0 28560 0 1 116285
box 0 0 1 1
use contact_33  contact_33_1415
timestamp 1624857261
transform 1 0 28424 0 1 116829
box 0 0 1 1
use contact_33  contact_33_1416
timestamp 1624857261
transform 1 0 28424 0 1 117101
box 0 0 1 1
use contact_33  contact_33_1486
timestamp 1624857261
transform 1 0 28560 0 1 117101
box 0 0 1 1
use contact_33  contact_33_5350
timestamp 1624857261
transform 1 0 1224 0 1 118053
box 0 0 1 1
use contact_13  contact_13_428
timestamp 1624857261
transform 1 0 1801 0 1 117267
box 0 0 1 1
use contact_13  contact_13_427
timestamp 1624857261
transform 1 0 1801 0 1 117603
box 0 0 1 1
use contact_19  contact_19_428
timestamp 1624857261
transform 1 0 1794 0 1 117276
box 0 0 1 1
use contact_14  contact_14_428
timestamp 1624857261
transform 1 0 1797 0 1 117275
box 0 0 1 1
use contact_13  contact_13_426
timestamp 1624857261
transform 1 0 1801 0 1 117939
box 0 0 1 1
use contact_19  contact_19_427
timestamp 1624857261
transform 1 0 1794 0 1 117612
box 0 0 1 1
use contact_14  contact_14_427
timestamp 1624857261
transform 1 0 1797 0 1 117611
box 0 0 1 1
use contact_7  contact_7_86
timestamp 1624857261
transform 1 0 1793 0 1 117943
box 0 0 1 1
use contact_13  contact_13_425
timestamp 1624857261
transform 1 0 1801 0 1 118275
box 0 0 1 1
use contact_19  contact_19_426
timestamp 1624857261
transform 1 0 1794 0 1 117948
box 0 0 1 1
use contact_19  contact_19_425
timestamp 1624857261
transform 1 0 1794 0 1 118284
box 0 0 1 1
use contact_14  contact_14_426
timestamp 1624857261
transform 1 0 1797 0 1 117947
box 0 0 1 1
use contact_14  contact_14_425
timestamp 1624857261
transform 1 0 1797 0 1 118283
box 0 0 1 1
use contact_13  contact_13_424
timestamp 1624857261
transform 1 0 1801 0 1 118611
box 0 0 1 1
use contact_19  contact_19_424
timestamp 1624857261
transform 1 0 1794 0 1 118620
box 0 0 1 1
use contact_14  contact_14_424
timestamp 1624857261
transform 1 0 1797 0 1 118619
box 0 0 1 1
use contact_33  contact_33_1929
timestamp 1624857261
transform 1 0 21896 0 1 117373
box 0 0 1 1
use contact_33  contact_33_2103
timestamp 1624857261
transform 1 0 21760 0 1 117509
box 0 0 1 1
use contact_33  contact_33_2104
timestamp 1624857261
transform 1 0 21760 0 1 117781
box 0 0 1 1
use contact_33  contact_33_1857
timestamp 1624857261
transform 1 0 22984 0 1 118189
box 0 0 1 1
use contact_33  contact_33_1858
timestamp 1624857261
transform 1 0 22984 0 1 118461
box 0 0 1 1
use contact_33  contact_33_1860
timestamp 1624857261
transform 1 0 22984 0 1 118597
box 0 0 1 1
use contact_33  contact_33_4890
timestamp 1624857261
transform 1 0 22576 0 1 118597
box 0 0 1 1
use contact_33  contact_33_5065
timestamp 1624857261
transform 1 0 22440 0 1 117373
box 0 0 1 1
use contact_33  contact_33_5076
timestamp 1624857261
transform 1 0 22168 0 1 117781
box 0 0 1 1
use contact_33  contact_33_5077
timestamp 1624857261
transform 1 0 22168 0 1 118053
box 0 0 1 1
use contact_33  contact_33_4675
timestamp 1624857261
transform 1 0 23392 0 1 118597
box 0 0 1 1
use contact_33  contact_33_4676
timestamp 1624857261
transform 1 0 23392 0 1 118189
box 0 0 1 1
use contact_33  contact_33_4677
timestamp 1624857261
transform 1 0 23392 0 1 118461
box 0 0 1 1
use contact_33  contact_33_1375
timestamp 1624857261
transform 1 0 28424 0 1 118053
box 0 0 1 1
use contact_33  contact_33_1376
timestamp 1624857261
transform 1 0 28424 0 1 118461
box 0 0 1 1
use contact_33  contact_33_1381
timestamp 1624857261
transform 1 0 28560 0 1 118461
box 0 0 1 1
use contact_33  contact_33_1383
timestamp 1624857261
transform 1 0 28424 0 1 117917
box 0 0 1 1
use contact_33  contact_33_1384
timestamp 1624857261
transform 1 0 28424 0 1 117645
box 0 0 1 1
use contact_33  contact_33_1485
timestamp 1624857261
transform 1 0 28560 0 1 117509
box 0 0 1 1
use contact_33  contact_33_5336
timestamp 1624857261
transform 1 0 1224 0 1 119685
box 0 0 1 1
use contact_13  contact_13_423
timestamp 1624857261
transform 1 0 1801 0 1 118947
box 0 0 1 1
use contact_19  contact_19_423
timestamp 1624857261
transform 1 0 1794 0 1 118956
box 0 0 1 1
use contact_14  contact_14_423
timestamp 1624857261
transform 1 0 1797 0 1 118955
box 0 0 1 1
use contact_13  contact_13_422
timestamp 1624857261
transform 1 0 1801 0 1 119283
box 0 0 1 1
use contact_19  contact_19_422
timestamp 1624857261
transform 1 0 1794 0 1 119292
box 0 0 1 1
use contact_14  contact_14_422
timestamp 1624857261
transform 1 0 1797 0 1 119291
box 0 0 1 1
use contact_13  contact_13_421
timestamp 1624857261
transform 1 0 1801 0 1 119619
box 0 0 1 1
use contact_19  contact_19_421
timestamp 1624857261
transform 1 0 1794 0 1 119628
box 0 0 1 1
use contact_14  contact_14_421
timestamp 1624857261
transform 1 0 1797 0 1 119627
box 0 0 1 1
use contact_7  contact_7_85
timestamp 1624857261
transform 1 0 1793 0 1 119623
box 0 0 1 1
use contact_13  contact_13_420
timestamp 1624857261
transform 1 0 1801 0 1 119955
box 0 0 1 1
use contact_19  contact_19_420
timestamp 1624857261
transform 1 0 1794 0 1 119964
box 0 0 1 1
use contact_14  contact_14_420
timestamp 1624857261
transform 1 0 1797 0 1 119963
box 0 0 1 1
use contact_33  contact_33_2071
timestamp 1624857261
transform 1 0 21760 0 1 119277
box 0 0 1 1
use contact_33  contact_33_2072
timestamp 1624857261
transform 1 0 21760 0 1 119005
box 0 0 1 1
use contact_33  contact_33_2137
timestamp 1624857261
transform 1 0 21896 0 1 119413
box 0 0 1 1
use contact_33  contact_33_2138
timestamp 1624857261
transform 1 0 21896 0 1 119685
box 0 0 1 1
use contact_33  contact_33_2140
timestamp 1624857261
transform 1 0 21760 0 1 119821
box 0 0 1 1
use contact_33  contact_33_5138
timestamp 1624857261
transform 1 0 22304 0 1 119005
box 0 0 1 1
use contact_33  contact_33_5136
timestamp 1624857261
transform 1 0 22440 0 1 119005
box 0 0 1 1
use contact_33  contact_33_4891
timestamp 1624857261
transform 1 0 22576 0 1 118869
box 0 0 1 1
use contact_33  contact_33_1859
timestamp 1624857261
transform 1 0 22984 0 1 118869
box 0 0 1 1
use contact_33  contact_33_1649
timestamp 1624857261
transform 1 0 23120 0 1 119005
box 0 0 1 1
use contact_33  contact_33_5139
timestamp 1624857261
transform 1 0 22304 0 1 119277
box 0 0 1 1
use contact_33  contact_33_5137
timestamp 1624857261
transform 1 0 22440 0 1 119277
box 0 0 1 1
use contact_33  contact_33_1650
timestamp 1624857261
transform 1 0 23120 0 1 119277
box 0 0 1 1
use contact_33  contact_33_1826
timestamp 1624857261
transform 1 0 22984 0 1 119685
box 0 0 1 1
use contact_33  contact_33_1825
timestamp 1624857261
transform 1 0 22984 0 1 119413
box 0 0 1 1
use contact_33  contact_33_4778
timestamp 1624857261
transform 1 0 22576 0 1 119821
box 0 0 1 1
use contact_33  contact_33_1828
timestamp 1624857261
transform 1 0 23120 0 1 119821
box 0 0 1 1
use contact_33  contact_33_4470
timestamp 1624857261
transform 1 0 23392 0 1 119005
box 0 0 1 1
use contact_33  contact_33_4471
timestamp 1624857261
transform 1 0 23392 0 1 119277
box 0 0 1 1
use contact_33  contact_33_4657
timestamp 1624857261
transform 1 0 23528 0 1 119821
box 0 0 1 1
use contact_33  contact_33_4658
timestamp 1624857261
transform 1 0 23392 0 1 119413
box 0 0 1 1
use contact_33  contact_33_4659
timestamp 1624857261
transform 1 0 23392 0 1 119685
box 0 0 1 1
use contact_33  contact_33_4674
timestamp 1624857261
transform 1 0 23392 0 1 118869
box 0 0 1 1
use contact_33  contact_33_1382
timestamp 1624857261
transform 1 0 28560 0 1 118733
box 0 0 1 1
use contact_13  contact_13_419
timestamp 1624857261
transform 1 0 1801 0 1 120291
box 0 0 1 1
use contact_19  contact_19_419
timestamp 1624857261
transform 1 0 1794 0 1 120300
box 0 0 1 1
use contact_14  contact_14_419
timestamp 1624857261
transform 1 0 1797 0 1 120299
box 0 0 1 1
use contact_13  contact_13_418
timestamp 1624857261
transform 1 0 1801 0 1 120627
box 0 0 1 1
use contact_19  contact_19_418
timestamp 1624857261
transform 1 0 1794 0 1 120636
box 0 0 1 1
use contact_14  contact_14_418
timestamp 1624857261
transform 1 0 1797 0 1 120635
box 0 0 1 1
use contact_13  contact_13_417
timestamp 1624857261
transform 1 0 1801 0 1 120963
box 0 0 1 1
use contact_19  contact_19_417
timestamp 1624857261
transform 1 0 1794 0 1 120972
box 0 0 1 1
use contact_14  contact_14_417
timestamp 1624857261
transform 1 0 1797 0 1 120971
box 0 0 1 1
use contact_13  contact_13_416
timestamp 1624857261
transform 1 0 1801 0 1 121299
box 0 0 1 1
use contact_19  contact_19_416
timestamp 1624857261
transform 1 0 1794 0 1 121308
box 0 0 1 1
use contact_14  contact_14_416
timestamp 1624857261
transform 1 0 1797 0 1 121307
box 0 0 1 1
use contact_7  contact_7_84
timestamp 1624857261
transform 1 0 1793 0 1 121303
box 0 0 1 1
use contact_33  contact_33_2051
timestamp 1624857261
transform 1 0 21760 0 1 120501
box 0 0 1 1
use contact_33  contact_33_2052
timestamp 1624857261
transform 1 0 21760 0 1 120229
box 0 0 1 1
use contact_33  contact_33_2139
timestamp 1624857261
transform 1 0 21760 0 1 120093
box 0 0 1 1
use contact_33  contact_33_1827
timestamp 1624857261
transform 1 0 23120 0 1 120093
box 0 0 1 1
use contact_33  contact_33_1847
timestamp 1624857261
transform 1 0 22984 0 1 120229
box 0 0 1 1
use contact_33  contact_33_1848
timestamp 1624857261
transform 1 0 22984 0 1 120501
box 0 0 1 1
use contact_33  contact_33_4776
timestamp 1624857261
transform 1 0 22576 0 1 120501
box 0 0 1 1
use contact_33  contact_33_4777
timestamp 1624857261
transform 1 0 22576 0 1 120229
box 0 0 1 1
use contact_33  contact_33_4779
timestamp 1624857261
transform 1 0 22576 0 1 120093
box 0 0 1 1
use contact_33  contact_33_5182
timestamp 1624857261
transform 1 0 22304 0 1 120229
box 0 0 1 1
use contact_33  contact_33_5183
timestamp 1624857261
transform 1 0 22304 0 1 120501
box 0 0 1 1
use contact_33  contact_33_4518
timestamp 1624857261
transform 1 0 23392 0 1 120229
box 0 0 1 1
use contact_33  contact_33_4519
timestamp 1624857261
transform 1 0 23392 0 1 120501
box 0 0 1 1
use contact_33  contact_33_4656
timestamp 1624857261
transform 1 0 23528 0 1 120093
box 0 0 1 1
use contact_33  contact_33_1484
timestamp 1624857261
transform 1 0 29920 0 1 121045
box 0 0 1 1
use contact_33  contact_33_5330
timestamp 1624857261
transform 1 0 1224 0 1 121453
box 0 0 1 1
use contact_13  contact_13_415
timestamp 1624857261
transform 1 0 1801 0 1 121635
box 0 0 1 1
use contact_19  contact_19_415
timestamp 1624857261
transform 1 0 1794 0 1 121644
box 0 0 1 1
use contact_14  contact_14_415
timestamp 1624857261
transform 1 0 1797 0 1 121643
box 0 0 1 1
use contact_13  contact_13_414
timestamp 1624857261
transform 1 0 1801 0 1 121971
box 0 0 1 1
use contact_19  contact_19_414
timestamp 1624857261
transform 1 0 1794 0 1 121980
box 0 0 1 1
use contact_14  contact_14_414
timestamp 1624857261
transform 1 0 1797 0 1 121979
box 0 0 1 1
use contact_13  contact_13_413
timestamp 1624857261
transform 1 0 1801 0 1 122307
box 0 0 1 1
use contact_19  contact_19_413
timestamp 1624857261
transform 1 0 1794 0 1 122316
box 0 0 1 1
use contact_14  contact_14_413
timestamp 1624857261
transform 1 0 1797 0 1 122315
box 0 0 1 1
use contact_13  contact_13_412
timestamp 1624857261
transform 1 0 1801 0 1 122643
box 0 0 1 1
use contact_19  contact_19_412
timestamp 1624857261
transform 1 0 1794 0 1 122652
box 0 0 1 1
use contact_14  contact_14_412
timestamp 1624857261
transform 1 0 1797 0 1 122651
box 0 0 1 1
use contact_33  contact_33_4304
timestamp 1624857261
transform 1 0 29648 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4305
timestamp 1624857261
transform 1 0 29648 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4288
timestamp 1624857261
transform 1 0 30464 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4289
timestamp 1624857261
transform 1 0 30464 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4302
timestamp 1624857261
transform 1 0 30328 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4303
timestamp 1624857261
transform 1 0 30328 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4280
timestamp 1624857261
transform 1 0 32776 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4281
timestamp 1624857261
transform 1 0 32776 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4282
timestamp 1624857261
transform 1 0 31688 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4283
timestamp 1624857261
transform 1 0 31688 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4254
timestamp 1624857261
transform 1 0 34136 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4255
timestamp 1624857261
transform 1 0 34136 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4260
timestamp 1624857261
transform 1 0 33456 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4261
timestamp 1624857261
transform 1 0 33456 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4236
timestamp 1624857261
transform 1 0 35360 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4237
timestamp 1624857261
transform 1 0 35360 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4250
timestamp 1624857261
transform 1 0 34680 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4251
timestamp 1624857261
transform 1 0 34680 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4226
timestamp 1624857261
transform 1 0 35904 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4227
timestamp 1624857261
transform 1 0 35904 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4220
timestamp 1624857261
transform 1 0 37128 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4221
timestamp 1624857261
transform 1 0 37128 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4192
timestamp 1624857261
transform 1 0 39576 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4193
timestamp 1624857261
transform 1 0 39576 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4196
timestamp 1624857261
transform 1 0 39168 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4197
timestamp 1624857261
transform 1 0 39168 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4204
timestamp 1624857261
transform 1 0 38488 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4205
timestamp 1624857261
transform 1 0 38488 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4176
timestamp 1624857261
transform 1 0 40936 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4177
timestamp 1624857261
transform 1 0 40936 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4182
timestamp 1624857261
transform 1 0 40392 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4183
timestamp 1624857261
transform 1 0 40392 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4170
timestamp 1624857261
transform 1 0 42160 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4171
timestamp 1624857261
transform 1 0 42160 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4152
timestamp 1624857261
transform 1 0 43384 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4153
timestamp 1624857261
transform 1 0 43384 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4154
timestamp 1624857261
transform 1 0 42840 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4155
timestamp 1624857261
transform 1 0 42840 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4138
timestamp 1624857261
transform 1 0 44608 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4139
timestamp 1624857261
transform 1 0 44608 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4144
timestamp 1624857261
transform 1 0 44064 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4145
timestamp 1624857261
transform 1 0 44064 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4148
timestamp 1624857261
transform 1 0 43928 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4149
timestamp 1624857261
transform 1 0 43928 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4128
timestamp 1624857261
transform 1 0 45696 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4129
timestamp 1624857261
transform 1 0 45696 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4118
timestamp 1624857261
transform 1 0 46648 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4119
timestamp 1624857261
transform 1 0 46648 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4090
timestamp 1624857261
transform 1 0 49096 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4091
timestamp 1624857261
transform 1 0 49096 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4096
timestamp 1624857261
transform 1 0 48416 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4097
timestamp 1624857261
transform 1 0 48416 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4100
timestamp 1624857261
transform 1 0 47872 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4101
timestamp 1624857261
transform 1 0 47872 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4072
timestamp 1624857261
transform 1 0 50320 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4073
timestamp 1624857261
transform 1 0 50320 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4084
timestamp 1624857261
transform 1 0 49232 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4085
timestamp 1624857261
transform 1 0 49232 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4068
timestamp 1624857261
transform 1 0 50864 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4069
timestamp 1624857261
transform 1 0 50864 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4046
timestamp 1624857261
transform 1 0 52904 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4047
timestamp 1624857261
transform 1 0 52904 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4060
timestamp 1624857261
transform 1 0 52224 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4061
timestamp 1624857261
transform 1 0 52224 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4040
timestamp 1624857261
transform 1 0 54128 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4041
timestamp 1624857261
transform 1 0 54128 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4042
timestamp 1624857261
transform 1 0 53312 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4043
timestamp 1624857261
transform 1 0 53312 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4016
timestamp 1624857261
transform 1 0 55352 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4017
timestamp 1624857261
transform 1 0 55352 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4032
timestamp 1624857261
transform 1 0 54672 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4033
timestamp 1624857261
transform 1 0 54672 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4004
timestamp 1624857261
transform 1 0 57120 0 1 121589
box 0 0 1 1
use contact_33  contact_33_4005
timestamp 1624857261
transform 1 0 57120 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4008
timestamp 1624857261
transform 1 0 56712 0 1 121997
box 0 0 1 1
use contact_33  contact_33_4009
timestamp 1624857261
transform 1 0 56712 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3984
timestamp 1624857261
transform 1 0 58072 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3985
timestamp 1624857261
transform 1 0 58072 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3978
timestamp 1624857261
transform 1 0 59160 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3979
timestamp 1624857261
transform 1 0 59160 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3960
timestamp 1624857261
transform 1 0 60928 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3961
timestamp 1624857261
transform 1 0 60928 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3948
timestamp 1624857261
transform 1 0 62152 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3949
timestamp 1624857261
transform 1 0 62152 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3954
timestamp 1624857261
transform 1 0 61608 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3955
timestamp 1624857261
transform 1 0 61608 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3926
timestamp 1624857261
transform 1 0 64056 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3927
timestamp 1624857261
transform 1 0 64056 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3928
timestamp 1624857261
transform 1 0 63376 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3929
timestamp 1624857261
transform 1 0 63376 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3932
timestamp 1624857261
transform 1 0 62832 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3933
timestamp 1624857261
transform 1 0 62832 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3916
timestamp 1624857261
transform 1 0 64600 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3917
timestamp 1624857261
transform 1 0 64600 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3904
timestamp 1624857261
transform 1 0 65688 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3905
timestamp 1624857261
transform 1 0 65688 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3896
timestamp 1624857261
transform 1 0 67184 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3897
timestamp 1624857261
transform 1 0 67184 0 1 121997
box 0 0 1 1
use contact_33  contact_33_5348
timestamp 1624857261
transform 1 0 1224 0 1 123085
box 0 0 1 1
use contact_13  contact_13_411
timestamp 1624857261
transform 1 0 1801 0 1 122979
box 0 0 1 1
use contact_19  contact_19_411
timestamp 1624857261
transform 1 0 1794 0 1 122988
box 0 0 1 1
use contact_14  contact_14_411
timestamp 1624857261
transform 1 0 1797 0 1 122987
box 0 0 1 1
use contact_7  contact_7_83
timestamp 1624857261
transform 1 0 1793 0 1 122983
box 0 0 1 1
use contact_13  contact_13_410
timestamp 1624857261
transform 1 0 1801 0 1 123315
box 0 0 1 1
use contact_19  contact_19_410
timestamp 1624857261
transform 1 0 1794 0 1 123324
box 0 0 1 1
use contact_14  contact_14_410
timestamp 1624857261
transform 1 0 1797 0 1 123323
box 0 0 1 1
use contact_13  contact_13_409
timestamp 1624857261
transform 1 0 1801 0 1 123651
box 0 0 1 1
use contact_19  contact_19_409
timestamp 1624857261
transform 1 0 1794 0 1 123660
box 0 0 1 1
use contact_14  contact_14_409
timestamp 1624857261
transform 1 0 1797 0 1 123659
box 0 0 1 1
use contact_13  contact_13_408
timestamp 1624857261
transform 1 0 1801 0 1 123987
box 0 0 1 1
use contact_19  contact_19_408
timestamp 1624857261
transform 1 0 1794 0 1 123996
box 0 0 1 1
use contact_14  contact_14_408
timestamp 1624857261
transform 1 0 1797 0 1 123995
box 0 0 1 1
use contact_33  contact_33_1347
timestamp 1624857261
transform 1 0 30056 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1483
timestamp 1624857261
transform 1 0 29920 0 1 123493
box 0 0 1 1
use contact_33  contact_33_1337
timestamp 1624857261
transform 1 0 32640 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1325
timestamp 1624857261
transform 1 0 35088 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1311
timestamp 1624857261
transform 1 0 37400 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1301
timestamp 1624857261
transform 1 0 40120 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1287
timestamp 1624857261
transform 1 0 42568 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1277
timestamp 1624857261
transform 1 0 44880 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1263
timestamp 1624857261
transform 1 0 47464 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1251
timestamp 1624857261
transform 1 0 50048 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1239
timestamp 1624857261
transform 1 0 52496 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1229
timestamp 1624857261
transform 1 0 55080 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1217
timestamp 1624857261
transform 1 0 57528 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1205
timestamp 1624857261
transform 1 0 59976 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1191
timestamp 1624857261
transform 1 0 62560 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1179
timestamp 1624857261
transform 1 0 64872 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1169
timestamp 1624857261
transform 1 0 67456 0 1 123765
box 0 0 1 1
use contact_33  contact_33_5354
timestamp 1624857261
transform 1 0 1224 0 1 124581
box 0 0 1 1
use contact_13  contact_13_407
timestamp 1624857261
transform 1 0 1801 0 1 124323
box 0 0 1 1
use contact_19  contact_19_407
timestamp 1624857261
transform 1 0 1794 0 1 124332
box 0 0 1 1
use contact_14  contact_14_407
timestamp 1624857261
transform 1 0 1797 0 1 124331
box 0 0 1 1
use contact_13  contact_13_406
timestamp 1624857261
transform 1 0 1801 0 1 124659
box 0 0 1 1
use contact_19  contact_19_406
timestamp 1624857261
transform 1 0 1794 0 1 124668
box 0 0 1 1
use contact_14  contact_14_406
timestamp 1624857261
transform 1 0 1797 0 1 124667
box 0 0 1 1
use contact_7  contact_7_82
timestamp 1624857261
transform 1 0 1793 0 1 124663
box 0 0 1 1
use contact_13  contact_13_405
timestamp 1624857261
transform 1 0 1801 0 1 124995
box 0 0 1 1
use contact_19  contact_19_405
timestamp 1624857261
transform 1 0 1794 0 1 125004
box 0 0 1 1
use contact_14  contact_14_405
timestamp 1624857261
transform 1 0 1797 0 1 125003
box 0 0 1 1
use contact_13  contact_13_404
timestamp 1624857261
transform 1 0 1801 0 1 125331
box 0 0 1 1
use contact_19  contact_19_404
timestamp 1624857261
transform 1 0 1794 0 1 125340
box 0 0 1 1
use contact_14  contact_14_404
timestamp 1624857261
transform 1 0 1797 0 1 125339
box 0 0 1 1
use contact_33  contact_33_5378
timestamp 1624857261
transform 1 0 1224 0 1 126349
box 0 0 1 1
use contact_13  contact_13_403
timestamp 1624857261
transform 1 0 1801 0 1 125667
box 0 0 1 1
use contact_19  contact_19_403
timestamp 1624857261
transform 1 0 1794 0 1 125676
box 0 0 1 1
use contact_14  contact_14_403
timestamp 1624857261
transform 1 0 1797 0 1 125675
box 0 0 1 1
use contact_13  contact_13_402
timestamp 1624857261
transform 1 0 1801 0 1 126003
box 0 0 1 1
use contact_19  contact_19_402
timestamp 1624857261
transform 1 0 1794 0 1 126012
box 0 0 1 1
use contact_14  contact_14_402
timestamp 1624857261
transform 1 0 1797 0 1 126011
box 0 0 1 1
use contact_13  contact_13_401
timestamp 1624857261
transform 1 0 1801 0 1 126339
box 0 0 1 1
use contact_19  contact_19_401
timestamp 1624857261
transform 1 0 1794 0 1 126348
box 0 0 1 1
use contact_14  contact_14_401
timestamp 1624857261
transform 1 0 1797 0 1 126347
box 0 0 1 1
use contact_7  contact_7_81
timestamp 1624857261
transform 1 0 1793 0 1 126343
box 0 0 1 1
use contact_13  contact_13_400
timestamp 1624857261
transform 1 0 1801 0 1 126675
box 0 0 1 1
use contact_19  contact_19_400
timestamp 1624857261
transform 1 0 1794 0 1 126684
box 0 0 1 1
use contact_14  contact_14_400
timestamp 1624857261
transform 1 0 1797 0 1 126683
box 0 0 1 1
use contact_33  contact_33_1348
timestamp 1624857261
transform 1 0 30056 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1353
timestamp 1624857261
transform 1 0 29920 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4297
timestamp 1624857261
transform 1 0 29784 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1338
timestamp 1624857261
transform 1 0 32640 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1341
timestamp 1624857261
transform 1 0 32504 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4269
timestamp 1624857261
transform 1 0 32368 0 1 126485
box 0 0 1 1
use contact_33  contact_33_4292
timestamp 1624857261
transform 1 0 32096 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1326
timestamp 1624857261
transform 1 0 35088 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1329
timestamp 1624857261
transform 1 0 34952 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4241
timestamp 1624857261
transform 1 0 34816 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1312
timestamp 1624857261
transform 1 0 37400 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1317
timestamp 1624857261
transform 1 0 37264 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4213
timestamp 1624857261
transform 1 0 37400 0 1 126485
box 0 0 1 1
use contact_33  contact_33_4239
timestamp 1624857261
transform 1 0 37128 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1302
timestamp 1624857261
transform 1 0 40120 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1303
timestamp 1624857261
transform 1 0 39984 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4187
timestamp 1624857261
transform 1 0 39848 0 1 126485
box 0 0 1 1
use contact_33  contact_33_4163
timestamp 1624857261
transform 1 0 42160 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1288
timestamp 1624857261
transform 1 0 42568 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1293
timestamp 1624857261
transform 1 0 42432 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1278
timestamp 1624857261
transform 1 0 44880 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1279
timestamp 1624857261
transform 1 0 44744 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4131
timestamp 1624857261
transform 1 0 44880 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1264
timestamp 1624857261
transform 1 0 47464 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1267
timestamp 1624857261
transform 1 0 47328 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4111
timestamp 1624857261
transform 1 0 47192 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1252
timestamp 1624857261
transform 1 0 50048 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1255
timestamp 1624857261
transform 1 0 49912 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4077
timestamp 1624857261
transform 1 0 49776 0 1 126485
box 0 0 1 1
use contact_33  contact_33_4106
timestamp 1624857261
transform 1 0 49504 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1240
timestamp 1624857261
transform 1 0 52496 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1243
timestamp 1624857261
transform 1 0 52360 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4053
timestamp 1624857261
transform 1 0 52224 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1230
timestamp 1624857261
transform 1 0 55080 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1231
timestamp 1624857261
transform 1 0 54944 0 1 125669
box 0 0 1 1
use contact_33  contact_33_4023
timestamp 1624857261
transform 1 0 54808 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3993
timestamp 1624857261
transform 1 0 57256 0 1 126485
box 0 0 1 1
use contact_33  contact_33_4021
timestamp 1624857261
transform 1 0 56984 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1218
timestamp 1624857261
transform 1 0 57528 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1219
timestamp 1624857261
transform 1 0 57392 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1206
timestamp 1624857261
transform 1 0 59976 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1207
timestamp 1624857261
transform 1 0 59704 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3965
timestamp 1624857261
transform 1 0 59840 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3991
timestamp 1624857261
transform 1 0 59568 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1192
timestamp 1624857261
transform 1 0 62560 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1195
timestamp 1624857261
transform 1 0 62424 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3941
timestamp 1624857261
transform 1 0 62288 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1180
timestamp 1624857261
transform 1 0 64872 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1183
timestamp 1624857261
transform 1 0 64736 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3911
timestamp 1624857261
transform 1 0 64872 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1170
timestamp 1624857261
transform 1 0 67456 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1171
timestamp 1624857261
transform 1 0 67320 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3889
timestamp 1624857261
transform 1 0 67184 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3906
timestamp 1624857261
transform 1 0 67048 0 1 126485
box 0 0 1 1
use contact_33  contact_33_5373
timestamp 1624857261
transform 1 0 1224 0 1 128117
box 0 0 1 1
use contact_13  contact_13_399
timestamp 1624857261
transform 1 0 1801 0 1 127011
box 0 0 1 1
use contact_19  contact_19_399
timestamp 1624857261
transform 1 0 1794 0 1 127020
box 0 0 1 1
use contact_14  contact_14_399
timestamp 1624857261
transform 1 0 1797 0 1 127019
box 0 0 1 1
use contact_13  contact_13_398
timestamp 1624857261
transform 1 0 1801 0 1 127347
box 0 0 1 1
use contact_19  contact_19_398
timestamp 1624857261
transform 1 0 1794 0 1 127356
box 0 0 1 1
use contact_14  contact_14_398
timestamp 1624857261
transform 1 0 1797 0 1 127355
box 0 0 1 1
use contact_13  contact_13_397
timestamp 1624857261
transform 1 0 1801 0 1 127683
box 0 0 1 1
use contact_19  contact_19_397
timestamp 1624857261
transform 1 0 1794 0 1 127692
box 0 0 1 1
use contact_14  contact_14_397
timestamp 1624857261
transform 1 0 1797 0 1 127691
box 0 0 1 1
use contact_13  contact_13_396
timestamp 1624857261
transform 1 0 1801 0 1 128019
box 0 0 1 1
use contact_19  contact_19_396
timestamp 1624857261
transform 1 0 1794 0 1 128028
box 0 0 1 1
use contact_14  contact_14_396
timestamp 1624857261
transform 1 0 1797 0 1 128027
box 0 0 1 1
use contact_7  contact_7_80
timestamp 1624857261
transform 1 0 1793 0 1 128023
box 0 0 1 1
use contact_7  contact_7_359
timestamp 1624857261
transform 1 0 29557 0 1 127542
box 0 0 1 1
use contact_19  contact_19_965
timestamp 1624857261
transform 1 0 29558 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1354
timestamp 1624857261
transform 1 0 29920 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4296
timestamp 1624857261
transform 1 0 29784 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5449
timestamp 1624857261
transform 1 0 29648 0 1 127573
box 0 0 1 1
use contact_7  contact_7_358
timestamp 1624857261
transform 1 0 32053 0 1 127542
box 0 0 1 1
use contact_19  contact_19_964
timestamp 1624857261
transform 1 0 32054 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1342
timestamp 1624857261
transform 1 0 32504 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4268
timestamp 1624857261
transform 1 0 32368 0 1 127165
box 0 0 1 1
use contact_33  contact_33_4293
timestamp 1624857261
transform 1 0 32096 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5448
timestamp 1624857261
transform 1 0 31960 0 1 127573
box 0 0 1 1
use contact_7  contact_7_357
timestamp 1624857261
transform 1 0 34549 0 1 127542
box 0 0 1 1
use contact_19  contact_19_963
timestamp 1624857261
transform 1 0 34550 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1330
timestamp 1624857261
transform 1 0 34952 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4240
timestamp 1624857261
transform 1 0 34816 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5447
timestamp 1624857261
transform 1 0 34544 0 1 127573
box 0 0 1 1
use contact_7  contact_7_356
timestamp 1624857261
transform 1 0 37045 0 1 127542
box 0 0 1 1
use contact_19  contact_19_962
timestamp 1624857261
transform 1 0 37046 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1318
timestamp 1624857261
transform 1 0 37264 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4212
timestamp 1624857261
transform 1 0 37400 0 1 127165
box 0 0 1 1
use contact_33  contact_33_4238
timestamp 1624857261
transform 1 0 37128 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5446
timestamp 1624857261
transform 1 0 36992 0 1 127573
box 0 0 1 1
use contact_7  contact_7_355
timestamp 1624857261
transform 1 0 39541 0 1 127542
box 0 0 1 1
use contact_19  contact_19_961
timestamp 1624857261
transform 1 0 39542 0 1 127547
box 0 0 1 1
use contact_33  contact_33_5445
timestamp 1624857261
transform 1 0 39576 0 1 127573
box 0 0 1 1
use contact_33  contact_33_1304
timestamp 1624857261
transform 1 0 39984 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4186
timestamp 1624857261
transform 1 0 39848 0 1 127165
box 0 0 1 1
use contact_7  contact_7_354
timestamp 1624857261
transform 1 0 42037 0 1 127542
box 0 0 1 1
use contact_19  contact_19_960
timestamp 1624857261
transform 1 0 42038 0 1 127547
box 0 0 1 1
use contact_33  contact_33_4162
timestamp 1624857261
transform 1 0 42160 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5444
timestamp 1624857261
transform 1 0 42024 0 1 127573
box 0 0 1 1
use contact_33  contact_33_1294
timestamp 1624857261
transform 1 0 42432 0 1 127437
box 0 0 1 1
use contact_7  contact_7_353
timestamp 1624857261
transform 1 0 44533 0 1 127542
box 0 0 1 1
use contact_19  contact_19_959
timestamp 1624857261
transform 1 0 44534 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1280
timestamp 1624857261
transform 1 0 44880 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4130
timestamp 1624857261
transform 1 0 44880 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5443
timestamp 1624857261
transform 1 0 44608 0 1 127573
box 0 0 1 1
use contact_7  contact_7_352
timestamp 1624857261
transform 1 0 47029 0 1 127542
box 0 0 1 1
use contact_19  contact_19_958
timestamp 1624857261
transform 1 0 47030 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1268
timestamp 1624857261
transform 1 0 47328 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4110
timestamp 1624857261
transform 1 0 47192 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5442
timestamp 1624857261
transform 1 0 47056 0 1 127573
box 0 0 1 1
use contact_7  contact_7_351
timestamp 1624857261
transform 1 0 49525 0 1 127542
box 0 0 1 1
use contact_19  contact_19_957
timestamp 1624857261
transform 1 0 49526 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1256
timestamp 1624857261
transform 1 0 49912 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4076
timestamp 1624857261
transform 1 0 49776 0 1 127165
box 0 0 1 1
use contact_33  contact_33_4107
timestamp 1624857261
transform 1 0 49504 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5441
timestamp 1624857261
transform 1 0 49504 0 1 127573
box 0 0 1 1
use contact_7  contact_7_350
timestamp 1624857261
transform 1 0 52021 0 1 127542
box 0 0 1 1
use contact_19  contact_19_956
timestamp 1624857261
transform 1 0 52022 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1244
timestamp 1624857261
transform 1 0 52360 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4052
timestamp 1624857261
transform 1 0 52224 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5440
timestamp 1624857261
transform 1 0 51952 0 1 127573
box 0 0 1 1
use contact_7  contact_7_349
timestamp 1624857261
transform 1 0 54517 0 1 127542
box 0 0 1 1
use contact_19  contact_19_955
timestamp 1624857261
transform 1 0 54518 0 1 127547
box 0 0 1 1
use contact_33  contact_33_5439
timestamp 1624857261
transform 1 0 54400 0 1 127573
box 0 0 1 1
use contact_33  contact_33_1232
timestamp 1624857261
transform 1 0 54944 0 1 127437
box 0 0 1 1
use contact_33  contact_33_4022
timestamp 1624857261
transform 1 0 54808 0 1 127165
box 0 0 1 1
use contact_7  contact_7_348
timestamp 1624857261
transform 1 0 57013 0 1 127542
box 0 0 1 1
use contact_19  contact_19_954
timestamp 1624857261
transform 1 0 57014 0 1 127547
box 0 0 1 1
use contact_33  contact_33_3992
timestamp 1624857261
transform 1 0 57256 0 1 127165
box 0 0 1 1
use contact_33  contact_33_4020
timestamp 1624857261
transform 1 0 56984 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5438
timestamp 1624857261
transform 1 0 56984 0 1 127573
box 0 0 1 1
use contact_33  contact_33_1220
timestamp 1624857261
transform 1 0 57392 0 1 127437
box 0 0 1 1
use contact_7  contact_7_347
timestamp 1624857261
transform 1 0 59509 0 1 127542
box 0 0 1 1
use contact_19  contact_19_953
timestamp 1624857261
transform 1 0 59510 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1208
timestamp 1624857261
transform 1 0 59840 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3964
timestamp 1624857261
transform 1 0 59840 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3990
timestamp 1624857261
transform 1 0 59568 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5437
timestamp 1624857261
transform 1 0 59568 0 1 127573
box 0 0 1 1
use contact_7  contact_7_346
timestamp 1624857261
transform 1 0 62005 0 1 127542
box 0 0 1 1
use contact_19  contact_19_952
timestamp 1624857261
transform 1 0 62006 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1196
timestamp 1624857261
transform 1 0 62424 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3940
timestamp 1624857261
transform 1 0 62288 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5436
timestamp 1624857261
transform 1 0 62016 0 1 127573
box 0 0 1 1
use contact_7  contact_7_345
timestamp 1624857261
transform 1 0 64501 0 1 127542
box 0 0 1 1
use contact_19  contact_19_951
timestamp 1624857261
transform 1 0 64502 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1184
timestamp 1624857261
transform 1 0 64736 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3910
timestamp 1624857261
transform 1 0 64872 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5435
timestamp 1624857261
transform 1 0 64600 0 1 127573
box 0 0 1 1
use contact_7  contact_7_344
timestamp 1624857261
transform 1 0 66997 0 1 127542
box 0 0 1 1
use contact_19  contact_19_950
timestamp 1624857261
transform 1 0 66998 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1172
timestamp 1624857261
transform 1 0 67320 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3888
timestamp 1624857261
transform 1 0 67184 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3907
timestamp 1624857261
transform 1 0 67048 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5434
timestamp 1624857261
transform 1 0 67048 0 1 127573
box 0 0 1 1
use contact_13  contact_13_395
timestamp 1624857261
transform 1 0 1801 0 1 128355
box 0 0 1 1
use contact_19  contact_19_395
timestamp 1624857261
transform 1 0 1794 0 1 128364
box 0 0 1 1
use contact_14  contact_14_395
timestamp 1624857261
transform 1 0 1797 0 1 128363
box 0 0 1 1
use contact_13  contact_13_394
timestamp 1624857261
transform 1 0 1801 0 1 128691
box 0 0 1 1
use contact_19  contact_19_394
timestamp 1624857261
transform 1 0 1794 0 1 128700
box 0 0 1 1
use contact_14  contact_14_394
timestamp 1624857261
transform 1 0 1797 0 1 128699
box 0 0 1 1
use contact_13  contact_13_393
timestamp 1624857261
transform 1 0 1801 0 1 129027
box 0 0 1 1
use contact_19  contact_19_393
timestamp 1624857261
transform 1 0 1794 0 1 129036
box 0 0 1 1
use contact_14  contact_14_393
timestamp 1624857261
transform 1 0 1797 0 1 129035
box 0 0 1 1
use contact_13  contact_13_392
timestamp 1624857261
transform 1 0 1801 0 1 129363
box 0 0 1 1
use contact_19  contact_19_392
timestamp 1624857261
transform 1 0 1794 0 1 129372
box 0 0 1 1
use contact_14  contact_14_392
timestamp 1624857261
transform 1 0 1797 0 1 129371
box 0 0 1 1
use contact_33  contact_33_5342
timestamp 1624857261
transform 1 0 1224 0 1 129749
box 0 0 1 1
use contact_13  contact_13_391
timestamp 1624857261
transform 1 0 1801 0 1 129699
box 0 0 1 1
use contact_19  contact_19_391
timestamp 1624857261
transform 1 0 1794 0 1 129708
box 0 0 1 1
use contact_14  contact_14_391
timestamp 1624857261
transform 1 0 1797 0 1 129707
box 0 0 1 1
use contact_7  contact_7_79
timestamp 1624857261
transform 1 0 1793 0 1 129703
box 0 0 1 1
use contact_13  contact_13_390
timestamp 1624857261
transform 1 0 1801 0 1 130035
box 0 0 1 1
use contact_19  contact_19_390
timestamp 1624857261
transform 1 0 1794 0 1 130044
box 0 0 1 1
use contact_14  contact_14_390
timestamp 1624857261
transform 1 0 1797 0 1 130043
box 0 0 1 1
use contact_13  contact_13_389
timestamp 1624857261
transform 1 0 1801 0 1 130371
box 0 0 1 1
use contact_19  contact_19_389
timestamp 1624857261
transform 1 0 1794 0 1 130380
box 0 0 1 1
use contact_14  contact_14_389
timestamp 1624857261
transform 1 0 1797 0 1 130379
box 0 0 1 1
use contact_13  contact_13_388
timestamp 1624857261
transform 1 0 1801 0 1 130707
box 0 0 1 1
use contact_19  contact_19_388
timestamp 1624857261
transform 1 0 1794 0 1 130716
box 0 0 1 1
use contact_14  contact_14_388
timestamp 1624857261
transform 1 0 1797 0 1 130715
box 0 0 1 1
use contact_13  contact_13_387
timestamp 1624857261
transform 1 0 1801 0 1 131043
box 0 0 1 1
use contact_19  contact_19_387
timestamp 1624857261
transform 1 0 1794 0 1 131052
box 0 0 1 1
use contact_14  contact_14_387
timestamp 1624857261
transform 1 0 1797 0 1 131051
box 0 0 1 1
use contact_13  contact_13_386
timestamp 1624857261
transform 1 0 1801 0 1 131379
box 0 0 1 1
use contact_19  contact_19_386
timestamp 1624857261
transform 1 0 1794 0 1 131388
box 0 0 1 1
use contact_14  contact_14_386
timestamp 1624857261
transform 1 0 1797 0 1 131387
box 0 0 1 1
use contact_7  contact_7_78
timestamp 1624857261
transform 1 0 1793 0 1 131383
box 0 0 1 1
use contact_33  contact_33_5370
timestamp 1624857261
transform 1 0 2040 0 1 131517
box 0 0 1 1
use contact_38  contact_38_0
timestamp 1624857261
transform 1 0 1730 0 1 131937
box 0 0 192 192
use contact_33  contact_33_5369
timestamp 1624857261
transform 1 0 2040 0 1 131925
box 0 0 1 1
use contact_33  contact_33_5293
timestamp 1624857261
transform 1 0 2176 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1172
timestamp 1624857261
transform 1 0 2137 0 1 131992
box 0 0 1 1
use contact_19  contact_19_852
timestamp 1624857261
transform 1 0 2130 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1172
timestamp 1624857261
transform 1 0 2133 0 1 132000
box 0 0 1 1
use contact_7  contact_7_236
timestamp 1624857261
transform 1 0 2129 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1171
timestamp 1624857261
transform 1 0 2473 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1171
timestamp 1624857261
transform 1 0 2469 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1170
timestamp 1624857261
transform 1 0 2809 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1170
timestamp 1624857261
transform 1 0 2805 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1169
timestamp 1624857261
transform 1 0 3145 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1169
timestamp 1624857261
transform 1 0 3141 0 1 132000
box 0 0 1 1
use contact_33  contact_33_5289
timestamp 1624857261
transform 1 0 3672 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1168
timestamp 1624857261
transform 1 0 3481 0 1 131992
box 0 0 1 1
use contact_19  contact_19_851
timestamp 1624857261
transform 1 0 3810 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1168
timestamp 1624857261
transform 1 0 3477 0 1 132000
box 0 0 1 1
use contact_7  contact_7_235
timestamp 1624857261
transform 1 0 3809 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1167
timestamp 1624857261
transform 1 0 3817 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1166
timestamp 1624857261
transform 1 0 4153 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1167
timestamp 1624857261
transform 1 0 3813 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1166
timestamp 1624857261
transform 1 0 4149 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1165
timestamp 1624857261
transform 1 0 4489 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1165
timestamp 1624857261
transform 1 0 4485 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1164
timestamp 1624857261
transform 1 0 4825 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1163
timestamp 1624857261
transform 1 0 5161 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1164
timestamp 1624857261
transform 1 0 4821 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1163
timestamp 1624857261
transform 1 0 5157 0 1 132000
box 0 0 1 1
use contact_33  contact_33_5287
timestamp 1624857261
transform 1 0 5440 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1162
timestamp 1624857261
transform 1 0 5497 0 1 131992
box 0 0 1 1
use contact_19  contact_19_850
timestamp 1624857261
transform 1 0 5490 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1162
timestamp 1624857261
transform 1 0 5493 0 1 132000
box 0 0 1 1
use contact_7  contact_7_234
timestamp 1624857261
transform 1 0 5489 0 1 131996
box 0 0 1 1
use contact_14  contact_14_1158
timestamp 1624857261
transform 1 0 6837 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1159
timestamp 1624857261
transform 1 0 6501 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1160
timestamp 1624857261
transform 1 0 6165 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1161
timestamp 1624857261
transform 1 0 5829 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1158
timestamp 1624857261
transform 1 0 6841 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1159
timestamp 1624857261
transform 1 0 6505 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1160
timestamp 1624857261
transform 1 0 6169 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1161
timestamp 1624857261
transform 1 0 5833 0 1 131992
box 0 0 1 1
use contact_33  contact_33_5281
timestamp 1624857261
transform 1 0 7208 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1157
timestamp 1624857261
transform 1 0 7177 0 1 131992
box 0 0 1 1
use contact_19  contact_19_849
timestamp 1624857261
transform 1 0 7170 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1157
timestamp 1624857261
transform 1 0 7173 0 1 132000
box 0 0 1 1
use contact_7  contact_7_233
timestamp 1624857261
transform 1 0 7169 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1156
timestamp 1624857261
transform 1 0 7513 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1155
timestamp 1624857261
transform 1 0 7849 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1156
timestamp 1624857261
transform 1 0 7509 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1155
timestamp 1624857261
transform 1 0 7845 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1154
timestamp 1624857261
transform 1 0 8185 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1154
timestamp 1624857261
transform 1 0 8181 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1153
timestamp 1624857261
transform 1 0 8521 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1153
timestamp 1624857261
transform 1 0 8517 0 1 132000
box 0 0 1 1
use contact_33  contact_33_5277
timestamp 1624857261
transform 1 0 8976 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1152
timestamp 1624857261
transform 1 0 8857 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1151
timestamp 1624857261
transform 1 0 9193 0 1 131992
box 0 0 1 1
use contact_19  contact_19_848
timestamp 1624857261
transform 1 0 8850 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1152
timestamp 1624857261
transform 1 0 8853 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1151
timestamp 1624857261
transform 1 0 9189 0 1 132000
box 0 0 1 1
use contact_7  contact_7_232
timestamp 1624857261
transform 1 0 8849 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1150
timestamp 1624857261
transform 1 0 9529 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1150
timestamp 1624857261
transform 1 0 9525 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1149
timestamp 1624857261
transform 1 0 9865 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1148
timestamp 1624857261
transform 1 0 10201 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1149
timestamp 1624857261
transform 1 0 9861 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1148
timestamp 1624857261
transform 1 0 10197 0 1 132000
box 0 0 1 1
use contact_33  contact_33_5273
timestamp 1624857261
transform 1 0 10472 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1147
timestamp 1624857261
transform 1 0 10537 0 1 131992
box 0 0 1 1
use contact_19  contact_19_847
timestamp 1624857261
transform 1 0 10530 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1147
timestamp 1624857261
transform 1 0 10533 0 1 132000
box 0 0 1 1
use contact_7  contact_7_231
timestamp 1624857261
transform 1 0 10529 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1146
timestamp 1624857261
transform 1 0 10873 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1146
timestamp 1624857261
transform 1 0 10869 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1145
timestamp 1624857261
transform 1 0 11209 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1144
timestamp 1624857261
transform 1 0 11545 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1145
timestamp 1624857261
transform 1 0 11205 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1144
timestamp 1624857261
transform 1 0 11541 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1143
timestamp 1624857261
transform 1 0 11881 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1143
timestamp 1624857261
transform 1 0 11877 0 1 132000
box 0 0 1 1
use contact_33  contact_33_5269
timestamp 1624857261
transform 1 0 12104 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1142
timestamp 1624857261
transform 1 0 12217 0 1 131992
box 0 0 1 1
use contact_19  contact_19_846
timestamp 1624857261
transform 1 0 12210 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1142
timestamp 1624857261
transform 1 0 12213 0 1 132000
box 0 0 1 1
use contact_7  contact_7_230
timestamp 1624857261
transform 1 0 12209 0 1 131996
box 0 0 1 1
use contact_14  contact_14_1138
timestamp 1624857261
transform 1 0 13557 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1139
timestamp 1624857261
transform 1 0 13221 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1140
timestamp 1624857261
transform 1 0 12885 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1141
timestamp 1624857261
transform 1 0 12549 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1138
timestamp 1624857261
transform 1 0 13561 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1139
timestamp 1624857261
transform 1 0 13225 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1140
timestamp 1624857261
transform 1 0 12889 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1141
timestamp 1624857261
transform 1 0 12553 0 1 131992
box 0 0 1 1
use contact_33  contact_33_5265
timestamp 1624857261
transform 1 0 13872 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1137
timestamp 1624857261
transform 1 0 13897 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1136
timestamp 1624857261
transform 1 0 14233 0 1 131992
box 0 0 1 1
use contact_19  contact_19_845
timestamp 1624857261
transform 1 0 13890 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1137
timestamp 1624857261
transform 1 0 13893 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1136
timestamp 1624857261
transform 1 0 14229 0 1 132000
box 0 0 1 1
use contact_7  contact_7_229
timestamp 1624857261
transform 1 0 13889 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1135
timestamp 1624857261
transform 1 0 14569 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1135
timestamp 1624857261
transform 1 0 14565 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1134
timestamp 1624857261
transform 1 0 14905 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1134
timestamp 1624857261
transform 1 0 14901 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1133
timestamp 1624857261
transform 1 0 15241 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1132
timestamp 1624857261
transform 1 0 15577 0 1 131992
box 0 0 1 1
use contact_7  contact_7_228
timestamp 1624857261
transform 1 0 15569 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1131
timestamp 1624857261
transform 1 0 15913 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1130
timestamp 1624857261
transform 1 0 16249 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1129
timestamp 1624857261
transform 1 0 16585 0 1 131992
box 0 0 1 1
use contact_19  contact_19_844
timestamp 1624857261
transform 1 0 15570 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1133
timestamp 1624857261
transform 1 0 15237 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1132
timestamp 1624857261
transform 1 0 15573 0 1 132000
box 0 0 1 1
use contact_33  contact_33_5245
timestamp 1624857261
transform 1 0 15640 0 1 132061
box 0 0 1 1
use contact_14  contact_14_1131
timestamp 1624857261
transform 1 0 15909 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1130
timestamp 1624857261
transform 1 0 16245 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1129
timestamp 1624857261
transform 1 0 16581 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1128
timestamp 1624857261
transform 1 0 16921 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1128
timestamp 1624857261
transform 1 0 16917 0 1 132000
box 0 0 1 1
use contact_33  contact_33_5239
timestamp 1624857261
transform 1 0 17136 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1127
timestamp 1624857261
transform 1 0 17257 0 1 131992
box 0 0 1 1
use contact_19  contact_19_843
timestamp 1624857261
transform 1 0 17250 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1127
timestamp 1624857261
transform 1 0 17253 0 1 132000
box 0 0 1 1
use contact_7  contact_7_227
timestamp 1624857261
transform 1 0 17249 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1126
timestamp 1624857261
transform 1 0 17593 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1126
timestamp 1624857261
transform 1 0 17589 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1125
timestamp 1624857261
transform 1 0 17929 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1125
timestamp 1624857261
transform 1 0 17925 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1124
timestamp 1624857261
transform 1 0 18265 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1124
timestamp 1624857261
transform 1 0 18261 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1123
timestamp 1624857261
transform 1 0 18601 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1123
timestamp 1624857261
transform 1 0 18597 0 1 132000
box 0 0 1 1
use contact_33  contact_33_5227
timestamp 1624857261
transform 1 0 18904 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1122
timestamp 1624857261
transform 1 0 18937 0 1 131992
box 0 0 1 1
use contact_19  contact_19_842
timestamp 1624857261
transform 1 0 18930 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1122
timestamp 1624857261
transform 1 0 18933 0 1 132000
box 0 0 1 1
use contact_7  contact_7_226
timestamp 1624857261
transform 1 0 18929 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1121
timestamp 1624857261
transform 1 0 19273 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1121
timestamp 1624857261
transform 1 0 19269 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1120
timestamp 1624857261
transform 1 0 19609 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1120
timestamp 1624857261
transform 1 0 19605 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1119
timestamp 1624857261
transform 1 0 19945 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1119
timestamp 1624857261
transform 1 0 19941 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1118
timestamp 1624857261
transform 1 0 20281 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1118
timestamp 1624857261
transform 1 0 20277 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1117
timestamp 1624857261
transform 1 0 20617 0 1 131992
box 0 0 1 1
use contact_19  contact_19_841
timestamp 1624857261
transform 1 0 20610 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1117
timestamp 1624857261
transform 1 0 20613 0 1 132000
box 0 0 1 1
use contact_7  contact_7_225
timestamp 1624857261
transform 1 0 20609 0 1 131996
box 0 0 1 1
use contact_14  contact_14_1113
timestamp 1624857261
transform 1 0 21957 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1114
timestamp 1624857261
transform 1 0 21621 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1115
timestamp 1624857261
transform 1 0 21285 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1116
timestamp 1624857261
transform 1 0 20949 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1113
timestamp 1624857261
transform 1 0 21961 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1114
timestamp 1624857261
transform 1 0 21625 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1115
timestamp 1624857261
transform 1 0 21289 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1116
timestamp 1624857261
transform 1 0 20953 0 1 131992
box 0 0 1 1
use contact_33  contact_33_5203
timestamp 1624857261
transform 1 0 20672 0 1 132061
box 0 0 1 1
use contact_33  contact_33_4903
timestamp 1624857261
transform 1 0 22168 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1112
timestamp 1624857261
transform 1 0 22297 0 1 131992
box 0 0 1 1
use contact_19  contact_19_840
timestamp 1624857261
transform 1 0 22290 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1112
timestamp 1624857261
transform 1 0 22293 0 1 132000
box 0 0 1 1
use contact_7  contact_7_224
timestamp 1624857261
transform 1 0 22289 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1111
timestamp 1624857261
transform 1 0 22633 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1111
timestamp 1624857261
transform 1 0 22629 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1110
timestamp 1624857261
transform 1 0 22969 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1110
timestamp 1624857261
transform 1 0 22965 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1109
timestamp 1624857261
transform 1 0 23305 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1109
timestamp 1624857261
transform 1 0 23301 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1108
timestamp 1624857261
transform 1 0 23641 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1108
timestamp 1624857261
transform 1 0 23637 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4325
timestamp 1624857261
transform 1 0 23936 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1107
timestamp 1624857261
transform 1 0 23977 0 1 131992
box 0 0 1 1
use contact_19  contact_19_839
timestamp 1624857261
transform 1 0 23970 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1107
timestamp 1624857261
transform 1 0 23973 0 1 132000
box 0 0 1 1
use contact_7  contact_7_223
timestamp 1624857261
transform 1 0 23969 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1106
timestamp 1624857261
transform 1 0 24313 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1106
timestamp 1624857261
transform 1 0 24309 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1105
timestamp 1624857261
transform 1 0 24649 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1105
timestamp 1624857261
transform 1 0 24645 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1104
timestamp 1624857261
transform 1 0 24985 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1104
timestamp 1624857261
transform 1 0 24981 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1103
timestamp 1624857261
transform 1 0 25321 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1103
timestamp 1624857261
transform 1 0 25317 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4321
timestamp 1624857261
transform 1 0 25704 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1102
timestamp 1624857261
transform 1 0 25657 0 1 131992
box 0 0 1 1
use contact_19  contact_19_838
timestamp 1624857261
transform 1 0 25650 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1102
timestamp 1624857261
transform 1 0 25653 0 1 132000
box 0 0 1 1
use contact_7  contact_7_222
timestamp 1624857261
transform 1 0 25649 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1101
timestamp 1624857261
transform 1 0 25993 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1101
timestamp 1624857261
transform 1 0 25989 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1100
timestamp 1624857261
transform 1 0 26329 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1100
timestamp 1624857261
transform 1 0 26325 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1099
timestamp 1624857261
transform 1 0 26665 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1099
timestamp 1624857261
transform 1 0 26661 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4317
timestamp 1624857261
transform 1 0 27200 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1098
timestamp 1624857261
transform 1 0 27001 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1097
timestamp 1624857261
transform 1 0 27337 0 1 131992
box 0 0 1 1
use contact_19  contact_19_837
timestamp 1624857261
transform 1 0 27330 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1098
timestamp 1624857261
transform 1 0 26997 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1097
timestamp 1624857261
transform 1 0 27333 0 1 132000
box 0 0 1 1
use contact_7  contact_7_221
timestamp 1624857261
transform 1 0 27329 0 1 131996
box 0 0 1 1
use contact_14  contact_14_1093
timestamp 1624857261
transform 1 0 28677 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1094
timestamp 1624857261
transform 1 0 28341 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1095
timestamp 1624857261
transform 1 0 28005 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1096
timestamp 1624857261
transform 1 0 27669 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1093
timestamp 1624857261
transform 1 0 28681 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1094
timestamp 1624857261
transform 1 0 28345 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1095
timestamp 1624857261
transform 1 0 28009 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1096
timestamp 1624857261
transform 1 0 27673 0 1 131992
box 0 0 1 1
use contact_33  contact_33_4309
timestamp 1624857261
transform 1 0 28968 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1092
timestamp 1624857261
transform 1 0 29017 0 1 131992
box 0 0 1 1
use contact_19  contact_19_836
timestamp 1624857261
transform 1 0 29010 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1092
timestamp 1624857261
transform 1 0 29013 0 1 132000
box 0 0 1 1
use contact_7  contact_7_220
timestamp 1624857261
transform 1 0 29009 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1091
timestamp 1624857261
transform 1 0 29353 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1091
timestamp 1624857261
transform 1 0 29349 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1090
timestamp 1624857261
transform 1 0 29689 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1089
timestamp 1624857261
transform 1 0 30025 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1090
timestamp 1624857261
transform 1 0 29685 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1089
timestamp 1624857261
transform 1 0 30021 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1088
timestamp 1624857261
transform 1 0 30361 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1088
timestamp 1624857261
transform 1 0 30357 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4287
timestamp 1624857261
transform 1 0 30736 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1087
timestamp 1624857261
transform 1 0 30697 0 1 131992
box 0 0 1 1
use contact_19  contact_19_835
timestamp 1624857261
transform 1 0 30690 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1087
timestamp 1624857261
transform 1 0 30693 0 1 132000
box 0 0 1 1
use contact_7  contact_7_219
timestamp 1624857261
transform 1 0 30689 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1086
timestamp 1624857261
transform 1 0 31033 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1085
timestamp 1624857261
transform 1 0 31369 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1086
timestamp 1624857261
transform 1 0 31029 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1085
timestamp 1624857261
transform 1 0 31365 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1084
timestamp 1624857261
transform 1 0 31705 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1084
timestamp 1624857261
transform 1 0 31701 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4265
timestamp 1624857261
transform 1 0 32232 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1083
timestamp 1624857261
transform 1 0 32041 0 1 131992
box 0 0 1 1
use contact_19  contact_19_834
timestamp 1624857261
transform 1 0 32370 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1083
timestamp 1624857261
transform 1 0 32037 0 1 132000
box 0 0 1 1
use contact_7  contact_7_218
timestamp 1624857261
transform 1 0 32369 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1082
timestamp 1624857261
transform 1 0 32377 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1081
timestamp 1624857261
transform 1 0 32713 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1082
timestamp 1624857261
transform 1 0 32373 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1081
timestamp 1624857261
transform 1 0 32709 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1080
timestamp 1624857261
transform 1 0 33049 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1080
timestamp 1624857261
transform 1 0 33045 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1079
timestamp 1624857261
transform 1 0 33385 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1078
timestamp 1624857261
transform 1 0 33721 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1079
timestamp 1624857261
transform 1 0 33381 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1078
timestamp 1624857261
transform 1 0 33717 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4257
timestamp 1624857261
transform 1 0 34136 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1077
timestamp 1624857261
transform 1 0 34057 0 1 131992
box 0 0 1 1
use contact_19  contact_19_833
timestamp 1624857261
transform 1 0 34050 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1077
timestamp 1624857261
transform 1 0 34053 0 1 132000
box 0 0 1 1
use contact_7  contact_7_217
timestamp 1624857261
transform 1 0 34049 0 1 131996
box 0 0 1 1
use contact_14  contact_14_1073
timestamp 1624857261
transform 1 0 35397 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1074
timestamp 1624857261
transform 1 0 35061 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1075
timestamp 1624857261
transform 1 0 34725 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1076
timestamp 1624857261
transform 1 0 34389 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1073
timestamp 1624857261
transform 1 0 35401 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1074
timestamp 1624857261
transform 1 0 35065 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1075
timestamp 1624857261
transform 1 0 34729 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1076
timestamp 1624857261
transform 1 0 34393 0 1 131992
box 0 0 1 1
use contact_33  contact_33_4229
timestamp 1624857261
transform 1 0 35632 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1072
timestamp 1624857261
transform 1 0 35737 0 1 131992
box 0 0 1 1
use contact_19  contact_19_832
timestamp 1624857261
transform 1 0 35730 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1072
timestamp 1624857261
transform 1 0 35733 0 1 132000
box 0 0 1 1
use contact_7  contact_7_216
timestamp 1624857261
transform 1 0 35729 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1071
timestamp 1624857261
transform 1 0 36073 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1070
timestamp 1624857261
transform 1 0 36409 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1071
timestamp 1624857261
transform 1 0 36069 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1070
timestamp 1624857261
transform 1 0 36405 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1069
timestamp 1624857261
transform 1 0 36745 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1069
timestamp 1624857261
transform 1 0 36741 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4209
timestamp 1624857261
transform 1 0 37400 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1068
timestamp 1624857261
transform 1 0 37081 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1068
timestamp 1624857261
transform 1 0 37077 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1067
timestamp 1624857261
transform 1 0 37417 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1066
timestamp 1624857261
transform 1 0 37753 0 1 131992
box 0 0 1 1
use contact_19  contact_19_831
timestamp 1624857261
transform 1 0 37410 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1067
timestamp 1624857261
transform 1 0 37413 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1066
timestamp 1624857261
transform 1 0 37749 0 1 132000
box 0 0 1 1
use contact_7  contact_7_215
timestamp 1624857261
transform 1 0 37409 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1065
timestamp 1624857261
transform 1 0 38089 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1065
timestamp 1624857261
transform 1 0 38085 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1064
timestamp 1624857261
transform 1 0 38425 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1063
timestamp 1624857261
transform 1 0 38761 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1064
timestamp 1624857261
transform 1 0 38421 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1063
timestamp 1624857261
transform 1 0 38757 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4203
timestamp 1624857261
transform 1 0 39168 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1062
timestamp 1624857261
transform 1 0 39097 0 1 131992
box 0 0 1 1
use contact_19  contact_19_830
timestamp 1624857261
transform 1 0 39090 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1062
timestamp 1624857261
transform 1 0 39093 0 1 132000
box 0 0 1 1
use contact_7  contact_7_214
timestamp 1624857261
transform 1 0 39089 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1061
timestamp 1624857261
transform 1 0 39433 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1061
timestamp 1624857261
transform 1 0 39429 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1060
timestamp 1624857261
transform 1 0 39769 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1059
timestamp 1624857261
transform 1 0 40105 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1060
timestamp 1624857261
transform 1 0 39765 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1059
timestamp 1624857261
transform 1 0 40101 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1058
timestamp 1624857261
transform 1 0 40441 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1058
timestamp 1624857261
transform 1 0 40437 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4181
timestamp 1624857261
transform 1 0 40664 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1057
timestamp 1624857261
transform 1 0 40777 0 1 131992
box 0 0 1 1
use contact_19  contact_19_829
timestamp 1624857261
transform 1 0 40770 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1057
timestamp 1624857261
transform 1 0 40773 0 1 132000
box 0 0 1 1
use contact_7  contact_7_213
timestamp 1624857261
transform 1 0 40769 0 1 131996
box 0 0 1 1
use contact_14  contact_14_1053
timestamp 1624857261
transform 1 0 42117 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1054
timestamp 1624857261
transform 1 0 41781 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1055
timestamp 1624857261
transform 1 0 41445 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1056
timestamp 1624857261
transform 1 0 41109 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1053
timestamp 1624857261
transform 1 0 42121 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1054
timestamp 1624857261
transform 1 0 41785 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1055
timestamp 1624857261
transform 1 0 41449 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1056
timestamp 1624857261
transform 1 0 41113 0 1 131992
box 0 0 1 1
use contact_33  contact_33_4159
timestamp 1624857261
transform 1 0 42432 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1052
timestamp 1624857261
transform 1 0 42457 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1051
timestamp 1624857261
transform 1 0 42793 0 1 131992
box 0 0 1 1
use contact_19  contact_19_828
timestamp 1624857261
transform 1 0 42450 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1052
timestamp 1624857261
transform 1 0 42453 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1051
timestamp 1624857261
transform 1 0 42789 0 1 132000
box 0 0 1 1
use contact_7  contact_7_212
timestamp 1624857261
transform 1 0 42449 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1050
timestamp 1624857261
transform 1 0 43129 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1050
timestamp 1624857261
transform 1 0 43125 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1049
timestamp 1624857261
transform 1 0 43465 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1049
timestamp 1624857261
transform 1 0 43461 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1048
timestamp 1624857261
transform 1 0 43801 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1047
timestamp 1624857261
transform 1 0 44137 0 1 131992
box 0 0 1 1
use contact_7  contact_7_211
timestamp 1624857261
transform 1 0 44129 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1046
timestamp 1624857261
transform 1 0 44473 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1045
timestamp 1624857261
transform 1 0 44809 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1044
timestamp 1624857261
transform 1 0 45145 0 1 131992
box 0 0 1 1
use contact_19  contact_19_827
timestamp 1624857261
transform 1 0 44130 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1048
timestamp 1624857261
transform 1 0 43797 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1047
timestamp 1624857261
transform 1 0 44133 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4143
timestamp 1624857261
transform 1 0 44200 0 1 132061
box 0 0 1 1
use contact_14  contact_14_1046
timestamp 1624857261
transform 1 0 44469 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1045
timestamp 1624857261
transform 1 0 44805 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1044
timestamp 1624857261
transform 1 0 45141 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1043
timestamp 1624857261
transform 1 0 45481 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1043
timestamp 1624857261
transform 1 0 45477 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4125
timestamp 1624857261
transform 1 0 45696 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1042
timestamp 1624857261
transform 1 0 45817 0 1 131992
box 0 0 1 1
use contact_19  contact_19_826
timestamp 1624857261
transform 1 0 45810 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1042
timestamp 1624857261
transform 1 0 45813 0 1 132000
box 0 0 1 1
use contact_7  contact_7_210
timestamp 1624857261
transform 1 0 45809 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1041
timestamp 1624857261
transform 1 0 46153 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1041
timestamp 1624857261
transform 1 0 46149 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1040
timestamp 1624857261
transform 1 0 46489 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1040
timestamp 1624857261
transform 1 0 46485 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1039
timestamp 1624857261
transform 1 0 46825 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1039
timestamp 1624857261
transform 1 0 46821 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1038
timestamp 1624857261
transform 1 0 47161 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1038
timestamp 1624857261
transform 1 0 47157 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4105
timestamp 1624857261
transform 1 0 47464 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1037
timestamp 1624857261
transform 1 0 47497 0 1 131992
box 0 0 1 1
use contact_19  contact_19_825
timestamp 1624857261
transform 1 0 47490 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1037
timestamp 1624857261
transform 1 0 47493 0 1 132000
box 0 0 1 1
use contact_7  contact_7_209
timestamp 1624857261
transform 1 0 47489 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1036
timestamp 1624857261
transform 1 0 47833 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1036
timestamp 1624857261
transform 1 0 47829 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1035
timestamp 1624857261
transform 1 0 48169 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1035
timestamp 1624857261
transform 1 0 48165 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1034
timestamp 1624857261
transform 1 0 48505 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1034
timestamp 1624857261
transform 1 0 48501 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4087
timestamp 1624857261
transform 1 0 49096 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1033
timestamp 1624857261
transform 1 0 48841 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1033
timestamp 1624857261
transform 1 0 48837 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1032
timestamp 1624857261
transform 1 0 49177 0 1 131992
box 0 0 1 1
use contact_19  contact_19_824
timestamp 1624857261
transform 1 0 49170 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1032
timestamp 1624857261
transform 1 0 49173 0 1 132000
box 0 0 1 1
use contact_7  contact_7_208
timestamp 1624857261
transform 1 0 49169 0 1 131996
box 0 0 1 1
use contact_14  contact_14_1028
timestamp 1624857261
transform 1 0 50517 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1029
timestamp 1624857261
transform 1 0 50181 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1030
timestamp 1624857261
transform 1 0 49845 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1031
timestamp 1624857261
transform 1 0 49509 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1028
timestamp 1624857261
transform 1 0 50521 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1029
timestamp 1624857261
transform 1 0 50185 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1030
timestamp 1624857261
transform 1 0 49849 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1031
timestamp 1624857261
transform 1 0 49513 0 1 131992
box 0 0 1 1
use contact_33  contact_33_4067
timestamp 1624857261
transform 1 0 50728 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1027
timestamp 1624857261
transform 1 0 50857 0 1 131992
box 0 0 1 1
use contact_19  contact_19_823
timestamp 1624857261
transform 1 0 50850 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1027
timestamp 1624857261
transform 1 0 50853 0 1 132000
box 0 0 1 1
use contact_7  contact_7_207
timestamp 1624857261
transform 1 0 50849 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1026
timestamp 1624857261
transform 1 0 51193 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1026
timestamp 1624857261
transform 1 0 51189 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1025
timestamp 1624857261
transform 1 0 51529 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1025
timestamp 1624857261
transform 1 0 51525 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1024
timestamp 1624857261
transform 1 0 51865 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1024
timestamp 1624857261
transform 1 0 51861 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1023
timestamp 1624857261
transform 1 0 52201 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1023
timestamp 1624857261
transform 1 0 52197 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4051
timestamp 1624857261
transform 1 0 52632 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1022
timestamp 1624857261
transform 1 0 52537 0 1 131992
box 0 0 1 1
use contact_19  contact_19_822
timestamp 1624857261
transform 1 0 52530 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1022
timestamp 1624857261
transform 1 0 52533 0 1 132000
box 0 0 1 1
use contact_7  contact_7_206
timestamp 1624857261
transform 1 0 52529 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1021
timestamp 1624857261
transform 1 0 52873 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1021
timestamp 1624857261
transform 1 0 52869 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1020
timestamp 1624857261
transform 1 0 53209 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1020
timestamp 1624857261
transform 1 0 53205 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1019
timestamp 1624857261
transform 1 0 53545 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1019
timestamp 1624857261
transform 1 0 53541 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4035
timestamp 1624857261
transform 1 0 54128 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1018
timestamp 1624857261
transform 1 0 53881 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1018
timestamp 1624857261
transform 1 0 53877 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1017
timestamp 1624857261
transform 1 0 54217 0 1 131992
box 0 0 1 1
use contact_19  contact_19_821
timestamp 1624857261
transform 1 0 54210 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1017
timestamp 1624857261
transform 1 0 54213 0 1 132000
box 0 0 1 1
use contact_7  contact_7_205
timestamp 1624857261
transform 1 0 54209 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1016
timestamp 1624857261
transform 1 0 54553 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1016
timestamp 1624857261
transform 1 0 54549 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1015
timestamp 1624857261
transform 1 0 54889 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1015
timestamp 1624857261
transform 1 0 54885 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1014
timestamp 1624857261
transform 1 0 55225 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1014
timestamp 1624857261
transform 1 0 55221 0 1 132000
box 0 0 1 1
use contact_33  contact_33_4011
timestamp 1624857261
transform 1 0 55896 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1013
timestamp 1624857261
transform 1 0 55561 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1012
timestamp 1624857261
transform 1 0 55897 0 1 131992
box 0 0 1 1
use contact_19  contact_19_820
timestamp 1624857261
transform 1 0 55890 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1013
timestamp 1624857261
transform 1 0 55557 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1012
timestamp 1624857261
transform 1 0 55893 0 1 132000
box 0 0 1 1
use contact_7  contact_7_204
timestamp 1624857261
transform 1 0 55889 0 1 131996
box 0 0 1 1
use contact_14  contact_14_1008
timestamp 1624857261
transform 1 0 57237 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1009
timestamp 1624857261
transform 1 0 56901 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1010
timestamp 1624857261
transform 1 0 56565 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1011
timestamp 1624857261
transform 1 0 56229 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1008
timestamp 1624857261
transform 1 0 57241 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1009
timestamp 1624857261
transform 1 0 56905 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1010
timestamp 1624857261
transform 1 0 56569 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1011
timestamp 1624857261
transform 1 0 56233 0 1 131992
box 0 0 1 1
use contact_33  contact_33_3989
timestamp 1624857261
transform 1 0 57664 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1007
timestamp 1624857261
transform 1 0 57577 0 1 131992
box 0 0 1 1
use contact_19  contact_19_819
timestamp 1624857261
transform 1 0 57570 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1007
timestamp 1624857261
transform 1 0 57573 0 1 132000
box 0 0 1 1
use contact_7  contact_7_203
timestamp 1624857261
transform 1 0 57569 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1006
timestamp 1624857261
transform 1 0 57913 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1006
timestamp 1624857261
transform 1 0 57909 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1005
timestamp 1624857261
transform 1 0 58249 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1004
timestamp 1624857261
transform 1 0 58585 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1005
timestamp 1624857261
transform 1 0 58245 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1004
timestamp 1624857261
transform 1 0 58581 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3977
timestamp 1624857261
transform 1 0 59160 0 1 132061
box 0 0 1 1
use contact_13  contact_13_1003
timestamp 1624857261
transform 1 0 58921 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1003
timestamp 1624857261
transform 1 0 58917 0 1 132000
box 0 0 1 1
use contact_13  contact_13_1002
timestamp 1624857261
transform 1 0 59257 0 1 131992
box 0 0 1 1
use contact_19  contact_19_818
timestamp 1624857261
transform 1 0 59250 0 1 132001
box 0 0 1 1
use contact_14  contact_14_1002
timestamp 1624857261
transform 1 0 59253 0 1 132000
box 0 0 1 1
use contact_7  contact_7_202
timestamp 1624857261
transform 1 0 59249 0 1 131996
box 0 0 1 1
use contact_13  contact_13_1001
timestamp 1624857261
transform 1 0 59593 0 1 131992
box 0 0 1 1
use contact_13  contact_13_1000
timestamp 1624857261
transform 1 0 59929 0 1 131992
box 0 0 1 1
use contact_14  contact_14_1001
timestamp 1624857261
transform 1 0 59589 0 1 132000
box 0 0 1 1
use contact_14  contact_14_1000
timestamp 1624857261
transform 1 0 59925 0 1 132000
box 0 0 1 1
use contact_13  contact_13_999
timestamp 1624857261
transform 1 0 60265 0 1 131992
box 0 0 1 1
use contact_14  contact_14_999
timestamp 1624857261
transform 1 0 60261 0 1 132000
box 0 0 1 1
use contact_13  contact_13_998
timestamp 1624857261
transform 1 0 60601 0 1 131992
box 0 0 1 1
use contact_19  contact_19_817
timestamp 1624857261
transform 1 0 60930 0 1 132001
box 0 0 1 1
use contact_14  contact_14_998
timestamp 1624857261
transform 1 0 60597 0 1 132000
box 0 0 1 1
use contact_7  contact_7_201
timestamp 1624857261
transform 1 0 60929 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3957
timestamp 1624857261
transform 1 0 61064 0 1 132061
box 0 0 1 1
use contact_13  contact_13_997
timestamp 1624857261
transform 1 0 60937 0 1 131992
box 0 0 1 1
use contact_13  contact_13_996
timestamp 1624857261
transform 1 0 61273 0 1 131992
box 0 0 1 1
use contact_14  contact_14_997
timestamp 1624857261
transform 1 0 60933 0 1 132000
box 0 0 1 1
use contact_14  contact_14_996
timestamp 1624857261
transform 1 0 61269 0 1 132000
box 0 0 1 1
use contact_13  contact_13_995
timestamp 1624857261
transform 1 0 61609 0 1 131992
box 0 0 1 1
use contact_14  contact_14_995
timestamp 1624857261
transform 1 0 61605 0 1 132000
box 0 0 1 1
use contact_13  contact_13_994
timestamp 1624857261
transform 1 0 61945 0 1 131992
box 0 0 1 1
use contact_13  contact_13_993
timestamp 1624857261
transform 1 0 62281 0 1 131992
box 0 0 1 1
use contact_14  contact_14_994
timestamp 1624857261
transform 1 0 61941 0 1 132000
box 0 0 1 1
use contact_14  contact_14_993
timestamp 1624857261
transform 1 0 62277 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3939
timestamp 1624857261
transform 1 0 62696 0 1 132061
box 0 0 1 1
use contact_13  contact_13_992
timestamp 1624857261
transform 1 0 62617 0 1 131992
box 0 0 1 1
use contact_19  contact_19_816
timestamp 1624857261
transform 1 0 62610 0 1 132001
box 0 0 1 1
use contact_14  contact_14_992
timestamp 1624857261
transform 1 0 62613 0 1 132000
box 0 0 1 1
use contact_7  contact_7_200
timestamp 1624857261
transform 1 0 62609 0 1 131996
box 0 0 1 1
use contact_14  contact_14_988
timestamp 1624857261
transform 1 0 63957 0 1 132000
box 0 0 1 1
use contact_14  contact_14_989
timestamp 1624857261
transform 1 0 63621 0 1 132000
box 0 0 1 1
use contact_14  contact_14_990
timestamp 1624857261
transform 1 0 63285 0 1 132000
box 0 0 1 1
use contact_14  contact_14_991
timestamp 1624857261
transform 1 0 62949 0 1 132000
box 0 0 1 1
use contact_13  contact_13_988
timestamp 1624857261
transform 1 0 63961 0 1 131992
box 0 0 1 1
use contact_13  contact_13_989
timestamp 1624857261
transform 1 0 63625 0 1 131992
box 0 0 1 1
use contact_13  contact_13_990
timestamp 1624857261
transform 1 0 63289 0 1 131992
box 0 0 1 1
use contact_13  contact_13_991
timestamp 1624857261
transform 1 0 62953 0 1 131992
box 0 0 1 1
use contact_33  contact_33_3923
timestamp 1624857261
transform 1 0 64192 0 1 132061
box 0 0 1 1
use contact_13  contact_13_987
timestamp 1624857261
transform 1 0 64297 0 1 131992
box 0 0 1 1
use contact_19  contact_19_815
timestamp 1624857261
transform 1 0 64290 0 1 132001
box 0 0 1 1
use contact_14  contact_14_987
timestamp 1624857261
transform 1 0 64293 0 1 132000
box 0 0 1 1
use contact_7  contact_7_199
timestamp 1624857261
transform 1 0 64289 0 1 131996
box 0 0 1 1
use contact_13  contact_13_986
timestamp 1624857261
transform 1 0 64633 0 1 131992
box 0 0 1 1
use contact_13  contact_13_985
timestamp 1624857261
transform 1 0 64969 0 1 131992
box 0 0 1 1
use contact_14  contact_14_986
timestamp 1624857261
transform 1 0 64629 0 1 132000
box 0 0 1 1
use contact_14  contact_14_985
timestamp 1624857261
transform 1 0 64965 0 1 132000
box 0 0 1 1
use contact_13  contact_13_984
timestamp 1624857261
transform 1 0 65305 0 1 131992
box 0 0 1 1
use contact_14  contact_14_984
timestamp 1624857261
transform 1 0 65301 0 1 132000
box 0 0 1 1
use contact_13  contact_13_983
timestamp 1624857261
transform 1 0 65641 0 1 131992
box 0 0 1 1
use contact_14  contact_14_983
timestamp 1624857261
transform 1 0 65637 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3899
timestamp 1624857261
transform 1 0 66096 0 1 132061
box 0 0 1 1
use contact_13  contact_13_982
timestamp 1624857261
transform 1 0 65977 0 1 131992
box 0 0 1 1
use contact_13  contact_13_981
timestamp 1624857261
transform 1 0 66313 0 1 131992
box 0 0 1 1
use contact_19  contact_19_814
timestamp 1624857261
transform 1 0 65970 0 1 132001
box 0 0 1 1
use contact_14  contact_14_982
timestamp 1624857261
transform 1 0 65973 0 1 132000
box 0 0 1 1
use contact_14  contact_14_981
timestamp 1624857261
transform 1 0 66309 0 1 132000
box 0 0 1 1
use contact_7  contact_7_198
timestamp 1624857261
transform 1 0 65969 0 1 131996
box 0 0 1 1
use contact_13  contact_13_980
timestamp 1624857261
transform 1 0 66649 0 1 131992
box 0 0 1 1
use contact_14  contact_14_980
timestamp 1624857261
transform 1 0 66645 0 1 132000
box 0 0 1 1
use contact_14  contact_14_978
timestamp 1624857261
transform 1 0 67317 0 1 132000
box 0 0 1 1
use contact_14  contact_14_979
timestamp 1624857261
transform 1 0 66981 0 1 132000
box 0 0 1 1
use contact_13  contact_13_978
timestamp 1624857261
transform 1 0 67321 0 1 131992
box 0 0 1 1
use contact_13  contact_13_979
timestamp 1624857261
transform 1 0 66985 0 1 131992
box 0 0 1 1
use contact_39  contact_39_67
timestamp 1624857261
transform 1 0 1088 0 1 132469
box 0 0 192 192
use contact_39  contact_39_54
timestamp 1624857261
transform 1 0 952 0 1 132469
box 0 0 192 192
use contact_39  contact_39_53
timestamp 1624857261
transform 1 0 1224 0 1 132469
box 0 0 192 192
use contact_39  contact_39_68
timestamp 1624857261
transform 1 0 1224 0 1 132741
box 0 0 192 192
use contact_39  contact_39_66
timestamp 1624857261
transform 1 0 1088 0 1 132605
box 0 0 192 192
use contact_39  contact_39_55
timestamp 1624857261
transform 1 0 952 0 1 132605
box 0 0 192 192
use contact_39  contact_39_46
timestamp 1624857261
transform 1 0 1224 0 1 132605
box 0 0 192 192
use contact_39  contact_39_43
timestamp 1624857261
transform 1 0 1088 0 1 132741
box 0 0 192 192
use contact_39  contact_39_38
timestamp 1624857261
transform 1 0 952 0 1 132741
box 0 0 192 192
use contact_39  contact_39_18
timestamp 1624857261
transform 1 0 408 0 1 133149
box 0 0 192 192
use contact_39  contact_39_15
timestamp 1624857261
transform 1 0 544 0 1 133149
box 0 0 192 192
use contact_39  contact_39_12
timestamp 1624857261
transform 1 0 272 0 1 133149
box 0 0 192 192
use contact_39  contact_39_33
timestamp 1624857261
transform 1 0 544 0 1 133285
box 0 0 192 192
use contact_39  contact_39_30
timestamp 1624857261
transform 1 0 544 0 1 133421
box 0 0 192 192
use contact_39  contact_39_25
timestamp 1624857261
transform 1 0 272 0 1 133285
box 0 0 192 192
use contact_39  contact_39_14
timestamp 1624857261
transform 1 0 272 0 1 133421
box 0 0 192 192
use contact_39  contact_39_4
timestamp 1624857261
transform 1 0 408 0 1 133421
box 0 0 192 192
use contact_39  contact_39_1
timestamp 1624857261
transform 1 0 408 0 1 133285
box 0 0 192 192
use contact_33  contact_33_5292
timestamp 1624857261
transform 1 0 2176 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5288
timestamp 1624857261
transform 1 0 3672 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5286
timestamp 1624857261
transform 1 0 5440 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5280
timestamp 1624857261
transform 1 0 7208 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5276
timestamp 1624857261
transform 1 0 8976 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5272
timestamp 1624857261
transform 1 0 10472 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5268
timestamp 1624857261
transform 1 0 12104 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5264
timestamp 1624857261
transform 1 0 13872 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5244
timestamp 1624857261
transform 1 0 15640 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5238
timestamp 1624857261
transform 1 0 17136 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5226
timestamp 1624857261
transform 1 0 18904 0 1 132469
box 0 0 1 1
use contact_33  contact_33_5202
timestamp 1624857261
transform 1 0 20672 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4902
timestamp 1624857261
transform 1 0 22168 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4324
timestamp 1624857261
transform 1 0 23936 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4320
timestamp 1624857261
transform 1 0 25704 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4316
timestamp 1624857261
transform 1 0 27200 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4308
timestamp 1624857261
transform 1 0 28968 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4286
timestamp 1624857261
transform 1 0 30736 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4264
timestamp 1624857261
transform 1 0 32232 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4256
timestamp 1624857261
transform 1 0 34136 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4228
timestamp 1624857261
transform 1 0 35632 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4208
timestamp 1624857261
transform 1 0 37400 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4202
timestamp 1624857261
transform 1 0 39168 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4180
timestamp 1624857261
transform 1 0 40664 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4158
timestamp 1624857261
transform 1 0 42432 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4142
timestamp 1624857261
transform 1 0 44200 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4124
timestamp 1624857261
transform 1 0 45696 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4104
timestamp 1624857261
transform 1 0 47464 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4086
timestamp 1624857261
transform 1 0 49096 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4066
timestamp 1624857261
transform 1 0 50728 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4050
timestamp 1624857261
transform 1 0 52632 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4034
timestamp 1624857261
transform 1 0 54128 0 1 132469
box 0 0 1 1
use contact_33  contact_33_4010
timestamp 1624857261
transform 1 0 55896 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3988
timestamp 1624857261
transform 1 0 57664 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3976
timestamp 1624857261
transform 1 0 59160 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3956
timestamp 1624857261
transform 1 0 61064 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3938
timestamp 1624857261
transform 1 0 62696 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3922
timestamp 1624857261
transform 1 0 64192 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3898
timestamp 1624857261
transform 1 0 66096 0 1 132469
box 0 0 1 1
use bank  bank_0
timestamp 1624857261
transform 1 0 15406 0 1 9422
box 0 0 67334 67312
use contact_33  contact_33_3868
timestamp 1624857261
transform 1 0 69224 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3842
timestamp 1624857261
transform 1 0 71128 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3824
timestamp 1624857261
transform 1 0 72624 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3810
timestamp 1624857261
transform 1 0 74256 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3782
timestamp 1624857261
transform 1 0 76024 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3760
timestamp 1624857261
transform 1 0 77656 0 1 1229
box 0 0 1 1
use contact_13  contact_13_1378
timestamp 1624857261
transform 1 0 67657 0 1 1683
box 0 0 1 1
use contact_19  contact_19_894
timestamp 1624857261
transform 1 0 67650 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1378
timestamp 1624857261
transform 1 0 67653 0 1 1691
box 0 0 1 1
use contact_7  contact_7_278
timestamp 1624857261
transform 1 0 67649 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1377
timestamp 1624857261
transform 1 0 67993 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1377
timestamp 1624857261
transform 1 0 67989 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1376
timestamp 1624857261
transform 1 0 68329 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1375
timestamp 1624857261
transform 1 0 68665 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1376
timestamp 1624857261
transform 1 0 68325 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1375
timestamp 1624857261
transform 1 0 68661 0 1 1691
box 0 0 1 1
use contact_7  contact_7_277
timestamp 1624857261
transform 1 0 69329 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1372
timestamp 1624857261
transform 1 0 69669 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1373
timestamp 1624857261
transform 1 0 69333 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1374
timestamp 1624857261
transform 1 0 68997 0 1 1691
box 0 0 1 1
use contact_19  contact_19_893
timestamp 1624857261
transform 1 0 69330 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1372
timestamp 1624857261
transform 1 0 69673 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1373
timestamp 1624857261
transform 1 0 69337 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1374
timestamp 1624857261
transform 1 0 69001 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3869
timestamp 1624857261
transform 1 0 69224 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1369
timestamp 1624857261
transform 1 0 70677 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1370
timestamp 1624857261
transform 1 0 70341 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1371
timestamp 1624857261
transform 1 0 70005 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1369
timestamp 1624857261
transform 1 0 70681 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1370
timestamp 1624857261
transform 1 0 70345 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1371
timestamp 1624857261
transform 1 0 70009 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3843
timestamp 1624857261
transform 1 0 71128 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1368
timestamp 1624857261
transform 1 0 71017 0 1 1683
box 0 0 1 1
use contact_19  contact_19_892
timestamp 1624857261
transform 1 0 71010 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1368
timestamp 1624857261
transform 1 0 71013 0 1 1691
box 0 0 1 1
use contact_7  contact_7_276
timestamp 1624857261
transform 1 0 71009 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1367
timestamp 1624857261
transform 1 0 71353 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1367
timestamp 1624857261
transform 1 0 71349 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1366
timestamp 1624857261
transform 1 0 71689 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1366
timestamp 1624857261
transform 1 0 71685 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1365
timestamp 1624857261
transform 1 0 72025 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1365
timestamp 1624857261
transform 1 0 72021 0 1 1691
box 0 0 1 1
use contact_7  contact_7_275
timestamp 1624857261
transform 1 0 72689 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1362
timestamp 1624857261
transform 1 0 73029 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1363
timestamp 1624857261
transform 1 0 72693 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1364
timestamp 1624857261
transform 1 0 72357 0 1 1691
box 0 0 1 1
use contact_19  contact_19_891
timestamp 1624857261
transform 1 0 72690 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1362
timestamp 1624857261
transform 1 0 73033 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1363
timestamp 1624857261
transform 1 0 72697 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1364
timestamp 1624857261
transform 1 0 72361 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3825
timestamp 1624857261
transform 1 0 72624 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1359
timestamp 1624857261
transform 1 0 74037 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1360
timestamp 1624857261
transform 1 0 73701 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1361
timestamp 1624857261
transform 1 0 73365 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1359
timestamp 1624857261
transform 1 0 74041 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1360
timestamp 1624857261
transform 1 0 73705 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1361
timestamp 1624857261
transform 1 0 73369 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3811
timestamp 1624857261
transform 1 0 74256 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1358
timestamp 1624857261
transform 1 0 74377 0 1 1683
box 0 0 1 1
use contact_19  contact_19_890
timestamp 1624857261
transform 1 0 74370 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1358
timestamp 1624857261
transform 1 0 74373 0 1 1691
box 0 0 1 1
use contact_7  contact_7_274
timestamp 1624857261
transform 1 0 74369 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1357
timestamp 1624857261
transform 1 0 74713 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1357
timestamp 1624857261
transform 1 0 74709 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1356
timestamp 1624857261
transform 1 0 75049 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1356
timestamp 1624857261
transform 1 0 75045 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1355
timestamp 1624857261
transform 1 0 75385 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1355
timestamp 1624857261
transform 1 0 75381 0 1 1691
box 0 0 1 1
use contact_7  contact_7_273
timestamp 1624857261
transform 1 0 76049 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1352
timestamp 1624857261
transform 1 0 76389 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1353
timestamp 1624857261
transform 1 0 76053 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1354
timestamp 1624857261
transform 1 0 75717 0 1 1691
box 0 0 1 1
use contact_19  contact_19_889
timestamp 1624857261
transform 1 0 76050 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1352
timestamp 1624857261
transform 1 0 76393 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1353
timestamp 1624857261
transform 1 0 76057 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1354
timestamp 1624857261
transform 1 0 75721 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3783
timestamp 1624857261
transform 1 0 76024 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1349
timestamp 1624857261
transform 1 0 77397 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1350
timestamp 1624857261
transform 1 0 77061 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1351
timestamp 1624857261
transform 1 0 76725 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1349
timestamp 1624857261
transform 1 0 77401 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1350
timestamp 1624857261
transform 1 0 77065 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1351
timestamp 1624857261
transform 1 0 76729 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3761
timestamp 1624857261
transform 1 0 77656 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1348
timestamp 1624857261
transform 1 0 77737 0 1 1683
box 0 0 1 1
use contact_19  contact_19_888
timestamp 1624857261
transform 1 0 77730 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1348
timestamp 1624857261
transform 1 0 77733 0 1 1691
box 0 0 1 1
use contact_7  contact_7_272
timestamp 1624857261
transform 1 0 77729 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1347
timestamp 1624857261
transform 1 0 78073 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1347
timestamp 1624857261
transform 1 0 78069 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1346
timestamp 1624857261
transform 1 0 78409 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1346
timestamp 1624857261
transform 1 0 78405 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1345
timestamp 1624857261
transform 1 0 78745 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1345
timestamp 1624857261
transform 1 0 78741 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1344
timestamp 1624857261
transform 1 0 79077 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1344
timestamp 1624857261
transform 1 0 79081 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3862
timestamp 1624857261
transform 1 0 69768 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3834
timestamp 1624857261
transform 1 0 72216 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3802
timestamp 1624857261
transform 1 0 74528 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3770
timestamp 1624857261
transform 1 0 77248 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3861
timestamp 1624857261
transform 1 0 69768 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3863
timestamp 1624857261
transform 1 0 69768 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1164
timestamp 1624857261
transform 1 0 69904 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1165
timestamp 1624857261
transform 1 0 69904 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1166
timestamp 1624857261
transform 1 0 69904 0 1 12245
box 0 0 1 1
use contact_33  contact_33_1152
timestamp 1624857261
transform 1 0 72488 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1153
timestamp 1624857261
transform 1 0 72488 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1154
timestamp 1624857261
transform 1 0 72488 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3833
timestamp 1624857261
transform 1 0 72352 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3835
timestamp 1624857261
transform 1 0 72216 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1140
timestamp 1624857261
transform 1 0 74936 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1141
timestamp 1624857261
transform 1 0 74664 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1142
timestamp 1624857261
transform 1 0 74664 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3801
timestamp 1624857261
transform 1 0 74800 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3803
timestamp 1624857261
transform 1 0 74528 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1128
timestamp 1624857261
transform 1 0 77248 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1129
timestamp 1624857261
transform 1 0 76976 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1130
timestamp 1624857261
transform 1 0 76976 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3769
timestamp 1624857261
transform 1 0 77112 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3771
timestamp 1624857261
transform 1 0 77248 0 1 11837
box 0 0 1 1
use contact_7  contact_7_391
timestamp 1624857261
transform 1 0 69493 0 1 13196
box 0 0 1 1
use contact_19  contact_19_981
timestamp 1624857261
transform 1 0 69494 0 1 13201
box 0 0 1 1
use contact_33  contact_33_3858
timestamp 1624857261
transform 1 0 69632 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3860
timestamp 1624857261
transform 1 0 69768 0 1 13605
box 0 0 1 1
use contact_33  contact_33_5398
timestamp 1624857261
transform 1 0 69496 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1162
timestamp 1624857261
transform 1 0 70040 0 1 12925
box 0 0 1 1
use contact_33  contact_33_1163
timestamp 1624857261
transform 1 0 69904 0 1 13061
box 0 0 1 1
use contact_7  contact_7_390
timestamp 1624857261
transform 1 0 71989 0 1 13196
box 0 0 1 1
use contact_19  contact_19_980
timestamp 1624857261
transform 1 0 71990 0 1 13201
box 0 0 1 1
use contact_33  contact_33_3855
timestamp 1624857261
transform 1 0 72080 0 1 13605
box 0 0 1 1
use contact_33  contact_33_5397
timestamp 1624857261
transform 1 0 71944 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1148
timestamp 1624857261
transform 1 0 72488 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1151
timestamp 1624857261
transform 1 0 72488 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3828
timestamp 1624857261
transform 1 0 72216 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3832
timestamp 1624857261
transform 1 0 72352 0 1 13469
box 0 0 1 1
use contact_7  contact_7_389
timestamp 1624857261
transform 1 0 74485 0 1 13196
box 0 0 1 1
use contact_19  contact_19_979
timestamp 1624857261
transform 1 0 74486 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1138
timestamp 1624857261
transform 1 0 74936 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1139
timestamp 1624857261
transform 1 0 74936 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3796
timestamp 1624857261
transform 1 0 74800 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3800
timestamp 1624857261
transform 1 0 74800 0 1 13469
box 0 0 1 1
use contact_33  contact_33_5396
timestamp 1624857261
transform 1 0 74392 0 1 13061
box 0 0 1 1
use contact_7  contact_7_388
timestamp 1624857261
transform 1 0 76981 0 1 13196
box 0 0 1 1
use contact_19  contact_19_978
timestamp 1624857261
transform 1 0 76982 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1126
timestamp 1624857261
transform 1 0 77384 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1127
timestamp 1624857261
transform 1 0 77248 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3762
timestamp 1624857261
transform 1 0 77248 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3768
timestamp 1624857261
transform 1 0 77112 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3794
timestamp 1624857261
transform 1 0 76976 0 1 13605
box 0 0 1 1
use contact_33  contact_33_5395
timestamp 1624857261
transform 1 0 76840 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3859
timestamp 1624857261
transform 1 0 69632 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3854
timestamp 1624857261
transform 1 0 72080 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3829
timestamp 1624857261
transform 1 0 72216 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3797
timestamp 1624857261
transform 1 0 74800 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3763
timestamp 1624857261
transform 1 0 77248 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3774
timestamp 1624857261
transform 1 0 77112 0 1 14421
box 0 0 1 1
use contact_33  contact_33_3795
timestamp 1624857261
transform 1 0 76976 0 1 14285
box 0 0 1 1
use contact_33  contact_33_1158
timestamp 1624857261
transform 1 0 69904 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1161
timestamp 1624857261
transform 1 0 70040 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1146
timestamp 1624857261
transform 1 0 72352 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1147
timestamp 1624857261
transform 1 0 72488 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1134
timestamp 1624857261
transform 1 0 75072 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1137
timestamp 1624857261
transform 1 0 74936 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1122
timestamp 1624857261
transform 1 0 77520 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1125
timestamp 1624857261
transform 1 0 77384 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1157
timestamp 1624857261
transform 1 0 69904 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1145
timestamp 1624857261
transform 1 0 72352 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1133
timestamp 1624857261
transform 1 0 75072 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1121
timestamp 1624857261
transform 1 0 77520 0 1 17005
box 0 0 1 1
use contact_33  contact_33_3775
timestamp 1624857261
transform 1 0 77112 0 1 18637
box 0 0 1 1
use contact_33  contact_33_3744
timestamp 1624857261
transform 1 0 79288 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3720
timestamp 1624857261
transform 1 0 81192 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3700
timestamp 1624857261
transform 1 0 82688 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3686
timestamp 1624857261
transform 1 0 84592 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3662
timestamp 1624857261
transform 1 0 86088 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3638
timestamp 1624857261
transform 1 0 87720 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3628
timestamp 1624857261
transform 1 0 89352 0 1 1229
box 0 0 1 1
use contact_7  contact_7_271
timestamp 1624857261
transform 1 0 79409 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1341
timestamp 1624857261
transform 1 0 80085 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1342
timestamp 1624857261
transform 1 0 79749 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1343
timestamp 1624857261
transform 1 0 79413 0 1 1691
box 0 0 1 1
use contact_19  contact_19_887
timestamp 1624857261
transform 1 0 79410 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1341
timestamp 1624857261
transform 1 0 80089 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1342
timestamp 1624857261
transform 1 0 79753 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1343
timestamp 1624857261
transform 1 0 79417 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3745
timestamp 1624857261
transform 1 0 79288 0 1 1637
box 0 0 1 1
use contact_7  contact_7_270
timestamp 1624857261
transform 1 0 81089 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1338
timestamp 1624857261
transform 1 0 81093 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1339
timestamp 1624857261
transform 1 0 80757 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1340
timestamp 1624857261
transform 1 0 80421 0 1 1691
box 0 0 1 1
use contact_19  contact_19_886
timestamp 1624857261
transform 1 0 81090 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1338
timestamp 1624857261
transform 1 0 81097 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1339
timestamp 1624857261
transform 1 0 80761 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1340
timestamp 1624857261
transform 1 0 80425 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3721
timestamp 1624857261
transform 1 0 81192 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1335
timestamp 1624857261
transform 1 0 82101 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1336
timestamp 1624857261
transform 1 0 81765 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1337
timestamp 1624857261
transform 1 0 81429 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1335
timestamp 1624857261
transform 1 0 82105 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1336
timestamp 1624857261
transform 1 0 81769 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1337
timestamp 1624857261
transform 1 0 81433 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3701
timestamp 1624857261
transform 1 0 82688 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1334
timestamp 1624857261
transform 1 0 82441 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1333
timestamp 1624857261
transform 1 0 82777 0 1 1683
box 0 0 1 1
use contact_7  contact_7_269
timestamp 1624857261
transform 1 0 82769 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1332
timestamp 1624857261
transform 1 0 83113 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1331
timestamp 1624857261
transform 1 0 83449 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1334
timestamp 1624857261
transform 1 0 82437 0 1 1691
box 0 0 1 1
use contact_19  contact_19_885
timestamp 1624857261
transform 1 0 82770 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1333
timestamp 1624857261
transform 1 0 82773 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1332
timestamp 1624857261
transform 1 0 83109 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1331
timestamp 1624857261
transform 1 0 83445 0 1 1691
box 0 0 1 1
use contact_7  contact_7_268
timestamp 1624857261
transform 1 0 84449 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1328
timestamp 1624857261
transform 1 0 84453 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1329
timestamp 1624857261
transform 1 0 84117 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1330
timestamp 1624857261
transform 1 0 83781 0 1 1691
box 0 0 1 1
use contact_19  contact_19_884
timestamp 1624857261
transform 1 0 84450 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1328
timestamp 1624857261
transform 1 0 84457 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1329
timestamp 1624857261
transform 1 0 84121 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1330
timestamp 1624857261
transform 1 0 83785 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1325
timestamp 1624857261
transform 1 0 85461 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1326
timestamp 1624857261
transform 1 0 85125 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1327
timestamp 1624857261
transform 1 0 84789 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1325
timestamp 1624857261
transform 1 0 85465 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1326
timestamp 1624857261
transform 1 0 85129 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1327
timestamp 1624857261
transform 1 0 84793 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3687
timestamp 1624857261
transform 1 0 84592 0 1 1637
box 0 0 1 1
use contact_7  contact_7_267
timestamp 1624857261
transform 1 0 86129 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1322
timestamp 1624857261
transform 1 0 86469 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1323
timestamp 1624857261
transform 1 0 86133 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1324
timestamp 1624857261
transform 1 0 85797 0 1 1691
box 0 0 1 1
use contact_19  contact_19_883
timestamp 1624857261
transform 1 0 86130 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1322
timestamp 1624857261
transform 1 0 86473 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1323
timestamp 1624857261
transform 1 0 86137 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1324
timestamp 1624857261
transform 1 0 85801 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3663
timestamp 1624857261
transform 1 0 86088 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1321
timestamp 1624857261
transform 1 0 86809 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1320
timestamp 1624857261
transform 1 0 87145 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1319
timestamp 1624857261
transform 1 0 87481 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3639
timestamp 1624857261
transform 1 0 87720 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1318
timestamp 1624857261
transform 1 0 87817 0 1 1683
box 0 0 1 1
use contact_7  contact_7_266
timestamp 1624857261
transform 1 0 87809 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1321
timestamp 1624857261
transform 1 0 86805 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1320
timestamp 1624857261
transform 1 0 87141 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1319
timestamp 1624857261
transform 1 0 87477 0 1 1691
box 0 0 1 1
use contact_19  contact_19_882
timestamp 1624857261
transform 1 0 87810 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1318
timestamp 1624857261
transform 1 0 87813 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1315
timestamp 1624857261
transform 1 0 88821 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1316
timestamp 1624857261
transform 1 0 88485 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1317
timestamp 1624857261
transform 1 0 88149 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1315
timestamp 1624857261
transform 1 0 88825 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1316
timestamp 1624857261
transform 1 0 88489 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1317
timestamp 1624857261
transform 1 0 88153 0 1 1683
box 0 0 1 1
use contact_7  contact_7_265
timestamp 1624857261
transform 1 0 89489 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1312
timestamp 1624857261
transform 1 0 89829 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1313
timestamp 1624857261
transform 1 0 89493 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1314
timestamp 1624857261
transform 1 0 89157 0 1 1691
box 0 0 1 1
use contact_19  contact_19_881
timestamp 1624857261
transform 1 0 89490 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1312
timestamp 1624857261
transform 1 0 89833 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1313
timestamp 1624857261
transform 1 0 89497 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1314
timestamp 1624857261
transform 1 0 89161 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3629
timestamp 1624857261
transform 1 0 89352 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1310
timestamp 1624857261
transform 1 0 90501 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1311
timestamp 1624857261
transform 1 0 90165 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1310
timestamp 1624857261
transform 1 0 90505 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1311
timestamp 1624857261
transform 1 0 90169 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3740
timestamp 1624857261
transform 1 0 79696 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3712
timestamp 1624857261
transform 1 0 82144 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3678
timestamp 1624857261
transform 1 0 84592 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3650
timestamp 1624857261
transform 1 0 87176 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3622
timestamp 1624857261
transform 1 0 89488 0 1 11021
box 0 0 1 1
use contact_33  contact_33_1117
timestamp 1624857261
transform 1 0 79968 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3739
timestamp 1624857261
transform 1 0 79832 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3741
timestamp 1624857261
transform 1 0 79696 0 1 11837
box 0 0 1 1
use contact_33  contact_33_3711
timestamp 1624857261
transform 1 0 82280 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3713
timestamp 1624857261
transform 1 0 82144 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1105
timestamp 1624857261
transform 1 0 82416 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1093
timestamp 1624857261
transform 1 0 84728 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3677
timestamp 1624857261
transform 1 0 84864 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3679
timestamp 1624857261
transform 1 0 84592 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1081
timestamp 1624857261
transform 1 0 87040 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3649
timestamp 1624857261
transform 1 0 87312 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3651
timestamp 1624857261
transform 1 0 87176 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1069
timestamp 1624857261
transform 1 0 89624 0 1 11701
box 0 0 1 1
use contact_33  contact_33_3621
timestamp 1624857261
transform 1 0 89760 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3623
timestamp 1624857261
transform 1 0 89488 0 1 11837
box 0 0 1 1
use contact_7  contact_7_387
timestamp 1624857261
transform 1 0 79477 0 1 13196
box 0 0 1 1
use contact_19  contact_19_977
timestamp 1624857261
transform 1 0 79478 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1114
timestamp 1624857261
transform 1 0 79968 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1115
timestamp 1624857261
transform 1 0 79968 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1116
timestamp 1624857261
transform 1 0 79968 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1118
timestamp 1624857261
transform 1 0 79968 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5394
timestamp 1624857261
transform 1 0 79424 0 1 13061
box 0 0 1 1
use contact_7  contact_7_386
timestamp 1624857261
transform 1 0 81973 0 1 13196
box 0 0 1 1
use contact_19  contact_19_976
timestamp 1624857261
transform 1 0 81974 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5393
timestamp 1624857261
transform 1 0 81872 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1100
timestamp 1624857261
transform 1 0 82416 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1103
timestamp 1624857261
transform 1 0 82416 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1104
timestamp 1624857261
transform 1 0 82416 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1106
timestamp 1624857261
transform 1 0 82416 0 1 12245
box 0 0 1 1
use contact_7  contact_7_385
timestamp 1624857261
transform 1 0 84469 0 1 13196
box 0 0 1 1
use contact_19  contact_19_975
timestamp 1624857261
transform 1 0 84470 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5392
timestamp 1624857261
transform 1 0 84320 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1088
timestamp 1624857261
transform 1 0 85000 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1091
timestamp 1624857261
transform 1 0 84728 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1092
timestamp 1624857261
transform 1 0 84728 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1094
timestamp 1624857261
transform 1 0 84728 0 1 12245
box 0 0 1 1
use contact_7  contact_7_384
timestamp 1624857261
transform 1 0 86965 0 1 13196
box 0 0 1 1
use contact_19  contact_19_974
timestamp 1624857261
transform 1 0 86966 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1078
timestamp 1624857261
transform 1 0 87448 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1079
timestamp 1624857261
transform 1 0 87448 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1080
timestamp 1624857261
transform 1 0 87448 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1082
timestamp 1624857261
transform 1 0 87040 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5391
timestamp 1624857261
transform 1 0 86904 0 1 13061
box 0 0 1 1
use contact_7  contact_7_383
timestamp 1624857261
transform 1 0 89461 0 1 13196
box 0 0 1 1
use contact_19  contact_19_973
timestamp 1624857261
transform 1 0 89462 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1066
timestamp 1624857261
transform 1 0 89896 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1067
timestamp 1624857261
transform 1 0 89896 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1068
timestamp 1624857261
transform 1 0 89896 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1070
timestamp 1624857261
transform 1 0 89624 0 1 12245
box 0 0 1 1
use contact_33  contact_33_5390
timestamp 1624857261
transform 1 0 89080 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3736
timestamp 1624857261
transform 1 0 79832 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3737
timestamp 1624857261
transform 1 0 79832 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3738
timestamp 1624857261
transform 1 0 79832 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3708
timestamp 1624857261
transform 1 0 82280 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3709
timestamp 1624857261
transform 1 0 82280 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3710
timestamp 1624857261
transform 1 0 82280 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3672
timestamp 1624857261
transform 1 0 84592 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3673
timestamp 1624857261
transform 1 0 84592 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3676
timestamp 1624857261
transform 1 0 84864 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3646
timestamp 1624857261
transform 1 0 87312 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3647
timestamp 1624857261
transform 1 0 87312 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3648
timestamp 1624857261
transform 1 0 87312 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3616
timestamp 1624857261
transform 1 0 89624 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3617
timestamp 1624857261
transform 1 0 89624 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3620
timestamp 1624857261
transform 1 0 89760 0 1 13469
box 0 0 1 1
use contact_33  contact_33_1110
timestamp 1624857261
transform 1 0 79832 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1113
timestamp 1624857261
transform 1 0 79968 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1098
timestamp 1624857261
transform 1 0 82552 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1099
timestamp 1624857261
transform 1 0 82416 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1084
timestamp 1624857261
transform 1 0 84864 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1087
timestamp 1624857261
transform 1 0 85000 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1074
timestamp 1624857261
transform 1 0 87312 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1077
timestamp 1624857261
transform 1 0 87448 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1065
timestamp 1624857261
transform 1 0 89896 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1060
timestamp 1624857261
transform 1 0 90032 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1109
timestamp 1624857261
transform 1 0 79832 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1097
timestamp 1624857261
transform 1 0 82552 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1083
timestamp 1624857261
transform 1 0 84864 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1073
timestamp 1624857261
transform 1 0 87312 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1059
timestamp 1624857261
transform 1 0 90032 0 1 17005
box 0 0 1 1
use contact_33  contact_33_3606
timestamp 1624857261
transform 1 0 91120 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3584
timestamp 1624857261
transform 1 0 92888 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3574
timestamp 1624857261
transform 1 0 94656 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3554
timestamp 1624857261
transform 1 0 96152 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3536
timestamp 1624857261
transform 1 0 97920 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3518
timestamp 1624857261
transform 1 0 99688 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3502
timestamp 1624857261
transform 1 0 101184 0 1 1229
box 0 0 1 1
use contact_7  contact_7_264
timestamp 1624857261
transform 1 0 91169 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1307
timestamp 1624857261
transform 1 0 91509 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1308
timestamp 1624857261
transform 1 0 91173 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1309
timestamp 1624857261
transform 1 0 90837 0 1 1691
box 0 0 1 1
use contact_19  contact_19_880
timestamp 1624857261
transform 1 0 91170 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1307
timestamp 1624857261
transform 1 0 91513 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1308
timestamp 1624857261
transform 1 0 91177 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1309
timestamp 1624857261
transform 1 0 90841 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3607
timestamp 1624857261
transform 1 0 91120 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1306
timestamp 1624857261
transform 1 0 91849 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1306
timestamp 1624857261
transform 1 0 91845 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1305
timestamp 1624857261
transform 1 0 92185 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1305
timestamp 1624857261
transform 1 0 92181 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1304
timestamp 1624857261
transform 1 0 92521 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1304
timestamp 1624857261
transform 1 0 92517 0 1 1691
box 0 0 1 1
use contact_33  contact_33_3585
timestamp 1624857261
transform 1 0 92888 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1303
timestamp 1624857261
transform 1 0 92857 0 1 1683
box 0 0 1 1
use contact_19  contact_19_879
timestamp 1624857261
transform 1 0 92850 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1303
timestamp 1624857261
transform 1 0 92853 0 1 1691
box 0 0 1 1
use contact_7  contact_7_263
timestamp 1624857261
transform 1 0 92849 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1300
timestamp 1624857261
transform 1 0 93861 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1301
timestamp 1624857261
transform 1 0 93525 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1302
timestamp 1624857261
transform 1 0 93189 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1300
timestamp 1624857261
transform 1 0 93865 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1301
timestamp 1624857261
transform 1 0 93529 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1302
timestamp 1624857261
transform 1 0 93193 0 1 1683
box 0 0 1 1
use contact_7  contact_7_262
timestamp 1624857261
transform 1 0 94529 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1297
timestamp 1624857261
transform 1 0 94869 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1298
timestamp 1624857261
transform 1 0 94533 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1299
timestamp 1624857261
transform 1 0 94197 0 1 1691
box 0 0 1 1
use contact_19  contact_19_878
timestamp 1624857261
transform 1 0 94530 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1297
timestamp 1624857261
transform 1 0 94873 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1298
timestamp 1624857261
transform 1 0 94537 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1299
timestamp 1624857261
transform 1 0 94201 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3575
timestamp 1624857261
transform 1 0 94656 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1296
timestamp 1624857261
transform 1 0 95209 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1296
timestamp 1624857261
transform 1 0 95205 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1295
timestamp 1624857261
transform 1 0 95545 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1295
timestamp 1624857261
transform 1 0 95541 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1294
timestamp 1624857261
transform 1 0 95881 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1294
timestamp 1624857261
transform 1 0 95877 0 1 1691
box 0 0 1 1
use contact_33  contact_33_3555
timestamp 1624857261
transform 1 0 96152 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1293
timestamp 1624857261
transform 1 0 96217 0 1 1683
box 0 0 1 1
use contact_19  contact_19_877
timestamp 1624857261
transform 1 0 96210 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1293
timestamp 1624857261
transform 1 0 96213 0 1 1691
box 0 0 1 1
use contact_7  contact_7_261
timestamp 1624857261
transform 1 0 96209 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1290
timestamp 1624857261
transform 1 0 97221 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1291
timestamp 1624857261
transform 1 0 96885 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1292
timestamp 1624857261
transform 1 0 96549 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1290
timestamp 1624857261
transform 1 0 97225 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1291
timestamp 1624857261
transform 1 0 96889 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1292
timestamp 1624857261
transform 1 0 96553 0 1 1683
box 0 0 1 1
use contact_7  contact_7_260
timestamp 1624857261
transform 1 0 97889 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1287
timestamp 1624857261
transform 1 0 98229 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1288
timestamp 1624857261
transform 1 0 97893 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1289
timestamp 1624857261
transform 1 0 97557 0 1 1691
box 0 0 1 1
use contact_19  contact_19_876
timestamp 1624857261
transform 1 0 97890 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1287
timestamp 1624857261
transform 1 0 98233 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1288
timestamp 1624857261
transform 1 0 97897 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1289
timestamp 1624857261
transform 1 0 97561 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3537
timestamp 1624857261
transform 1 0 97920 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1286
timestamp 1624857261
transform 1 0 98569 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1286
timestamp 1624857261
transform 1 0 98565 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1285
timestamp 1624857261
transform 1 0 98905 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1285
timestamp 1624857261
transform 1 0 98901 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1284
timestamp 1624857261
transform 1 0 99241 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1284
timestamp 1624857261
transform 1 0 99237 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1283
timestamp 1624857261
transform 1 0 99577 0 1 1683
box 0 0 1 1
use contact_19  contact_19_875
timestamp 1624857261
transform 1 0 99570 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1283
timestamp 1624857261
transform 1 0 99573 0 1 1691
box 0 0 1 1
use contact_7  contact_7_259
timestamp 1624857261
transform 1 0 99569 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1280
timestamp 1624857261
transform 1 0 100581 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1281
timestamp 1624857261
transform 1 0 100245 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1282
timestamp 1624857261
transform 1 0 99909 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1280
timestamp 1624857261
transform 1 0 100585 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1281
timestamp 1624857261
transform 1 0 100249 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1282
timestamp 1624857261
transform 1 0 99913 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3519
timestamp 1624857261
transform 1 0 99688 0 1 1637
box 0 0 1 1
use contact_7  contact_7_258
timestamp 1624857261
transform 1 0 101249 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1277
timestamp 1624857261
transform 1 0 101589 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1278
timestamp 1624857261
transform 1 0 101253 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1279
timestamp 1624857261
transform 1 0 100917 0 1 1691
box 0 0 1 1
use contact_19  contact_19_874
timestamp 1624857261
transform 1 0 101250 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1277
timestamp 1624857261
transform 1 0 101593 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1278
timestamp 1624857261
transform 1 0 101257 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1279
timestamp 1624857261
transform 1 0 100921 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3503
timestamp 1624857261
transform 1 0 101184 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1276
timestamp 1624857261
transform 1 0 101925 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1276
timestamp 1624857261
transform 1 0 101929 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3598
timestamp 1624857261
transform 1 0 92208 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3570
timestamp 1624857261
transform 1 0 94656 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3548
timestamp 1624857261
transform 1 0 97104 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3516
timestamp 1624857261
transform 1 0 99552 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3492
timestamp 1624857261
transform 1 0 102136 0 1 11021
box 0 0 1 1
use contact_33  contact_33_1056
timestamp 1624857261
transform 1 0 92208 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1057
timestamp 1624857261
transform 1 0 92480 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1058
timestamp 1624857261
transform 1 0 92480 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3597
timestamp 1624857261
transform 1 0 92344 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3599
timestamp 1624857261
transform 1 0 92208 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1044
timestamp 1624857261
transform 1 0 94928 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1045
timestamp 1624857261
transform 1 0 94928 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1046
timestamp 1624857261
transform 1 0 94928 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3569
timestamp 1624857261
transform 1 0 94792 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3571
timestamp 1624857261
transform 1 0 94656 0 1 11837
box 0 0 1 1
use contact_33  contact_33_3547
timestamp 1624857261
transform 1 0 97240 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3549
timestamp 1624857261
transform 1 0 97104 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1032
timestamp 1624857261
transform 1 0 97376 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1033
timestamp 1624857261
transform 1 0 97376 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1034
timestamp 1624857261
transform 1 0 97376 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3517
timestamp 1624857261
transform 1 0 99552 0 1 11837
box 0 0 1 1
use contact_33  contact_33_1020
timestamp 1624857261
transform 1 0 99688 0 1 12517
box 0 0 1 1
use contact_33  contact_33_1021
timestamp 1624857261
transform 1 0 99688 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1022
timestamp 1624857261
transform 1 0 99688 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3515
timestamp 1624857261
transform 1 0 99824 0 1 11973
box 0 0 1 1
use contact_33  contact_33_1009
timestamp 1624857261
transform 1 0 102000 0 1 11701
box 0 0 1 1
use contact_33  contact_33_1010
timestamp 1624857261
transform 1 0 102000 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3493
timestamp 1624857261
transform 1 0 102136 0 1 11837
box 0 0 1 1
use contact_7  contact_7_382
timestamp 1624857261
transform 1 0 91957 0 1 13196
box 0 0 1 1
use contact_19  contact_19_972
timestamp 1624857261
transform 1 0 91958 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1052
timestamp 1624857261
transform 1 0 92480 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1055
timestamp 1624857261
transform 1 0 92208 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3594
timestamp 1624857261
transform 1 0 92208 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3596
timestamp 1624857261
transform 1 0 92344 0 1 13469
box 0 0 1 1
use contact_33  contact_33_5389
timestamp 1624857261
transform 1 0 91936 0 1 13061
box 0 0 1 1
use contact_7  contact_7_381
timestamp 1624857261
transform 1 0 94453 0 1 13196
box 0 0 1 1
use contact_19  contact_19_971
timestamp 1624857261
transform 1 0 94454 0 1 13201
box 0 0 1 1
use contact_33  contact_33_1042
timestamp 1624857261
transform 1 0 94928 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1043
timestamp 1624857261
transform 1 0 94928 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3566
timestamp 1624857261
transform 1 0 94656 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3568
timestamp 1624857261
transform 1 0 94792 0 1 13469
box 0 0 1 1
use contact_33  contact_33_5388
timestamp 1624857261
transform 1 0 94384 0 1 13061
box 0 0 1 1
use contact_7  contact_7_380
timestamp 1624857261
transform 1 0 96949 0 1 13196
box 0 0 1 1
use contact_19  contact_19_970
timestamp 1624857261
transform 1 0 96950 0 1 13201
box 0 0 1 1
use contact_33  contact_33_3544
timestamp 1624857261
transform 1 0 97240 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3546
timestamp 1624857261
transform 1 0 97240 0 1 13469
box 0 0 1 1
use contact_33  contact_33_5387
timestamp 1624857261
transform 1 0 96832 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1030
timestamp 1624857261
transform 1 0 97376 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1031
timestamp 1624857261
transform 1 0 97376 0 1 13061
box 0 0 1 1
use contact_7  contact_7_379
timestamp 1624857261
transform 1 0 99445 0 1 13196
box 0 0 1 1
use contact_19  contact_19_969
timestamp 1624857261
transform 1 0 99446 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5386
timestamp 1624857261
transform 1 0 99416 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1018
timestamp 1624857261
transform 1 0 99960 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1019
timestamp 1624857261
transform 1 0 99688 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3512
timestamp 1624857261
transform 1 0 99688 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3514
timestamp 1624857261
transform 1 0 99824 0 1 13469
box 0 0 1 1
use contact_7  contact_7_378
timestamp 1624857261
transform 1 0 101941 0 1 13196
box 0 0 1 1
use contact_19  contact_19_968
timestamp 1624857261
transform 1 0 101942 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5385
timestamp 1624857261
transform 1 0 101864 0 1 13061
box 0 0 1 1
use contact_33  contact_33_3595
timestamp 1624857261
transform 1 0 92208 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3567
timestamp 1624857261
transform 1 0 94656 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3545
timestamp 1624857261
transform 1 0 97240 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3513
timestamp 1624857261
transform 1 0 99688 0 1 14285
box 0 0 1 1
use contact_33  contact_33_1048
timestamp 1624857261
transform 1 0 92344 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1051
timestamp 1624857261
transform 1 0 92480 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1036
timestamp 1624857261
transform 1 0 94792 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1041
timestamp 1624857261
transform 1 0 94928 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1024
timestamp 1624857261
transform 1 0 97512 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1029
timestamp 1624857261
transform 1 0 97376 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1012
timestamp 1624857261
transform 1 0 99824 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1017
timestamp 1624857261
transform 1 0 99960 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1047
timestamp 1624857261
transform 1 0 92344 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1035
timestamp 1624857261
transform 1 0 94928 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1023
timestamp 1624857261
transform 1 0 97512 0 1 17005
box 0 0 1 1
use contact_33  contact_33_1011
timestamp 1624857261
transform 1 0 99824 0 1 17005
box 0 0 1 1
use contact_33  contact_33_3482
timestamp 1624857261
transform 1 0 102952 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3460
timestamp 1624857261
transform 1 0 104584 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3448
timestamp 1624857261
transform 1 0 106216 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3424
timestamp 1624857261
transform 1 0 107848 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3414
timestamp 1624857261
transform 1 0 109616 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3410
timestamp 1624857261
transform 1 0 111384 0 1 1229
box 0 0 1 1
use contact_33  contact_33_3406
timestamp 1624857261
transform 1 0 112880 0 1 1229
box 0 0 1 1
use contact_13  contact_13_1275
timestamp 1624857261
transform 1 0 102265 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1275
timestamp 1624857261
transform 1 0 102261 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1274
timestamp 1624857261
transform 1 0 102601 0 1 1683
box 0 0 1 1
use contact_19  contact_19_873
timestamp 1624857261
transform 1 0 102930 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1274
timestamp 1624857261
transform 1 0 102597 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1273
timestamp 1624857261
transform 1 0 102933 0 1 1691
box 0 0 1 1
use contact_7  contact_7_257
timestamp 1624857261
transform 1 0 102929 0 1 1687
box 0 0 1 1
use contact_33  contact_33_3483
timestamp 1624857261
transform 1 0 102952 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1273
timestamp 1624857261
transform 1 0 102937 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1272
timestamp 1624857261
transform 1 0 103273 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1272
timestamp 1624857261
transform 1 0 103269 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1271
timestamp 1624857261
transform 1 0 103609 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1271
timestamp 1624857261
transform 1 0 103605 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1270
timestamp 1624857261
transform 1 0 103945 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1270
timestamp 1624857261
transform 1 0 103941 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1269
timestamp 1624857261
transform 1 0 104281 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1269
timestamp 1624857261
transform 1 0 104277 0 1 1691
box 0 0 1 1
use contact_33  contact_33_3461
timestamp 1624857261
transform 1 0 104584 0 1 1637
box 0 0 1 1
use contact_19  contact_19_872
timestamp 1624857261
transform 1 0 104610 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1268
timestamp 1624857261
transform 1 0 104613 0 1 1691
box 0 0 1 1
use contact_7  contact_7_256
timestamp 1624857261
transform 1 0 104609 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1265
timestamp 1624857261
transform 1 0 105621 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1266
timestamp 1624857261
transform 1 0 105285 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1267
timestamp 1624857261
transform 1 0 104949 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1265
timestamp 1624857261
transform 1 0 105625 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1266
timestamp 1624857261
transform 1 0 105289 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1267
timestamp 1624857261
transform 1 0 104953 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1268
timestamp 1624857261
transform 1 0 104617 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1264
timestamp 1624857261
transform 1 0 105961 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1264
timestamp 1624857261
transform 1 0 105957 0 1 1691
box 0 0 1 1
use contact_33  contact_33_3449
timestamp 1624857261
transform 1 0 106216 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1263
timestamp 1624857261
transform 1 0 106297 0 1 1683
box 0 0 1 1
use contact_19  contact_19_871
timestamp 1624857261
transform 1 0 106290 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1263
timestamp 1624857261
transform 1 0 106293 0 1 1691
box 0 0 1 1
use contact_7  contact_7_255
timestamp 1624857261
transform 1 0 106289 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1262
timestamp 1624857261
transform 1 0 106633 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1262
timestamp 1624857261
transform 1 0 106629 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1261
timestamp 1624857261
transform 1 0 106969 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1261
timestamp 1624857261
transform 1 0 106965 0 1 1691
box 0 0 1 1
use contact_7  contact_7_254
timestamp 1624857261
transform 1 0 107969 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1258
timestamp 1624857261
transform 1 0 107973 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1259
timestamp 1624857261
transform 1 0 107637 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1260
timestamp 1624857261
transform 1 0 107301 0 1 1691
box 0 0 1 1
use contact_19  contact_19_870
timestamp 1624857261
transform 1 0 107970 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1258
timestamp 1624857261
transform 1 0 107977 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1259
timestamp 1624857261
transform 1 0 107641 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1260
timestamp 1624857261
transform 1 0 107305 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3425
timestamp 1624857261
transform 1 0 107848 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1254
timestamp 1624857261
transform 1 0 109317 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1255
timestamp 1624857261
transform 1 0 108981 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1256
timestamp 1624857261
transform 1 0 108645 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1257
timestamp 1624857261
transform 1 0 108309 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1254
timestamp 1624857261
transform 1 0 109321 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1255
timestamp 1624857261
transform 1 0 108985 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1256
timestamp 1624857261
transform 1 0 108649 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1257
timestamp 1624857261
transform 1 0 108313 0 1 1683
box 0 0 1 1
use contact_7  contact_7_253
timestamp 1624857261
transform 1 0 109649 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1251
timestamp 1624857261
transform 1 0 110325 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1252
timestamp 1624857261
transform 1 0 109989 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1253
timestamp 1624857261
transform 1 0 109653 0 1 1691
box 0 0 1 1
use contact_19  contact_19_869
timestamp 1624857261
transform 1 0 109650 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1251
timestamp 1624857261
transform 1 0 110329 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1252
timestamp 1624857261
transform 1 0 109993 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1253
timestamp 1624857261
transform 1 0 109657 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3415
timestamp 1624857261
transform 1 0 109616 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1250
timestamp 1624857261
transform 1 0 110665 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1250
timestamp 1624857261
transform 1 0 110661 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1249
timestamp 1624857261
transform 1 0 110997 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1249
timestamp 1624857261
transform 1 0 111001 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1248
timestamp 1624857261
transform 1 0 111337 0 1 1683
box 0 0 1 1
use contact_19  contact_19_868
timestamp 1624857261
transform 1 0 111330 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1248
timestamp 1624857261
transform 1 0 111333 0 1 1691
box 0 0 1 1
use contact_7  contact_7_252
timestamp 1624857261
transform 1 0 111329 0 1 1687
box 0 0 1 1
use contact_33  contact_33_3411
timestamp 1624857261
transform 1 0 111384 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1247
timestamp 1624857261
transform 1 0 111673 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1247
timestamp 1624857261
transform 1 0 111669 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1246
timestamp 1624857261
transform 1 0 112009 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1246
timestamp 1624857261
transform 1 0 112005 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1245
timestamp 1624857261
transform 1 0 112345 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1245
timestamp 1624857261
transform 1 0 112341 0 1 1691
box 0 0 1 1
use contact_33  contact_33_3407
timestamp 1624857261
transform 1 0 112880 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1244
timestamp 1624857261
transform 1 0 112681 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1244
timestamp 1624857261
transform 1 0 112677 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1243
timestamp 1624857261
transform 1 0 113017 0 1 1683
box 0 0 1 1
use contact_19  contact_19_867
timestamp 1624857261
transform 1 0 113010 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1243
timestamp 1624857261
transform 1 0 113013 0 1 1691
box 0 0 1 1
use contact_7  contact_7_251
timestamp 1624857261
transform 1 0 113009 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1241
timestamp 1624857261
transform 1 0 113685 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1242
timestamp 1624857261
transform 1 0 113349 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1241
timestamp 1624857261
transform 1 0 113689 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1242
timestamp 1624857261
transform 1 0 113353 0 1 1683
box 0 0 1 1
use contact_33  contact_33_985
timestamp 1624857261
transform 1 0 109344 0 1 9525
box 0 0 1 1
use contact_33  contact_33_3466
timestamp 1624857261
transform 1 0 104584 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3438
timestamp 1624857261
transform 1 0 107168 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3434
timestamp 1624857261
transform 1 0 109208 0 1 10613
box 0 0 1 1
use contact_33  contact_33_3435
timestamp 1624857261
transform 1 0 109208 0 1 11021
box 0 0 1 1
use contact_33  contact_33_3491
timestamp 1624857261
transform 1 0 102272 0 1 11973
box 0 0 1 1
use contact_33  contact_33_997
timestamp 1624857261
transform 1 0 104448 0 1 11701
box 0 0 1 1
use contact_33  contact_33_998
timestamp 1624857261
transform 1 0 104448 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3467
timestamp 1624857261
transform 1 0 104584 0 1 11837
box 0 0 1 1
use contact_33  contact_33_3465
timestamp 1624857261
transform 1 0 104720 0 1 11973
box 0 0 1 1
use contact_33  contact_33_983
timestamp 1624857261
transform 1 0 107440 0 1 11701
box 0 0 1 1
use contact_33  contact_33_984
timestamp 1624857261
transform 1 0 107440 0 1 12245
box 0 0 1 1
use contact_33  contact_33_3437
timestamp 1624857261
transform 1 0 107304 0 1 11973
box 0 0 1 1
use contact_33  contact_33_3439
timestamp 1624857261
transform 1 0 107168 0 1 11837
box 0 0 1 1
use contact_33  contact_33_986
timestamp 1624857261
transform 1 0 109344 0 1 11293
box 0 0 1 1
use contact_33  contact_33_1004
timestamp 1624857261
transform 1 0 102408 0 1 13197
box 0 0 1 1
use contact_33  contact_33_1007
timestamp 1624857261
transform 1 0 102408 0 1 13061
box 0 0 1 1
use contact_33  contact_33_1008
timestamp 1624857261
transform 1 0 102408 0 1 12517
box 0 0 1 1
use contact_33  contact_33_3490
timestamp 1624857261
transform 1 0 102272 0 1 13469
box 0 0 1 1
use contact_7  contact_7_377
timestamp 1624857261
transform 1 0 104437 0 1 13196
box 0 0 1 1
use contact_19  contact_19_967
timestamp 1624857261
transform 1 0 104438 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5384
timestamp 1624857261
transform 1 0 104312 0 1 13061
box 0 0 1 1
use contact_33  contact_33_994
timestamp 1624857261
transform 1 0 104856 0 1 13197
box 0 0 1 1
use contact_33  contact_33_995
timestamp 1624857261
transform 1 0 104856 0 1 13061
box 0 0 1 1
use contact_33  contact_33_996
timestamp 1624857261
transform 1 0 104856 0 1 12517
box 0 0 1 1
use contact_33  contact_33_3464
timestamp 1624857261
transform 1 0 104720 0 1 13469
box 0 0 1 1
use contact_7  contact_7_376
timestamp 1624857261
transform 1 0 106933 0 1 13196
box 0 0 1 1
use contact_19  contact_19_966
timestamp 1624857261
transform 1 0 106934 0 1 13201
box 0 0 1 1
use contact_33  contact_33_5383
timestamp 1624857261
transform 1 0 106896 0 1 13061
box 0 0 1 1
use contact_33  contact_33_978
timestamp 1624857261
transform 1 0 107440 0 1 13197
box 0 0 1 1
use contact_33  contact_33_981
timestamp 1624857261
transform 1 0 107440 0 1 13061
box 0 0 1 1
use contact_33  contact_33_982
timestamp 1624857261
transform 1 0 107440 0 1 12517
box 0 0 1 1
use contact_33  contact_33_3436
timestamp 1624857261
transform 1 0 107304 0 1 13469
box 0 0 1 1
use contact_33  contact_33_3488
timestamp 1624857261
transform 1 0 102272 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3489
timestamp 1624857261
transform 1 0 102272 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3458
timestamp 1624857261
transform 1 0 104720 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3459
timestamp 1624857261
transform 1 0 104720 0 1 14285
box 0 0 1 1
use contact_33  contact_33_3432
timestamp 1624857261
transform 1 0 107304 0 1 13605
box 0 0 1 1
use contact_33  contact_33_3433
timestamp 1624857261
transform 1 0 107304 0 1 14285
box 0 0 1 1
use contact_33  contact_33_1000
timestamp 1624857261
transform 1 0 102272 0 1 15101
box 0 0 1 1
use contact_33  contact_33_1003
timestamp 1624857261
transform 1 0 102408 0 1 15101
box 0 0 1 1
use contact_33  contact_33_988
timestamp 1624857261
transform 1 0 104992 0 1 15101
box 0 0 1 1
use contact_33  contact_33_993
timestamp 1624857261
transform 1 0 104856 0 1 15101
box 0 0 1 1
use contact_33  contact_33_974
timestamp 1624857261
transform 1 0 107304 0 1 15101
box 0 0 1 1
use contact_33  contact_33_977
timestamp 1624857261
transform 1 0 107440 0 1 15101
box 0 0 1 1
use contact_33  contact_33_999
timestamp 1624857261
transform 1 0 102408 0 1 17005
box 0 0 1 1
use contact_33  contact_33_987
timestamp 1624857261
transform 1 0 104992 0 1 17005
box 0 0 1 1
use contact_33  contact_33_973
timestamp 1624857261
transform 1 0 107304 0 1 17005
box 0 0 1 1
use contact_33  contact_33_972
timestamp 1624857261
transform 1 0 110160 0 1 17141
box 0 0 1 1
use contact_33  contact_33_3402
timestamp 1624857261
transform 1 0 114648 0 1 1229
box 0 0 1 1
use contact_14  contact_14_1240
timestamp 1624857261
transform 1 0 114021 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1240
timestamp 1624857261
transform 1 0 114025 0 1 1683
box 0 0 1 1
use contact_7  contact_7_250
timestamp 1624857261
transform 1 0 114689 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1238
timestamp 1624857261
transform 1 0 114693 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1239
timestamp 1624857261
transform 1 0 114357 0 1 1691
box 0 0 1 1
use contact_19  contact_19_866
timestamp 1624857261
transform 1 0 114690 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1238
timestamp 1624857261
transform 1 0 114697 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1239
timestamp 1624857261
transform 1 0 114361 0 1 1683
box 0 0 1 1
use contact_33  contact_33_3403
timestamp 1624857261
transform 1 0 114648 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1234
timestamp 1624857261
transform 1 0 116037 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1235
timestamp 1624857261
transform 1 0 115701 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1236
timestamp 1624857261
transform 1 0 115365 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1237
timestamp 1624857261
transform 1 0 115029 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1234
timestamp 1624857261
transform 1 0 116041 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1235
timestamp 1624857261
transform 1 0 115705 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1236
timestamp 1624857261
transform 1 0 115369 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1237
timestamp 1624857261
transform 1 0 115033 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2690
timestamp 1624857261
transform 1 0 116280 0 1 1229
box 0 0 1 1
use contact_7  contact_7_249
timestamp 1624857261
transform 1 0 116369 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1233
timestamp 1624857261
transform 1 0 116373 0 1 1691
box 0 0 1 1
use contact_19  contact_19_865
timestamp 1624857261
transform 1 0 116370 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1233
timestamp 1624857261
transform 1 0 116377 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2691
timestamp 1624857261
transform 1 0 116280 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1232
timestamp 1624857261
transform 1 0 116709 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1232
timestamp 1624857261
transform 1 0 116713 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1230
timestamp 1624857261
transform 1 0 117381 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1231
timestamp 1624857261
transform 1 0 117045 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1230
timestamp 1624857261
transform 1 0 117385 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1231
timestamp 1624857261
transform 1 0 117049 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2528
timestamp 1624857261
transform 1 0 118048 0 1 1229
box 0 0 1 1
use contact_14  contact_14_1229
timestamp 1624857261
transform 1 0 117717 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1229
timestamp 1624857261
transform 1 0 117721 0 1 1683
box 0 0 1 1
use contact_7  contact_7_248
timestamp 1624857261
transform 1 0 118049 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1227
timestamp 1624857261
transform 1 0 118389 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1228
timestamp 1624857261
transform 1 0 118053 0 1 1691
box 0 0 1 1
use contact_19  contact_19_864
timestamp 1624857261
transform 1 0 118050 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1227
timestamp 1624857261
transform 1 0 118393 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1228
timestamp 1624857261
transform 1 0 118057 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2529
timestamp 1624857261
transform 1 0 118048 0 1 1637
box 0 0 1 1
use contact_33  contact_33_2508
timestamp 1624857261
transform 1 0 119680 0 1 1229
box 0 0 1 1
use contact_14  contact_14_1225
timestamp 1624857261
transform 1 0 119061 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1226
timestamp 1624857261
transform 1 0 118725 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1225
timestamp 1624857261
transform 1 0 119065 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1226
timestamp 1624857261
transform 1 0 118729 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1224
timestamp 1624857261
transform 1 0 119397 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1224
timestamp 1624857261
transform 1 0 119401 0 1 1683
box 0 0 1 1
use contact_7  contact_7_247
timestamp 1624857261
transform 1 0 119729 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1223
timestamp 1624857261
transform 1 0 119733 0 1 1691
box 0 0 1 1
use contact_19  contact_19_863
timestamp 1624857261
transform 1 0 119730 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1223
timestamp 1624857261
transform 1 0 119737 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2509
timestamp 1624857261
transform 1 0 119680 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1219
timestamp 1624857261
transform 1 0 121077 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1220
timestamp 1624857261
transform 1 0 120741 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1221
timestamp 1624857261
transform 1 0 120405 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1222
timestamp 1624857261
transform 1 0 120069 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1219
timestamp 1624857261
transform 1 0 121081 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1220
timestamp 1624857261
transform 1 0 120745 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1221
timestamp 1624857261
transform 1 0 120409 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1222
timestamp 1624857261
transform 1 0 120073 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2486
timestamp 1624857261
transform 1 0 121448 0 1 1229
box 0 0 1 1
use contact_7  contact_7_246
timestamp 1624857261
transform 1 0 121409 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1218
timestamp 1624857261
transform 1 0 121413 0 1 1691
box 0 0 1 1
use contact_19  contact_19_862
timestamp 1624857261
transform 1 0 121410 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1218
timestamp 1624857261
transform 1 0 121417 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2487
timestamp 1624857261
transform 1 0 121448 0 1 1637
box 0 0 1 1
use contact_14  contact_14_1217
timestamp 1624857261
transform 1 0 121749 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1217
timestamp 1624857261
transform 1 0 121753 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1216
timestamp 1624857261
transform 1 0 122085 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1216
timestamp 1624857261
transform 1 0 122089 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1215
timestamp 1624857261
transform 1 0 122421 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1215
timestamp 1624857261
transform 1 0 122425 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2488
timestamp 1624857261
transform 1 0 121312 0 1 18501
box 0 0 1 1
use contact_33  contact_33_2480
timestamp 1624857261
transform 1 0 122944 0 1 1229
box 0 0 1 1
use contact_33  contact_33_2481
timestamp 1624857261
transform 1 0 122944 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1214
timestamp 1624857261
transform 1 0 122761 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1214
timestamp 1624857261
transform 1 0 122757 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1213
timestamp 1624857261
transform 1 0 123097 0 1 1683
box 0 0 1 1
use contact_19  contact_19_861
timestamp 1624857261
transform 1 0 123090 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1213
timestamp 1624857261
transform 1 0 123093 0 1 1691
box 0 0 1 1
use contact_7  contact_7_245
timestamp 1624857261
transform 1 0 123089 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1212
timestamp 1624857261
transform 1 0 123433 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1212
timestamp 1624857261
transform 1 0 123429 0 1 1691
box 0 0 1 1
use contact_7  contact_7_443
timestamp 1624857261
transform 1 0 122766 0 1 9132
box 0 0 1 1
use contact_7  contact_7_444
timestamp 1624857261
transform 1 0 123664 0 1 9132
box 0 0 1 1
use contact_19  contact_19_998
timestamp 1624857261
transform 1 0 122767 0 1 9137
box 0 0 1 1
use contact_7  contact_7_445
timestamp 1624857261
transform 1 0 122846 0 1 10690
box 0 0 1 1
use contact_7  contact_7_446
timestamp 1624857261
transform 1 0 123664 0 1 10690
box 0 0 1 1
use contact_19  contact_19_999
timestamp 1624857261
transform 1 0 122847 0 1 10695
box 0 0 1 1
use contact_7  contact_7_447
timestamp 1624857261
transform 1 0 122926 0 1 11960
box 0 0 1 1
use contact_7  contact_7_448
timestamp 1624857261
transform 1 0 123664 0 1 11960
box 0 0 1 1
use contact_19  contact_19_1000
timestamp 1624857261
transform 1 0 122927 0 1 11965
box 0 0 1 1
use contact_7  contact_7_449
timestamp 1624857261
transform 1 0 123006 0 1 13518
box 0 0 1 1
use contact_7  contact_7_450
timestamp 1624857261
transform 1 0 123664 0 1 13518
box 0 0 1 1
use contact_19  contact_19_1001
timestamp 1624857261
transform 1 0 123007 0 1 13523
box 0 0 1 1
use contact_7  contact_7_451
timestamp 1624857261
transform 1 0 123086 0 1 14788
box 0 0 1 1
use contact_7  contact_7_452
timestamp 1624857261
transform 1 0 123664 0 1 14788
box 0 0 1 1
use contact_19  contact_19_1002
timestamp 1624857261
transform 1 0 123087 0 1 14793
box 0 0 1 1
use contact_7  contact_7_453
timestamp 1624857261
transform 1 0 123166 0 1 16346
box 0 0 1 1
use contact_7  contact_7_454
timestamp 1624857261
transform 1 0 123664 0 1 16346
box 0 0 1 1
use contact_19  contact_19_1003
timestamp 1624857261
transform 1 0 123167 0 1 16351
box 0 0 1 1
use contact_7  contact_7_455
timestamp 1624857261
transform 1 0 123246 0 1 17616
box 0 0 1 1
use contact_7  contact_7_456
timestamp 1624857261
transform 1 0 123664 0 1 17616
box 0 0 1 1
use contact_19  contact_19_1004
timestamp 1624857261
transform 1 0 123247 0 1 17621
box 0 0 1 1
use row_addr_dff  row_addr_dff_0
timestamp 1624857261
transform -1 0 124812 0 -1 19846
box -36 -49 1204 9951
use contact_14  contact_14_1211
timestamp 1624857261
transform 1 0 123765 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1211
timestamp 1624857261
transform 1 0 123769 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1210
timestamp 1624857261
transform 1 0 124101 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1210
timestamp 1624857261
transform 1 0 124105 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1209
timestamp 1624857261
transform 1 0 124437 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1209
timestamp 1624857261
transform 1 0 124441 0 1 1683
box 0 0 1 1
use contact_7  contact_7_244
timestamp 1624857261
transform 1 0 124769 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1208
timestamp 1624857261
transform 1 0 124773 0 1 1691
box 0 0 1 1
use contact_19  contact_19_860
timestamp 1624857261
transform 1 0 124770 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1208
timestamp 1624857261
transform 1 0 124777 0 1 1683
box 0 0 1 1
use contact_33  contact_33_12
timestamp 1624857261
transform 1 0 124168 0 1 8573
box 0 0 1 1
use contact_33  contact_33_5417
timestamp 1624857261
transform 1 0 124712 0 1 8981
box 0 0 1 1
use contact_7  contact_7_318
timestamp 1624857261
transform 1 0 124609 0 1 9061
box 0 0 1 1
use contact_33  contact_33_2470
timestamp 1624857261
transform 1 0 124304 0 1 9933
box 0 0 1 1
use contact_33  contact_33_5416
timestamp 1624857261
transform 1 0 124576 0 1 10749
box 0 0 1 1
use contact_7  contact_7_319
timestamp 1624857261
transform 1 0 124609 0 1 10761
box 0 0 1 1
use contact_33  contact_33_13
timestamp 1624857261
transform 1 0 124168 0 1 11429
box 0 0 1 1
use contact_33  contact_33_11
timestamp 1624857261
transform 1 0 124168 0 1 11293
box 0 0 1 1
use contact_33  contact_33_5415
timestamp 1624857261
transform 1 0 124440 0 1 11837
box 0 0 1 1
use contact_7  contact_7_320
timestamp 1624857261
transform 1 0 124609 0 1 11889
box 0 0 1 1
use contact_33  contact_33_2471
timestamp 1624857261
transform 1 0 124304 0 1 12653
box 0 0 1 1
use contact_33  contact_33_2473
timestamp 1624857261
transform 1 0 124304 0 1 12789
box 0 0 1 1
use contact_33  contact_33_5382
timestamp 1624857261
transform 1 0 124848 0 1 13469
box 0 0 1 1
use contact_7  contact_7_321
timestamp 1624857261
transform 1 0 124609 0 1 13589
box 0 0 1 1
use contact_33  contact_33_16
timestamp 1624857261
transform 1 0 124440 0 1 14285
box 0 0 1 1
use contact_33  contact_33_14
timestamp 1624857261
transform 1 0 124168 0 1 14013
box 0 0 1 1
use contact_7  contact_7_322
timestamp 1624857261
transform 1 0 124609 0 1 14717
box 0 0 1 1
use contact_33  contact_33_2474
timestamp 1624857261
transform 1 0 124168 0 1 15645
box 0 0 1 1
use contact_33  contact_33_2472
timestamp 1624857261
transform 1 0 124304 0 1 15509
box 0 0 1 1
use contact_7  contact_7_323
timestamp 1624857261
transform 1 0 124609 0 1 16417
box 0 0 1 1
use contact_33  contact_33_15
timestamp 1624857261
transform 1 0 124440 0 1 16869
box 0 0 1 1
use contact_33  contact_33_10
timestamp 1624857261
transform 1 0 124304 0 1 17005
box 0 0 1 1
use contact_7  contact_7_324
timestamp 1624857261
transform 1 0 124609 0 1 17545
box 0 0 1 1
use contact_33  contact_33_2475
timestamp 1624857261
transform 1 0 124168 0 1 18365
box 0 0 1 1
use contact_14  contact_14_1207
timestamp 1624857261
transform 1 0 125109 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1207
timestamp 1624857261
transform 1 0 125113 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2468
timestamp 1624857261
transform 1 0 125120 0 1 1229
box 0 0 1 1
use contact_33  contact_33_2469
timestamp 1624857261
transform 1 0 125120 0 1 1637
box 0 0 1 1
use contact_33  contact_33_2462
timestamp 1624857261
transform 1 0 126344 0 1 1229
box 0 0 1 1
use contact_13  contact_13_1206
timestamp 1624857261
transform 1 0 125449 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1206
timestamp 1624857261
transform 1 0 125445 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1205
timestamp 1624857261
transform 1 0 125785 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1204
timestamp 1624857261
transform 1 0 126121 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1205
timestamp 1624857261
transform 1 0 125781 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1204
timestamp 1624857261
transform 1 0 126117 0 1 1691
box 0 0 1 1
use contact_33  contact_33_2463
timestamp 1624857261
transform 1 0 126344 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1203
timestamp 1624857261
transform 1 0 126457 0 1 1683
box 0 0 1 1
use contact_19  contact_19_859
timestamp 1624857261
transform 1 0 126450 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1203
timestamp 1624857261
transform 1 0 126453 0 1 1691
box 0 0 1 1
use contact_7  contact_7_243
timestamp 1624857261
transform 1 0 126449 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1202
timestamp 1624857261
transform 1 0 126793 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1202
timestamp 1624857261
transform 1 0 126789 0 1 1691
box 0 0 1 1
use contact_33  contact_33_2458
timestamp 1624857261
transform 1 0 128112 0 1 1229
box 0 0 1 1
use contact_13  contact_13_1201
timestamp 1624857261
transform 1 0 127129 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1201
timestamp 1624857261
transform 1 0 127125 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1200
timestamp 1624857261
transform 1 0 127465 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1200
timestamp 1624857261
transform 1 0 127461 0 1 1691
box 0 0 1 1
use contact_33  contact_33_2459
timestamp 1624857261
transform 1 0 128112 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1199
timestamp 1624857261
transform 1 0 127801 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1198
timestamp 1624857261
transform 1 0 128137 0 1 1683
box 0 0 1 1
use contact_19  contact_19_858
timestamp 1624857261
transform 1 0 128130 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1199
timestamp 1624857261
transform 1 0 127797 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1198
timestamp 1624857261
transform 1 0 128133 0 1 1691
box 0 0 1 1
use contact_7  contact_7_242
timestamp 1624857261
transform 1 0 128129 0 1 1687
box 0 0 1 1
use contact_13  contact_13_1197
timestamp 1624857261
transform 1 0 128473 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1197
timestamp 1624857261
transform 1 0 128469 0 1 1691
box 0 0 1 1
use contact_33  contact_33_2455
timestamp 1624857261
transform 1 0 129880 0 1 1637
box 0 0 1 1
use contact_33  contact_33_2454
timestamp 1624857261
transform 1 0 129880 0 1 1229
box 0 0 1 1
use contact_13  contact_13_1196
timestamp 1624857261
transform 1 0 128809 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1196
timestamp 1624857261
transform 1 0 128805 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1195
timestamp 1624857261
transform 1 0 129145 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1195
timestamp 1624857261
transform 1 0 129141 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1194
timestamp 1624857261
transform 1 0 129481 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1193
timestamp 1624857261
transform 1 0 129817 0 1 1683
box 0 0 1 1
use contact_19  contact_19_857
timestamp 1624857261
transform 1 0 129810 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1194
timestamp 1624857261
transform 1 0 129477 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1193
timestamp 1624857261
transform 1 0 129813 0 1 1691
box 0 0 1 1
use contact_7  contact_7_241
timestamp 1624857261
transform 1 0 129809 0 1 1687
box 0 0 1 1
use contact_33  contact_33_2452
timestamp 1624857261
transform 1 0 131376 0 1 1229
box 0 0 1 1
use contact_13  contact_13_1192
timestamp 1624857261
transform 1 0 130153 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1191
timestamp 1624857261
transform 1 0 130489 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1192
timestamp 1624857261
transform 1 0 130149 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1191
timestamp 1624857261
transform 1 0 130485 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1190
timestamp 1624857261
transform 1 0 130825 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1190
timestamp 1624857261
transform 1 0 130821 0 1 1691
box 0 0 1 1
use contact_33  contact_33_2453
timestamp 1624857261
transform 1 0 131376 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1189
timestamp 1624857261
transform 1 0 131161 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1189
timestamp 1624857261
transform 1 0 131157 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1188
timestamp 1624857261
transform 1 0 131497 0 1 1683
box 0 0 1 1
use contact_19  contact_19_856
timestamp 1624857261
transform 1 0 131490 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1188
timestamp 1624857261
transform 1 0 131493 0 1 1691
box 0 0 1 1
use contact_7  contact_7_240
timestamp 1624857261
transform 1 0 131489 0 1 1687
box 0 0 1 1
use contact_33  contact_33_2446
timestamp 1624857261
transform 1 0 133144 0 1 1229
box 0 0 1 1
use contact_13  contact_13_1187
timestamp 1624857261
transform 1 0 131833 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1187
timestamp 1624857261
transform 1 0 131829 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1186
timestamp 1624857261
transform 1 0 132169 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1185
timestamp 1624857261
transform 1 0 132505 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1186
timestamp 1624857261
transform 1 0 132165 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1185
timestamp 1624857261
transform 1 0 132501 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1184
timestamp 1624857261
transform 1 0 132841 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1184
timestamp 1624857261
transform 1 0 132837 0 1 1691
box 0 0 1 1
use contact_33  contact_33_2447
timestamp 1624857261
transform 1 0 133144 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1183
timestamp 1624857261
transform 1 0 133177 0 1 1683
box 0 0 1 1
use contact_19  contact_19_855
timestamp 1624857261
transform 1 0 133170 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1183
timestamp 1624857261
transform 1 0 133173 0 1 1691
box 0 0 1 1
use contact_7  contact_7_239
timestamp 1624857261
transform 1 0 133169 0 1 1687
box 0 0 1 1
use contact_33  contact_33_2442
timestamp 1624857261
transform 1 0 134776 0 1 1229
box 0 0 1 1
use contact_13  contact_13_1182
timestamp 1624857261
transform 1 0 133513 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1182
timestamp 1624857261
transform 1 0 133509 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1181
timestamp 1624857261
transform 1 0 133849 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1180
timestamp 1624857261
transform 1 0 134185 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1181
timestamp 1624857261
transform 1 0 133845 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1180
timestamp 1624857261
transform 1 0 134181 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1179
timestamp 1624857261
transform 1 0 134521 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1179
timestamp 1624857261
transform 1 0 134517 0 1 1691
box 0 0 1 1
use contact_33  contact_33_2443
timestamp 1624857261
transform 1 0 134776 0 1 1637
box 0 0 1 1
use contact_13  contact_13_1178
timestamp 1624857261
transform 1 0 134857 0 1 1683
box 0 0 1 1
use contact_19  contact_19_854
timestamp 1624857261
transform 1 0 134850 0 1 1692
box 0 0 1 1
use contact_14  contact_14_1178
timestamp 1624857261
transform 1 0 134853 0 1 1691
box 0 0 1 1
use contact_7  contact_7_238
timestamp 1624857261
transform 1 0 134849 0 1 1687
box 0 0 1 1
use contact_33  contact_33_3870
timestamp 1624857261
transform 1 0 69088 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3871
timestamp 1624857261
transform 1 0 69088 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3874
timestamp 1624857261
transform 1 0 68408 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3875
timestamp 1624857261
transform 1 0 68408 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3880
timestamp 1624857261
transform 1 0 67864 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3881
timestamp 1624857261
transform 1 0 67864 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3840
timestamp 1624857261
transform 1 0 71536 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3841
timestamp 1624857261
transform 1 0 71536 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3846
timestamp 1624857261
transform 1 0 70856 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3847
timestamp 1624857261
transform 1 0 70856 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3850
timestamp 1624857261
transform 1 0 70312 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3851
timestamp 1624857261
transform 1 0 70312 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3792
timestamp 1624857261
transform 1 0 75344 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3793
timestamp 1624857261
transform 1 0 75344 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3804
timestamp 1624857261
transform 1 0 75208 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3805
timestamp 1624857261
transform 1 0 75208 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3806
timestamp 1624857261
transform 1 0 74664 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3807
timestamp 1624857261
transform 1 0 74664 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3818
timestamp 1624857261
transform 1 0 73304 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3819
timestamp 1624857261
transform 1 0 73304 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3754
timestamp 1624857261
transform 1 0 77928 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3755
timestamp 1624857261
transform 1 0 77928 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3776
timestamp 1624857261
transform 1 0 77112 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3777
timestamp 1624857261
transform 1 0 77112 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3780
timestamp 1624857261
transform 1 0 76568 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3781
timestamp 1624857261
transform 1 0 76568 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3788
timestamp 1624857261
transform 1 0 75888 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3789
timestamp 1624857261
transform 1 0 75888 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3752
timestamp 1624857261
transform 1 0 78336 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3753
timestamp 1624857261
transform 1 0 78336 0 1 18909
box 0 0 1 1
use contact_33  contact_33_3716
timestamp 1624857261
transform 1 0 81600 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3717
timestamp 1624857261
transform 1 0 81600 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3724
timestamp 1624857261
transform 1 0 81464 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3725
timestamp 1624857261
transform 1 0 81464 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3728
timestamp 1624857261
transform 1 0 80512 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3729
timestamp 1624857261
transform 1 0 80512 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3748
timestamp 1624857261
transform 1 0 79152 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3749
timestamp 1624857261
transform 1 0 79152 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3688
timestamp 1624857261
transform 1 0 84048 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3689
timestamp 1624857261
transform 1 0 84048 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3694
timestamp 1624857261
transform 1 0 83368 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3695
timestamp 1624857261
transform 1 0 83368 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3698
timestamp 1624857261
transform 1 0 82824 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3699
timestamp 1624857261
transform 1 0 82824 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3714
timestamp 1624857261
transform 1 0 82008 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3715
timestamp 1624857261
transform 1 0 82008 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3683
timestamp 1624857261
transform 1 0 84592 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3682
timestamp 1624857261
transform 1 0 84592 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3671
timestamp 1624857261
transform 1 0 85272 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3670
timestamp 1624857261
transform 1 0 85272 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3667
timestamp 1624857261
transform 1 0 85816 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3666
timestamp 1624857261
transform 1 0 85816 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3659
timestamp 1624857261
transform 1 0 86496 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3658
timestamp 1624857261
transform 1 0 86496 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3655
timestamp 1624857261
transform 1 0 86768 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3654
timestamp 1624857261
transform 1 0 86768 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3640
timestamp 1624857261
transform 1 0 88128 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3641
timestamp 1624857261
transform 1 0 88128 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3614
timestamp 1624857261
transform 1 0 90304 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3615
timestamp 1624857261
transform 1 0 90304 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3624
timestamp 1624857261
transform 1 0 89624 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3625
timestamp 1624857261
transform 1 0 89624 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3590
timestamp 1624857261
transform 1 0 92752 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3591
timestamp 1624857261
transform 1 0 92752 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3600
timestamp 1624857261
transform 1 0 92072 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3601
timestamp 1624857261
transform 1 0 92072 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3610
timestamp 1624857261
transform 1 0 90848 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3611
timestamp 1624857261
transform 1 0 90848 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3558
timestamp 1624857261
transform 1 0 95744 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3559
timestamp 1624857261
transform 1 0 95744 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3562
timestamp 1624857261
transform 1 0 95336 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3563
timestamp 1624857261
transform 1 0 95336 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3578
timestamp 1624857261
transform 1 0 94248 0 1 19317
box 0 0 1 1
use contact_33  contact_33_3579
timestamp 1624857261
transform 1 0 94248 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3580
timestamp 1624857261
transform 1 0 94384 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3581
timestamp 1624857261
transform 1 0 94384 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3532
timestamp 1624857261
transform 1 0 98328 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3533
timestamp 1624857261
transform 1 0 98328 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3552
timestamp 1624857261
transform 1 0 96560 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3553
timestamp 1624857261
transform 1 0 96560 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3500
timestamp 1624857261
transform 1 0 101592 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3501
timestamp 1624857261
transform 1 0 101592 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3508
timestamp 1624857261
transform 1 0 100368 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3509
timestamp 1624857261
transform 1 0 100368 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3522
timestamp 1624857261
transform 1 0 99552 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3523
timestamp 1624857261
transform 1 0 99552 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3528
timestamp 1624857261
transform 1 0 99144 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3529
timestamp 1624857261
transform 1 0 99144 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3494
timestamp 1624857261
transform 1 0 102000 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3495
timestamp 1624857261
transform 1 0 102000 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3474
timestamp 1624857261
transform 1 0 104040 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3475
timestamp 1624857261
transform 1 0 104040 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3484
timestamp 1624857261
transform 1 0 102952 0 1 19317
box 0 0 1 1
use contact_33  contact_33_3485
timestamp 1624857261
transform 1 0 102952 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3452
timestamp 1624857261
transform 1 0 105808 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3453
timestamp 1624857261
transform 1 0 105808 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3454
timestamp 1624857261
transform 1 0 105264 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3455
timestamp 1624857261
transform 1 0 105264 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3470
timestamp 1624857261
transform 1 0 104584 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3471
timestamp 1624857261
transform 1 0 104584 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3422
timestamp 1624857261
transform 1 0 108256 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3423
timestamp 1624857261
transform 1 0 108256 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3442
timestamp 1624857261
transform 1 0 107032 0 1 19181
box 0 0 1 1
use contact_33  contact_33_3443
timestamp 1624857261
transform 1 0 107032 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3444
timestamp 1624857261
transform 1 0 106624 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3445
timestamp 1624857261
transform 1 0 106624 0 1 19181
box 0 0 1 1
use contact_33  contact_33_971
timestamp 1624857261
transform 1 0 110160 0 1 19725
box 0 0 1 1
use contact_33  contact_33_3420
timestamp 1624857261
transform 1 0 109072 0 1 18773
box 0 0 1 1
use contact_33  contact_33_3421
timestamp 1624857261
transform 1 0 109072 0 1 19181
box 0 0 1 1
use contact_33  contact_33_923
timestamp 1624857261
transform 1 0 110160 0 1 22445
box 0 0 1 1
use contact_33  contact_33_924
timestamp 1624857261
transform 1 0 110160 0 1 22717
box 0 0 1 1
use contact_33  contact_33_926
timestamp 1624857261
transform 1 0 110432 0 1 22853
box 0 0 1 1
use contact_33  contact_33_837
timestamp 1624857261
transform 1 0 110432 0 1 23669
box 0 0 1 1
use contact_33  contact_33_838
timestamp 1624857261
transform 1 0 110432 0 1 23941
box 0 0 1 1
use contact_33  contact_33_925
timestamp 1624857261
transform 1 0 110432 0 1 23125
box 0 0 1 1
use contact_33  contact_33_839
timestamp 1624857261
transform 1 0 110432 0 1 26253
box 0 0 1 1
use contact_33  contact_33_840
timestamp 1624857261
transform 1 0 110432 0 1 25981
box 0 0 1 1
use contact_33  contact_33_935
timestamp 1624857261
transform 1 0 110296 0 1 26389
box 0 0 1 1
use contact_33  contact_33_936
timestamp 1624857261
transform 1 0 110296 0 1 26661
box 0 0 1 1
use contact_33  contact_33_937
timestamp 1624857261
transform 1 0 110296 0 1 27069
box 0 0 1 1
use contact_33  contact_33_938
timestamp 1624857261
transform 1 0 110296 0 1 26797
box 0 0 1 1
use contact_33  contact_33_953
timestamp 1624857261
transform 1 0 110160 0 1 27341
box 0 0 1 1
use contact_33  contact_33_954
timestamp 1624857261
transform 1 0 110160 0 1 27069
box 0 0 1 1
use contact_33  contact_33_831
timestamp 1624857261
transform 1 0 110160 0 1 31557
box 0 0 1 1
use contact_33  contact_33_931
timestamp 1624857261
transform 1 0 110432 0 1 30333
box 0 0 1 1
use contact_33  contact_33_932
timestamp 1624857261
transform 1 0 110432 0 1 30605
box 0 0 1 1
use contact_33  contact_33_967
timestamp 1624857261
transform 1 0 110160 0 1 30197
box 0 0 1 1
use contact_33  contact_33_968
timestamp 1624857261
transform 1 0 110160 0 1 29925
box 0 0 1 1
use contact_33  contact_33_832
timestamp 1624857261
transform 1 0 110160 0 1 31829
box 0 0 1 1
use contact_33  contact_33_889
timestamp 1624857261
transform 1 0 110160 0 1 34413
box 0 0 1 1
use contact_33  contact_33_890
timestamp 1624857261
transform 1 0 110160 0 1 34685
box 0 0 1 1
use contact_33  contact_33_899
timestamp 1624857261
transform 1 0 110296 0 1 35773
box 0 0 1 1
use contact_33  contact_33_900
timestamp 1624857261
transform 1 0 110296 0 1 35501
box 0 0 1 1
use contact_33  contact_33_957
timestamp 1624857261
transform 1 0 110432 0 1 34685
box 0 0 1 1
use contact_33  contact_33_958
timestamp 1624857261
transform 1 0 110432 0 1 34957
box 0 0 1 1
use contact_32  contact_32_1
timestamp 1624857261
transform 1 0 123527 0 1 19501
box 0 0 1 1
use contact_7  contact_7_457
timestamp 1624857261
transform 1 0 123326 0 1 19174
box 0 0 1 1
use contact_7  contact_7_458
timestamp 1624857261
transform 1 0 123664 0 1 19174
box 0 0 1 1
use contact_19  contact_19_1005
timestamp 1624857261
transform 1 0 123327 0 1 19179
box 0 0 1 1
use contact_7  contact_7_325
timestamp 1624857261
transform 1 0 124609 0 1 19245
box 0 0 1 1
use contact_33  contact_33_3221
timestamp 1624857261
transform 1 0 115192 0 1 20269
box 0 0 1 1
use contact_33  contact_33_764
timestamp 1624857261
transform 1 0 115600 0 1 20269
box 0 0 1 1
use contact_33  contact_33_2830
timestamp 1624857261
transform 1 0 116008 0 1 20269
box 0 0 1 1
use contact_33  contact_33_246
timestamp 1624857261
transform 1 0 116960 0 1 20269
box 0 0 1 1
use contact_33  contact_33_2515
timestamp 1624857261
transform 1 0 118864 0 1 20269
box 0 0 1 1
use contact_33  contact_33_45
timestamp 1624857261
transform 1 0 119408 0 1 20269
box 0 0 1 1
use contact_33  contact_33_2507
timestamp 1624857261
transform 1 0 119816 0 1 20269
box 0 0 1 1
use contact_33  contact_33_2489
timestamp 1624857261
transform 1 0 121312 0 1 20133
box 0 0 1 1
use contact_33  contact_33_9
timestamp 1624857261
transform 1 0 124304 0 1 19725
box 0 0 1 1
use contact_33  contact_33_25
timestamp 1624857261
transform 1 0 124168 0 1 19861
box 0 0 1 1
use contact_33  contact_33_26
timestamp 1624857261
transform 1 0 124168 0 1 20133
box 0 0 1 1
use contact_33  contact_33_3098
timestamp 1624857261
transform 1 0 115192 0 1 20949
box 0 0 1 1
use contact_33  contact_33_3099
timestamp 1624857261
transform 1 0 115192 0 1 20677
box 0 0 1 1
use contact_33  contact_33_3220
timestamp 1624857261
transform 1 0 115192 0 1 20541
box 0 0 1 1
use contact_33  contact_33_651
timestamp 1624857261
transform 1 0 115600 0 1 20949
box 0 0 1 1
use contact_33  contact_33_652
timestamp 1624857261
transform 1 0 115600 0 1 20677
box 0 0 1 1
use contact_33  contact_33_763
timestamp 1624857261
transform 1 0 115600 0 1 20541
box 0 0 1 1
use contact_33  contact_33_767
timestamp 1624857261
transform 1 0 115600 0 1 21085
box 0 0 1 1
use contact_33  contact_33_2725
timestamp 1624857261
transform 1 0 116008 0 1 21085
box 0 0 1 1
use contact_33  contact_33_2828
timestamp 1624857261
transform 1 0 116008 0 1 20949
box 0 0 1 1
use contact_33  contact_33_2829
timestamp 1624857261
transform 1 0 116008 0 1 20677
box 0 0 1 1
use contact_33  contact_33_2831
timestamp 1624857261
transform 1 0 116008 0 1 20541
box 0 0 1 1
use contact_33  contact_33_3047
timestamp 1624857261
transform 1 0 115328 0 1 21085
box 0 0 1 1
use contact_33  contact_33_127
timestamp 1624857261
transform 1 0 116824 0 1 20677
box 0 0 1 1
use contact_33  contact_33_128
timestamp 1624857261
transform 1 0 116824 0 1 20949
box 0 0 1 1
use contact_33  contact_33_245
timestamp 1624857261
transform 1 0 116960 0 1 20541
box 0 0 1 1
use contact_33  contact_33_329
timestamp 1624857261
transform 1 0 116960 0 1 21085
box 0 0 1 1
use contact_33  contact_33_2514
timestamp 1624857261
transform 1 0 118864 0 1 20949
box 0 0 1 1
use contact_33  contact_33_2520
timestamp 1624857261
transform 1 0 119000 0 1 21085
box 0 0 1 1
use contact_33  contact_33_46
timestamp 1624857261
transform 1 0 119408 0 1 20949
box 0 0 1 1
use contact_33  contact_33_2506
timestamp 1624857261
transform 1 0 119816 0 1 20949
box 0 0 1 1
use contact_33  contact_33_42
timestamp 1624857261
transform 1 0 120496 0 1 21085
box 0 0 1 1
use contact_33  contact_33_3022
timestamp 1624857261
transform 1 0 115192 0 1 21493
box 0 0 1 1
use contact_33  contact_33_3023
timestamp 1624857261
transform 1 0 115192 0 1 21765
box 0 0 1 1
use contact_33  contact_33_765
timestamp 1624857261
transform 1 0 115600 0 1 21765
box 0 0 1 1
use contact_33  contact_33_766
timestamp 1624857261
transform 1 0 115600 0 1 21493
box 0 0 1 1
use contact_33  contact_33_768
timestamp 1624857261
transform 1 0 115600 0 1 21357
box 0 0 1 1
use contact_33  contact_33_2724
timestamp 1624857261
transform 1 0 116008 0 1 21357
box 0 0 1 1
use contact_33  contact_33_3046
timestamp 1624857261
transform 1 0 115328 0 1 21357
box 0 0 1 1
use contact_33  contact_33_2588
timestamp 1624857261
transform 1 0 116552 0 1 21765
box 0 0 1 1
use contact_33  contact_33_2589
timestamp 1624857261
transform 1 0 116552 0 1 21493
box 0 0 1 1
use contact_33  contact_33_330
timestamp 1624857261
transform 1 0 116960 0 1 21357
box 0 0 1 1
use contact_33  contact_33_331
timestamp 1624857261
transform 1 0 116960 0 1 21765
box 0 0 1 1
use contact_33  contact_33_332
timestamp 1624857261
transform 1 0 116960 0 1 21493
box 0 0 1 1
use contact_33  contact_33_171
timestamp 1624857261
transform 1 0 116824 0 1 22581
box 0 0 1 1
use contact_33  contact_33_172
timestamp 1624857261
transform 1 0 116824 0 1 22309
box 0 0 1 1
use contact_33  contact_33_173
timestamp 1624857261
transform 1 0 116824 0 1 21901
box 0 0 1 1
use contact_33  contact_33_174
timestamp 1624857261
transform 1 0 116824 0 1 22173
box 0 0 1 1
use contact_33  contact_33_2812
timestamp 1624857261
transform 1 0 116280 0 1 22309
box 0 0 1 1
use contact_33  contact_33_2813
timestamp 1624857261
transform 1 0 116280 0 1 22581
box 0 0 1 1
use contact_33  contact_33_2521
timestamp 1624857261
transform 1 0 119000 0 1 22445
box 0 0 1 1
use contact_33  contact_33_41
timestamp 1624857261
transform 1 0 120496 0 1 22581
box 0 0 1 1
use contact_33  contact_33_638
timestamp 1624857261
transform 1 0 115736 0 1 23397
box 0 0 1 1
use contact_33  contact_33_693
timestamp 1624857261
transform 1 0 115736 0 1 23261
box 0 0 1 1
use contact_33  contact_33_694
timestamp 1624857261
transform 1 0 115736 0 1 22989
box 0 0 1 1
use contact_33  contact_33_3037
timestamp 1624857261
transform 1 0 115328 0 1 23397
box 0 0 1 1
use contact_33  contact_33_3228
timestamp 1624857261
transform 1 0 115328 0 1 23261
box 0 0 1 1
use contact_33  contact_33_3229
timestamp 1624857261
transform 1 0 115328 0 1 22989
box 0 0 1 1
use contact_33  contact_33_191
timestamp 1624857261
transform 1 0 116824 0 1 22717
box 0 0 1 1
use contact_33  contact_33_192
timestamp 1624857261
transform 1 0 116824 0 1 22989
box 0 0 1 1
use contact_33  contact_33_2848
timestamp 1624857261
transform 1 0 116280 0 1 23261
box 0 0 1 1
use contact_33  contact_33_2849
timestamp 1624857261
transform 1 0 116280 0 1 22989
box 0 0 1 1
use contact_33  contact_33_2523
timestamp 1624857261
transform 1 0 119000 0 1 23397
box 0 0 1 1
use contact_33  contact_33_2524
timestamp 1624857261
transform 1 0 119000 0 1 22717
box 0 0 1 1
use contact_33  contact_33_2525
timestamp 1624857261
transform 1 0 119000 0 1 23261
box 0 0 1 1
use contact_33  contact_33_58
timestamp 1624857261
transform 1 0 119272 0 1 23397
box 0 0 1 1
use contact_33  contact_33_59
timestamp 1624857261
transform 1 0 119272 0 1 22717
box 0 0 1 1
use contact_33  contact_33_60
timestamp 1624857261
transform 1 0 119272 0 1 23261
box 0 0 1 1
use contact_33  contact_33_2496
timestamp 1624857261
transform 1 0 119680 0 1 22717
box 0 0 1 1
use contact_33  contact_33_2497
timestamp 1624857261
transform 1 0 119680 0 1 23261
box 0 0 1 1
use contact_33  contact_33_35
timestamp 1624857261
transform 1 0 120632 0 1 23261
box 0 0 1 1
use contact_33  contact_33_36
timestamp 1624857261
transform 1 0 120632 0 1 22717
box 0 0 1 1
use contact_33  contact_33_3276
timestamp 1624857261
transform 1 0 115192 0 1 24213
box 0 0 1 1
use contact_33  contact_33_469
timestamp 1624857261
transform 1 0 115736 0 1 23805
box 0 0 1 1
use contact_33  contact_33_470
timestamp 1624857261
transform 1 0 115736 0 1 24077
box 0 0 1 1
use contact_33  contact_33_637
timestamp 1624857261
transform 1 0 115736 0 1 23669
box 0 0 1 1
use contact_33  contact_33_657
timestamp 1624857261
transform 1 0 115736 0 1 24213
box 0 0 1 1
use contact_33  contact_33_2976
timestamp 1624857261
transform 1 0 116008 0 1 24213
box 0 0 1 1
use contact_33  contact_33_3036
timestamp 1624857261
transform 1 0 115328 0 1 23669
box 0 0 1 1
use contact_33  contact_33_3148
timestamp 1624857261
transform 1 0 115328 0 1 23805
box 0 0 1 1
use contact_33  contact_33_3149
timestamp 1624857261
transform 1 0 115328 0 1 24077
box 0 0 1 1
use contact_33  contact_33_72
timestamp 1624857261
transform 1 0 116824 0 1 24213
box 0 0 1 1
use contact_33  contact_33_2648
timestamp 1624857261
transform 1 0 116552 0 1 24077
box 0 0 1 1
use contact_33  contact_33_2649
timestamp 1624857261
transform 1 0 116552 0 1 23805
box 0 0 1 1
use contact_33  contact_33_2852
timestamp 1624857261
transform 1 0 116144 0 1 23805
box 0 0 1 1
use contact_33  contact_33_2853
timestamp 1624857261
transform 1 0 116144 0 1 24077
box 0 0 1 1
use contact_33  contact_33_2517
timestamp 1624857261
transform 1 0 119000 0 1 24213
box 0 0 1 1
use contact_33  contact_33_2522
timestamp 1624857261
transform 1 0 119000 0 1 24077
box 0 0 1 1
use contact_33  contact_33_52
timestamp 1624857261
transform 1 0 119408 0 1 24213
box 0 0 1 1
use contact_33  contact_33_57
timestamp 1624857261
transform 1 0 119272 0 1 24077
box 0 0 1 1
use contact_33  contact_33_2498
timestamp 1624857261
transform 1 0 119680 0 1 23533
box 0 0 1 1
use contact_33  contact_33_2499
timestamp 1624857261
transform 1 0 119680 0 1 24077
box 0 0 1 1
use contact_33  contact_33_37
timestamp 1624857261
transform 1 0 120632 0 1 23533
box 0 0 1 1
use contact_33  contact_33_38
timestamp 1624857261
transform 1 0 120632 0 1 24077
box 0 0 1 1
use contact_33  contact_33_39
timestamp 1624857261
transform 1 0 120632 0 1 24213
box 0 0 1 1
use contact_33  contact_33_49
timestamp 1624857261
transform 1 0 120496 0 1 23533
box 0 0 1 1
use contact_33  contact_33_50
timestamp 1624857261
transform 1 0 120496 0 1 23941
box 0 0 1 1
use contact_33  contact_33_2495
timestamp 1624857261
transform 1 0 120088 0 1 24213
box 0 0 1 1
use contact_33  contact_33_3277
timestamp 1624857261
transform 1 0 115192 0 1 24485
box 0 0 1 1
use contact_33  contact_33_3348
timestamp 1624857261
transform 1 0 115192 0 1 24621
box 0 0 1 1
use contact_33  contact_33_3349
timestamp 1624857261
transform 1 0 115192 0 1 24893
box 0 0 1 1
use contact_33  contact_33_658
timestamp 1624857261
transform 1 0 115736 0 1 24485
box 0 0 1 1
use contact_33  contact_33_659
timestamp 1624857261
transform 1 0 115600 0 1 24893
box 0 0 1 1
use contact_33  contact_33_660
timestamp 1624857261
transform 1 0 115600 0 1 24621
box 0 0 1 1
use contact_33  contact_33_2977
timestamp 1624857261
transform 1 0 116008 0 1 24485
box 0 0 1 1
use contact_33  contact_33_71
timestamp 1624857261
transform 1 0 116824 0 1 24485
box 0 0 1 1
use contact_33  contact_33_2974
timestamp 1624857261
transform 1 0 116144 0 1 24893
box 0 0 1 1
use contact_33  contact_33_2975
timestamp 1624857261
transform 1 0 116144 0 1 24621
box 0 0 1 1
use contact_33  contact_33_237
timestamp 1624857261
transform 1 0 116960 0 1 24621
box 0 0 1 1
use contact_33  contact_33_238
timestamp 1624857261
transform 1 0 116960 0 1 24893
box 0 0 1 1
use contact_33  contact_33_2516
timestamp 1624857261
transform 1 0 119000 0 1 24893
box 0 0 1 1
use contact_33  contact_33_51
timestamp 1624857261
transform 1 0 119408 0 1 24893
box 0 0 1 1
use contact_33  contact_33_40
timestamp 1624857261
transform 1 0 120632 0 1 24893
box 0 0 1 1
use contact_33  contact_33_2494
timestamp 1624857261
transform 1 0 120088 0 1 24893
box 0 0 1 1
use contact_33  contact_33_3346
timestamp 1624857261
transform 1 0 115192 0 1 25301
box 0 0 1 1
use contact_33  contact_33_3347
timestamp 1624857261
transform 1 0 115192 0 1 25029
box 0 0 1 1
use contact_33  contact_33_743
timestamp 1624857261
transform 1 0 115736 0 1 25029
box 0 0 1 1
use contact_33  contact_33_744
timestamp 1624857261
transform 1 0 115736 0 1 25301
box 0 0 1 1
use contact_33  contact_33_745
timestamp 1624857261
transform 1 0 115736 0 1 25709
box 0 0 1 1
use contact_33  contact_33_746
timestamp 1624857261
transform 1 0 115736 0 1 25437
box 0 0 1 1
use contact_33  contact_33_3092
timestamp 1624857261
transform 1 0 115328 0 1 25709
box 0 0 1 1
use contact_33  contact_33_3093
timestamp 1624857261
transform 1 0 115328 0 1 25437
box 0 0 1 1
use contact_33  contact_33_2584
timestamp 1624857261
transform 1 0 116416 0 1 25709
box 0 0 1 1
use contact_33  contact_33_2585
timestamp 1624857261
transform 1 0 116416 0 1 25437
box 0 0 1 1
use contact_33  contact_33_2594
timestamp 1624857261
transform 1 0 116552 0 1 25301
box 0 0 1 1
use contact_33  contact_33_2595
timestamp 1624857261
transform 1 0 116552 0 1 25029
box 0 0 1 1
use contact_33  contact_33_2846
timestamp 1624857261
transform 1 0 116280 0 1 25709
box 0 0 1 1
use contact_33  contact_33_2847
timestamp 1624857261
transform 1 0 116280 0 1 25437
box 0 0 1 1
use contact_33  contact_33_117
timestamp 1624857261
transform 1 0 116960 0 1 25437
box 0 0 1 1
use contact_33  contact_33_118
timestamp 1624857261
transform 1 0 116960 0 1 25709
box 0 0 1 1
use contact_33  contact_33_239
timestamp 1624857261
transform 1 0 116960 0 1 25301
box 0 0 1 1
use contact_33  contact_33_240
timestamp 1624857261
transform 1 0 116960 0 1 25029
box 0 0 1 1
use contact_33  contact_33_44
timestamp 1624857261
transform 1 0 119408 0 1 25029
box 0 0 1 1
use contact_33  contact_33_115
timestamp 1624857261
transform 1 0 119272 0 1 25029
box 0 0 1 1
use contact_33  contact_33_116
timestamp 1624857261
transform 1 0 119272 0 1 25709
box 0 0 1 1
use contact_33  contact_33_2505
timestamp 1624857261
transform 1 0 119816 0 1 25029
box 0 0 1 1
use contact_33  contact_33_3132
timestamp 1624857261
transform 1 0 115192 0 1 25845
box 0 0 1 1
use contact_33  contact_33_3133
timestamp 1624857261
transform 1 0 115192 0 1 26117
box 0 0 1 1
use contact_33  contact_33_633
timestamp 1624857261
transform 1 0 115600 0 1 26117
box 0 0 1 1
use contact_33  contact_33_634
timestamp 1624857261
transform 1 0 115600 0 1 25845
box 0 0 1 1
use contact_33  contact_33_2806
timestamp 1624857261
transform 1 0 116008 0 1 26253
box 0 0 1 1
use contact_33  contact_33_2807
timestamp 1624857261
transform 1 0 116008 0 1 26525
box 0 0 1 1
use contact_33  contact_33_223
timestamp 1624857261
transform 1 0 116824 0 1 26253
box 0 0 1 1
use contact_33  contact_33_224
timestamp 1624857261
transform 1 0 116824 0 1 26525
box 0 0 1 1
use contact_33  contact_33_119
timestamp 1624857261
transform 1 0 116960 0 1 25845
box 0 0 1 1
use contact_33  contact_33_120
timestamp 1624857261
transform 1 0 116960 0 1 26117
box 0 0 1 1
use contact_33  contact_33_43
timestamp 1624857261
transform 1 0 119408 0 1 26389
box 0 0 1 1
use contact_33  contact_33_2504
timestamp 1624857261
transform 1 0 119816 0 1 26525
box 0 0 1 1
use contact_33  contact_33_787
timestamp 1624857261
transform 1 0 115736 0 1 27341
box 0 0 1 1
use contact_33  contact_33_3321
timestamp 1624857261
transform 1 0 115328 0 1 27341
box 0 0 1 1
use contact_33  contact_33_221
timestamp 1624857261
transform 1 0 116824 0 1 26933
box 0 0 1 1
use contact_33  contact_33_222
timestamp 1624857261
transform 1 0 116824 0 1 26661
box 0 0 1 1
use contact_33  contact_33_2570
timestamp 1624857261
transform 1 0 116552 0 1 27205
box 0 0 1 1
use contact_33  contact_33_2571
timestamp 1624857261
transform 1 0 116552 0 1 26933
box 0 0 1 1
use contact_33  contact_33_2519
timestamp 1624857261
transform 1 0 119000 0 1 27341
box 0 0 1 1
use contact_33  contact_33_53
timestamp 1624857261
transform 1 0 119272 0 1 26661
box 0 0 1 1
use contact_33  contact_33_54
timestamp 1624857261
transform 1 0 119272 0 1 27205
box 0 0 1 1
use contact_33  contact_33_56
timestamp 1624857261
transform 1 0 119408 0 1 27341
box 0 0 1 1
use contact_33  contact_33_31
timestamp 1624857261
transform 1 0 120496 0 1 27205
box 0 0 1 1
use contact_33  contact_33_32
timestamp 1624857261
transform 1 0 120496 0 1 26661
box 0 0 1 1
use contact_33  contact_33_2492
timestamp 1624857261
transform 1 0 120088 0 1 27205
box 0 0 1 1
use contact_33  contact_33_2493
timestamp 1624857261
transform 1 0 120088 0 1 26661
box 0 0 1 1
use contact_33  contact_33_788
timestamp 1624857261
transform 1 0 115736 0 1 27613
box 0 0 1 1
use contact_33  contact_33_789
timestamp 1624857261
transform 1 0 115736 0 1 28021
box 0 0 1 1
use contact_33  contact_33_790
timestamp 1624857261
transform 1 0 115736 0 1 27749
box 0 0 1 1
use contact_33  contact_33_2898
timestamp 1624857261
transform 1 0 116008 0 1 28021
box 0 0 1 1
use contact_33  contact_33_2899
timestamp 1624857261
transform 1 0 116008 0 1 27749
box 0 0 1 1
use contact_33  contact_33_3058
timestamp 1624857261
transform 1 0 115328 0 1 28021
box 0 0 1 1
use contact_33  contact_33_3059
timestamp 1624857261
transform 1 0 115328 0 1 27749
box 0 0 1 1
use contact_33  contact_33_3320
timestamp 1624857261
transform 1 0 115328 0 1 27613
box 0 0 1 1
use contact_33  contact_33_2518
timestamp 1624857261
transform 1 0 119000 0 1 28021
box 0 0 1 1
use contact_33  contact_33_55
timestamp 1624857261
transform 1 0 119408 0 1 28021
box 0 0 1 1
use contact_33  contact_33_2500
timestamp 1624857261
transform 1 0 119952 0 1 27477
box 0 0 1 1
use contact_33  contact_33_2501
timestamp 1624857261
transform 1 0 119952 0 1 28021
box 0 0 1 1
use contact_33  contact_33_29
timestamp 1624857261
transform 1 0 120632 0 1 27477
box 0 0 1 1
use contact_33  contact_33_30
timestamp 1624857261
transform 1 0 120632 0 1 28021
box 0 0 1 1
use contact_33  contact_33_3208
timestamp 1624857261
transform 1 0 115328 0 1 28157
box 0 0 1 1
use contact_33  contact_33_793
timestamp 1624857261
transform 1 0 115736 0 1 28157
box 0 0 1 1
use contact_33  contact_33_3211
timestamp 1624857261
transform 1 0 115328 0 1 28565
box 0 0 1 1
use contact_33  contact_33_3209
timestamp 1624857261
transform 1 0 115328 0 1 28429
box 0 0 1 1
use contact_33  contact_33_794
timestamp 1624857261
transform 1 0 115736 0 1 28429
box 0 0 1 1
use contact_33  contact_33_792
timestamp 1624857261
transform 1 0 115736 0 1 28565
box 0 0 1 1
use contact_33  contact_33_2966
timestamp 1624857261
transform 1 0 116008 0 1 28565
box 0 0 1 1
use contact_33  contact_33_3210
timestamp 1624857261
transform 1 0 115328 0 1 28837
box 0 0 1 1
use contact_33  contact_33_791
timestamp 1624857261
transform 1 0 115736 0 1 28837
box 0 0 1 1
use contact_33  contact_33_2967
timestamp 1624857261
transform 1 0 116008 0 1 28837
box 0 0 1 1
use contact_33  contact_33_213
timestamp 1624857261
transform 1 0 116824 0 1 28565
box 0 0 1 1
use contact_33  contact_33_214
timestamp 1624857261
transform 1 0 116824 0 1 28837
box 0 0 1 1
use contact_33  contact_33_165
timestamp 1624857261
transform 1 0 116960 0 1 28429
box 0 0 1 1
use contact_33  contact_33_166
timestamp 1624857261
transform 1 0 116960 0 1 28157
box 0 0 1 1
use contact_33  contact_33_2526
timestamp 1624857261
transform 1 0 119000 0 1 28157
box 0 0 1 1
use contact_33  contact_33_2527
timestamp 1624857261
transform 1 0 119000 0 1 28837
box 0 0 1 1
use contact_33  contact_33_47
timestamp 1624857261
transform 1 0 119272 0 1 28837
box 0 0 1 1
use contact_33  contact_33_48
timestamp 1624857261
transform 1 0 119272 0 1 28157
box 0 0 1 1
use contact_33  contact_33_2502
timestamp 1624857261
transform 1 0 119952 0 1 28837
box 0 0 1 1
use contact_33  contact_33_2503
timestamp 1624857261
transform 1 0 119952 0 1 28157
box 0 0 1 1
use contact_33  contact_33_33
timestamp 1624857261
transform 1 0 120496 0 1 28157
box 0 0 1 1
use contact_33  contact_33_34
timestamp 1624857261
transform 1 0 120496 0 1 28837
box 0 0 1 1
use contact_33  contact_33_3372
timestamp 1624857261
transform 1 0 115192 0 1 28973
box 0 0 1 1
use contact_33  contact_33_3373
timestamp 1624857261
transform 1 0 115192 0 1 29245
box 0 0 1 1
use contact_33  contact_33_3374
timestamp 1624857261
transform 1 0 115192 0 1 29653
box 0 0 1 1
use contact_33  contact_33_3375
timestamp 1624857261
transform 1 0 115192 0 1 29381
box 0 0 1 1
use contact_33  contact_33_797
timestamp 1624857261
transform 1 0 115600 0 1 28973
box 0 0 1 1
use contact_33  contact_33_798
timestamp 1624857261
transform 1 0 115600 0 1 29245
box 0 0 1 1
use contact_33  contact_33_799
timestamp 1624857261
transform 1 0 115600 0 1 29653
box 0 0 1 1
use contact_33  contact_33_800
timestamp 1624857261
transform 1 0 115600 0 1 29381
box 0 0 1 1
use contact_33  contact_33_2710
timestamp 1624857261
transform 1 0 116008 0 1 29381
box 0 0 1 1
use contact_33  contact_33_2711
timestamp 1624857261
transform 1 0 116008 0 1 29653
box 0 0 1 1
use contact_33  contact_33_2964
timestamp 1624857261
transform 1 0 116144 0 1 29245
box 0 0 1 1
use contact_33  contact_33_2965
timestamp 1624857261
transform 1 0 116144 0 1 28973
box 0 0 1 1
use contact_33  contact_33_105
timestamp 1624857261
transform 1 0 116960 0 1 29653
box 0 0 1 1
use contact_33  contact_33_106
timestamp 1624857261
transform 1 0 116960 0 1 29381
box 0 0 1 1
use contact_33  contact_33_215
timestamp 1624857261
transform 1 0 116960 0 1 29245
box 0 0 1 1
use contact_33  contact_33_216
timestamp 1624857261
transform 1 0 116960 0 1 28973
box 0 0 1 1
use contact_33  contact_33_757
timestamp 1624857261
transform 1 0 115736 0 1 30061
box 0 0 1 1
use contact_33  contact_33_758
timestamp 1624857261
transform 1 0 115736 0 1 29789
box 0 0 1 1
use contact_33  contact_33_3306
timestamp 1624857261
transform 1 0 115328 0 1 30061
box 0 0 1 1
use contact_33  contact_33_3307
timestamp 1624857261
transform 1 0 115328 0 1 29789
box 0 0 1 1
use contact_33  contact_33_2698
timestamp 1624857261
transform 1 0 116280 0 1 30197
box 0 0 1 1
use contact_33  contact_33_2699
timestamp 1624857261
transform 1 0 116280 0 1 30469
box 0 0 1 1
use contact_33  contact_33_341
timestamp 1624857261
transform 1 0 116960 0 1 29789
box 0 0 1 1
use contact_33  contact_33_342
timestamp 1624857261
transform 1 0 116960 0 1 30061
box 0 0 1 1
use contact_33  contact_33_343
timestamp 1624857261
transform 1 0 116960 0 1 30469
box 0 0 1 1
use contact_33  contact_33_344
timestamp 1624857261
transform 1 0 116960 0 1 30197
box 0 0 1 1
use contact_33  contact_33_3029
timestamp 1624857261
transform 1 0 115192 0 1 31285
box 0 0 1 1
use contact_33  contact_33_523
timestamp 1624857261
transform 1 0 115600 0 1 31285
box 0 0 1 1
use contact_33  contact_33_2928
timestamp 1624857261
transform 1 0 116008 0 1 31149
box 0 0 1 1
use contact_33  contact_33_2929
timestamp 1624857261
transform 1 0 116008 0 1 30877
box 0 0 1 1
use contact_33  contact_33_367
timestamp 1624857261
transform 1 0 116824 0 1 30605
box 0 0 1 1
use contact_33  contact_33_368
timestamp 1624857261
transform 1 0 116824 0 1 30877
box 0 0 1 1
use contact_33  contact_33_3028
timestamp 1624857261
transform 1 0 115192 0 1 31557
box 0 0 1 1
use contact_33  contact_33_521
timestamp 1624857261
transform 1 0 115736 0 1 31965
box 0 0 1 1
use contact_33  contact_33_522
timestamp 1624857261
transform 1 0 115736 0 1 31693
box 0 0 1 1
use contact_33  contact_33_524
timestamp 1624857261
transform 1 0 115600 0 1 31557
box 0 0 1 1
use contact_33  contact_33_3020
timestamp 1624857261
transform 1 0 115328 0 1 31965
box 0 0 1 1
use contact_33  contact_33_3021
timestamp 1624857261
transform 1 0 115328 0 1 31693
box 0 0 1 1
use contact_33  contact_33_423
timestamp 1624857261
transform 1 0 116824 0 1 31421
box 0 0 1 1
use contact_33  contact_33_424
timestamp 1624857261
transform 1 0 116824 0 1 31693
box 0 0 1 1
use contact_33  contact_33_2694
timestamp 1624857261
transform 1 0 116416 0 1 31693
box 0 0 1 1
use contact_33  contact_33_2695
timestamp 1624857261
transform 1 0 116144 0 1 31693
box 0 0 1 1
use contact_33  contact_33_2696
timestamp 1624857261
transform 1 0 116416 0 1 31421
box 0 0 1 1
use contact_33  contact_33_2697
timestamp 1624857261
transform 1 0 116280 0 1 31693
box 0 0 1 1
use contact_33  contact_33_3174
timestamp 1624857261
transform 1 0 115192 0 1 32101
box 0 0 1 1
use contact_33  contact_33_3175
timestamp 1624857261
transform 1 0 115192 0 1 32373
box 0 0 1 1
use contact_33  contact_33_805
timestamp 1624857261
transform 1 0 115600 0 1 32101
box 0 0 1 1
use contact_33  contact_33_3001
timestamp 1624857261
transform 1 0 116008 0 1 32101
box 0 0 1 1
use contact_33  contact_33_3218
timestamp 1624857261
transform 1 0 115328 0 1 32509
box 0 0 1 1
use contact_33  contact_33_808
timestamp 1624857261
transform 1 0 115600 0 1 32509
box 0 0 1 1
use contact_33  contact_33_806
timestamp 1624857261
transform 1 0 115600 0 1 32373
box 0 0 1 1
use contact_33  contact_33_3000
timestamp 1624857261
transform 1 0 116008 0 1 32373
box 0 0 1 1
use contact_33  contact_33_2857
timestamp 1624857261
transform 1 0 116008 0 1 32509
box 0 0 1 1
use contact_33  contact_33_3219
timestamp 1624857261
transform 1 0 115328 0 1 32781
box 0 0 1 1
use contact_33  contact_33_807
timestamp 1624857261
transform 1 0 115600 0 1 32781
box 0 0 1 1
use contact_33  contact_33_2856
timestamp 1624857261
transform 1 0 116008 0 1 32781
box 0 0 1 1
use contact_33  contact_33_153
timestamp 1624857261
transform 1 0 116824 0 1 32509
box 0 0 1 1
use contact_33  contact_33_154
timestamp 1624857261
transform 1 0 116824 0 1 32781
box 0 0 1 1
use contact_33  contact_33_2792
timestamp 1624857261
transform 1 0 116280 0 1 32509
box 0 0 1 1
use contact_33  contact_33_2793
timestamp 1624857261
transform 1 0 116280 0 1 32781
box 0 0 1 1
use contact_33  contact_33_2854
timestamp 1624857261
transform 1 0 116280 0 1 32101
box 0 0 1 1
use contact_33  contact_33_2855
timestamp 1624857261
transform 1 0 116280 0 1 32373
box 0 0 1 1
use contact_33  contact_33_143
timestamp 1624857261
transform 1 0 116960 0 1 32101
box 0 0 1 1
use contact_33  contact_33_144
timestamp 1624857261
transform 1 0 116960 0 1 32373
box 0 0 1 1
use contact_33  contact_33_3054
timestamp 1624857261
transform 1 0 115192 0 1 33597
box 0 0 1 1
use contact_33  contact_33_3055
timestamp 1624857261
transform 1 0 115192 0 1 33325
box 0 0 1 1
use contact_33  contact_33_597
timestamp 1624857261
transform 1 0 115600 0 1 33597
box 0 0 1 1
use contact_33  contact_33_598
timestamp 1624857261
transform 1 0 115600 0 1 33325
box 0 0 1 1
use contact_33  contact_33_599
timestamp 1624857261
transform 1 0 115736 0 1 32917
box 0 0 1 1
use contact_33  contact_33_600
timestamp 1624857261
transform 1 0 115736 0 1 33189
box 0 0 1 1
use contact_33  contact_33_3216
timestamp 1624857261
transform 1 0 115328 0 1 33189
box 0 0 1 1
use contact_33  contact_33_3217
timestamp 1624857261
transform 1 0 115328 0 1 32917
box 0 0 1 1
use contact_33  contact_33_177
timestamp 1624857261
transform 1 0 116824 0 1 32917
box 0 0 1 1
use contact_33  contact_33_178
timestamp 1624857261
transform 1 0 116824 0 1 33189
box 0 0 1 1
use contact_33  contact_33_2580
timestamp 1624857261
transform 1 0 116416 0 1 32917
box 0 0 1 1
use contact_33  contact_33_2581
timestamp 1624857261
transform 1 0 116416 0 1 33189
box 0 0 1 1
use contact_33  contact_33_2752
timestamp 1624857261
transform 1 0 116144 0 1 33597
box 0 0 1 1
use contact_33  contact_33_2753
timestamp 1624857261
transform 1 0 116144 0 1 33325
box 0 0 1 1
use contact_33  contact_33_2794
timestamp 1624857261
transform 1 0 116144 0 1 33189
box 0 0 1 1
use contact_33  contact_33_2795
timestamp 1624857261
transform 1 0 116144 0 1 32917
box 0 0 1 1
use contact_33  contact_33_175
timestamp 1624857261
transform 1 0 116960 0 1 33597
box 0 0 1 1
use contact_33  contact_33_176
timestamp 1624857261
transform 1 0 116960 0 1 33325
box 0 0 1 1
use contact_33  contact_33_3264
timestamp 1624857261
transform 1 0 115328 0 1 33733
box 0 0 1 1
use contact_33  contact_33_466
timestamp 1624857261
transform 1 0 115600 0 1 33733
box 0 0 1 1
use contact_33  contact_33_3265
timestamp 1624857261
transform 1 0 115328 0 1 34005
box 0 0 1 1
use contact_33  contact_33_465
timestamp 1624857261
transform 1 0 115600 0 1 34005
box 0 0 1 1
use contact_33  contact_33_3267
timestamp 1624857261
transform 1 0 115328 0 1 34141
box 0 0 1 1
use contact_33  contact_33_519
timestamp 1624857261
transform 1 0 115600 0 1 34141
box 0 0 1 1
use contact_33  contact_33_3015
timestamp 1624857261
transform 1 0 116008 0 1 34141
box 0 0 1 1
use contact_33  contact_33_3266
timestamp 1624857261
transform 1 0 115328 0 1 34413
box 0 0 1 1
use contact_33  contact_33_520
timestamp 1624857261
transform 1 0 115600 0 1 34413
box 0 0 1 1
use contact_33  contact_33_3014
timestamp 1624857261
transform 1 0 116008 0 1 34413
box 0 0 1 1
use contact_33  contact_33_99
timestamp 1624857261
transform 1 0 116824 0 1 33733
box 0 0 1 1
use contact_33  contact_33_100
timestamp 1624857261
transform 1 0 116824 0 1 34005
box 0 0 1 1
use contact_33  contact_33_2626
timestamp 1624857261
transform 1 0 116552 0 1 34005
box 0 0 1 1
use contact_33  contact_33_2627
timestamp 1624857261
transform 1 0 116552 0 1 33733
box 0 0 1 1
use contact_33  contact_33_2712
timestamp 1624857261
transform 1 0 116280 0 1 34005
box 0 0 1 1
use contact_33  contact_33_2713
timestamp 1624857261
transform 1 0 116280 0 1 33733
box 0 0 1 1
use contact_33  contact_33_147
timestamp 1624857261
transform 1 0 116960 0 1 34141
box 0 0 1 1
use contact_33  contact_33_148
timestamp 1624857261
transform 1 0 116960 0 1 34413
box 0 0 1 1
use contact_33  contact_33_66
timestamp 1624857261
transform 1 0 116824 0 1 34957
box 0 0 1 1
use contact_33  contact_33_2647
timestamp 1624857261
transform 1 0 116552 0 1 34821
box 0 0 1 1
use contact_33  contact_33_145
timestamp 1624857261
transform 1 0 116960 0 1 34821
box 0 0 1 1
use contact_33  contact_33_146
timestamp 1624857261
transform 1 0 116960 0 1 34549
box 0 0 1 1
use contact_33  contact_33_635
timestamp 1624857261
transform 1 0 115600 0 1 35909
box 0 0 1 1
use contact_33  contact_33_636
timestamp 1624857261
transform 1 0 115600 0 1 35637
box 0 0 1 1
use contact_33  contact_33_3094
timestamp 1624857261
transform 1 0 115328 0 1 35637
box 0 0 1 1
use contact_33  contact_33_3095
timestamp 1624857261
transform 1 0 115328 0 1 35909
box 0 0 1 1
use contact_33  contact_33_65
timestamp 1624857261
transform 1 0 116824 0 1 35229
box 0 0 1 1
use contact_33  contact_33_2540
timestamp 1624857261
transform 1 0 116552 0 1 35637
box 0 0 1 1
use contact_33  contact_33_2541
timestamp 1624857261
transform 1 0 116552 0 1 35909
box 0 0 1 1
use contact_33  contact_33_2646
timestamp 1624857261
transform 1 0 116552 0 1 35229
box 0 0 1 1
use contact_33  contact_33_2766
timestamp 1624857261
transform 1 0 116280 0 1 35365
box 0 0 1 1
use contact_33  contact_33_2767
timestamp 1624857261
transform 1 0 116280 0 1 35637
box 0 0 1 1
use contact_33  contact_33_111
timestamp 1624857261
transform 1 0 116960 0 1 35365
box 0 0 1 1
use contact_33  contact_33_112
timestamp 1624857261
transform 1 0 116960 0 1 35637
box 0 0 1 1
use contact_33  contact_33_3274
timestamp 1624857261
transform 1 0 115192 0 1 36453
box 0 0 1 1
use contact_33  contact_33_3275
timestamp 1624857261
transform 1 0 115192 0 1 36725
box 0 0 1 1
use contact_33  contact_33_505
timestamp 1624857261
transform 1 0 115736 0 1 36045
box 0 0 1 1
use contact_33  contact_33_506
timestamp 1624857261
transform 1 0 115736 0 1 36317
box 0 0 1 1
use contact_33  contact_33_573
timestamp 1624857261
transform 1 0 115600 0 1 36453
box 0 0 1 1
use contact_33  contact_33_574
timestamp 1624857261
transform 1 0 115600 0 1 36725
box 0 0 1 1
use contact_33  contact_33_2804
timestamp 1624857261
transform 1 0 116008 0 1 36453
box 0 0 1 1
use contact_33  contact_33_2805
timestamp 1624857261
transform 1 0 116008 0 1 36725
box 0 0 1 1
use contact_33  contact_33_3096
timestamp 1624857261
transform 1 0 115328 0 1 36317
box 0 0 1 1
use contact_33  contact_33_3097
timestamp 1624857261
transform 1 0 115328 0 1 36045
box 0 0 1 1
use contact_33  contact_33_2732
timestamp 1624857261
transform 1 0 116280 0 1 36317
box 0 0 1 1
use contact_33  contact_33_2733
timestamp 1624857261
transform 1 0 116280 0 1 36045
box 0 0 1 1
use contact_33  contact_33_2802
timestamp 1624857261
transform 1 0 116280 0 1 36453
box 0 0 1 1
use contact_33  contact_33_2803
timestamp 1624857261
transform 1 0 116280 0 1 36725
box 0 0 1 1
use contact_33  contact_33_393
timestamp 1624857261
transform 1 0 116960 0 1 36317
box 0 0 1 1
use contact_33  contact_33_394
timestamp 1624857261
transform 1 0 116960 0 1 36045
box 0 0 1 1
use contact_33  contact_33_575
timestamp 1624857261
transform 1 0 115600 0 1 37133
box 0 0 1 1
use contact_33  contact_33_576
timestamp 1624857261
transform 1 0 115600 0 1 36861
box 0 0 1 1
use contact_33  contact_33_3370
timestamp 1624857261
transform 1 0 115328 0 1 36861
box 0 0 1 1
use contact_33  contact_33_3371
timestamp 1624857261
transform 1 0 115328 0 1 37133
box 0 0 1 1
use contact_33  contact_33_369
timestamp 1624857261
transform 1 0 116824 0 1 36861
box 0 0 1 1
use contact_33  contact_33_370
timestamp 1624857261
transform 1 0 116824 0 1 37133
box 0 0 1 1
use contact_33  contact_33_2614
timestamp 1624857261
transform 1 0 116552 0 1 37133
box 0 0 1 1
use contact_33  contact_33_2615
timestamp 1624857261
transform 1 0 116552 0 1 36861
box 0 0 1 1
use contact_33  contact_33_2958
timestamp 1624857261
transform 1 0 116280 0 1 36861
box 0 0 1 1
use contact_33  contact_33_2959
timestamp 1624857261
transform 1 0 116280 0 1 37133
box 0 0 1 1
use contact_33  contact_33_2962
timestamp 1624857261
transform 1 0 116144 0 1 36861
box 0 0 1 1
use contact_33  contact_33_2963
timestamp 1624857261
transform 1 0 116144 0 1 37133
box 0 0 1 1
use contact_33  contact_33_841
timestamp 1624857261
transform 1 0 110432 0 1 39037
box 0 0 1 1
use contact_33  contact_33_842
timestamp 1624857261
transform 1 0 110432 0 1 39309
box 0 0 1 1
use contact_33  contact_33_885
timestamp 1624857261
transform 1 0 110160 0 1 38357
box 0 0 1 1
use contact_33  contact_33_886
timestamp 1624857261
transform 1 0 110160 0 1 38629
box 0 0 1 1
use contact_33  contact_33_927
timestamp 1624857261
transform 1 0 110432 0 1 42029
box 0 0 1 1
use contact_33  contact_33_928
timestamp 1624857261
transform 1 0 110432 0 1 41757
box 0 0 1 1
use contact_33  contact_33_933
timestamp 1624857261
transform 1 0 110160 0 1 40261
box 0 0 1 1
use contact_33  contact_33_934
timestamp 1624857261
transform 1 0 110160 0 1 40533
box 0 0 1 1
use contact_33  contact_33_865
timestamp 1624857261
transform 1 0 110432 0 1 43661
box 0 0 1 1
use contact_33  contact_33_866
timestamp 1624857261
transform 1 0 110432 0 1 43389
box 0 0 1 1
use contact_33  contact_33_917
timestamp 1624857261
transform 1 0 110160 0 1 43253
box 0 0 1 1
use contact_33  contact_33_918
timestamp 1624857261
transform 1 0 110160 0 1 42981
box 0 0 1 1
use contact_33  contact_33_929
timestamp 1624857261
transform 1 0 110160 0 1 44205
box 0 0 1 1
use contact_33  contact_33_930
timestamp 1624857261
transform 1 0 110160 0 1 44477
box 0 0 1 1
use contact_33  contact_33_843
timestamp 1624857261
transform 1 0 110296 0 1 46925
box 0 0 1 1
use contact_33  contact_33_844
timestamp 1624857261
transform 1 0 110296 0 1 47197
box 0 0 1 1
use contact_33  contact_33_845
timestamp 1624857261
transform 1 0 110160 0 1 47605
box 0 0 1 1
use contact_33  contact_33_846
timestamp 1624857261
transform 1 0 110160 0 1 47333
box 0 0 1 1
use contact_33  contact_33_951
timestamp 1624857261
transform 1 0 110432 0 1 46789
box 0 0 1 1
use contact_33  contact_33_952
timestamp 1624857261
transform 1 0 110432 0 1 46517
box 0 0 1 1
use contact_33  contact_33_897
timestamp 1624857261
transform 1 0 110432 0 1 50733
box 0 0 1 1
use contact_33  contact_33_898
timestamp 1624857261
transform 1 0 110432 0 1 50461
box 0 0 1 1
use contact_33  contact_33_921
timestamp 1624857261
transform 1 0 110432 0 1 52093
box 0 0 1 1
use contact_33  contact_33_922
timestamp 1624857261
transform 1 0 110432 0 1 52365
box 0 0 1 1
use contact_33  contact_33_836
timestamp 1624857261
transform 1 0 110432 0 1 55629
box 0 0 1 1
use contact_33  contact_33_867
timestamp 1624857261
transform 1 0 110432 0 1 55493
box 0 0 1 1
use contact_33  contact_33_868
timestamp 1624857261
transform 1 0 110432 0 1 55221
box 0 0 1 1
use contact_33  contact_33_3130
timestamp 1624857261
transform 1 0 115192 0 1 37949
box 0 0 1 1
use contact_33  contact_33_3131
timestamp 1624857261
transform 1 0 115192 0 1 37677
box 0 0 1 1
use contact_33  contact_33_3368
timestamp 1624857261
transform 1 0 115328 0 1 37541
box 0 0 1 1
use contact_33  contact_33_3369
timestamp 1624857261
transform 1 0 115328 0 1 37269
box 0 0 1 1
use contact_33  contact_33_481
timestamp 1624857261
transform 1 0 115600 0 1 37949
box 0 0 1 1
use contact_33  contact_33_482
timestamp 1624857261
transform 1 0 115600 0 1 37677
box 0 0 1 1
use contact_33  contact_33_529
timestamp 1624857261
transform 1 0 115736 0 1 37541
box 0 0 1 1
use contact_33  contact_33_530
timestamp 1624857261
transform 1 0 115736 0 1 37269
box 0 0 1 1
use contact_33  contact_33_2780
timestamp 1624857261
transform 1 0 116008 0 1 37677
box 0 0 1 1
use contact_33  contact_33_2781
timestamp 1624857261
transform 1 0 116008 0 1 37949
box 0 0 1 1
use contact_33  contact_33_2960
timestamp 1624857261
transform 1 0 116144 0 1 37541
box 0 0 1 1
use contact_33  contact_33_2961
timestamp 1624857261
transform 1 0 116144 0 1 37269
box 0 0 1 1
use contact_33  contact_33_259
timestamp 1624857261
transform 1 0 116960 0 1 37677
box 0 0 1 1
use contact_33  contact_33_260
timestamp 1624857261
transform 1 0 116960 0 1 37949
box 0 0 1 1
use contact_33  contact_33_371
timestamp 1624857261
transform 1 0 116824 0 1 37541
box 0 0 1 1
use contact_33  contact_33_372
timestamp 1624857261
transform 1 0 116824 0 1 37269
box 0 0 1 1
use contact_33  contact_33_2956
timestamp 1624857261
transform 1 0 116280 0 1 37541
box 0 0 1 1
use contact_33  contact_33_2957
timestamp 1624857261
transform 1 0 116280 0 1 37269
box 0 0 1 1
use contact_33  contact_33_3182
timestamp 1624857261
transform 1 0 115328 0 1 38085
box 0 0 1 1
use contact_33  contact_33_3183
timestamp 1624857261
transform 1 0 115328 0 1 38357
box 0 0 1 1
use contact_33  contact_33_717
timestamp 1624857261
transform 1 0 115736 0 1 38085
box 0 0 1 1
use contact_33  contact_33_718
timestamp 1624857261
transform 1 0 115736 0 1 38357
box 0 0 1 1
use contact_33  contact_33_2916
timestamp 1624857261
transform 1 0 116008 0 1 38085
box 0 0 1 1
use contact_33  contact_33_2917
timestamp 1624857261
transform 1 0 116008 0 1 38357
box 0 0 1 1
use contact_33  contact_33_293
timestamp 1624857261
transform 1 0 116824 0 1 38085
box 0 0 1 1
use contact_33  contact_33_294
timestamp 1624857261
transform 1 0 116824 0 1 38357
box 0 0 1 1
use contact_33  contact_33_323
timestamp 1624857261
transform 1 0 116960 0 1 38493
box 0 0 1 1
use contact_33  contact_33_324
timestamp 1624857261
transform 1 0 116960 0 1 38765
box 0 0 1 1
use contact_33  contact_33_3060
timestamp 1624857261
transform 1 0 115192 0 1 39581
box 0 0 1 1
use contact_33  contact_33_533
timestamp 1624857261
transform 1 0 115600 0 1 39581
box 0 0 1 1
use contact_33  contact_33_205
timestamp 1624857261
transform 1 0 116824 0 1 39581
box 0 0 1 1
use contact_33  contact_33_206
timestamp 1624857261
transform 1 0 116824 0 1 39309
box 0 0 1 1
use contact_33  contact_33_321
timestamp 1624857261
transform 1 0 116960 0 1 39173
box 0 0 1 1
use contact_33  contact_33_322
timestamp 1624857261
transform 1 0 116960 0 1 38901
box 0 0 1 1
use contact_33  contact_33_2578
timestamp 1624857261
transform 1 0 116552 0 1 38901
box 0 0 1 1
use contact_33  contact_33_2579
timestamp 1624857261
transform 1 0 116552 0 1 39173
box 0 0 1 1
use contact_33  contact_33_2611
timestamp 1624857261
transform 1 0 116416 0 1 39581
box 0 0 1 1
use contact_33  contact_33_3061
timestamp 1624857261
transform 1 0 115192 0 1 39853
box 0 0 1 1
use contact_33  contact_33_3171
timestamp 1624857261
transform 1 0 115192 0 1 40397
box 0 0 1 1
use contact_33  contact_33_3172
timestamp 1624857261
transform 1 0 115192 0 1 39989
box 0 0 1 1
use contact_33  contact_33_3173
timestamp 1624857261
transform 1 0 115192 0 1 40261
box 0 0 1 1
use contact_33  contact_33_531
timestamp 1624857261
transform 1 0 115600 0 1 40261
box 0 0 1 1
use contact_33  contact_33_532
timestamp 1624857261
transform 1 0 115600 0 1 39989
box 0 0 1 1
use contact_33  contact_33_534
timestamp 1624857261
transform 1 0 115600 0 1 39853
box 0 0 1 1
use contact_33  contact_33_759
timestamp 1624857261
transform 1 0 115736 0 1 40397
box 0 0 1 1
use contact_33  contact_33_2876
timestamp 1624857261
transform 1 0 116008 0 1 40397
box 0 0 1 1
use contact_33  contact_33_2610
timestamp 1624857261
transform 1 0 116416 0 1 39853
box 0 0 1 1
use contact_33  contact_33_3170
timestamp 1624857261
transform 1 0 115192 0 1 40669
box 0 0 1 1
use contact_33  contact_33_3242
timestamp 1624857261
transform 1 0 115192 0 1 40805
box 0 0 1 1
use contact_33  contact_33_3243
timestamp 1624857261
transform 1 0 115192 0 1 41077
box 0 0 1 1
use contact_33  contact_33_3245
timestamp 1624857261
transform 1 0 115192 0 1 41213
box 0 0 1 1
use contact_33  contact_33_514
timestamp 1624857261
transform 1 0 115600 0 1 41213
box 0 0 1 1
use contact_33  contact_33_760
timestamp 1624857261
transform 1 0 115736 0 1 40669
box 0 0 1 1
use contact_33  contact_33_761
timestamp 1624857261
transform 1 0 115736 0 1 41077
box 0 0 1 1
use contact_33  contact_33_762
timestamp 1624857261
transform 1 0 115736 0 1 40805
box 0 0 1 1
use contact_33  contact_33_2737
timestamp 1624857261
transform 1 0 116008 0 1 41213
box 0 0 1 1
use contact_33  contact_33_2874
timestamp 1624857261
transform 1 0 116008 0 1 41077
box 0 0 1 1
use contact_33  contact_33_2875
timestamp 1624857261
transform 1 0 116008 0 1 40805
box 0 0 1 1
use contact_33  contact_33_2877
timestamp 1624857261
transform 1 0 116008 0 1 40669
box 0 0 1 1
use contact_33  contact_33_360
timestamp 1624857261
transform 1 0 116960 0 1 41213
box 0 0 1 1
use contact_33  contact_33_361
timestamp 1624857261
transform 1 0 116960 0 1 40805
box 0 0 1 1
use contact_33  contact_33_362
timestamp 1624857261
transform 1 0 116960 0 1 41077
box 0 0 1 1
use contact_33  contact_33_2621
timestamp 1624857261
transform 1 0 116552 0 1 41213
box 0 0 1 1
use contact_33  contact_33_2735
timestamp 1624857261
transform 1 0 116280 0 1 41213
box 0 0 1 1
use contact_33  contact_33_3069
timestamp 1624857261
transform 1 0 115192 0 1 42029
box 0 0 1 1
use contact_33  contact_33_3128
timestamp 1624857261
transform 1 0 115328 0 1 41893
box 0 0 1 1
use contact_33  contact_33_3129
timestamp 1624857261
transform 1 0 115328 0 1 41621
box 0 0 1 1
use contact_33  contact_33_3244
timestamp 1624857261
transform 1 0 115192 0 1 41485
box 0 0 1 1
use contact_33  contact_33_513
timestamp 1624857261
transform 1 0 115600 0 1 41485
box 0 0 1 1
use contact_33  contact_33_611
timestamp 1624857261
transform 1 0 115736 0 1 41621
box 0 0 1 1
use contact_33  contact_33_612
timestamp 1624857261
transform 1 0 115736 0 1 41893
box 0 0 1 1
use contact_33  contact_33_783
timestamp 1624857261
transform 1 0 115600 0 1 42029
box 0 0 1 1
use contact_33  contact_33_2736
timestamp 1624857261
transform 1 0 116008 0 1 41485
box 0 0 1 1
use contact_33  contact_33_2796
timestamp 1624857261
transform 1 0 116008 0 1 41621
box 0 0 1 1
use contact_33  contact_33_2797
timestamp 1624857261
transform 1 0 116008 0 1 41893
box 0 0 1 1
use contact_33  contact_33_2799
timestamp 1624857261
transform 1 0 116144 0 1 42029
box 0 0 1 1
use contact_33  contact_33_255
timestamp 1624857261
transform 1 0 116824 0 1 41893
box 0 0 1 1
use contact_33  contact_33_256
timestamp 1624857261
transform 1 0 116824 0 1 41621
box 0 0 1 1
use contact_33  contact_33_313
timestamp 1624857261
transform 1 0 116960 0 1 42029
box 0 0 1 1
use contact_33  contact_33_359
timestamp 1624857261
transform 1 0 116960 0 1 41485
box 0 0 1 1
use contact_33  contact_33_2576
timestamp 1624857261
transform 1 0 116416 0 1 41621
box 0 0 1 1
use contact_33  contact_33_2577
timestamp 1624857261
transform 1 0 116416 0 1 41893
box 0 0 1 1
use contact_33  contact_33_2620
timestamp 1624857261
transform 1 0 116552 0 1 41485
box 0 0 1 1
use contact_33  contact_33_2734
timestamp 1624857261
transform 1 0 116280 0 1 41485
box 0 0 1 1
use contact_33  contact_33_3068
timestamp 1624857261
transform 1 0 115192 0 1 42301
box 0 0 1 1
use contact_33  contact_33_3192
timestamp 1624857261
transform 1 0 115328 0 1 42437
box 0 0 1 1
use contact_33  contact_33_3193
timestamp 1624857261
transform 1 0 115328 0 1 42709
box 0 0 1 1
use contact_33  contact_33_784
timestamp 1624857261
transform 1 0 115600 0 1 42301
box 0 0 1 1
use contact_33  contact_33_785
timestamp 1624857261
transform 1 0 115600 0 1 42709
box 0 0 1 1
use contact_33  contact_33_786
timestamp 1624857261
transform 1 0 115600 0 1 42437
box 0 0 1 1
use contact_33  contact_33_2798
timestamp 1624857261
transform 1 0 116144 0 1 42301
box 0 0 1 1
use contact_33  contact_33_295
timestamp 1624857261
transform 1 0 116960 0 1 42845
box 0 0 1 1
use contact_33  contact_33_311
timestamp 1624857261
transform 1 0 116960 0 1 42709
box 0 0 1 1
use contact_33  contact_33_312
timestamp 1624857261
transform 1 0 116960 0 1 42437
box 0 0 1 1
use contact_33  contact_33_314
timestamp 1624857261
transform 1 0 116960 0 1 42301
box 0 0 1 1
use contact_33  contact_33_3120
timestamp 1624857261
transform 1 0 115192 0 1 43797
box 0 0 1 1
use contact_33  contact_33_3121
timestamp 1624857261
transform 1 0 115192 0 1 43525
box 0 0 1 1
use contact_33  contact_33_455
timestamp 1624857261
transform 1 0 115600 0 1 43797
box 0 0 1 1
use contact_33  contact_33_456
timestamp 1624857261
transform 1 0 115600 0 1 43525
box 0 0 1 1
use contact_33  contact_33_2888
timestamp 1624857261
transform 1 0 116008 0 1 43797
box 0 0 1 1
use contact_33  contact_33_2889
timestamp 1624857261
transform 1 0 116008 0 1 43525
box 0 0 1 1
use contact_33  contact_33_296
timestamp 1624857261
transform 1 0 116960 0 1 43117
box 0 0 1 1
use contact_33  contact_33_297
timestamp 1624857261
transform 1 0 116960 0 1 43525
box 0 0 1 1
use contact_33  contact_33_298
timestamp 1624857261
transform 1 0 116960 0 1 43253
box 0 0 1 1
use contact_33  contact_33_2596
timestamp 1624857261
transform 1 0 116552 0 1 43797
box 0 0 1 1
use contact_33  contact_33_2597
timestamp 1624857261
transform 1 0 116552 0 1 43525
box 0 0 1 1
use contact_33  contact_33_3184
timestamp 1624857261
transform 1 0 115192 0 1 43933
box 0 0 1 1
use contact_33  contact_33_3185
timestamp 1624857261
transform 1 0 115192 0 1 44205
box 0 0 1 1
use contact_33  contact_33_3186
timestamp 1624857261
transform 1 0 115192 0 1 44613
box 0 0 1 1
use contact_33  contact_33_3187
timestamp 1624857261
transform 1 0 115192 0 1 44341
box 0 0 1 1
use contact_33  contact_33_451
timestamp 1624857261
transform 1 0 115600 0 1 43933
box 0 0 1 1
use contact_33  contact_33_452
timestamp 1624857261
transform 1 0 115600 0 1 44205
box 0 0 1 1
use contact_33  contact_33_453
timestamp 1624857261
transform 1 0 115600 0 1 44613
box 0 0 1 1
use contact_33  contact_33_454
timestamp 1624857261
transform 1 0 115600 0 1 44341
box 0 0 1 1
use contact_33  contact_33_2542
timestamp 1624857261
transform 1 0 116552 0 1 44613
box 0 0 1 1
use contact_33  contact_33_2543
timestamp 1624857261
transform 1 0 116552 0 1 44341
box 0 0 1 1
use contact_33  contact_33_2882
timestamp 1624857261
transform 1 0 116280 0 1 44069
box 0 0 1 1
use contact_33  contact_33_2883
timestamp 1624857261
transform 1 0 116280 0 1 44341
box 0 0 1 1
use contact_33  contact_33_3252
timestamp 1624857261
transform 1 0 115328 0 1 44749
box 0 0 1 1
use contact_33  contact_33_3253
timestamp 1624857261
transform 1 0 115328 0 1 45021
box 0 0 1 1
use contact_33  contact_33_3254
timestamp 1624857261
transform 1 0 115328 0 1 45429
box 0 0 1 1
use contact_33  contact_33_3255
timestamp 1624857261
transform 1 0 115328 0 1 45157
box 0 0 1 1
use contact_33  contact_33_495
timestamp 1624857261
transform 1 0 115736 0 1 44749
box 0 0 1 1
use contact_33  contact_33_496
timestamp 1624857261
transform 1 0 115736 0 1 45021
box 0 0 1 1
use contact_33  contact_33_497
timestamp 1624857261
transform 1 0 115736 0 1 45429
box 0 0 1 1
use contact_33  contact_33_498
timestamp 1624857261
transform 1 0 115736 0 1 45157
box 0 0 1 1
use contact_33  contact_33_3012
timestamp 1624857261
transform 1 0 116144 0 1 45157
box 0 0 1 1
use contact_33  contact_33_3013
timestamp 1624857261
transform 1 0 116144 0 1 45429
box 0 0 1 1
use contact_33  contact_33_123
timestamp 1624857261
transform 1 0 116960 0 1 45157
box 0 0 1 1
use contact_33  contact_33_124
timestamp 1624857261
transform 1 0 116960 0 1 45429
box 0 0 1 1
use contact_33  contact_33_199
timestamp 1624857261
transform 1 0 116824 0 1 45021
box 0 0 1 1
use contact_33  contact_33_200
timestamp 1624857261
transform 1 0 116824 0 1 44749
box 0 0 1 1
use contact_33  contact_33_2592
timestamp 1624857261
transform 1 0 116416 0 1 44749
box 0 0 1 1
use contact_33  contact_33_2593
timestamp 1624857261
transform 1 0 116416 0 1 45021
box 0 0 1 1
use contact_33  contact_33_3010
timestamp 1624857261
transform 1 0 116280 0 1 45157
box 0 0 1 1
use contact_33  contact_33_3011
timestamp 1624857261
transform 1 0 116280 0 1 45429
box 0 0 1 1
use contact_33  contact_33_3050
timestamp 1624857261
transform 1 0 115328 0 1 46245
box 0 0 1 1
use contact_33  contact_33_3051
timestamp 1624857261
transform 1 0 115328 0 1 45973
box 0 0 1 1
use contact_33  contact_33_3086
timestamp 1624857261
transform 1 0 115192 0 1 45837
box 0 0 1 1
use contact_33  contact_33_3087
timestamp 1624857261
transform 1 0 115192 0 1 45565
box 0 0 1 1
use contact_33  contact_33_471
timestamp 1624857261
transform 1 0 115600 0 1 45837
box 0 0 1 1
use contact_33  contact_33_472
timestamp 1624857261
transform 1 0 115600 0 1 45565
box 0 0 1 1
use contact_33  contact_33_499
timestamp 1624857261
transform 1 0 115736 0 1 45973
box 0 0 1 1
use contact_33  contact_33_500
timestamp 1624857261
transform 1 0 115736 0 1 46245
box 0 0 1 1
use contact_33  contact_33_2748
timestamp 1624857261
transform 1 0 116008 0 1 45973
box 0 0 1 1
use contact_33  contact_33_2749
timestamp 1624857261
transform 1 0 116008 0 1 46245
box 0 0 1 1
use contact_33  contact_33_93
timestamp 1624857261
transform 1 0 116824 0 1 46245
box 0 0 1 1
use contact_33  contact_33_94
timestamp 1624857261
transform 1 0 116824 0 1 45973
box 0 0 1 1
use contact_33  contact_33_125
timestamp 1624857261
transform 1 0 116960 0 1 45837
box 0 0 1 1
use contact_33  contact_33_126
timestamp 1624857261
transform 1 0 116960 0 1 45565
box 0 0 1 1
use contact_33  contact_33_2658
timestamp 1624857261
transform 1 0 116416 0 1 45565
box 0 0 1 1
use contact_33  contact_33_2659
timestamp 1624857261
transform 1 0 116416 0 1 45837
box 0 0 1 1
use contact_33  contact_33_3384
timestamp 1624857261
transform 1 0 115192 0 1 46381
box 0 0 1 1
use contact_33  contact_33_3385
timestamp 1624857261
transform 1 0 115192 0 1 46653
box 0 0 1 1
use contact_33  contact_33_703
timestamp 1624857261
transform 1 0 115600 0 1 46381
box 0 0 1 1
use contact_33  contact_33_704
timestamp 1624857261
transform 1 0 115600 0 1 46653
box 0 0 1 1
use contact_33  contact_33_2818
timestamp 1624857261
transform 1 0 116144 0 1 46789
box 0 0 1 1
use contact_33  contact_33_2819
timestamp 1624857261
transform 1 0 116144 0 1 47061
box 0 0 1 1
use contact_33  contact_33_67
timestamp 1624857261
transform 1 0 116824 0 1 46653
box 0 0 1 1
use contact_33  contact_33_68
timestamp 1624857261
transform 1 0 116824 0 1 46381
box 0 0 1 1
use contact_33  contact_33_73
timestamp 1624857261
transform 1 0 116824 0 1 46789
box 0 0 1 1
use contact_33  contact_33_74
timestamp 1624857261
transform 1 0 116824 0 1 47061
box 0 0 1 1
use contact_33  contact_33_2816
timestamp 1624857261
transform 1 0 116280 0 1 46789
box 0 0 1 1
use contact_33  contact_33_2817
timestamp 1624857261
transform 1 0 116280 0 1 47061
box 0 0 1 1
use contact_33  contact_33_3395
timestamp 1624857261
transform 1 0 115192 0 1 47877
box 0 0 1 1
use contact_33  contact_33_673
timestamp 1624857261
transform 1 0 115736 0 1 47877
box 0 0 1 1
use contact_33  contact_33_133
timestamp 1624857261
transform 1 0 116960 0 1 47197
box 0 0 1 1
use contact_33  contact_33_134
timestamp 1624857261
transform 1 0 116960 0 1 47469
box 0 0 1 1
use contact_33  contact_33_2544
timestamp 1624857261
transform 1 0 116552 0 1 47469
box 0 0 1 1
use contact_33  contact_33_2545
timestamp 1624857261
transform 1 0 116552 0 1 47741
box 0 0 1 1
use contact_33  contact_33_3140
timestamp 1624857261
transform 1 0 115328 0 1 48557
box 0 0 1 1
use contact_33  contact_33_3141
timestamp 1624857261
transform 1 0 115328 0 1 48285
box 0 0 1 1
use contact_33  contact_33_3162
timestamp 1624857261
transform 1 0 115192 0 1 48693
box 0 0 1 1
use contact_33  contact_33_3394
timestamp 1624857261
transform 1 0 115192 0 1 48149
box 0 0 1 1
use contact_33  contact_33_494
timestamp 1624857261
transform 1 0 115600 0 1 48693
box 0 0 1 1
use contact_33  contact_33_674
timestamp 1624857261
transform 1 0 115736 0 1 48149
box 0 0 1 1
use contact_33  contact_33_675
timestamp 1624857261
transform 1 0 115736 0 1 48557
box 0 0 1 1
use contact_33  contact_33_676
timestamp 1624857261
transform 1 0 115736 0 1 48285
box 0 0 1 1
use contact_33  contact_33_2837
timestamp 1624857261
transform 1 0 116144 0 1 48149
box 0 0 1 1
use contact_33  contact_33_2924
timestamp 1624857261
transform 1 0 116144 0 1 48285
box 0 0 1 1
use contact_33  contact_33_2925
timestamp 1624857261
transform 1 0 116144 0 1 48557
box 0 0 1 1
use contact_33  contact_33_155
timestamp 1624857261
transform 1 0 116960 0 1 48693
box 0 0 1 1
use contact_33  contact_33_181
timestamp 1624857261
transform 1 0 116824 0 1 48013
box 0 0 1 1
use contact_33  contact_33_182
timestamp 1624857261
transform 1 0 116824 0 1 48285
box 0 0 1 1
use contact_33  contact_33_2669
timestamp 1624857261
transform 1 0 116552 0 1 48693
box 0 0 1 1
use contact_33  contact_33_2836
timestamp 1624857261
transform 1 0 116280 0 1 48013
box 0 0 1 1
use contact_33  contact_33_2838
timestamp 1624857261
transform 1 0 116280 0 1 48557
box 0 0 1 1
use contact_33  contact_33_2839
timestamp 1624857261
transform 1 0 116280 0 1 48285
box 0 0 1 1
use contact_33  contact_33_3163
timestamp 1624857261
transform 1 0 115192 0 1 48965
box 0 0 1 1
use contact_33  contact_33_3246
timestamp 1624857261
transform 1 0 115328 0 1 49101
box 0 0 1 1
use contact_33  contact_33_3247
timestamp 1624857261
transform 1 0 115328 0 1 49373
box 0 0 1 1
use contact_33  contact_33_3249
timestamp 1624857261
transform 1 0 115328 0 1 49509
box 0 0 1 1
use contact_33  contact_33_493
timestamp 1624857261
transform 1 0 115600 0 1 48965
box 0 0 1 1
use contact_33  contact_33_647
timestamp 1624857261
transform 1 0 115736 0 1 49101
box 0 0 1 1
use contact_33  contact_33_648
timestamp 1624857261
transform 1 0 115736 0 1 49373
box 0 0 1 1
use contact_33  contact_33_650
timestamp 1624857261
transform 1 0 115736 0 1 49509
box 0 0 1 1
use contact_33  contact_33_2744
timestamp 1624857261
transform 1 0 116008 0 1 49509
box 0 0 1 1
use contact_33  contact_33_156
timestamp 1624857261
transform 1 0 116960 0 1 48965
box 0 0 1 1
use contact_33  contact_33_157
timestamp 1624857261
transform 1 0 116824 0 1 49373
box 0 0 1 1
use contact_33  contact_33_158
timestamp 1624857261
transform 1 0 116824 0 1 49101
box 0 0 1 1
use contact_33  contact_33_403
timestamp 1624857261
transform 1 0 116960 0 1 49509
box 0 0 1 1
use contact_33  contact_33_2564
timestamp 1624857261
transform 1 0 116416 0 1 49101
box 0 0 1 1
use contact_33  contact_33_2565
timestamp 1624857261
transform 1 0 116416 0 1 49373
box 0 0 1 1
use contact_33  contact_33_2668
timestamp 1624857261
transform 1 0 116552 0 1 48965
box 0 0 1 1
use contact_33  contact_33_3248
timestamp 1624857261
transform 1 0 115328 0 1 49781
box 0 0 1 1
use contact_33  contact_33_3293
timestamp 1624857261
transform 1 0 115328 0 1 50325
box 0 0 1 1
use contact_33  contact_33_3294
timestamp 1624857261
transform 1 0 115328 0 1 49917
box 0 0 1 1
use contact_33  contact_33_3295
timestamp 1624857261
transform 1 0 115328 0 1 50189
box 0 0 1 1
use contact_33  contact_33_591
timestamp 1624857261
transform 1 0 115600 0 1 50189
box 0 0 1 1
use contact_33  contact_33_592
timestamp 1624857261
transform 1 0 115600 0 1 49917
box 0 0 1 1
use contact_33  contact_33_649
timestamp 1624857261
transform 1 0 115736 0 1 49781
box 0 0 1 1
use contact_33  contact_33_701
timestamp 1624857261
transform 1 0 115736 0 1 50325
box 0 0 1 1
use contact_33  contact_33_2745
timestamp 1624857261
transform 1 0 116008 0 1 49781
box 0 0 1 1
use contact_33  contact_33_2746
timestamp 1624857261
transform 1 0 116144 0 1 50189
box 0 0 1 1
use contact_33  contact_33_2747
timestamp 1624857261
transform 1 0 116144 0 1 49917
box 0 0 1 1
use contact_33  contact_33_2764
timestamp 1624857261
transform 1 0 116008 0 1 50325
box 0 0 1 1
use contact_33  contact_33_91
timestamp 1624857261
transform 1 0 116824 0 1 50325
box 0 0 1 1
use contact_33  contact_33_401
timestamp 1624857261
transform 1 0 116960 0 1 50189
box 0 0 1 1
use contact_33  contact_33_402
timestamp 1624857261
transform 1 0 116960 0 1 49917
box 0 0 1 1
use contact_33  contact_33_404
timestamp 1624857261
transform 1 0 116960 0 1 49781
box 0 0 1 1
use contact_33  contact_33_2684
timestamp 1624857261
transform 1 0 116416 0 1 50325
box 0 0 1 1
use contact_33  contact_33_2742
timestamp 1624857261
transform 1 0 116280 0 1 50189
box 0 0 1 1
use contact_33  contact_33_2743
timestamp 1624857261
transform 1 0 116280 0 1 49917
box 0 0 1 1
use contact_33  contact_33_3180
timestamp 1624857261
transform 1 0 115192 0 1 51005
box 0 0 1 1
use contact_33  contact_33_3181
timestamp 1624857261
transform 1 0 115192 0 1 50733
box 0 0 1 1
use contact_33  contact_33_3292
timestamp 1624857261
transform 1 0 115328 0 1 50597
box 0 0 1 1
use contact_33  contact_33_702
timestamp 1624857261
transform 1 0 115736 0 1 50597
box 0 0 1 1
use contact_33  contact_33_781
timestamp 1624857261
transform 1 0 115600 0 1 50733
box 0 0 1 1
use contact_33  contact_33_782
timestamp 1624857261
transform 1 0 115600 0 1 51005
box 0 0 1 1
use contact_33  contact_33_2765
timestamp 1624857261
transform 1 0 116008 0 1 50597
box 0 0 1 1
use contact_33  contact_33_89
timestamp 1624857261
transform 1 0 116824 0 1 51005
box 0 0 1 1
use contact_33  contact_33_90
timestamp 1624857261
transform 1 0 116824 0 1 50733
box 0 0 1 1
use contact_33  contact_33_92
timestamp 1624857261
transform 1 0 116824 0 1 50597
box 0 0 1 1
use contact_33  contact_33_211
timestamp 1624857261
transform 1 0 116824 0 1 51141
box 0 0 1 1
use contact_33  contact_33_2682
timestamp 1624857261
transform 1 0 116552 0 1 51005
box 0 0 1 1
use contact_33  contact_33_2683
timestamp 1624857261
transform 1 0 116552 0 1 50733
box 0 0 1 1
use contact_33  contact_33_2685
timestamp 1624857261
transform 1 0 116416 0 1 50597
box 0 0 1 1
use contact_33  contact_33_3103
timestamp 1624857261
transform 1 0 115192 0 1 51821
box 0 0 1 1
use contact_33  contact_33_553
timestamp 1624857261
transform 1 0 115600 0 1 51821
box 0 0 1 1
use contact_33  contact_33_2972
timestamp 1624857261
transform 1 0 116008 0 1 51413
box 0 0 1 1
use contact_33  contact_33_2973
timestamp 1624857261
transform 1 0 116008 0 1 51685
box 0 0 1 1
use contact_33  contact_33_179
timestamp 1624857261
transform 1 0 116960 0 1 51957
box 0 0 1 1
use contact_33  contact_33_212
timestamp 1624857261
transform 1 0 116824 0 1 51413
box 0 0 1 1
use contact_33  contact_33_2568
timestamp 1624857261
transform 1 0 116416 0 1 51413
box 0 0 1 1
use contact_33  contact_33_2569
timestamp 1624857261
transform 1 0 116416 0 1 51685
box 0 0 1 1
use contact_33  contact_33_3102
timestamp 1624857261
transform 1 0 115192 0 1 52093
box 0 0 1 1
use contact_33  contact_33_3177
timestamp 1624857261
transform 1 0 115328 0 1 52637
box 0 0 1 1
use contact_33  contact_33_3178
timestamp 1624857261
transform 1 0 115328 0 1 52229
box 0 0 1 1
use contact_33  contact_33_3179
timestamp 1624857261
transform 1 0 115328 0 1 52501
box 0 0 1 1
use contact_33  contact_33_554
timestamp 1624857261
transform 1 0 115600 0 1 52093
box 0 0 1 1
use contact_33  contact_33_802
timestamp 1624857261
transform 1 0 115736 0 1 52637
box 0 0 1 1
use contact_33  contact_33_803
timestamp 1624857261
transform 1 0 115736 0 1 52229
box 0 0 1 1
use contact_33  contact_33_804
timestamp 1624857261
transform 1 0 115736 0 1 52501
box 0 0 1 1
use contact_33  contact_33_2730
timestamp 1624857261
transform 1 0 116008 0 1 52501
box 0 0 1 1
use contact_33  contact_33_2731
timestamp 1624857261
transform 1 0 116008 0 1 52229
box 0 0 1 1
use contact_33  contact_33_2988
timestamp 1624857261
transform 1 0 116144 0 1 52637
box 0 0 1 1
use contact_33  contact_33_180
timestamp 1624857261
transform 1 0 116960 0 1 52229
box 0 0 1 1
use contact_33  contact_33_258
timestamp 1624857261
transform 1 0 116824 0 1 52637
box 0 0 1 1
use contact_33  contact_33_2657
timestamp 1624857261
transform 1 0 116416 0 1 52637
box 0 0 1 1
use contact_33  contact_33_2706
timestamp 1624857261
transform 1 0 116280 0 1 52229
box 0 0 1 1
use contact_33  contact_33_2707
timestamp 1624857261
transform 1 0 116280 0 1 52501
box 0 0 1 1
use contact_33  contact_33_2986
timestamp 1624857261
transform 1 0 116280 0 1 52637
box 0 0 1 1
use contact_33  contact_33_3088
timestamp 1624857261
transform 1 0 115192 0 1 53317
box 0 0 1 1
use contact_33  contact_33_3089
timestamp 1624857261
transform 1 0 115192 0 1 53045
box 0 0 1 1
use contact_33  contact_33_3176
timestamp 1624857261
transform 1 0 115328 0 1 52909
box 0 0 1 1
use contact_33  contact_33_3198
timestamp 1624857261
transform 1 0 115328 0 1 53453
box 0 0 1 1
use contact_33  contact_33_538
timestamp 1624857261
transform 1 0 115736 0 1 53453
box 0 0 1 1
use contact_33  contact_33_539
timestamp 1624857261
transform 1 0 115600 0 1 53045
box 0 0 1 1
use contact_33  contact_33_540
timestamp 1624857261
transform 1 0 115600 0 1 53317
box 0 0 1 1
use contact_33  contact_33_801
timestamp 1624857261
transform 1 0 115736 0 1 52909
box 0 0 1 1
use contact_33  contact_33_2989
timestamp 1624857261
transform 1 0 116144 0 1 52909
box 0 0 1 1
use contact_33  contact_33_257
timestamp 1624857261
transform 1 0 116824 0 1 52909
box 0 0 1 1
use contact_33  contact_33_429
timestamp 1624857261
transform 1 0 116824 0 1 53453
box 0 0 1 1
use contact_33  contact_33_2622
timestamp 1624857261
transform 1 0 116552 0 1 53045
box 0 0 1 1
use contact_33  contact_33_2623
timestamp 1624857261
transform 1 0 116552 0 1 53317
box 0 0 1 1
use contact_33  contact_33_2656
timestamp 1624857261
transform 1 0 116416 0 1 52909
box 0 0 1 1
use contact_33  contact_33_2777
timestamp 1624857261
transform 1 0 116280 0 1 53453
box 0 0 1 1
use contact_33  contact_33_2987
timestamp 1624857261
transform 1 0 116280 0 1 52909
box 0 0 1 1
use contact_33  contact_33_3078
timestamp 1624857261
transform 1 0 115328 0 1 54269
box 0 0 1 1
use contact_33  contact_33_3196
timestamp 1624857261
transform 1 0 115328 0 1 54133
box 0 0 1 1
use contact_33  contact_33_3197
timestamp 1624857261
transform 1 0 115328 0 1 53861
box 0 0 1 1
use contact_33  contact_33_3199
timestamp 1624857261
transform 1 0 115328 0 1 53725
box 0 0 1 1
use contact_33  contact_33_527
timestamp 1624857261
transform 1 0 115600 0 1 53861
box 0 0 1 1
use contact_33  contact_33_528
timestamp 1624857261
transform 1 0 115600 0 1 54133
box 0 0 1 1
use contact_33  contact_33_537
timestamp 1624857261
transform 1 0 115736 0 1 53725
box 0 0 1 1
use contact_33  contact_33_545
timestamp 1624857261
transform 1 0 115736 0 1 54269
box 0 0 1 1
use contact_33  contact_33_2790
timestamp 1624857261
transform 1 0 116008 0 1 54133
box 0 0 1 1
use contact_33  contact_33_2791
timestamp 1624857261
transform 1 0 116008 0 1 53861
box 0 0 1 1
use contact_33  contact_33_2990
timestamp 1624857261
transform 1 0 116144 0 1 54269
box 0 0 1 1
use contact_33  contact_33_319
timestamp 1624857261
transform 1 0 116824 0 1 54269
box 0 0 1 1
use contact_33  contact_33_427
timestamp 1624857261
transform 1 0 116824 0 1 54133
box 0 0 1 1
use contact_33  contact_33_428
timestamp 1624857261
transform 1 0 116824 0 1 53861
box 0 0 1 1
use contact_33  contact_33_430
timestamp 1624857261
transform 1 0 116824 0 1 53725
box 0 0 1 1
use contact_33  contact_33_2688
timestamp 1624857261
transform 1 0 116416 0 1 54133
box 0 0 1 1
use contact_33  contact_33_2689
timestamp 1624857261
transform 1 0 116416 0 1 53861
box 0 0 1 1
use contact_33  contact_33_2773
timestamp 1624857261
transform 1 0 116280 0 1 54269
box 0 0 1 1
use contact_33  contact_33_2776
timestamp 1624857261
transform 1 0 116280 0 1 53725
box 0 0 1 1
use contact_33  contact_33_3079
timestamp 1624857261
transform 1 0 115328 0 1 54541
box 0 0 1 1
use contact_33  contact_33_3256
timestamp 1624857261
transform 1 0 115192 0 1 54677
box 0 0 1 1
use contact_33  contact_33_3257
timestamp 1624857261
transform 1 0 115192 0 1 54949
box 0 0 1 1
use contact_33  contact_33_546
timestamp 1624857261
transform 1 0 115736 0 1 54541
box 0 0 1 1
use contact_33  contact_33_671
timestamp 1624857261
transform 1 0 115736 0 1 54677
box 0 0 1 1
use contact_33  contact_33_672
timestamp 1624857261
transform 1 0 115736 0 1 54949
box 0 0 1 1
use contact_33  contact_33_2991
timestamp 1624857261
transform 1 0 116144 0 1 54541
box 0 0 1 1
use contact_33  contact_33_193
timestamp 1624857261
transform 1 0 116960 0 1 55085
box 0 0 1 1
use contact_33  contact_33_317
timestamp 1624857261
transform 1 0 116824 0 1 54949
box 0 0 1 1
use contact_33  contact_33_318
timestamp 1624857261
transform 1 0 116824 0 1 54677
box 0 0 1 1
use contact_33  contact_33_320
timestamp 1624857261
transform 1 0 116824 0 1 54541
box 0 0 1 1
use contact_33  contact_33_2722
timestamp 1624857261
transform 1 0 116280 0 1 54677
box 0 0 1 1
use contact_33  contact_33_2723
timestamp 1624857261
transform 1 0 116280 0 1 54949
box 0 0 1 1
use contact_33  contact_33_2772
timestamp 1624857261
transform 1 0 116280 0 1 54541
box 0 0 1 1
use contact_33  contact_33_194
timestamp 1624857261
transform 1 0 116960 0 1 55357
box 0 0 1 1
use contact_33  contact_33_196
timestamp 1624857261
transform 1 0 116960 0 1 55493
box 0 0 1 1
use contact_33  contact_33_2677
timestamp 1624857261
transform 1 0 116552 0 1 55493
box 0 0 1 1
use contact_33  contact_33_835
timestamp 1624857261
transform 1 0 110432 0 1 55901
box 0 0 1 1
use contact_33  contact_33_875
timestamp 1624857261
transform 1 0 110432 0 1 56037
box 0 0 1 1
use contact_33  contact_33_876
timestamp 1624857261
transform 1 0 110432 0 1 56309
box 0 0 1 1
use contact_33  contact_33_910
timestamp 1624857261
transform 1 0 110432 0 1 58349
box 0 0 1 1
use contact_33  contact_33_827
timestamp 1624857261
transform 1 0 110160 0 1 59573
box 0 0 1 1
use contact_33  contact_33_828
timestamp 1624857261
transform 1 0 110160 0 1 59845
box 0 0 1 1
use contact_33  contact_33_907
timestamp 1624857261
transform 1 0 110432 0 1 59437
box 0 0 1 1
use contact_33  contact_33_908
timestamp 1624857261
transform 1 0 110432 0 1 59165
box 0 0 1 1
use contact_33  contact_33_909
timestamp 1624857261
transform 1 0 110432 0 1 58621
box 0 0 1 1
use contact_33  contact_33_913
timestamp 1624857261
transform 1 0 110432 0 1 61069
box 0 0 1 1
use contact_33  contact_33_914
timestamp 1624857261
transform 1 0 110432 0 1 60797
box 0 0 1 1
use contact_33  contact_33_873
timestamp 1624857261
transform 1 0 110160 0 1 63925
box 0 0 1 1
use contact_33  contact_33_895
timestamp 1624857261
transform 1 0 110160 0 1 62565
box 0 0 1 1
use contact_33  contact_33_896
timestamp 1624857261
transform 1 0 110160 0 1 62293
box 0 0 1 1
use contact_33  contact_33_939
timestamp 1624857261
transform 1 0 110432 0 1 63789
box 0 0 1 1
use contact_33  contact_33_940
timestamp 1624857261
transform 1 0 110432 0 1 63517
box 0 0 1 1
use contact_33  contact_33_874
timestamp 1624857261
transform 1 0 110160 0 1 64197
box 0 0 1 1
use contact_33  contact_33_863
timestamp 1624857261
transform 1 0 110432 0 1 68957
box 0 0 1 1
use contact_33  contact_33_864
timestamp 1624857261
transform 1 0 110432 0 1 68685
box 0 0 1 1
use contact_33  contact_33_887
timestamp 1624857261
transform 1 0 110296 0 1 67053
box 0 0 1 1
use contact_33  contact_33_888
timestamp 1624857261
transform 1 0 110296 0 1 67325
box 0 0 1 1
use contact_33  contact_33_945
timestamp 1624857261
transform 1 0 110432 0 1 68141
box 0 0 1 1
use contact_33  contact_33_946
timestamp 1624857261
transform 1 0 110432 0 1 67869
box 0 0 1 1
use contact_33  contact_33_920
timestamp 1624857261
transform 1 0 113288 0 1 69637
box 0 0 1 1
use contact_33  contact_33_829
timestamp 1624857261
transform 1 0 110432 0 1 72493
box 0 0 1 1
use contact_33  contact_33_830
timestamp 1624857261
transform 1 0 110432 0 1 72221
box 0 0 1 1
use contact_33  contact_33_919
timestamp 1624857261
transform 1 0 113288 0 1 70317
box 0 0 1 1
use contact_33  contact_33_3108
timestamp 1624857261
transform 1 0 115192 0 1 56445
box 0 0 1 1
use contact_33  contact_33_3109
timestamp 1624857261
transform 1 0 115192 0 1 56173
box 0 0 1 1
use contact_33  contact_33_747
timestamp 1624857261
transform 1 0 115600 0 1 56173
box 0 0 1 1
use contact_33  contact_33_748
timestamp 1624857261
transform 1 0 115600 0 1 56445
box 0 0 1 1
use contact_33  contact_33_163
timestamp 1624857261
transform 1 0 116960 0 1 55901
box 0 0 1 1
use contact_33  contact_33_164
timestamp 1624857261
transform 1 0 116960 0 1 56173
box 0 0 1 1
use contact_33  contact_33_195
timestamp 1624857261
transform 1 0 116960 0 1 55765
box 0 0 1 1
use contact_33  contact_33_2554
timestamp 1624857261
transform 1 0 116552 0 1 56173
box 0 0 1 1
use contact_33  contact_33_2555
timestamp 1624857261
transform 1 0 116552 0 1 56445
box 0 0 1 1
use contact_33  contact_33_2676
timestamp 1624857261
transform 1 0 116552 0 1 55765
box 0 0 1 1
use contact_33  contact_33_3030
timestamp 1624857261
transform 1 0 115328 0 1 57261
box 0 0 1 1
use contact_33  contact_33_3031
timestamp 1624857261
transform 1 0 115328 0 1 56989
box 0 0 1 1
use contact_33  contact_33_3104
timestamp 1624857261
transform 1 0 115192 0 1 56853
box 0 0 1 1
use contact_33  contact_33_3105
timestamp 1624857261
transform 1 0 115192 0 1 56581
box 0 0 1 1
use contact_33  contact_33_3322
timestamp 1624857261
transform 1 0 115192 0 1 57397
box 0 0 1 1
use contact_33  contact_33_625
timestamp 1624857261
transform 1 0 115600 0 1 57397
box 0 0 1 1
use contact_33  contact_33_687
timestamp 1624857261
transform 1 0 115736 0 1 57261
box 0 0 1 1
use contact_33  contact_33_688
timestamp 1624857261
transform 1 0 115736 0 1 56989
box 0 0 1 1
use contact_33  contact_33_749
timestamp 1624857261
transform 1 0 115600 0 1 56853
box 0 0 1 1
use contact_33  contact_33_750
timestamp 1624857261
transform 1 0 115600 0 1 56581
box 0 0 1 1
use contact_33  contact_33_2738
timestamp 1624857261
transform 1 0 116280 0 1 56989
box 0 0 1 1
use contact_33  contact_33_2739
timestamp 1624857261
transform 1 0 116280 0 1 57261
box 0 0 1 1
use contact_33  contact_33_2740
timestamp 1624857261
transform 1 0 116144 0 1 56989
box 0 0 1 1
use contact_33  contact_33_2741
timestamp 1624857261
transform 1 0 116144 0 1 57261
box 0 0 1 1
use contact_33  contact_33_236
timestamp 1624857261
transform 1 0 116960 0 1 57397
box 0 0 1 1
use contact_33  contact_33_2672
timestamp 1624857261
transform 1 0 116552 0 1 57397
box 0 0 1 1
use contact_33  contact_33_3298
timestamp 1624857261
transform 1 0 115192 0 1 58213
box 0 0 1 1
use contact_33  contact_33_3323
timestamp 1624857261
transform 1 0 115192 0 1 57669
box 0 0 1 1
use contact_33  contact_33_3324
timestamp 1624857261
transform 1 0 115192 0 1 58077
box 0 0 1 1
use contact_33  contact_33_3325
timestamp 1624857261
transform 1 0 115192 0 1 57805
box 0 0 1 1
use contact_33  contact_33_490
timestamp 1624857261
transform 1 0 115736 0 1 58213
box 0 0 1 1
use contact_33  contact_33_626
timestamp 1624857261
transform 1 0 115600 0 1 57669
box 0 0 1 1
use contact_33  contact_33_627
timestamp 1624857261
transform 1 0 115736 0 1 58077
box 0 0 1 1
use contact_33  contact_33_628
timestamp 1624857261
transform 1 0 115736 0 1 57805
box 0 0 1 1
use contact_33  contact_33_2885
timestamp 1624857261
transform 1 0 116008 0 1 58213
box 0 0 1 1
use contact_33  contact_33_235
timestamp 1624857261
transform 1 0 116960 0 1 57669
box 0 0 1 1
use contact_33  contact_33_377
timestamp 1624857261
transform 1 0 116824 0 1 57805
box 0 0 1 1
use contact_33  contact_33_378
timestamp 1624857261
transform 1 0 116824 0 1 58077
box 0 0 1 1
use contact_33  contact_33_380
timestamp 1624857261
transform 1 0 116824 0 1 58213
box 0 0 1 1
use contact_33  contact_33_2673
timestamp 1624857261
transform 1 0 116552 0 1 57669
box 0 0 1 1
use contact_33  contact_33_3273
timestamp 1624857261
transform 1 0 115328 0 1 59029
box 0 0 1 1
use contact_33  contact_33_3299
timestamp 1624857261
transform 1 0 115192 0 1 58485
box 0 0 1 1
use contact_33  contact_33_3300
timestamp 1624857261
transform 1 0 115192 0 1 58893
box 0 0 1 1
use contact_33  contact_33_3301
timestamp 1624857261
transform 1 0 115192 0 1 58621
box 0 0 1 1
use contact_33  contact_33_489
timestamp 1624857261
transform 1 0 115736 0 1 58485
box 0 0 1 1
use contact_33  contact_33_606
timestamp 1624857261
transform 1 0 115736 0 1 59029
box 0 0 1 1
use contact_33  contact_33_607
timestamp 1624857261
transform 1 0 115736 0 1 58621
box 0 0 1 1
use contact_33  contact_33_608
timestamp 1624857261
transform 1 0 115736 0 1 58893
box 0 0 1 1
use contact_33  contact_33_2884
timestamp 1624857261
transform 1 0 116008 0 1 58485
box 0 0 1 1
use contact_33  contact_33_2906
timestamp 1624857261
transform 1 0 116144 0 1 58621
box 0 0 1 1
use contact_33  contact_33_2907
timestamp 1624857261
transform 1 0 116144 0 1 58893
box 0 0 1 1
use contact_33  contact_33_379
timestamp 1624857261
transform 1 0 116824 0 1 58485
box 0 0 1 1
use contact_33  contact_33_439
timestamp 1624857261
transform 1 0 116824 0 1 58621
box 0 0 1 1
use contact_33  contact_33_440
timestamp 1624857261
transform 1 0 116824 0 1 58893
box 0 0 1 1
use contact_33  contact_33_442
timestamp 1624857261
transform 1 0 116824 0 1 59029
box 0 0 1 1
use contact_33  contact_33_2608
timestamp 1624857261
transform 1 0 116552 0 1 58893
box 0 0 1 1
use contact_33  contact_33_2609
timestamp 1624857261
transform 1 0 116552 0 1 58621
box 0 0 1 1
use contact_33  contact_33_3272
timestamp 1624857261
transform 1 0 115328 0 1 59301
box 0 0 1 1
use contact_33  contact_33_605
timestamp 1624857261
transform 1 0 115736 0 1 59301
box 0 0 1 1
use contact_33  contact_33_149
timestamp 1624857261
transform 1 0 116824 0 1 59845
box 0 0 1 1
use contact_33  contact_33_335
timestamp 1624857261
transform 1 0 116960 0 1 59709
box 0 0 1 1
use contact_33  contact_33_336
timestamp 1624857261
transform 1 0 116960 0 1 59437
box 0 0 1 1
use contact_33  contact_33_441
timestamp 1624857261
transform 1 0 116824 0 1 59301
box 0 0 1 1
use contact_33  contact_33_2634
timestamp 1624857261
transform 1 0 116552 0 1 59437
box 0 0 1 1
use contact_33  contact_33_2635
timestamp 1624857261
transform 1 0 116552 0 1 59709
box 0 0 1 1
use contact_33  contact_33_3110
timestamp 1624857261
transform 1 0 115192 0 1 60525
box 0 0 1 1
use contact_33  contact_33_3111
timestamp 1624857261
transform 1 0 115192 0 1 60797
box 0 0 1 1
use contact_33  contact_33_3134
timestamp 1624857261
transform 1 0 115328 0 1 60389
box 0 0 1 1
use contact_33  contact_33_3135
timestamp 1624857261
transform 1 0 115328 0 1 60117
box 0 0 1 1
use contact_33  contact_33_725
timestamp 1624857261
transform 1 0 115600 0 1 60797
box 0 0 1 1
use contact_33  contact_33_726
timestamp 1624857261
transform 1 0 115600 0 1 60525
box 0 0 1 1
use contact_33  contact_33_729
timestamp 1624857261
transform 1 0 115736 0 1 60389
box 0 0 1 1
use contact_33  contact_33_730
timestamp 1624857261
transform 1 0 115736 0 1 60117
box 0 0 1 1
use contact_33  contact_33_2940
timestamp 1624857261
transform 1 0 116008 0 1 60117
box 0 0 1 1
use contact_33  contact_33_2941
timestamp 1624857261
transform 1 0 116008 0 1 60389
box 0 0 1 1
use contact_33  contact_33_150
timestamp 1624857261
transform 1 0 116824 0 1 60117
box 0 0 1 1
use contact_33  contact_33_2628
timestamp 1624857261
transform 1 0 116416 0 1 60117
box 0 0 1 1
use contact_33  contact_33_2629
timestamp 1624857261
transform 1 0 116416 0 1 60389
box 0 0 1 1
use contact_33  contact_33_3064
timestamp 1624857261
transform 1 0 115328 0 1 61613
box 0 0 1 1
use contact_33  contact_33_3065
timestamp 1624857261
transform 1 0 115328 0 1 61341
box 0 0 1 1
use contact_33  contact_33_3112
timestamp 1624857261
transform 1 0 115192 0 1 61205
box 0 0 1 1
use contact_33  contact_33_3113
timestamp 1624857261
transform 1 0 115192 0 1 60933
box 0 0 1 1
use contact_33  contact_33_541
timestamp 1624857261
transform 1 0 115736 0 1 61613
box 0 0 1 1
use contact_33  contact_33_542
timestamp 1624857261
transform 1 0 115736 0 1 61341
box 0 0 1 1
use contact_33  contact_33_543
timestamp 1624857261
transform 1 0 115736 0 1 60933
box 0 0 1 1
use contact_33  contact_33_544
timestamp 1624857261
transform 1 0 115736 0 1 61205
box 0 0 1 1
use contact_33  contact_33_2760
timestamp 1624857261
transform 1 0 116008 0 1 60933
box 0 0 1 1
use contact_33  contact_33_2761
timestamp 1624857261
transform 1 0 116008 0 1 61205
box 0 0 1 1
use contact_33  contact_33_3006
timestamp 1624857261
transform 1 0 116144 0 1 61341
box 0 0 1 1
use contact_33  contact_33_3007
timestamp 1624857261
transform 1 0 116144 0 1 61613
box 0 0 1 1
use contact_33  contact_33_207
timestamp 1624857261
transform 1 0 116824 0 1 61613
box 0 0 1 1
use contact_33  contact_33_208
timestamp 1624857261
transform 1 0 116824 0 1 61341
box 0 0 1 1
use contact_33  contact_33_2556
timestamp 1624857261
transform 1 0 116552 0 1 61205
box 0 0 1 1
use contact_33  contact_33_2557
timestamp 1624857261
transform 1 0 116552 0 1 60933
box 0 0 1 1
use contact_33  contact_33_3026
timestamp 1624857261
transform 1 0 115192 0 1 61749
box 0 0 1 1
use contact_33  contact_33_3027
timestamp 1624857261
transform 1 0 115192 0 1 62021
box 0 0 1 1
use contact_33  contact_33_3056
timestamp 1624857261
transform 1 0 115328 0 1 62157
box 0 0 1 1
use contact_33  contact_33_3057
timestamp 1624857261
transform 1 0 115328 0 1 62429
box 0 0 1 1
use contact_33  contact_33_3082
timestamp 1624857261
transform 1 0 115192 0 1 62565
box 0 0 1 1
use contact_33  contact_33_665
timestamp 1624857261
transform 1 0 115600 0 1 62565
box 0 0 1 1
use contact_33  contact_33_719
timestamp 1624857261
transform 1 0 115600 0 1 61749
box 0 0 1 1
use contact_33  contact_33_720
timestamp 1624857261
transform 1 0 115600 0 1 62021
box 0 0 1 1
use contact_33  contact_33_721
timestamp 1624857261
transform 1 0 115736 0 1 62429
box 0 0 1 1
use contact_33  contact_33_722
timestamp 1624857261
transform 1 0 115736 0 1 62157
box 0 0 1 1
use contact_33  contact_33_2726
timestamp 1624857261
transform 1 0 116280 0 1 62565
box 0 0 1 1
use contact_33  contact_33_2728
timestamp 1624857261
transform 1 0 116144 0 1 62565
box 0 0 1 1
use contact_33  contact_33_241
timestamp 1624857261
transform 1 0 116824 0 1 62429
box 0 0 1 1
use contact_33  contact_33_242
timestamp 1624857261
transform 1 0 116824 0 1 62157
box 0 0 1 1
use contact_33  contact_33_243
timestamp 1624857261
transform 1 0 116960 0 1 61749
box 0 0 1 1
use contact_33  contact_33_244
timestamp 1624857261
transform 1 0 116960 0 1 62021
box 0 0 1 1
use contact_33  contact_33_271
timestamp 1624857261
transform 1 0 116960 0 1 62565
box 0 0 1 1
use contact_33  contact_33_2562
timestamp 1624857261
transform 1 0 116416 0 1 62157
box 0 0 1 1
use contact_33  contact_33_2563
timestamp 1624857261
transform 1 0 116416 0 1 62429
box 0 0 1 1
use contact_33  contact_33_2624
timestamp 1624857261
transform 1 0 116552 0 1 62021
box 0 0 1 1
use contact_33  contact_33_2625
timestamp 1624857261
transform 1 0 116552 0 1 61749
box 0 0 1 1
use contact_33  contact_33_3080
timestamp 1624857261
transform 1 0 115192 0 1 63245
box 0 0 1 1
use contact_33  contact_33_3081
timestamp 1624857261
transform 1 0 115192 0 1 62973
box 0 0 1 1
use contact_33  contact_33_3083
timestamp 1624857261
transform 1 0 115192 0 1 62837
box 0 0 1 1
use contact_33  contact_33_666
timestamp 1624857261
transform 1 0 115600 0 1 62837
box 0 0 1 1
use contact_33  contact_33_667
timestamp 1624857261
transform 1 0 115600 0 1 63245
box 0 0 1 1
use contact_33  contact_33_668
timestamp 1624857261
transform 1 0 115600 0 1 62973
box 0 0 1 1
use contact_33  contact_33_2705
timestamp 1624857261
transform 1 0 116280 0 1 63381
box 0 0 1 1
use contact_33  contact_33_2727
timestamp 1624857261
transform 1 0 116280 0 1 62837
box 0 0 1 1
use contact_33  contact_33_2729
timestamp 1624857261
transform 1 0 116144 0 1 62837
box 0 0 1 1
use contact_33  contact_33_140
timestamp 1624857261
transform 1 0 116824 0 1 63381
box 0 0 1 1
use contact_33  contact_33_272
timestamp 1624857261
transform 1 0 116960 0 1 62837
box 0 0 1 1
use contact_33  contact_33_273
timestamp 1624857261
transform 1 0 116960 0 1 63245
box 0 0 1 1
use contact_33  contact_33_274
timestamp 1624857261
transform 1 0 116960 0 1 62973
box 0 0 1 1
use contact_33  contact_33_2704
timestamp 1624857261
transform 1 0 116280 0 1 63653
box 0 0 1 1
use contact_33  contact_33_2843
timestamp 1624857261
transform 1 0 116008 0 1 64061
box 0 0 1 1
use contact_33  contact_33_131
timestamp 1624857261
transform 1 0 116824 0 1 64061
box 0 0 1 1
use contact_33  contact_33_132
timestamp 1624857261
transform 1 0 116824 0 1 63789
box 0 0 1 1
use contact_33  contact_33_139
timestamp 1624857261
transform 1 0 116824 0 1 63653
box 0 0 1 1
use contact_33  contact_33_2603
timestamp 1624857261
transform 1 0 116552 0 1 64061
box 0 0 1 1
use contact_33  contact_33_3214
timestamp 1624857261
transform 1 0 115192 0 1 64877
box 0 0 1 1
use contact_33  contact_33_3318
timestamp 1624857261
transform 1 0 115328 0 1 64741
box 0 0 1 1
use contact_33  contact_33_3319
timestamp 1624857261
transform 1 0 115328 0 1 64469
box 0 0 1 1
use contact_33  contact_33_640
timestamp 1624857261
transform 1 0 115600 0 1 64877
box 0 0 1 1
use contact_33  contact_33_641
timestamp 1624857261
transform 1 0 115736 0 1 64469
box 0 0 1 1
use contact_33  contact_33_642
timestamp 1624857261
transform 1 0 115736 0 1 64741
box 0 0 1 1
use contact_33  contact_33_2842
timestamp 1624857261
transform 1 0 116008 0 1 64333
box 0 0 1 1
use contact_33  contact_33_2921
timestamp 1624857261
transform 1 0 116144 0 1 64877
box 0 0 1 1
use contact_33  contact_33_2602
timestamp 1624857261
transform 1 0 116552 0 1 64333
box 0 0 1 1
use contact_33  contact_33_3212
timestamp 1624857261
transform 1 0 115192 0 1 65557
box 0 0 1 1
use contact_33  contact_33_3213
timestamp 1624857261
transform 1 0 115192 0 1 65285
box 0 0 1 1
use contact_33  contact_33_3215
timestamp 1624857261
transform 1 0 115192 0 1 65149
box 0 0 1 1
use contact_33  contact_33_3362
timestamp 1624857261
transform 1 0 115192 0 1 65693
box 0 0 1 1
use contact_33  contact_33_3363
timestamp 1624857261
transform 1 0 115192 0 1 65965
box 0 0 1 1
use contact_33  contact_33_639
timestamp 1624857261
transform 1 0 115600 0 1 65149
box 0 0 1 1
use contact_33  contact_33_460
timestamp 1624857261
transform 1 0 115600 0 1 65285
box 0 0 1 1
use contact_33  contact_33_2920
timestamp 1624857261
transform 1 0 116144 0 1 65149
box 0 0 1 1
use contact_33  contact_33_2787
timestamp 1624857261
transform 1 0 116008 0 1 65285
box 0 0 1 1
use contact_33  contact_33_459
timestamp 1624857261
transform 1 0 115600 0 1 65557
box 0 0 1 1
use contact_33  contact_33_2786
timestamp 1624857261
transform 1 0 116008 0 1 65557
box 0 0 1 1
use contact_33  contact_33_517
timestamp 1624857261
transform 1 0 115600 0 1 65693
box 0 0 1 1
use contact_33  contact_33_2862
timestamp 1624857261
transform 1 0 116144 0 1 65693
box 0 0 1 1
use contact_33  contact_33_518
timestamp 1624857261
transform 1 0 115600 0 1 65965
box 0 0 1 1
use contact_33  contact_33_2863
timestamp 1624857261
transform 1 0 116144 0 1 65965
box 0 0 1 1
use contact_33  contact_33_275
timestamp 1624857261
transform 1 0 116824 0 1 65965
box 0 0 1 1
use contact_33  contact_33_276
timestamp 1624857261
transform 1 0 116824 0 1 65693
box 0 0 1 1
use contact_33  contact_33_277
timestamp 1624857261
transform 1 0 116824 0 1 65285
box 0 0 1 1
use contact_33  contact_33_278
timestamp 1624857261
transform 1 0 116824 0 1 65557
box 0 0 1 1
use contact_33  contact_33_2686
timestamp 1624857261
transform 1 0 116416 0 1 65965
box 0 0 1 1
use contact_33  contact_33_2687
timestamp 1624857261
transform 1 0 116416 0 1 65693
box 0 0 1 1
use contact_33  contact_33_3066
timestamp 1624857261
transform 1 0 115328 0 1 66509
box 0 0 1 1
use contact_33  contact_33_3067
timestamp 1624857261
transform 1 0 115328 0 1 66781
box 0 0 1 1
use contact_33  contact_33_3360
timestamp 1624857261
transform 1 0 115192 0 1 66373
box 0 0 1 1
use contact_33  contact_33_3361
timestamp 1624857261
transform 1 0 115192 0 1 66101
box 0 0 1 1
use contact_33  contact_33_449
timestamp 1624857261
transform 1 0 115736 0 1 66509
box 0 0 1 1
use contact_33  contact_33_450
timestamp 1624857261
transform 1 0 115736 0 1 66781
box 0 0 1 1
use contact_33  contact_33_515
timestamp 1624857261
transform 1 0 115600 0 1 66373
box 0 0 1 1
use contact_33  contact_33_516
timestamp 1624857261
transform 1 0 115600 0 1 66101
box 0 0 1 1
use contact_33  contact_33_2750
timestamp 1624857261
transform 1 0 116280 0 1 66781
box 0 0 1 1
use contact_33  contact_33_2751
timestamp 1624857261
transform 1 0 116280 0 1 66509
box 0 0 1 1
use contact_33  contact_33_69
timestamp 1624857261
transform 1 0 116824 0 1 66509
box 0 0 1 1
use contact_33  contact_33_70
timestamp 1624857261
transform 1 0 116824 0 1 66781
box 0 0 1 1
use contact_33  contact_33_79
timestamp 1624857261
transform 1 0 116960 0 1 66373
box 0 0 1 1
use contact_33  contact_33_80
timestamp 1624857261
transform 1 0 116960 0 1 66101
box 0 0 1 1
use contact_33  contact_33_2558
timestamp 1624857261
transform 1 0 116552 0 1 66373
box 0 0 1 1
use contact_33  contact_33_2559
timestamp 1624857261
transform 1 0 116552 0 1 66101
box 0 0 1 1
use contact_33  contact_33_3146
timestamp 1624857261
transform 1 0 115192 0 1 66917
box 0 0 1 1
use contact_33  contact_33_3147
timestamp 1624857261
transform 1 0 115192 0 1 67189
box 0 0 1 1
use contact_33  contact_33_815
timestamp 1624857261
transform 1 0 115600 0 1 66917
box 0 0 1 1
use contact_33  contact_33_816
timestamp 1624857261
transform 1 0 115600 0 1 67189
box 0 0 1 1
use contact_33  contact_33_305
timestamp 1624857261
transform 1 0 116960 0 1 66917
box 0 0 1 1
use contact_33  contact_33_306
timestamp 1624857261
transform 1 0 116960 0 1 67189
box 0 0 1 1
use contact_33  contact_33_365
timestamp 1624857261
transform 1 0 116824 0 1 67325
box 0 0 1 1
use contact_33  contact_33_366
timestamp 1624857261
transform 1 0 116824 0 1 67597
box 0 0 1 1
use contact_33  contact_33_2652
timestamp 1624857261
transform 1 0 116552 0 1 67597
box 0 0 1 1
use contact_33  contact_33_2653
timestamp 1624857261
transform 1 0 116552 0 1 67325
box 0 0 1 1
use contact_33  contact_33_3310
timestamp 1624857261
transform 1 0 115328 0 1 68413
box 0 0 1 1
use contact_33  contact_33_751
timestamp 1624857261
transform 1 0 115736 0 1 68413
box 0 0 1 1
use contact_33  contact_33_2886
timestamp 1624857261
transform 1 0 116008 0 1 68277
box 0 0 1 1
use contact_33  contact_33_2887
timestamp 1624857261
transform 1 0 116008 0 1 68005
box 0 0 1 1
use contact_33  contact_33_350
timestamp 1624857261
transform 1 0 116960 0 1 68549
box 0 0 1 1
use contact_33  contact_33_363
timestamp 1624857261
transform 1 0 116824 0 1 68005
box 0 0 1 1
use contact_33  contact_33_364
timestamp 1624857261
transform 1 0 116824 0 1 67733
box 0 0 1 1
use contact_33  contact_33_3297
timestamp 1624857261
transform 1 0 115192 0 1 69229
box 0 0 1 1
use contact_33  contact_33_3311
timestamp 1624857261
transform 1 0 115328 0 1 68685
box 0 0 1 1
use contact_33  contact_33_3312
timestamp 1624857261
transform 1 0 115328 0 1 69093
box 0 0 1 1
use contact_33  contact_33_3313
timestamp 1624857261
transform 1 0 115328 0 1 68821
box 0 0 1 1
use contact_33  contact_33_731
timestamp 1624857261
transform 1 0 115600 0 1 69229
box 0 0 1 1
use contact_33  contact_33_752
timestamp 1624857261
transform 1 0 115736 0 1 68685
box 0 0 1 1
use contact_33  contact_33_753
timestamp 1624857261
transform 1 0 115736 0 1 69093
box 0 0 1 1
use contact_33  contact_33_754
timestamp 1624857261
transform 1 0 115736 0 1 68821
box 0 0 1 1
use contact_33  contact_33_2870
timestamp 1624857261
transform 1 0 116280 0 1 68821
box 0 0 1 1
use contact_33  contact_33_2871
timestamp 1624857261
transform 1 0 116280 0 1 69093
box 0 0 1 1
use contact_33  contact_33_2873
timestamp 1624857261
transform 1 0 116144 0 1 69229
box 0 0 1 1
use contact_33  contact_33_287
timestamp 1624857261
transform 1 0 116824 0 1 69229
box 0 0 1 1
use contact_33  contact_33_349
timestamp 1624857261
transform 1 0 116960 0 1 68821
box 0 0 1 1
use contact_33  contact_33_3024
timestamp 1624857261
transform 1 0 115192 0 1 69909
box 0 0 1 1
use contact_33  contact_33_3025
timestamp 1624857261
transform 1 0 115192 0 1 69637
box 0 0 1 1
use contact_33  contact_33_3122
timestamp 1624857261
transform 1 0 115192 0 1 70045
box 0 0 1 1
use contact_33  contact_33_3296
timestamp 1624857261
transform 1 0 115192 0 1 69501
box 0 0 1 1
use contact_33  contact_33_632
timestamp 1624857261
transform 1 0 115736 0 1 70045
box 0 0 1 1
use contact_33  contact_33_732
timestamp 1624857261
transform 1 0 115600 0 1 69501
box 0 0 1 1
use contact_33  contact_33_733
timestamp 1624857261
transform 1 0 115600 0 1 69909
box 0 0 1 1
use contact_33  contact_33_734
timestamp 1624857261
transform 1 0 115600 0 1 69637
box 0 0 1 1
use contact_33  contact_33_2868
timestamp 1624857261
transform 1 0 116008 0 1 69909
box 0 0 1 1
use contact_33  contact_33_2869
timestamp 1624857261
transform 1 0 116008 0 1 69637
box 0 0 1 1
use contact_33  contact_33_2872
timestamp 1624857261
transform 1 0 116144 0 1 69501
box 0 0 1 1
use contact_33  contact_33_2982
timestamp 1624857261
transform 1 0 116144 0 1 70045
box 0 0 1 1
use contact_33  contact_33_197
timestamp 1624857261
transform 1 0 116960 0 1 70045
box 0 0 1 1
use contact_33  contact_33_288
timestamp 1624857261
transform 1 0 116824 0 1 69501
box 0 0 1 1
use contact_33  contact_33_2546
timestamp 1624857261
transform 1 0 116552 0 1 69909
box 0 0 1 1
use contact_33  contact_33_2547
timestamp 1624857261
transform 1 0 116552 0 1 69637
box 0 0 1 1
use contact_33  contact_33_3123
timestamp 1624857261
transform 1 0 115192 0 1 70317
box 0 0 1 1
use contact_33  contact_33_3124
timestamp 1624857261
transform 1 0 115192 0 1 70725
box 0 0 1 1
use contact_33  contact_33_3125
timestamp 1624857261
transform 1 0 115192 0 1 70453
box 0 0 1 1
use contact_33  contact_33_3226
timestamp 1624857261
transform 1 0 115328 0 1 70861
box 0 0 1 1
use contact_33  contact_33_3227
timestamp 1624857261
transform 1 0 115328 0 1 71133
box 0 0 1 1
use contact_33  contact_33_579
timestamp 1624857261
transform 1 0 115600 0 1 70725
box 0 0 1 1
use contact_33  contact_33_580
timestamp 1624857261
transform 1 0 115600 0 1 70453
box 0 0 1 1
use contact_33  contact_33_631
timestamp 1624857261
transform 1 0 115736 0 1 70317
box 0 0 1 1
use contact_33  contact_33_661
timestamp 1624857261
transform 1 0 115736 0 1 70861
box 0 0 1 1
use contact_33  contact_33_662
timestamp 1624857261
transform 1 0 115736 0 1 71133
box 0 0 1 1
use contact_33  contact_33_2784
timestamp 1624857261
transform 1 0 116280 0 1 71133
box 0 0 1 1
use contact_33  contact_33_2785
timestamp 1624857261
transform 1 0 116280 0 1 70861
box 0 0 1 1
use contact_33  contact_33_2983
timestamp 1624857261
transform 1 0 116144 0 1 70317
box 0 0 1 1
use contact_33  contact_33_198
timestamp 1624857261
transform 1 0 116960 0 1 70317
box 0 0 1 1
use contact_33  contact_33_209
timestamp 1624857261
transform 1 0 116960 0 1 70453
box 0 0 1 1
use contact_33  contact_33_210
timestamp 1624857261
transform 1 0 116960 0 1 70725
box 0 0 1 1
use contact_33  contact_33_433
timestamp 1624857261
transform 1 0 116824 0 1 70861
box 0 0 1 1
use contact_33  contact_33_434
timestamp 1624857261
transform 1 0 116824 0 1 71133
box 0 0 1 1
use contact_33  contact_33_2536
timestamp 1624857261
transform 1 0 116552 0 1 70725
box 0 0 1 1
use contact_33  contact_33_2537
timestamp 1624857261
transform 1 0 116552 0 1 70453
box 0 0 1 1
use contact_33  contact_33_3290
timestamp 1624857261
transform 1 0 115192 0 1 71269
box 0 0 1 1
use contact_33  contact_33_3291
timestamp 1624857261
transform 1 0 115192 0 1 71541
box 0 0 1 1
use contact_33  contact_33_663
timestamp 1624857261
transform 1 0 115736 0 1 71541
box 0 0 1 1
use contact_33  contact_33_664
timestamp 1624857261
transform 1 0 115736 0 1 71269
box 0 0 1 1
use contact_33  contact_33_2708
timestamp 1624857261
transform 1 0 116280 0 1 71269
box 0 0 1 1
use contact_33  contact_33_2709
timestamp 1624857261
transform 1 0 116280 0 1 71541
box 0 0 1 1
use contact_33  contact_33_3016
timestamp 1624857261
transform 1 0 116008 0 1 71541
box 0 0 1 1
use contact_33  contact_33_3017
timestamp 1624857261
transform 1 0 116008 0 1 71269
box 0 0 1 1
use contact_33  contact_33_159
timestamp 1624857261
transform 1 0 116824 0 1 71677
box 0 0 1 1
use contact_33  contact_33_160
timestamp 1624857261
transform 1 0 116824 0 1 71949
box 0 0 1 1
use contact_33  contact_33_431
timestamp 1624857261
transform 1 0 116824 0 1 71541
box 0 0 1 1
use contact_33  contact_33_432
timestamp 1624857261
transform 1 0 116824 0 1 71269
box 0 0 1 1
use contact_33  contact_33_3034
timestamp 1624857261
transform 1 0 115328 0 1 72765
box 0 0 1 1
use contact_33  contact_33_737
timestamp 1624857261
transform 1 0 115736 0 1 72765
box 0 0 1 1
use contact_33  contact_33_2867
timestamp 1624857261
transform 1 0 116008 0 1 72765
box 0 0 1 1
use contact_33  contact_33_3004
timestamp 1624857261
transform 1 0 116008 0 1 72085
box 0 0 1 1
use contact_33  contact_33_3005
timestamp 1624857261
transform 1 0 116008 0 1 72357
box 0 0 1 1
use contact_33  contact_33_249
timestamp 1624857261
transform 1 0 116824 0 1 72085
box 0 0 1 1
use contact_33  contact_33_250
timestamp 1624857261
transform 1 0 116824 0 1 72357
box 0 0 1 1
use contact_33  contact_33_443
timestamp 1624857261
transform 1 0 116960 0 1 72493
box 0 0 1 1
use contact_33  contact_33_444
timestamp 1624857261
transform 1 0 116960 0 1 72765
box 0 0 1 1
use contact_33  contact_33_2606
timestamp 1624857261
transform 1 0 116416 0 1 72765
box 0 0 1 1
use contact_33  contact_33_3035
timestamp 1624857261
transform 1 0 115328 0 1 73037
box 0 0 1 1
use contact_33  contact_33_3336
timestamp 1624857261
transform 1 0 115328 0 1 73173
box 0 0 1 1
use contact_33  contact_33_3337
timestamp 1624857261
transform 1 0 115328 0 1 73445
box 0 0 1 1
use contact_33  contact_33_3339
timestamp 1624857261
transform 1 0 115192 0 1 73581
box 0 0 1 1
use contact_33  contact_33_567
timestamp 1624857261
transform 1 0 115600 0 1 73581
box 0 0 1 1
use contact_33  contact_33_735
timestamp 1624857261
transform 1 0 115736 0 1 73445
box 0 0 1 1
use contact_33  contact_33_736
timestamp 1624857261
transform 1 0 115736 0 1 73173
box 0 0 1 1
use contact_33  contact_33_738
timestamp 1624857261
transform 1 0 115736 0 1 73037
box 0 0 1 1
use contact_33  contact_33_2866
timestamp 1624857261
transform 1 0 116008 0 1 73037
box 0 0 1 1
use contact_33  contact_33_2948
timestamp 1624857261
transform 1 0 116008 0 1 73173
box 0 0 1 1
use contact_33  contact_33_2949
timestamp 1624857261
transform 1 0 116008 0 1 73445
box 0 0 1 1
use contact_33  contact_33_2951
timestamp 1624857261
transform 1 0 116144 0 1 73581
box 0 0 1 1
use contact_33  contact_33_161
timestamp 1624857261
transform 1 0 116824 0 1 73445
box 0 0 1 1
use contact_33  contact_33_162
timestamp 1624857261
transform 1 0 116824 0 1 73173
box 0 0 1 1
use contact_33  contact_33_2607
timestamp 1624857261
transform 1 0 116416 0 1 73037
box 0 0 1 1
use contact_33  contact_33_3207
timestamp 1624857261
transform 1 0 115192 0 1 73989
box 0 0 1 1
use contact_33  contact_33_3338
timestamp 1624857261
transform 1 0 115192 0 1 73853
box 0 0 1 1
use contact_33  contact_33_568
timestamp 1624857261
transform 1 0 115600 0 1 73853
box 0 0 1 1
use contact_33  contact_33_570
timestamp 1624857261
transform 1 0 115600 0 1 73989
box 0 0 1 1
use contact_33  contact_33_2860
timestamp 1624857261
transform 1 0 116008 0 1 73989
box 0 0 1 1
use contact_33  contact_33_2950
timestamp 1624857261
transform 1 0 116144 0 1 73853
box 0 0 1 1
use contact_33  contact_33_104
timestamp 1624857261
transform 1 0 116960 0 1 73989
box 0 0 1 1
use cr_5  cr_5_0
timestamp 1624857261
transform 1 0 15406 0 1 9422
box 61024 65420 64083 68762
use contact_33  contact_33_891
timestamp 1624857261
transform 1 0 110432 0 1 76845
box 0 0 1 1
use contact_33  contact_33_892
timestamp 1624857261
transform 1 0 110432 0 1 76573
box 0 0 1 1
use contact_33  contact_33_893
timestamp 1624857261
transform 1 0 110296 0 1 76165
box 0 0 1 1
use contact_33  contact_33_894
timestamp 1624857261
transform 1 0 110296 0 1 76437
box 0 0 1 1
use contact_33  contact_33_856
timestamp 1624857261
transform 1 0 110432 0 1 80109
box 0 0 1 1
use contact_33  contact_33_881
timestamp 1624857261
transform 1 0 110432 0 1 77661
box 0 0 1 1
use contact_33  contact_33_882
timestamp 1624857261
transform 1 0 110432 0 1 77389
box 0 0 1 1
use contact_33  contact_33_903
timestamp 1624857261
transform 1 0 110160 0 1 79973
box 0 0 1 1
use contact_33  contact_33_904
timestamp 1624857261
transform 1 0 110160 0 1 79701
box 0 0 1 1
use contact_33  contact_33_855
timestamp 1624857261
transform 1 0 110432 0 1 80381
box 0 0 1 1
use contact_33  contact_33_861
timestamp 1624857261
transform 1 0 110160 0 1 84325
box 0 0 1 1
use contact_33  contact_33_862
timestamp 1624857261
transform 1 0 110160 0 1 84053
box 0 0 1 1
use contact_33  contact_33_955
timestamp 1624857261
transform 1 0 110160 0 1 85277
box 0 0 1 1
use contact_33  contact_33_956
timestamp 1624857261
transform 1 0 110160 0 1 85549
box 0 0 1 1
use contact_33  contact_33_853
timestamp 1624857261
transform 1 0 110160 0 1 88677
box 0 0 1 1
use contact_33  contact_33_854
timestamp 1624857261
transform 1 0 110160 0 1 88949
box 0 0 1 1
use contact_33  contact_33_869
timestamp 1624857261
transform 1 0 110296 0 1 88405
box 0 0 1 1
use contact_33  contact_33_870
timestamp 1624857261
transform 1 0 110296 0 1 88677
box 0 0 1 1
use contact_33  contact_33_915
timestamp 1624857261
transform 1 0 110432 0 1 88405
box 0 0 1 1
use contact_33  contact_33_916
timestamp 1624857261
transform 1 0 110432 0 1 88133
box 0 0 1 1
use contact_33  contact_33_857
timestamp 1624857261
transform 1 0 110432 0 1 91805
box 0 0 1 1
use contact_33  contact_33_858
timestamp 1624857261
transform 1 0 110432 0 1 91533
box 0 0 1 1
use contact_33  contact_33_947
timestamp 1624857261
transform 1 0 110296 0 1 92349
box 0 0 1 1
use contact_33  contact_33_948
timestamp 1624857261
transform 1 0 110296 0 1 92621
box 0 0 1 1
use contact_33  contact_33_3206
timestamp 1624857261
transform 1 0 115192 0 1 74261
box 0 0 1 1
use contact_33  contact_33_3326
timestamp 1624857261
transform 1 0 115192 0 1 74397
box 0 0 1 1
use contact_33  contact_33_3327
timestamp 1624857261
transform 1 0 115192 0 1 74669
box 0 0 1 1
use contact_33  contact_33_3329
timestamp 1624857261
transform 1 0 115192 0 1 74805
box 0 0 1 1
use contact_33  contact_33_569
timestamp 1624857261
transform 1 0 115600 0 1 74261
box 0 0 1 1
use contact_33  contact_33_653
timestamp 1624857261
transform 1 0 115600 0 1 74397
box 0 0 1 1
use contact_33  contact_33_654
timestamp 1624857261
transform 1 0 115600 0 1 74669
box 0 0 1 1
use contact_33  contact_33_656
timestamp 1624857261
transform 1 0 115600 0 1 74805
box 0 0 1 1
use contact_33  contact_33_2858
timestamp 1624857261
transform 1 0 116008 0 1 74669
box 0 0 1 1
use contact_33  contact_33_2859
timestamp 1624857261
transform 1 0 116008 0 1 74397
box 0 0 1 1
use contact_33  contact_33_2861
timestamp 1624857261
transform 1 0 116008 0 1 74261
box 0 0 1 1
use contact_33  contact_33_103
timestamp 1624857261
transform 1 0 116960 0 1 74261
box 0 0 1 1
use contact_33  contact_33_373
timestamp 1624857261
transform 1 0 116960 0 1 74397
box 0 0 1 1
use contact_33  contact_33_374
timestamp 1624857261
transform 1 0 116960 0 1 74669
box 0 0 1 1
use contact_33  contact_33_376
timestamp 1624857261
transform 1 0 116960 0 1 74805
box 0 0 1 1
use contact_33  contact_33_2573
timestamp 1624857261
transform 1 0 116552 0 1 74805
box 0 0 1 1
use contact_33  contact_33_3328
timestamp 1624857261
transform 1 0 115192 0 1 75077
box 0 0 1 1
use contact_33  contact_33_3330
timestamp 1624857261
transform 1 0 115328 0 1 75213
box 0 0 1 1
use contact_33  contact_33_3331
timestamp 1624857261
transform 1 0 115328 0 1 75485
box 0 0 1 1
use contact_33  contact_33_619
timestamp 1624857261
transform 1 0 115736 0 1 75213
box 0 0 1 1
use contact_33  contact_33_620
timestamp 1624857261
transform 1 0 115736 0 1 75485
box 0 0 1 1
use contact_33  contact_33_655
timestamp 1624857261
transform 1 0 115600 0 1 75077
box 0 0 1 1
use contact_33  contact_33_2926
timestamp 1624857261
transform 1 0 116144 0 1 75485
box 0 0 1 1
use contact_33  contact_33_2927
timestamp 1624857261
transform 1 0 116144 0 1 75213
box 0 0 1 1
use contact_33  contact_33_375
timestamp 1624857261
transform 1 0 116960 0 1 75077
box 0 0 1 1
use contact_33  contact_33_419
timestamp 1624857261
transform 1 0 116824 0 1 75213
box 0 0 1 1
use contact_33  contact_33_420
timestamp 1624857261
transform 1 0 116824 0 1 75485
box 0 0 1 1
use contact_33  contact_33_422
timestamp 1624857261
transform 1 0 116824 0 1 75621
box 0 0 1 1
use contact_33  contact_33_2572
timestamp 1624857261
transform 1 0 116552 0 1 75077
box 0 0 1 1
use contact_33  contact_33_2666
timestamp 1624857261
transform 1 0 116416 0 1 75213
box 0 0 1 1
use contact_33  contact_33_2667
timestamp 1624857261
transform 1 0 116416 0 1 75485
box 0 0 1 1
use contact_33  contact_33_3063
timestamp 1624857261
transform 1 0 115328 0 1 76709
box 0 0 1 1
use contact_33  contact_33_712
timestamp 1624857261
transform 1 0 115736 0 1 76709
box 0 0 1 1
use contact_33  contact_33_2763
timestamp 1624857261
transform 1 0 116008 0 1 76709
box 0 0 1 1
use contact_33  contact_33_2954
timestamp 1624857261
transform 1 0 116144 0 1 76029
box 0 0 1 1
use contact_33  contact_33_2955
timestamp 1624857261
transform 1 0 116144 0 1 76301
box 0 0 1 1
use contact_33  contact_33_121
timestamp 1624857261
transform 1 0 116824 0 1 76709
box 0 0 1 1
use contact_33  contact_33_122
timestamp 1624857261
transform 1 0 116824 0 1 76437
box 0 0 1 1
use contact_33  contact_33_299
timestamp 1624857261
transform 1 0 116960 0 1 76301
box 0 0 1 1
use contact_33  contact_33_300
timestamp 1624857261
transform 1 0 116960 0 1 76029
box 0 0 1 1
use contact_33  contact_33_421
timestamp 1624857261
transform 1 0 116824 0 1 75893
box 0 0 1 1
use contact_33  contact_33_2680
timestamp 1624857261
transform 1 0 116552 0 1 76301
box 0 0 1 1
use contact_33  contact_33_2681
timestamp 1624857261
transform 1 0 116552 0 1 76029
box 0 0 1 1
use contact_33  contact_33_3044
timestamp 1624857261
transform 1 0 115328 0 1 77117
box 0 0 1 1
use contact_33  contact_33_3045
timestamp 1624857261
transform 1 0 115328 0 1 77389
box 0 0 1 1
use contact_33  contact_33_3062
timestamp 1624857261
transform 1 0 115328 0 1 76981
box 0 0 1 1
use contact_33  contact_33_3142
timestamp 1624857261
transform 1 0 115328 0 1 77525
box 0 0 1 1
use contact_33  contact_33_571
timestamp 1624857261
transform 1 0 115600 0 1 77389
box 0 0 1 1
use contact_33  contact_33_572
timestamp 1624857261
transform 1 0 115600 0 1 77117
box 0 0 1 1
use contact_33  contact_33_679
timestamp 1624857261
transform 1 0 115736 0 1 77525
box 0 0 1 1
use contact_33  contact_33_711
timestamp 1624857261
transform 1 0 115736 0 1 76981
box 0 0 1 1
use contact_33  contact_33_2762
timestamp 1624857261
transform 1 0 116008 0 1 76981
box 0 0 1 1
use contact_33  contact_33_2714
timestamp 1624857261
transform 1 0 116280 0 1 77525
box 0 0 1 1
use contact_33  contact_33_3143
timestamp 1624857261
transform 1 0 115328 0 1 77797
box 0 0 1 1
use contact_33  contact_33_3144
timestamp 1624857261
transform 1 0 115328 0 1 78205
box 0 0 1 1
use contact_33  contact_33_3145
timestamp 1624857261
transform 1 0 115328 0 1 77933
box 0 0 1 1
use contact_33  contact_33_3232
timestamp 1624857261
transform 1 0 115328 0 1 78341
box 0 0 1 1
use contact_33  contact_33_680
timestamp 1624857261
transform 1 0 115736 0 1 77797
box 0 0 1 1
use contact_33  contact_33_681
timestamp 1624857261
transform 1 0 115600 0 1 78205
box 0 0 1 1
use contact_33  contact_33_682
timestamp 1624857261
transform 1 0 115600 0 1 77933
box 0 0 1 1
use contact_33  contact_33_739
timestamp 1624857261
transform 1 0 115736 0 1 78341
box 0 0 1 1
use contact_33  contact_33_2944
timestamp 1624857261
transform 1 0 116008 0 1 77933
box 0 0 1 1
use contact_33  contact_33_2945
timestamp 1624857261
transform 1 0 116008 0 1 78205
box 0 0 1 1
use contact_33  contact_33_2947
timestamp 1624857261
transform 1 0 116008 0 1 78341
box 0 0 1 1
use contact_33  contact_33_82
timestamp 1624857261
transform 1 0 116960 0 1 78341
box 0 0 1 1
use contact_33  contact_33_315
timestamp 1624857261
transform 1 0 116960 0 1 78205
box 0 0 1 1
use contact_33  contact_33_316
timestamp 1624857261
transform 1 0 116960 0 1 77933
box 0 0 1 1
use contact_33  contact_33_2715
timestamp 1624857261
transform 1 0 116280 0 1 77797
box 0 0 1 1
use contact_33  contact_33_3233
timestamp 1624857261
transform 1 0 115328 0 1 78613
box 0 0 1 1
use contact_33  contact_33_3355
timestamp 1624857261
transform 1 0 115192 0 1 79157
box 0 0 1 1
use contact_33  contact_33_3356
timestamp 1624857261
transform 1 0 115192 0 1 78749
box 0 0 1 1
use contact_33  contact_33_3357
timestamp 1624857261
transform 1 0 115192 0 1 79021
box 0 0 1 1
use contact_33  contact_33_610
timestamp 1624857261
transform 1 0 115600 0 1 79157
box 0 0 1 1
use contact_33  contact_33_740
timestamp 1624857261
transform 1 0 115736 0 1 78613
box 0 0 1 1
use contact_33  contact_33_741
timestamp 1624857261
transform 1 0 115736 0 1 79021
box 0 0 1 1
use contact_33  contact_33_742
timestamp 1624857261
transform 1 0 115736 0 1 78749
box 0 0 1 1
use contact_33  contact_33_2908
timestamp 1624857261
transform 1 0 116008 0 1 79021
box 0 0 1 1
use contact_33  contact_33_2909
timestamp 1624857261
transform 1 0 116008 0 1 78749
box 0 0 1 1
use contact_33  contact_33_2946
timestamp 1624857261
transform 1 0 116008 0 1 78613
box 0 0 1 1
use contact_33  contact_33_77
timestamp 1624857261
transform 1 0 116960 0 1 78749
box 0 0 1 1
use contact_33  contact_33_78
timestamp 1624857261
transform 1 0 116960 0 1 79021
box 0 0 1 1
use contact_33  contact_33_81
timestamp 1624857261
transform 1 0 116960 0 1 78613
box 0 0 1 1
use contact_33  contact_33_409
timestamp 1624857261
transform 1 0 116960 0 1 79157
box 0 0 1 1
use contact_33  contact_33_2661
timestamp 1624857261
transform 1 0 116552 0 1 79157
box 0 0 1 1
use contact_33  contact_33_3262
timestamp 1624857261
transform 1 0 115328 0 1 79565
box 0 0 1 1
use contact_33  contact_33_3263
timestamp 1624857261
transform 1 0 115328 0 1 79837
box 0 0 1 1
use contact_33  contact_33_3354
timestamp 1624857261
transform 1 0 115192 0 1 79429
box 0 0 1 1
use contact_33  contact_33_609
timestamp 1624857261
transform 1 0 115600 0 1 79429
box 0 0 1 1
use contact_33  contact_33_723
timestamp 1624857261
transform 1 0 115736 0 1 79565
box 0 0 1 1
use contact_33  contact_33_724
timestamp 1624857261
transform 1 0 115736 0 1 79837
box 0 0 1 1
use contact_33  contact_33_2824
timestamp 1624857261
transform 1 0 116008 0 1 79973
box 0 0 1 1
use contact_33  contact_33_186
timestamp 1624857261
transform 1 0 116824 0 1 79973
box 0 0 1 1
use contact_33  contact_33_410
timestamp 1624857261
transform 1 0 116960 0 1 79429
box 0 0 1 1
use contact_33  contact_33_411
timestamp 1624857261
transform 1 0 116824 0 1 79837
box 0 0 1 1
use contact_33  contact_33_412
timestamp 1624857261
transform 1 0 116824 0 1 79565
box 0 0 1 1
use contact_33  contact_33_2660
timestamp 1624857261
transform 1 0 116552 0 1 79429
box 0 0 1 1
use contact_33  contact_33_2720
timestamp 1624857261
transform 1 0 116280 0 1 79701
box 0 0 1 1
use contact_33  contact_33_2721
timestamp 1624857261
transform 1 0 116280 0 1 79429
box 0 0 1 1
use contact_33  contact_33_2822
timestamp 1624857261
transform 1 0 116280 0 1 79973
box 0 0 1 1
use contact_33  contact_33_2825
timestamp 1624857261
transform 1 0 116008 0 1 80245
box 0 0 1 1
use contact_33  contact_33_2912
timestamp 1624857261
transform 1 0 116144 0 1 80925
box 0 0 1 1
use contact_33  contact_33_2913
timestamp 1624857261
transform 1 0 116144 0 1 80653
box 0 0 1 1
use contact_33  contact_33_185
timestamp 1624857261
transform 1 0 116824 0 1 80245
box 0 0 1 1
use contact_33  contact_33_233
timestamp 1624857261
transform 1 0 116824 0 1 80381
box 0 0 1 1
use contact_33  contact_33_234
timestamp 1624857261
transform 1 0 116824 0 1 80653
box 0 0 1 1
use contact_33  contact_33_2823
timestamp 1624857261
transform 1 0 116280 0 1 80245
box 0 0 1 1
use contact_33  contact_33_3302
timestamp 1624857261
transform 1 0 115192 0 1 81061
box 0 0 1 1
use contact_33  contact_33_3303
timestamp 1624857261
transform 1 0 115192 0 1 81333
box 0 0 1 1
use contact_33  contact_33_3304
timestamp 1624857261
transform 1 0 115192 0 1 81741
box 0 0 1 1
use contact_33  contact_33_3305
timestamp 1624857261
transform 1 0 115192 0 1 81469
box 0 0 1 1
use contact_33  contact_33_697
timestamp 1624857261
transform 1 0 115600 0 1 81061
box 0 0 1 1
use contact_33  contact_33_698
timestamp 1624857261
transform 1 0 115600 0 1 81333
box 0 0 1 1
use contact_33  contact_33_699
timestamp 1624857261
transform 1 0 115600 0 1 81741
box 0 0 1 1
use contact_33  contact_33_700
timestamp 1624857261
transform 1 0 115600 0 1 81469
box 0 0 1 1
use contact_33  contact_33_2768
timestamp 1624857261
transform 1 0 116280 0 1 81469
box 0 0 1 1
use contact_33  contact_33_2769
timestamp 1624857261
transform 1 0 116280 0 1 81741
box 0 0 1 1
use contact_33  contact_33_3070
timestamp 1624857261
transform 1 0 115328 0 1 82149
box 0 0 1 1
use contact_33  contact_33_3071
timestamp 1624857261
transform 1 0 115328 0 1 81877
box 0 0 1 1
use contact_33  contact_33_3342
timestamp 1624857261
transform 1 0 115192 0 1 82285
box 0 0 1 1
use contact_33  contact_33_3343
timestamp 1624857261
transform 1 0 115192 0 1 82557
box 0 0 1 1
use contact_33  contact_33_559
timestamp 1624857261
transform 1 0 115600 0 1 82557
box 0 0 1 1
use contact_33  contact_33_560
timestamp 1624857261
transform 1 0 115600 0 1 82285
box 0 0 1 1
use contact_33  contact_33_561
timestamp 1624857261
transform 1 0 115736 0 1 81877
box 0 0 1 1
use contact_33  contact_33_562
timestamp 1624857261
transform 1 0 115736 0 1 82149
box 0 0 1 1
use contact_33  contact_33_2810
timestamp 1624857261
transform 1 0 116008 0 1 81877
box 0 0 1 1
use contact_33  contact_33_2811
timestamp 1624857261
transform 1 0 116008 0 1 82149
box 0 0 1 1
use contact_33  contact_33_2992
timestamp 1624857261
transform 1 0 116008 0 1 82285
box 0 0 1 1
use contact_33  contact_33_2993
timestamp 1624857261
transform 1 0 116008 0 1 82557
box 0 0 1 1
use contact_33  contact_33_101
timestamp 1624857261
transform 1 0 116824 0 1 81877
box 0 0 1 1
use contact_33  contact_33_102
timestamp 1624857261
transform 1 0 116824 0 1 82149
box 0 0 1 1
use contact_33  contact_33_129
timestamp 1624857261
transform 1 0 116960 0 1 82285
box 0 0 1 1
use contact_33  contact_33_130
timestamp 1624857261
transform 1 0 116960 0 1 82557
box 0 0 1 1
use contact_33  contact_33_2636
timestamp 1624857261
transform 1 0 116416 0 1 81877
box 0 0 1 1
use contact_33  contact_33_2637
timestamp 1624857261
transform 1 0 116416 0 1 82149
box 0 0 1 1
use contact_33  contact_33_3032
timestamp 1624857261
transform 1 0 115192 0 1 83101
box 0 0 1 1
use contact_33  contact_33_3033
timestamp 1624857261
transform 1 0 115192 0 1 83373
box 0 0 1 1
use contact_33  contact_33_3340
timestamp 1624857261
transform 1 0 115192 0 1 82965
box 0 0 1 1
use contact_33  contact_33_3341
timestamp 1624857261
transform 1 0 115192 0 1 82693
box 0 0 1 1
use contact_33  contact_33_773
timestamp 1624857261
transform 1 0 115736 0 1 83373
box 0 0 1 1
use contact_33  contact_33_774
timestamp 1624857261
transform 1 0 115736 0 1 83101
box 0 0 1 1
use contact_33  contact_33_775
timestamp 1624857261
transform 1 0 115736 0 1 82693
box 0 0 1 1
use contact_33  contact_33_776
timestamp 1624857261
transform 1 0 115736 0 1 82965
box 0 0 1 1
use contact_33  contact_33_2850
timestamp 1624857261
transform 1 0 116008 0 1 83373
box 0 0 1 1
use contact_33  contact_33_2851
timestamp 1624857261
transform 1 0 116008 0 1 83101
box 0 0 1 1
use contact_33  contact_33_2994
timestamp 1624857261
transform 1 0 116008 0 1 82965
box 0 0 1 1
use contact_33  contact_33_2995
timestamp 1624857261
transform 1 0 116008 0 1 82693
box 0 0 1 1
use contact_33  contact_33_183
timestamp 1624857261
transform 1 0 116824 0 1 82693
box 0 0 1 1
use contact_33  contact_33_184
timestamp 1624857261
transform 1 0 116824 0 1 82965
box 0 0 1 1
use contact_33  contact_33_309
timestamp 1624857261
transform 1 0 116960 0 1 83101
box 0 0 1 1
use contact_33  contact_33_310
timestamp 1624857261
transform 1 0 116960 0 1 83373
box 0 0 1 1
use contact_33  contact_33_2632
timestamp 1624857261
transform 1 0 116416 0 1 83373
box 0 0 1 1
use contact_33  contact_33_2633
timestamp 1624857261
transform 1 0 116416 0 1 83101
box 0 0 1 1
use contact_33  contact_33_3358
timestamp 1624857261
transform 1 0 115192 0 1 83509
box 0 0 1 1
use contact_33  contact_33_3359
timestamp 1624857261
transform 1 0 115192 0 1 83781
box 0 0 1 1
use contact_33  contact_33_795
timestamp 1624857261
transform 1 0 115600 0 1 83509
box 0 0 1 1
use contact_33  contact_33_796
timestamp 1624857261
transform 1 0 115600 0 1 83781
box 0 0 1 1
use contact_33  contact_33_83
timestamp 1624857261
transform 1 0 116824 0 1 83917
box 0 0 1 1
use contact_33  contact_33_84
timestamp 1624857261
transform 1 0 116824 0 1 84189
box 0 0 1 1
use contact_33  contact_33_201
timestamp 1624857261
transform 1 0 116960 0 1 84325
box 0 0 1 1
use contact_33  contact_33_307
timestamp 1624857261
transform 1 0 116960 0 1 83781
box 0 0 1 1
use contact_33  contact_33_308
timestamp 1624857261
transform 1 0 116960 0 1 83509
box 0 0 1 1
use contact_33  contact_33_3157
timestamp 1624857261
transform 1 0 115328 0 1 85005
box 0 0 1 1
use contact_33  contact_33_669
timestamp 1624857261
transform 1 0 115736 0 1 85005
box 0 0 1 1
use contact_33  contact_33_202
timestamp 1624857261
transform 1 0 116960 0 1 84597
box 0 0 1 1
use contact_33  contact_33_426
timestamp 1624857261
transform 1 0 116960 0 1 85141
box 0 0 1 1
use contact_33  contact_33_2560
timestamp 1624857261
transform 1 0 116552 0 1 84869
box 0 0 1 1
use contact_33  contact_33_2561
timestamp 1624857261
transform 1 0 116552 0 1 84597
box 0 0 1 1
use contact_33  contact_33_3072
timestamp 1624857261
transform 1 0 115328 0 1 85821
box 0 0 1 1
use contact_33  contact_33_3100
timestamp 1624857261
transform 1 0 115328 0 1 85685
box 0 0 1 1
use contact_33  contact_33_3101
timestamp 1624857261
transform 1 0 115328 0 1 85413
box 0 0 1 1
use contact_33  contact_33_3156
timestamp 1624857261
transform 1 0 115328 0 1 85277
box 0 0 1 1
use contact_33  contact_33_670
timestamp 1624857261
transform 1 0 115736 0 1 85277
box 0 0 1 1
use contact_33  contact_33_818
timestamp 1624857261
transform 1 0 115600 0 1 85821
box 0 0 1 1
use contact_33  contact_33_819
timestamp 1624857261
transform 1 0 115600 0 1 85413
box 0 0 1 1
use contact_33  contact_33_820
timestamp 1624857261
transform 1 0 115600 0 1 85685
box 0 0 1 1
use contact_33  contact_33_2820
timestamp 1624857261
transform 1 0 116008 0 1 85685
box 0 0 1 1
use contact_33  contact_33_2821
timestamp 1624857261
transform 1 0 116008 0 1 85413
box 0 0 1 1
use contact_33  contact_33_325
timestamp 1624857261
transform 1 0 116824 0 1 85821
box 0 0 1 1
use contact_33  contact_33_425
timestamp 1624857261
transform 1 0 116960 0 1 85413
box 0 0 1 1
use contact_33  contact_33_3073
timestamp 1624857261
transform 1 0 115328 0 1 86093
box 0 0 1 1
use contact_33  contact_33_3074
timestamp 1624857261
transform 1 0 115328 0 1 86501
box 0 0 1 1
use contact_33  contact_33_3075
timestamp 1624857261
transform 1 0 115328 0 1 86229
box 0 0 1 1
use contact_33  contact_33_3314
timestamp 1624857261
transform 1 0 115192 0 1 86637
box 0 0 1 1
use contact_33  contact_33_564
timestamp 1624857261
transform 1 0 115600 0 1 86637
box 0 0 1 1
use contact_33  contact_33_565
timestamp 1624857261
transform 1 0 115736 0 1 86229
box 0 0 1 1
use contact_33  contact_33_566
timestamp 1624857261
transform 1 0 115736 0 1 86501
box 0 0 1 1
use contact_33  contact_33_817
timestamp 1624857261
transform 1 0 115600 0 1 86093
box 0 0 1 1
use contact_33  contact_33_2996
timestamp 1624857261
transform 1 0 116008 0 1 86229
box 0 0 1 1
use contact_33  contact_33_2997
timestamp 1624857261
transform 1 0 116008 0 1 86501
box 0 0 1 1
use contact_33  contact_33_2999
timestamp 1624857261
transform 1 0 116144 0 1 86637
box 0 0 1 1
use contact_33  contact_33_326
timestamp 1624857261
transform 1 0 116824 0 1 86093
box 0 0 1 1
use contact_33  contact_33_327
timestamp 1624857261
transform 1 0 116824 0 1 86501
box 0 0 1 1
use contact_33  contact_33_328
timestamp 1624857261
transform 1 0 116824 0 1 86229
box 0 0 1 1
use contact_33  contact_33_437
timestamp 1624857261
transform 1 0 116960 0 1 86637
box 0 0 1 1
use contact_33  contact_33_2654
timestamp 1624857261
transform 1 0 116416 0 1 86229
box 0 0 1 1
use contact_33  contact_33_2655
timestamp 1624857261
transform 1 0 116416 0 1 86501
box 0 0 1 1
use contact_33  contact_33_3309
timestamp 1624857261
transform 1 0 115328 0 1 87453
box 0 0 1 1
use contact_33  contact_33_3315
timestamp 1624857261
transform 1 0 115192 0 1 86909
box 0 0 1 1
use contact_33  contact_33_3316
timestamp 1624857261
transform 1 0 115192 0 1 87317
box 0 0 1 1
use contact_33  contact_33_3317
timestamp 1624857261
transform 1 0 115192 0 1 87045
box 0 0 1 1
use contact_33  contact_33_502
timestamp 1624857261
transform 1 0 115736 0 1 87453
box 0 0 1 1
use contact_33  contact_33_503
timestamp 1624857261
transform 1 0 115736 0 1 87045
box 0 0 1 1
use contact_33  contact_33_504
timestamp 1624857261
transform 1 0 115736 0 1 87317
box 0 0 1 1
use contact_33  contact_33_563
timestamp 1624857261
transform 1 0 115600 0 1 86909
box 0 0 1 1
use contact_33  contact_33_2878
timestamp 1624857261
transform 1 0 116144 0 1 87453
box 0 0 1 1
use contact_33  contact_33_2900
timestamp 1624857261
transform 1 0 116008 0 1 87317
box 0 0 1 1
use contact_33  contact_33_2901
timestamp 1624857261
transform 1 0 116008 0 1 87045
box 0 0 1 1
use contact_33  contact_33_2998
timestamp 1624857261
transform 1 0 116144 0 1 86909
box 0 0 1 1
use contact_33  contact_33_415
timestamp 1624857261
transform 1 0 116960 0 1 87453
box 0 0 1 1
use contact_33  contact_33_435
timestamp 1624857261
transform 1 0 116960 0 1 87317
box 0 0 1 1
use contact_33  contact_33_436
timestamp 1624857261
transform 1 0 116960 0 1 87045
box 0 0 1 1
use contact_33  contact_33_438
timestamp 1624857261
transform 1 0 116960 0 1 86909
box 0 0 1 1
use contact_33  contact_33_2583
timestamp 1624857261
transform 1 0 116416 0 1 87453
box 0 0 1 1
use contact_33  contact_33_2700
timestamp 1624857261
transform 1 0 116280 0 1 87045
box 0 0 1 1
use contact_33  contact_33_2701
timestamp 1624857261
transform 1 0 116280 0 1 87317
box 0 0 1 1
use contact_33  contact_33_2703
timestamp 1624857261
transform 1 0 116280 0 1 87453
box 0 0 1 1
use contact_33  contact_33_3288
timestamp 1624857261
transform 1 0 115192 0 1 88133
box 0 0 1 1
use contact_33  contact_33_3289
timestamp 1624857261
transform 1 0 115192 0 1 87861
box 0 0 1 1
use contact_33  contact_33_3308
timestamp 1624857261
transform 1 0 115328 0 1 87725
box 0 0 1 1
use contact_33  contact_33_501
timestamp 1624857261
transform 1 0 115736 0 1 87725
box 0 0 1 1
use contact_33  contact_33_511
timestamp 1624857261
transform 1 0 115600 0 1 87861
box 0 0 1 1
use contact_33  contact_33_512
timestamp 1624857261
transform 1 0 115600 0 1 88133
box 0 0 1 1
use contact_33  contact_33_2879
timestamp 1624857261
transform 1 0 116144 0 1 87725
box 0 0 1 1
use contact_33  contact_33_2702
timestamp 1624857261
transform 1 0 116280 0 1 87725
box 0 0 1 1
use contact_33  contact_33_2582
timestamp 1624857261
transform 1 0 116416 0 1 87725
box 0 0 1 1
use contact_33  contact_33_2575
timestamp 1624857261
transform 1 0 116552 0 1 87861
box 0 0 1 1
use contact_33  contact_33_418
timestamp 1624857261
transform 1 0 116960 0 1 87861
box 0 0 1 1
use contact_33  contact_33_416
timestamp 1624857261
transform 1 0 116960 0 1 87725
box 0 0 1 1
use contact_33  contact_33_2779
timestamp 1624857261
transform 1 0 116280 0 1 88133
box 0 0 1 1
use contact_33  contact_33_2574
timestamp 1624857261
transform 1 0 116552 0 1 88133
box 0 0 1 1
use contact_33  contact_33_417
timestamp 1624857261
transform 1 0 116960 0 1 88133
box 0 0 1 1
use contact_33  contact_33_2778
timestamp 1624857261
transform 1 0 116280 0 1 88405
box 0 0 1 1
use contact_33  contact_33_291
timestamp 1624857261
transform 1 0 116824 0 1 88269
box 0 0 1 1
use contact_33  contact_33_2586
timestamp 1624857261
transform 1 0 116552 0 1 88541
box 0 0 1 1
use contact_33  contact_33_292
timestamp 1624857261
transform 1 0 116824 0 1 88541
box 0 0 1 1
use contact_33  contact_33_3169
timestamp 1624857261
transform 1 0 115192 0 1 89357
box 0 0 1 1
use contact_33  contact_33_756
timestamp 1624857261
transform 1 0 115736 0 1 89357
box 0 0 1 1
use contact_33  contact_33_141
timestamp 1624857261
transform 1 0 116960 0 1 89357
box 0 0 1 1
use contact_33  contact_33_142
timestamp 1624857261
transform 1 0 116960 0 1 89085
box 0 0 1 1
use contact_33  contact_33_289
timestamp 1624857261
transform 1 0 116824 0 1 88949
box 0 0 1 1
use contact_33  contact_33_290
timestamp 1624857261
transform 1 0 116824 0 1 88677
box 0 0 1 1
use contact_33  contact_33_2587
timestamp 1624857261
transform 1 0 116552 0 1 88949
box 0 0 1 1
use contact_33  contact_33_3106
timestamp 1624857261
transform 1 0 115192 0 1 89765
box 0 0 1 1
use contact_33  contact_33_3107
timestamp 1624857261
transform 1 0 115192 0 1 90037
box 0 0 1 1
use contact_33  contact_33_3168
timestamp 1624857261
transform 1 0 115192 0 1 89629
box 0 0 1 1
use contact_33  contact_33_3234
timestamp 1624857261
transform 1 0 115328 0 1 90173
box 0 0 1 1
use contact_33  contact_33_477
timestamp 1624857261
transform 1 0 115736 0 1 90037
box 0 0 1 1
use contact_33  contact_33_478
timestamp 1624857261
transform 1 0 115736 0 1 89765
box 0 0 1 1
use contact_33  contact_33_689
timestamp 1624857261
transform 1 0 115736 0 1 90173
box 0 0 1 1
use contact_33  contact_33_755
timestamp 1624857261
transform 1 0 115736 0 1 89629
box 0 0 1 1
use contact_33  contact_33_2826
timestamp 1624857261
transform 1 0 116008 0 1 90037
box 0 0 1 1
use contact_33  contact_33_2827
timestamp 1624857261
transform 1 0 116008 0 1 89765
box 0 0 1 1
use contact_33  contact_33_3018
timestamp 1624857261
transform 1 0 116144 0 1 90173
box 0 0 1 1
use contact_33  contact_33_445
timestamp 1624857261
transform 1 0 116824 0 1 90037
box 0 0 1 1
use contact_33  contact_33_446
timestamp 1624857261
transform 1 0 116824 0 1 89765
box 0 0 1 1
use contact_33  contact_33_2716
timestamp 1624857261
transform 1 0 116280 0 1 89765
box 0 0 1 1
use contact_33  contact_33_2717
timestamp 1624857261
transform 1 0 116280 0 1 90037
box 0 0 1 1
use contact_33  contact_33_2719
timestamp 1624857261
transform 1 0 116280 0 1 90173
box 0 0 1 1
use contact_33  contact_33_3235
timestamp 1624857261
transform 1 0 115328 0 1 90445
box 0 0 1 1
use contact_33  contact_33_3236
timestamp 1624857261
transform 1 0 115328 0 1 90581
box 0 0 1 1
use contact_33  contact_33_3237
timestamp 1624857261
transform 1 0 115328 0 1 90853
box 0 0 1 1
use contact_33  contact_33_3250
timestamp 1624857261
transform 1 0 115192 0 1 90989
box 0 0 1 1
use contact_33  contact_33_690
timestamp 1624857261
transform 1 0 115736 0 1 90445
box 0 0 1 1
use contact_33  contact_33_691
timestamp 1624857261
transform 1 0 115736 0 1 90853
box 0 0 1 1
use contact_33  contact_33_692
timestamp 1624857261
transform 1 0 115736 0 1 90581
box 0 0 1 1
use contact_33  contact_33_709
timestamp 1624857261
transform 1 0 115600 0 1 90989
box 0 0 1 1
use contact_33  contact_33_2953
timestamp 1624857261
transform 1 0 116144 0 1 90989
box 0 0 1 1
use contact_33  contact_33_3019
timestamp 1624857261
transform 1 0 116144 0 1 90445
box 0 0 1 1
use contact_33  contact_33_151
timestamp 1624857261
transform 1 0 116824 0 1 90853
box 0 0 1 1
use contact_33  contact_33_152
timestamp 1624857261
transform 1 0 116824 0 1 90581
box 0 0 1 1
use contact_33  contact_33_189
timestamp 1624857261
transform 1 0 116960 0 1 90989
box 0 0 1 1
use contact_33  contact_33_2674
timestamp 1624857261
transform 1 0 116416 0 1 90581
box 0 0 1 1
use contact_33  contact_33_2675
timestamp 1624857261
transform 1 0 116416 0 1 90853
box 0 0 1 1
use contact_33  contact_33_2718
timestamp 1624857261
transform 1 0 116280 0 1 90445
box 0 0 1 1
use contact_33  contact_33_3251
timestamp 1624857261
transform 1 0 115192 0 1 91261
box 0 0 1 1
use contact_33  contact_33_3259
timestamp 1624857261
transform 1 0 115328 0 1 91805
box 0 0 1 1
use contact_33  contact_33_3260
timestamp 1624857261
transform 1 0 115328 0 1 91397
box 0 0 1 1
use contact_33  contact_33_3261
timestamp 1624857261
transform 1 0 115328 0 1 91669
box 0 0 1 1
use contact_33  contact_33_551
timestamp 1624857261
transform 1 0 115600 0 1 91805
box 0 0 1 1
use contact_33  contact_33_707
timestamp 1624857261
transform 1 0 115600 0 1 91669
box 0 0 1 1
use contact_33  contact_33_708
timestamp 1624857261
transform 1 0 115600 0 1 91397
box 0 0 1 1
use contact_33  contact_33_710
timestamp 1624857261
transform 1 0 115600 0 1 91261
box 0 0 1 1
use contact_33  contact_33_2910
timestamp 1624857261
transform 1 0 116144 0 1 91397
box 0 0 1 1
use contact_33  contact_33_2911
timestamp 1624857261
transform 1 0 116144 0 1 91669
box 0 0 1 1
use contact_33  contact_33_2952
timestamp 1624857261
transform 1 0 116144 0 1 91261
box 0 0 1 1
use contact_33  contact_33_187
timestamp 1624857261
transform 1 0 116960 0 1 91669
box 0 0 1 1
use contact_33  contact_33_188
timestamp 1624857261
transform 1 0 116960 0 1 91397
box 0 0 1 1
use contact_33  contact_33_190
timestamp 1624857261
transform 1 0 116960 0 1 91261
box 0 0 1 1
use contact_33  contact_33_389
timestamp 1624857261
transform 1 0 116960 0 1 91805
box 0 0 1 1
use contact_33  contact_33_2770
timestamp 1624857261
transform 1 0 116280 0 1 91805
box 0 0 1 1
use contact_33  contact_33_3258
timestamp 1624857261
transform 1 0 115328 0 1 92077
box 0 0 1 1
use contact_33  contact_33_552
timestamp 1624857261
transform 1 0 115600 0 1 92077
box 0 0 1 1
use contact_33  contact_33_385
timestamp 1624857261
transform 1 0 116824 0 1 92621
box 0 0 1 1
use contact_33  contact_33_390
timestamp 1624857261
transform 1 0 116960 0 1 92077
box 0 0 1 1
use contact_33  contact_33_391
timestamp 1624857261
transform 1 0 116960 0 1 92485
box 0 0 1 1
use contact_33  contact_33_392
timestamp 1624857261
transform 1 0 116960 0 1 92213
box 0 0 1 1
use contact_33  contact_33_2638
timestamp 1624857261
transform 1 0 116416 0 1 92621
box 0 0 1 1
use contact_33  contact_33_2771
timestamp 1624857261
transform 1 0 116280 0 1 92077
box 0 0 1 1
use contact_33  contact_33_825
timestamp 1624857261
transform 1 0 110160 0 1 93981
box 0 0 1 1
use contact_33  contact_33_826
timestamp 1624857261
transform 1 0 110160 0 1 94253
box 0 0 1 1
use contact_33  contact_33_905
timestamp 1624857261
transform 1 0 110160 0 1 95477
box 0 0 1 1
use contact_33  contact_33_959
timestamp 1624857261
transform 1 0 110296 0 1 92757
box 0 0 1 1
use contact_33  contact_33_960
timestamp 1624857261
transform 1 0 110296 0 1 93029
box 0 0 1 1
use contact_33  contact_33_877
timestamp 1624857261
transform 1 0 110160 0 1 97381
box 0 0 1 1
use contact_33  contact_33_878
timestamp 1624857261
transform 1 0 110160 0 1 97109
box 0 0 1 1
use contact_33  contact_33_879
timestamp 1624857261
transform 1 0 110296 0 1 96701
box 0 0 1 1
use contact_33  contact_33_880
timestamp 1624857261
transform 1 0 110296 0 1 96973
box 0 0 1 1
use contact_33  contact_33_906
timestamp 1624857261
transform 1 0 110160 0 1 95749
box 0 0 1 1
use contact_33  contact_33_872
timestamp 1624857261
transform 1 0 110160 0 1 101053
box 0 0 1 1
use contact_33  contact_33_941
timestamp 1624857261
transform 1 0 110296 0 1 100237
box 0 0 1 1
use contact_33  contact_33_942
timestamp 1624857261
transform 1 0 110296 0 1 100509
box 0 0 1 1
use contact_33  contact_33_943
timestamp 1624857261
transform 1 0 110296 0 1 100917
box 0 0 1 1
use contact_33  contact_33_944
timestamp 1624857261
transform 1 0 110296 0 1 100645
box 0 0 1 1
use contact_33  contact_33_871
timestamp 1624857261
transform 1 0 110160 0 1 101325
box 0 0 1 1
use contact_33  contact_33_859
timestamp 1624857261
transform 1 0 110296 0 1 105813
box 0 0 1 1
use contact_33  contact_33_860
timestamp 1624857261
transform 1 0 110296 0 1 106085
box 0 0 1 1
use contact_33  contact_33_949
timestamp 1624857261
transform 1 0 110432 0 1 109213
box 0 0 1 1
use contact_33  contact_33_950
timestamp 1624857261
transform 1 0 110432 0 1 108941
box 0 0 1 1
use contact_33  contact_33_961
timestamp 1624857261
transform 1 0 110296 0 1 109213
box 0 0 1 1
use contact_33  contact_33_962
timestamp 1624857261
transform 1 0 110296 0 1 109621
box 0 0 1 1
use contact_33  contact_33_964
timestamp 1624857261
transform 1 0 110160 0 1 109757
box 0 0 1 1
use contact_33  contact_33_965
timestamp 1624857261
transform 1 0 110160 0 1 109349
box 0 0 1 1
use contact_33  contact_33_966
timestamp 1624857261
transform 1 0 110160 0 1 109621
box 0 0 1 1
use contact_33  contact_33_963
timestamp 1624857261
transform 1 0 110160 0 1 110029
box 0 0 1 1
use contact_33  contact_33_3090
timestamp 1624857261
transform 1 0 115192 0 1 93301
box 0 0 1 1
use contact_33  contact_33_814
timestamp 1624857261
transform 1 0 115600 0 1 93301
box 0 0 1 1
use contact_33  contact_33_386
timestamp 1624857261
transform 1 0 116824 0 1 92893
box 0 0 1 1
use contact_33  contact_33_387
timestamp 1624857261
transform 1 0 116824 0 1 93301
box 0 0 1 1
use contact_33  contact_33_388
timestamp 1624857261
transform 1 0 116824 0 1 93029
box 0 0 1 1
use contact_33  contact_33_2639
timestamp 1624857261
transform 1 0 116416 0 1 92893
box 0 0 1 1
use contact_33  contact_33_2670
timestamp 1624857261
transform 1 0 116416 0 1 93301
box 0 0 1 1
use contact_33  contact_33_3091
timestamp 1624857261
transform 1 0 115192 0 1 93573
box 0 0 1 1
use contact_33  contact_33_3188
timestamp 1624857261
transform 1 0 115328 0 1 94389
box 0 0 1 1
use contact_33  contact_33_3189
timestamp 1624857261
transform 1 0 115328 0 1 94117
box 0 0 1 1
use contact_33  contact_33_3190
timestamp 1624857261
transform 1 0 115328 0 1 93709
box 0 0 1 1
use contact_33  contact_33_3191
timestamp 1624857261
transform 1 0 115328 0 1 93981
box 0 0 1 1
use contact_33  contact_33_615
timestamp 1624857261
transform 1 0 115600 0 1 94117
box 0 0 1 1
use contact_33  contact_33_616
timestamp 1624857261
transform 1 0 115600 0 1 94389
box 0 0 1 1
use contact_33  contact_33_629
timestamp 1624857261
transform 1 0 115736 0 1 93981
box 0 0 1 1
use contact_33  contact_33_630
timestamp 1624857261
transform 1 0 115736 0 1 93709
box 0 0 1 1
use contact_33  contact_33_813
timestamp 1624857261
transform 1 0 115600 0 1 93573
box 0 0 1 1
use contact_33  contact_33_2890
timestamp 1624857261
transform 1 0 116280 0 1 94117
box 0 0 1 1
use contact_33  contact_33_2891
timestamp 1624857261
transform 1 0 116280 0 1 94389
box 0 0 1 1
use contact_33  contact_33_2892
timestamp 1624857261
transform 1 0 116008 0 1 94117
box 0 0 1 1
use contact_33  contact_33_2893
timestamp 1624857261
transform 1 0 116008 0 1 94389
box 0 0 1 1
use contact_33  contact_33_2671
timestamp 1624857261
transform 1 0 116416 0 1 93573
box 0 0 1 1
use contact_33  contact_33_3042
timestamp 1624857261
transform 1 0 115328 0 1 95205
box 0 0 1 1
use contact_33  contact_33_3043
timestamp 1624857261
transform 1 0 115328 0 1 94933
box 0 0 1 1
use contact_33  contact_33_3084
timestamp 1624857261
transform 1 0 115192 0 1 94797
box 0 0 1 1
use contact_33  contact_33_3085
timestamp 1624857261
transform 1 0 115192 0 1 94525
box 0 0 1 1
use contact_33  contact_33_547
timestamp 1624857261
transform 1 0 115736 0 1 94933
box 0 0 1 1
use contact_33  contact_33_548
timestamp 1624857261
transform 1 0 115736 0 1 95205
box 0 0 1 1
use contact_33  contact_33_613
timestamp 1624857261
transform 1 0 115600 0 1 94797
box 0 0 1 1
use contact_33  contact_33_614
timestamp 1624857261
transform 1 0 115600 0 1 94525
box 0 0 1 1
use contact_33  contact_33_2932
timestamp 1624857261
transform 1 0 116008 0 1 94933
box 0 0 1 1
use contact_33  contact_33_2933
timestamp 1624857261
transform 1 0 116008 0 1 95205
box 0 0 1 1
use contact_33  contact_33_351
timestamp 1624857261
transform 1 0 116824 0 1 94525
box 0 0 1 1
use contact_33  contact_33_352
timestamp 1624857261
transform 1 0 116824 0 1 94797
box 0 0 1 1
use contact_33  contact_33_353
timestamp 1624857261
transform 1 0 116824 0 1 95205
box 0 0 1 1
use contact_33  contact_33_354
timestamp 1624857261
transform 1 0 116824 0 1 94933
box 0 0 1 1
use contact_33  contact_33_2566
timestamp 1624857261
transform 1 0 116416 0 1 94933
box 0 0 1 1
use contact_33  contact_33_2567
timestamp 1624857261
transform 1 0 116416 0 1 95205
box 0 0 1 1
use contact_33  contact_33_3364
timestamp 1624857261
transform 1 0 115192 0 1 95341
box 0 0 1 1
use contact_33  contact_33_3365
timestamp 1624857261
transform 1 0 115192 0 1 95613
box 0 0 1 1
use contact_33  contact_33_3378
timestamp 1624857261
transform 1 0 115328 0 1 95749
box 0 0 1 1
use contact_33  contact_33_3379
timestamp 1624857261
transform 1 0 115328 0 1 96021
box 0 0 1 1
use contact_33  contact_33_549
timestamp 1624857261
transform 1 0 115600 0 1 95613
box 0 0 1 1
use contact_33  contact_33_550
timestamp 1624857261
transform 1 0 115600 0 1 95341
box 0 0 1 1
use contact_33  contact_33_809
timestamp 1624857261
transform 1 0 115736 0 1 95749
box 0 0 1 1
use contact_33  contact_33_810
timestamp 1624857261
transform 1 0 115736 0 1 96021
box 0 0 1 1
use contact_33  contact_33_2930
timestamp 1624857261
transform 1 0 116144 0 1 95613
box 0 0 1 1
use contact_33  contact_33_2931
timestamp 1624857261
transform 1 0 116144 0 1 95341
box 0 0 1 1
use contact_33  contact_33_397
timestamp 1624857261
transform 1 0 116960 0 1 96021
box 0 0 1 1
use contact_33  contact_33_398
timestamp 1624857261
transform 1 0 116960 0 1 95749
box 0 0 1 1
use contact_33  contact_33_399
timestamp 1624857261
transform 1 0 116960 0 1 95341
box 0 0 1 1
use contact_33  contact_33_400
timestamp 1624857261
transform 1 0 116960 0 1 95613
box 0 0 1 1
use contact_33  contact_33_2548
timestamp 1624857261
transform 1 0 116552 0 1 96021
box 0 0 1 1
use contact_33  contact_33_2549
timestamp 1624857261
transform 1 0 116552 0 1 95749
box 0 0 1 1
use contact_33  contact_33_3376
timestamp 1624857261
transform 1 0 115328 0 1 96429
box 0 0 1 1
use contact_33  contact_33_3377
timestamp 1624857261
transform 1 0 115328 0 1 96157
box 0 0 1 1
use contact_33  contact_33_811
timestamp 1624857261
transform 1 0 115736 0 1 96429
box 0 0 1 1
use contact_33  contact_33_812
timestamp 1624857261
transform 1 0 115736 0 1 96157
box 0 0 1 1
use contact_33  contact_33_2902
timestamp 1624857261
transform 1 0 116280 0 1 96157
box 0 0 1 1
use contact_33  contact_33_2903
timestamp 1624857261
transform 1 0 116280 0 1 96429
box 0 0 1 1
use contact_33  contact_33_251
timestamp 1624857261
transform 1 0 116960 0 1 96157
box 0 0 1 1
use contact_33  contact_33_252
timestamp 1624857261
transform 1 0 116960 0 1 96429
box 0 0 1 1
use contact_33  contact_33_253
timestamp 1624857261
transform 1 0 116960 0 1 96837
box 0 0 1 1
use contact_33  contact_33_254
timestamp 1624857261
transform 1 0 116960 0 1 96565
box 0 0 1 1
use contact_33  contact_33_2664
timestamp 1624857261
transform 1 0 116552 0 1 96837
box 0 0 1 1
use contact_33  contact_33_2665
timestamp 1624857261
transform 1 0 116552 0 1 96565
box 0 0 1 1
use contact_33  contact_33_3038
timestamp 1624857261
transform 1 0 115192 0 1 97653
box 0 0 1 1
use contact_33  contact_33_3204
timestamp 1624857261
transform 1 0 115328 0 1 97517
box 0 0 1 1
use contact_33  contact_33_3205
timestamp 1624857261
transform 1 0 115328 0 1 97245
box 0 0 1 1
use contact_33  contact_33_475
timestamp 1624857261
transform 1 0 115600 0 1 97653
box 0 0 1 1
use contact_33  contact_33_727
timestamp 1624857261
transform 1 0 115736 0 1 97517
box 0 0 1 1
use contact_33  contact_33_728
timestamp 1624857261
transform 1 0 115736 0 1 97245
box 0 0 1 1
use contact_33  contact_33_2788
timestamp 1624857261
transform 1 0 116280 0 1 97245
box 0 0 1 1
use contact_33  contact_33_2789
timestamp 1624857261
transform 1 0 116280 0 1 97517
box 0 0 1 1
use contact_33  contact_33_225
timestamp 1624857261
transform 1 0 116824 0 1 97245
box 0 0 1 1
use contact_33  contact_33_226
timestamp 1624857261
transform 1 0 116824 0 1 96973
box 0 0 1 1
use contact_33  contact_33_3039
timestamp 1624857261
transform 1 0 115192 0 1 97925
box 0 0 1 1
use contact_33  contact_33_3040
timestamp 1624857261
transform 1 0 115328 0 1 98333
box 0 0 1 1
use contact_33  contact_33_3041
timestamp 1624857261
transform 1 0 115328 0 1 98061
box 0 0 1 1
use contact_33  contact_33_3270
timestamp 1624857261
transform 1 0 115192 0 1 98469
box 0 0 1 1
use contact_33  contact_33_473
timestamp 1624857261
transform 1 0 115736 0 1 98333
box 0 0 1 1
use contact_33  contact_33_474
timestamp 1624857261
transform 1 0 115736 0 1 98061
box 0 0 1 1
use contact_33  contact_33_476
timestamp 1624857261
transform 1 0 115600 0 1 97925
box 0 0 1 1
use contact_33  contact_33_603
timestamp 1624857261
transform 1 0 115600 0 1 98469
box 0 0 1 1
use contact_33  contact_33_2969
timestamp 1624857261
transform 1 0 116008 0 1 98469
box 0 0 1 1
use contact_33  contact_33_2970
timestamp 1624857261
transform 1 0 116008 0 1 98061
box 0 0 1 1
use contact_33  contact_33_2971
timestamp 1624857261
transform 1 0 116008 0 1 98333
box 0 0 1 1
use contact_33  contact_33_303
timestamp 1624857261
transform 1 0 116960 0 1 98469
box 0 0 1 1
use contact_33  contact_33_2590
timestamp 1624857261
transform 1 0 116416 0 1 98061
box 0 0 1 1
use contact_33  contact_33_2591
timestamp 1624857261
transform 1 0 116416 0 1 98333
box 0 0 1 1
use contact_33  contact_33_3268
timestamp 1624857261
transform 1 0 115192 0 1 99149
box 0 0 1 1
use contact_33  contact_33_3269
timestamp 1624857261
transform 1 0 115192 0 1 98877
box 0 0 1 1
use contact_33  contact_33_3271
timestamp 1624857261
transform 1 0 115192 0 1 98741
box 0 0 1 1
use contact_33  contact_33_3352
timestamp 1624857261
transform 1 0 115192 0 1 99285
box 0 0 1 1
use contact_33  contact_33_595
timestamp 1624857261
transform 1 0 115736 0 1 99285
box 0 0 1 1
use contact_33  contact_33_601
timestamp 1624857261
transform 1 0 115600 0 1 99149
box 0 0 1 1
use contact_33  contact_33_602
timestamp 1624857261
transform 1 0 115600 0 1 98877
box 0 0 1 1
use contact_33  contact_33_604
timestamp 1624857261
transform 1 0 115600 0 1 98741
box 0 0 1 1
use contact_33  contact_33_2800
timestamp 1624857261
transform 1 0 116280 0 1 99285
box 0 0 1 1
use contact_33  contact_33_2904
timestamp 1624857261
transform 1 0 116144 0 1 98877
box 0 0 1 1
use contact_33  contact_33_2905
timestamp 1624857261
transform 1 0 116144 0 1 99149
box 0 0 1 1
use contact_33  contact_33_2968
timestamp 1624857261
transform 1 0 116008 0 1 98741
box 0 0 1 1
use contact_33  contact_33_265
timestamp 1624857261
transform 1 0 116824 0 1 99285
box 0 0 1 1
use contact_33  contact_33_301
timestamp 1624857261
transform 1 0 116960 0 1 99149
box 0 0 1 1
use contact_33  contact_33_302
timestamp 1624857261
transform 1 0 116960 0 1 98877
box 0 0 1 1
use contact_33  contact_33_304
timestamp 1624857261
transform 1 0 116960 0 1 98741
box 0 0 1 1
use contact_33  contact_33_2616
timestamp 1624857261
transform 1 0 116416 0 1 99285
box 0 0 1 1
use contact_33  contact_33_2650
timestamp 1624857261
transform 1 0 116552 0 1 99149
box 0 0 1 1
use contact_33  contact_33_2651
timestamp 1624857261
transform 1 0 116552 0 1 98877
box 0 0 1 1
use contact_33  contact_33_3126
timestamp 1624857261
transform 1 0 115328 0 1 100101
box 0 0 1 1
use contact_33  contact_33_3127
timestamp 1624857261
transform 1 0 115328 0 1 100373
box 0 0 1 1
use contact_33  contact_33_3350
timestamp 1624857261
transform 1 0 115192 0 1 99965
box 0 0 1 1
use contact_33  contact_33_3351
timestamp 1624857261
transform 1 0 115192 0 1 99693
box 0 0 1 1
use contact_33  contact_33_3353
timestamp 1624857261
transform 1 0 115192 0 1 99557
box 0 0 1 1
use contact_33  contact_33_593
timestamp 1624857261
transform 1 0 115600 0 1 99965
box 0 0 1 1
use contact_33  contact_33_594
timestamp 1624857261
transform 1 0 115600 0 1 99693
box 0 0 1 1
use contact_33  contact_33_596
timestamp 1624857261
transform 1 0 115736 0 1 99557
box 0 0 1 1
use contact_33  contact_33_677
timestamp 1624857261
transform 1 0 115736 0 1 100101
box 0 0 1 1
use contact_33  contact_33_678
timestamp 1624857261
transform 1 0 115736 0 1 100373
box 0 0 1 1
use contact_33  contact_33_2801
timestamp 1624857261
transform 1 0 116280 0 1 99557
box 0 0 1 1
use contact_33  contact_33_2914
timestamp 1624857261
transform 1 0 116008 0 1 99693
box 0 0 1 1
use contact_33  contact_33_2915
timestamp 1624857261
transform 1 0 116008 0 1 99965
box 0 0 1 1
use contact_33  contact_33_169
timestamp 1624857261
transform 1 0 116960 0 1 100373
box 0 0 1 1
use contact_33  contact_33_170
timestamp 1624857261
transform 1 0 116960 0 1 100101
box 0 0 1 1
use contact_33  contact_33_266
timestamp 1624857261
transform 1 0 116824 0 1 99557
box 0 0 1 1
use contact_33  contact_33_267
timestamp 1624857261
transform 1 0 116824 0 1 99965
box 0 0 1 1
use contact_33  contact_33_268
timestamp 1624857261
transform 1 0 116824 0 1 99693
box 0 0 1 1
use contact_33  contact_33_2617
timestamp 1624857261
transform 1 0 116416 0 1 99557
box 0 0 1 1
use contact_33  contact_33_2865
timestamp 1624857261
transform 1 0 116280 0 1 101189
box 0 0 1 1
use contact_33  contact_33_2922
timestamp 1624857261
transform 1 0 116144 0 1 100509
box 0 0 1 1
use contact_33  contact_33_2923
timestamp 1624857261
transform 1 0 116144 0 1 100781
box 0 0 1 1
use contact_33  contact_33_355
timestamp 1624857261
transform 1 0 116960 0 1 100509
box 0 0 1 1
use contact_33  contact_33_356
timestamp 1624857261
transform 1 0 116960 0 1 100781
box 0 0 1 1
use contact_33  contact_33_357
timestamp 1624857261
transform 1 0 116960 0 1 101189
box 0 0 1 1
use contact_33  contact_33_358
timestamp 1624857261
transform 1 0 116960 0 1 100917
box 0 0 1 1
use contact_33  contact_33_2618
timestamp 1624857261
transform 1 0 116416 0 1 100781
box 0 0 1 1
use contact_33  contact_33_2619
timestamp 1624857261
transform 1 0 116416 0 1 100509
box 0 0 1 1
use contact_33  contact_33_3387
timestamp 1624857261
transform 1 0 115192 0 1 102005
box 0 0 1 1
use contact_33  contact_33_3388
timestamp 1624857261
transform 1 0 115192 0 1 101597
box 0 0 1 1
use contact_33  contact_33_3389
timestamp 1624857261
transform 1 0 115192 0 1 101869
box 0 0 1 1
use contact_33  contact_33_622
timestamp 1624857261
transform 1 0 115600 0 1 102005
box 0 0 1 1
use contact_33  contact_33_623
timestamp 1624857261
transform 1 0 115600 0 1 101597
box 0 0 1 1
use contact_33  contact_33_624
timestamp 1624857261
transform 1 0 115600 0 1 101869
box 0 0 1 1
use contact_33  contact_33_2864
timestamp 1624857261
transform 1 0 116280 0 1 101461
box 0 0 1 1
use contact_33  contact_33_203
timestamp 1624857261
transform 1 0 116960 0 1 102005
box 0 0 1 1
use contact_33  contact_33_204
timestamp 1624857261
transform 1 0 116960 0 1 101733
box 0 0 1 1
use contact_33  contact_33_2539
timestamp 1624857261
transform 1 0 116552 0 1 102005
box 0 0 1 1
use contact_33  contact_33_3077
timestamp 1624857261
transform 1 0 115328 0 1 102821
box 0 0 1 1
use contact_33  contact_33_3202
timestamp 1624857261
transform 1 0 115192 0 1 102685
box 0 0 1 1
use contact_33  contact_33_3203
timestamp 1624857261
transform 1 0 115192 0 1 102413
box 0 0 1 1
use contact_33  contact_33_3386
timestamp 1624857261
transform 1 0 115192 0 1 102277
box 0 0 1 1
use contact_33  contact_33_588
timestamp 1624857261
transform 1 0 115736 0 1 102821
box 0 0 1 1
use contact_33  contact_33_589
timestamp 1624857261
transform 1 0 115736 0 1 102413
box 0 0 1 1
use contact_33  contact_33_590
timestamp 1624857261
transform 1 0 115736 0 1 102685
box 0 0 1 1
use contact_33  contact_33_621
timestamp 1624857261
transform 1 0 115600 0 1 102277
box 0 0 1 1
use contact_33  contact_33_2834
timestamp 1624857261
transform 1 0 116144 0 1 102685
box 0 0 1 1
use contact_33  contact_33_2835
timestamp 1624857261
transform 1 0 116144 0 1 102413
box 0 0 1 1
use contact_33  contact_33_75
timestamp 1624857261
transform 1 0 116824 0 1 102685
box 0 0 1 1
use contact_33  contact_33_76
timestamp 1624857261
transform 1 0 116824 0 1 102413
box 0 0 1 1
use contact_33  contact_33_85
timestamp 1624857261
transform 1 0 116960 0 1 102821
box 0 0 1 1
use contact_33  contact_33_2538
timestamp 1624857261
transform 1 0 116552 0 1 102277
box 0 0 1 1
use contact_33  contact_33_2552
timestamp 1624857261
transform 1 0 116416 0 1 102413
box 0 0 1 1
use contact_33  contact_33_2553
timestamp 1624857261
transform 1 0 116416 0 1 102685
box 0 0 1 1
use contact_33  contact_33_3076
timestamp 1624857261
transform 1 0 115328 0 1 103093
box 0 0 1 1
use contact_33  contact_33_3116
timestamp 1624857261
transform 1 0 115328 0 1 103229
box 0 0 1 1
use contact_33  contact_33_3117
timestamp 1624857261
transform 1 0 115328 0 1 103501
box 0 0 1 1
use contact_33  contact_33_3119
timestamp 1624857261
transform 1 0 115328 0 1 103637
box 0 0 1 1
use contact_33  contact_33_461
timestamp 1624857261
transform 1 0 115736 0 1 103229
box 0 0 1 1
use contact_33  contact_33_462
timestamp 1624857261
transform 1 0 115736 0 1 103501
box 0 0 1 1
use contact_33  contact_33_535
timestamp 1624857261
transform 1 0 115736 0 1 103637
box 0 0 1 1
use contact_33  contact_33_587
timestamp 1624857261
transform 1 0 115736 0 1 103093
box 0 0 1 1
use contact_33  contact_33_2774
timestamp 1624857261
transform 1 0 116280 0 1 103229
box 0 0 1 1
use contact_33  contact_33_2775
timestamp 1624857261
transform 1 0 116280 0 1 103501
box 0 0 1 1
use contact_33  contact_33_2978
timestamp 1624857261
transform 1 0 116008 0 1 103637
box 0 0 1 1
use contact_33  contact_33_86
timestamp 1624857261
transform 1 0 116960 0 1 103093
box 0 0 1 1
use contact_33  contact_33_95
timestamp 1624857261
transform 1 0 116824 0 1 103229
box 0 0 1 1
use contact_33  contact_33_96
timestamp 1624857261
transform 1 0 116824 0 1 103501
box 0 0 1 1
use contact_33  contact_33_227
timestamp 1624857261
transform 1 0 116824 0 1 103637
box 0 0 1 1
use contact_33  contact_33_3049
timestamp 1624857261
transform 1 0 115192 0 1 104453
box 0 0 1 1
use contact_33  contact_33_3114
timestamp 1624857261
transform 1 0 115192 0 1 104317
box 0 0 1 1
use contact_33  contact_33_3115
timestamp 1624857261
transform 1 0 115192 0 1 104045
box 0 0 1 1
use contact_33  contact_33_3118
timestamp 1624857261
transform 1 0 115328 0 1 103909
box 0 0 1 1
use contact_33  contact_33_536
timestamp 1624857261
transform 1 0 115736 0 1 103909
box 0 0 1 1
use contact_33  contact_33_643
timestamp 1624857261
transform 1 0 115600 0 1 104045
box 0 0 1 1
use contact_33  contact_33_644
timestamp 1624857261
transform 1 0 115600 0 1 104317
box 0 0 1 1
use contact_33  contact_33_646
timestamp 1624857261
transform 1 0 115600 0 1 104453
box 0 0 1 1
use contact_33  contact_33_2918
timestamp 1624857261
transform 1 0 116008 0 1 104453
box 0 0 1 1
use contact_33  contact_33_2979
timestamp 1624857261
transform 1 0 116008 0 1 103909
box 0 0 1 1
use contact_33  contact_33_2980
timestamp 1624857261
transform 1 0 116144 0 1 104317
box 0 0 1 1
use contact_33  contact_33_2981
timestamp 1624857261
transform 1 0 116144 0 1 104045
box 0 0 1 1
use contact_33  contact_33_228
timestamp 1624857261
transform 1 0 116824 0 1 103909
box 0 0 1 1
use contact_33  contact_33_338
timestamp 1624857261
transform 1 0 116960 0 1 104453
box 0 0 1 1
use contact_33  contact_33_339
timestamp 1624857261
transform 1 0 116960 0 1 104045
box 0 0 1 1
use contact_33  contact_33_340
timestamp 1624857261
transform 1 0 116960 0 1 104317
box 0 0 1 1
use contact_33  contact_33_3048
timestamp 1624857261
transform 1 0 115192 0 1 104725
box 0 0 1 1
use contact_33  contact_33_645
timestamp 1624857261
transform 1 0 115600 0 1 104725
box 0 0 1 1
use contact_33  contact_33_2919
timestamp 1624857261
transform 1 0 116008 0 1 104725
box 0 0 1 1
use contact_33  contact_33_333
timestamp 1624857261
transform 1 0 116960 0 1 104861
box 0 0 1 1
use contact_33  contact_33_334
timestamp 1624857261
transform 1 0 116960 0 1 105133
box 0 0 1 1
use contact_33  contact_33_337
timestamp 1624857261
transform 1 0 116960 0 1 104725
box 0 0 1 1
use contact_33  contact_33_2600
timestamp 1624857261
transform 1 0 116416 0 1 105133
box 0 0 1 1
use contact_33  contact_33_2601
timestamp 1624857261
transform 1 0 116416 0 1 105405
box 0 0 1 1
use contact_33  contact_33_3158
timestamp 1624857261
transform 1 0 115328 0 1 105541
box 0 0 1 1
use contact_33  contact_33_3159
timestamp 1624857261
transform 1 0 115328 0 1 105813
box 0 0 1 1
use contact_33  contact_33_3160
timestamp 1624857261
transform 1 0 115328 0 1 106221
box 0 0 1 1
use contact_33  contact_33_3161
timestamp 1624857261
transform 1 0 115328 0 1 105949
box 0 0 1 1
use contact_33  contact_33_3332
timestamp 1624857261
transform 1 0 115192 0 1 106357
box 0 0 1 1
use contact_33  contact_33_584
timestamp 1624857261
transform 1 0 115600 0 1 106357
box 0 0 1 1
use contact_33  contact_33_821
timestamp 1624857261
transform 1 0 115736 0 1 106221
box 0 0 1 1
use contact_33  contact_33_822
timestamp 1624857261
transform 1 0 115736 0 1 105949
box 0 0 1 1
use contact_33  contact_33_823
timestamp 1624857261
transform 1 0 115736 0 1 105541
box 0 0 1 1
use contact_33  contact_33_824
timestamp 1624857261
transform 1 0 115736 0 1 105813
box 0 0 1 1
use contact_33  contact_33_168
timestamp 1624857261
transform 1 0 116960 0 1 106357
box 0 0 1 1
use contact_33  contact_33_269
timestamp 1624857261
transform 1 0 116824 0 1 105677
box 0 0 1 1
use contact_33  contact_33_270
timestamp 1624857261
transform 1 0 116824 0 1 105949
box 0 0 1 1
use contact_33  contact_33_2641
timestamp 1624857261
transform 1 0 116552 0 1 106357
box 0 0 1 1
use contact_33  contact_33_3238
timestamp 1624857261
transform 1 0 115192 0 1 107173
box 0 0 1 1
use contact_33  contact_33_3333
timestamp 1624857261
transform 1 0 115192 0 1 106629
box 0 0 1 1
use contact_33  contact_33_3334
timestamp 1624857261
transform 1 0 115192 0 1 107037
box 0 0 1 1
use contact_33  contact_33_3335
timestamp 1624857261
transform 1 0 115192 0 1 106765
box 0 0 1 1
use contact_33  contact_33_491
timestamp 1624857261
transform 1 0 115736 0 1 106765
box 0 0 1 1
use contact_33  contact_33_492
timestamp 1624857261
transform 1 0 115736 0 1 107037
box 0 0 1 1
use contact_33  contact_33_583
timestamp 1624857261
transform 1 0 115600 0 1 106629
box 0 0 1 1
use contact_33  contact_33_771
timestamp 1624857261
transform 1 0 115600 0 1 107173
box 0 0 1 1
use contact_33  contact_33_2894
timestamp 1624857261
transform 1 0 116008 0 1 106765
box 0 0 1 1
use contact_33  contact_33_2895
timestamp 1624857261
transform 1 0 116008 0 1 107037
box 0 0 1 1
use contact_33  contact_33_2897
timestamp 1624857261
transform 1 0 116008 0 1 107173
box 0 0 1 1
use contact_33  contact_33_167
timestamp 1624857261
transform 1 0 116960 0 1 106629
box 0 0 1 1
use contact_33  contact_33_383
timestamp 1624857261
transform 1 0 116960 0 1 107173
box 0 0 1 1
use contact_33  contact_33_2640
timestamp 1624857261
transform 1 0 116552 0 1 106629
box 0 0 1 1
use contact_33  contact_33_3231
timestamp 1624857261
transform 1 0 115328 0 1 107989
box 0 0 1 1
use contact_33  contact_33_3239
timestamp 1624857261
transform 1 0 115192 0 1 107445
box 0 0 1 1
use contact_33  contact_33_3240
timestamp 1624857261
transform 1 0 115192 0 1 107853
box 0 0 1 1
use contact_33  contact_33_3241
timestamp 1624857261
transform 1 0 115192 0 1 107581
box 0 0 1 1
use contact_33  contact_33_483
timestamp 1624857261
transform 1 0 115736 0 1 107989
box 0 0 1 1
use contact_33  contact_33_769
timestamp 1624857261
transform 1 0 115600 0 1 107853
box 0 0 1 1
use contact_33  contact_33_770
timestamp 1624857261
transform 1 0 115600 0 1 107581
box 0 0 1 1
use contact_33  contact_33_772
timestamp 1624857261
transform 1 0 115600 0 1 107445
box 0 0 1 1
use contact_33  contact_33_2832
timestamp 1624857261
transform 1 0 116280 0 1 107989
box 0 0 1 1
use contact_33  contact_33_2896
timestamp 1624857261
transform 1 0 116008 0 1 107445
box 0 0 1 1
use contact_33  contact_33_3002
timestamp 1624857261
transform 1 0 116144 0 1 107581
box 0 0 1 1
use contact_33  contact_33_3003
timestamp 1624857261
transform 1 0 116144 0 1 107853
box 0 0 1 1
use contact_33  contact_33_136
timestamp 1624857261
transform 1 0 116824 0 1 107989
box 0 0 1 1
use contact_33  contact_33_381
timestamp 1624857261
transform 1 0 116960 0 1 107853
box 0 0 1 1
use contact_33  contact_33_382
timestamp 1624857261
transform 1 0 116960 0 1 107581
box 0 0 1 1
use contact_33  contact_33_384
timestamp 1624857261
transform 1 0 116960 0 1 107445
box 0 0 1 1
use contact_33  contact_33_2662
timestamp 1624857261
transform 1 0 116416 0 1 107581
box 0 0 1 1
use contact_33  contact_33_2663
timestamp 1624857261
transform 1 0 116416 0 1 107853
box 0 0 1 1
use contact_33  contact_33_3200
timestamp 1624857261
transform 1 0 115192 0 1 108669
box 0 0 1 1
use contact_33  contact_33_3201
timestamp 1624857261
transform 1 0 115192 0 1 108397
box 0 0 1 1
use contact_33  contact_33_3230
timestamp 1624857261
transform 1 0 115328 0 1 108261
box 0 0 1 1
use contact_33  contact_33_484
timestamp 1624857261
transform 1 0 115736 0 1 108261
box 0 0 1 1
use contact_33  contact_33_581
timestamp 1624857261
transform 1 0 115600 0 1 108397
box 0 0 1 1
use contact_33  contact_33_582
timestamp 1624857261
transform 1 0 115600 0 1 108669
box 0 0 1 1
use contact_33  contact_33_2833
timestamp 1624857261
transform 1 0 116280 0 1 108261
box 0 0 1 1
use contact_33  contact_33_2934
timestamp 1624857261
transform 1 0 116008 0 1 108397
box 0 0 1 1
use contact_33  contact_33_2935
timestamp 1624857261
transform 1 0 116008 0 1 108669
box 0 0 1 1
use contact_33  contact_33_135
timestamp 1624857261
transform 1 0 116824 0 1 108261
box 0 0 1 1
use contact_33  contact_33_217
timestamp 1624857261
transform 1 0 116960 0 1 108397
box 0 0 1 1
use contact_33  contact_33_218
timestamp 1624857261
transform 1 0 116960 0 1 108669
box 0 0 1 1
use contact_33  contact_33_220
timestamp 1624857261
transform 1 0 116960 0 1 108805
box 0 0 1 1
use contact_33  contact_33_2936
timestamp 1624857261
transform 1 0 116280 0 1 109213
box 0 0 1 1
use contact_33  contact_33_2937
timestamp 1624857261
transform 1 0 116280 0 1 109485
box 0 0 1 1
use contact_33  contact_33_2938
timestamp 1624857261
transform 1 0 116144 0 1 109213
box 0 0 1 1
use contact_33  contact_33_2939
timestamp 1624857261
transform 1 0 116144 0 1 109485
box 0 0 1 1
use contact_33  contact_33_109
timestamp 1624857261
transform 1 0 116960 0 1 109213
box 0 0 1 1
use contact_33  contact_33_110
timestamp 1624857261
transform 1 0 116960 0 1 109485
box 0 0 1 1
use contact_33  contact_33_219
timestamp 1624857261
transform 1 0 116960 0 1 109077
box 0 0 1 1
use contact_33  contact_33_413
timestamp 1624857261
transform 1 0 116960 0 1 109621
box 0 0 1 1
use contact_33  contact_33_3224
timestamp 1624857261
transform 1 0 115192 0 1 110301
box 0 0 1 1
use contact_33  contact_33_3225
timestamp 1624857261
transform 1 0 115192 0 1 110573
box 0 0 1 1
use contact_33  contact_33_3366
timestamp 1624857261
transform 1 0 115192 0 1 110165
box 0 0 1 1
use contact_33  contact_33_3367
timestamp 1624857261
transform 1 0 115192 0 1 109893
box 0 0 1 1
use contact_33  contact_33_555
timestamp 1624857261
transform 1 0 115736 0 1 109893
box 0 0 1 1
use contact_33  contact_33_556
timestamp 1624857261
transform 1 0 115736 0 1 110165
box 0 0 1 1
use contact_33  contact_33_557
timestamp 1624857261
transform 1 0 115736 0 1 110573
box 0 0 1 1
use contact_33  contact_33_558
timestamp 1624857261
transform 1 0 115736 0 1 110301
box 0 0 1 1
use contact_33  contact_33_2756
timestamp 1624857261
transform 1 0 116008 0 1 110165
box 0 0 1 1
use contact_33  contact_33_2757
timestamp 1624857261
transform 1 0 116008 0 1 109893
box 0 0 1 1
use contact_33  contact_33_414
timestamp 1624857261
transform 1 0 116960 0 1 109893
box 0 0 1 1
use contact_33  contact_33_3222
timestamp 1624857261
transform 1 0 115192 0 1 110981
box 0 0 1 1
use contact_33  contact_33_3223
timestamp 1624857261
transform 1 0 115192 0 1 110709
box 0 0 1 1
use contact_33  contact_33_3280
timestamp 1624857261
transform 1 0 115328 0 1 111117
box 0 0 1 1
use contact_33  contact_33_463
timestamp 1624857261
transform 1 0 115600 0 1 110981
box 0 0 1 1
use contact_33  contact_33_464
timestamp 1624857261
transform 1 0 115600 0 1 110709
box 0 0 1 1
use contact_33  contact_33_479
timestamp 1624857261
transform 1 0 115736 0 1 111117
box 0 0 1 1
use contact_33  contact_33_114
timestamp 1624857261
transform 1 0 116824 0 1 111117
box 0 0 1 1
use contact_33  contact_33_2550
timestamp 1624857261
transform 1 0 116552 0 1 110981
box 0 0 1 1
use contact_33  contact_33_2551
timestamp 1624857261
transform 1 0 116552 0 1 110709
box 0 0 1 1
use contact_33  contact_33_2598
timestamp 1624857261
transform 1 0 116416 0 1 111117
box 0 0 1 1
use contact_33  contact_33_3872
timestamp 1624857261
transform 1 0 69088 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3873
timestamp 1624857261
transform 1 0 69088 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3876
timestamp 1624857261
transform 1 0 68408 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3877
timestamp 1624857261
transform 1 0 68408 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3878
timestamp 1624857261
transform 1 0 67864 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3879
timestamp 1624857261
transform 1 0 67864 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3848
timestamp 1624857261
transform 1 0 70856 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3849
timestamp 1624857261
transform 1 0 70856 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3852
timestamp 1624857261
transform 1 0 70312 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3853
timestamp 1624857261
transform 1 0 70312 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3864
timestamp 1624857261
transform 1 0 69632 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3865
timestamp 1624857261
transform 1 0 69632 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3838
timestamp 1624857261
transform 1 0 72080 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3839
timestamp 1624857261
transform 1 0 72080 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3814
timestamp 1624857261
transform 1 0 74120 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3815
timestamp 1624857261
transform 1 0 74120 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3816
timestamp 1624857261
transform 1 0 73304 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3817
timestamp 1624857261
transform 1 0 73304 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3820
timestamp 1624857261
transform 1 0 72896 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3821
timestamp 1624857261
transform 1 0 72896 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3836
timestamp 1624857261
transform 1 0 72760 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3837
timestamp 1624857261
transform 1 0 72760 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3786
timestamp 1624857261
transform 1 0 75888 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3787
timestamp 1624857261
transform 1 0 75888 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3790
timestamp 1624857261
transform 1 0 75344 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3791
timestamp 1624857261
transform 1 0 75344 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3808
timestamp 1624857261
transform 1 0 75208 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3809
timestamp 1624857261
transform 1 0 75208 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3772
timestamp 1624857261
transform 1 0 77112 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3773
timestamp 1624857261
transform 1 0 77112 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3778
timestamp 1624857261
transform 1 0 76568 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3779
timestamp 1624857261
transform 1 0 76568 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3750
timestamp 1624857261
transform 1 0 78336 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3751
timestamp 1624857261
transform 1 0 78336 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3756
timestamp 1624857261
transform 1 0 77792 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3757
timestamp 1624857261
transform 1 0 77792 0 1 121589
box 0 0 1 1
use contact_33  contact_33_1155
timestamp 1624857261
transform 1 0 69904 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1143
timestamp 1624857261
transform 1 0 72488 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1131
timestamp 1624857261
transform 1 0 75072 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1119
timestamp 1624857261
transform 1 0 77520 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1156
timestamp 1624857261
transform 1 0 69904 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1159
timestamp 1624857261
transform 1 0 69768 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1144
timestamp 1624857261
transform 1 0 72488 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1149
timestamp 1624857261
transform 1 0 72352 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1132
timestamp 1624857261
transform 1 0 75072 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1135
timestamp 1624857261
transform 1 0 74936 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1120
timestamp 1624857261
transform 1 0 77520 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1123
timestamp 1624857261
transform 1 0 77384 0 1 125669
box 0 0 1 1
use contact_7  contact_7_343
timestamp 1624857261
transform 1 0 69493 0 1 127542
box 0 0 1 1
use contact_19  contact_19_949
timestamp 1624857261
transform 1 0 69494 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1160
timestamp 1624857261
transform 1 0 69768 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3856
timestamp 1624857261
transform 1 0 69632 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3857
timestamp 1624857261
transform 1 0 69632 0 1 126485
box 0 0 1 1
use contact_33  contact_33_5433
timestamp 1624857261
transform 1 0 69360 0 1 127573
box 0 0 1 1
use contact_7  contact_7_342
timestamp 1624857261
transform 1 0 71989 0 1 127542
box 0 0 1 1
use contact_19  contact_19_948
timestamp 1624857261
transform 1 0 71990 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1150
timestamp 1624857261
transform 1 0 72352 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3830
timestamp 1624857261
transform 1 0 72216 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3831
timestamp 1624857261
transform 1 0 72216 0 1 126485
box 0 0 1 1
use contact_33  contact_33_5432
timestamp 1624857261
transform 1 0 72080 0 1 127573
box 0 0 1 1
use contact_33  contact_33_5431
timestamp 1624857261
transform 1 0 74392 0 1 127573
box 0 0 1 1
use contact_7  contact_7_341
timestamp 1624857261
transform 1 0 74485 0 1 127542
box 0 0 1 1
use contact_19  contact_19_947
timestamp 1624857261
transform 1 0 74486 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1136
timestamp 1624857261
transform 1 0 74936 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3798
timestamp 1624857261
transform 1 0 74800 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3799
timestamp 1624857261
transform 1 0 74800 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3826
timestamp 1624857261
transform 1 0 74528 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3827
timestamp 1624857261
transform 1 0 74528 0 1 127165
box 0 0 1 1
use contact_7  contact_7_340
timestamp 1624857261
transform 1 0 76981 0 1 127542
box 0 0 1 1
use contact_19  contact_19_946
timestamp 1624857261
transform 1 0 76982 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1124
timestamp 1624857261
transform 1 0 77384 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3766
timestamp 1624857261
transform 1 0 77248 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3767
timestamp 1624857261
transform 1 0 77248 0 1 126485
box 0 0 1 1
use contact_33  contact_33_5430
timestamp 1624857261
transform 1 0 76976 0 1 127573
box 0 0 1 1
use contact_33  contact_33_3730
timestamp 1624857261
transform 1 0 80512 0 1 121453
box 0 0 1 1
use contact_33  contact_33_3731
timestamp 1624857261
transform 1 0 80512 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3742
timestamp 1624857261
transform 1 0 79560 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3743
timestamp 1624857261
transform 1 0 79560 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3718
timestamp 1624857261
transform 1 0 81600 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3719
timestamp 1624857261
transform 1 0 81600 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3726
timestamp 1624857261
transform 1 0 81464 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3727
timestamp 1624857261
transform 1 0 81464 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3692
timestamp 1624857261
transform 1 0 83368 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3693
timestamp 1624857261
transform 1 0 83368 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3696
timestamp 1624857261
transform 1 0 82824 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3697
timestamp 1624857261
transform 1 0 82824 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3668
timestamp 1624857261
transform 1 0 85408 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3669
timestamp 1624857261
transform 1 0 85408 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3680
timestamp 1624857261
transform 1 0 84592 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3681
timestamp 1624857261
transform 1 0 84592 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3690
timestamp 1624857261
transform 1 0 84048 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3691
timestamp 1624857261
transform 1 0 84048 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3652
timestamp 1624857261
transform 1 0 87040 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3653
timestamp 1624857261
transform 1 0 87040 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3656
timestamp 1624857261
transform 1 0 86496 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3657
timestamp 1624857261
transform 1 0 86496 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3664
timestamp 1624857261
transform 1 0 85816 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3665
timestamp 1624857261
transform 1 0 85816 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3634
timestamp 1624857261
transform 1 0 88400 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3635
timestamp 1624857261
transform 1 0 88400 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3642
timestamp 1624857261
transform 1 0 87856 0 1 122133
box 0 0 1 1
use contact_33  contact_33_3630
timestamp 1624857261
transform 1 0 89216 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3631
timestamp 1624857261
transform 1 0 89216 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3632
timestamp 1624857261
transform 1 0 89080 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3633
timestamp 1624857261
transform 1 0 89080 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3612
timestamp 1624857261
transform 1 0 90304 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3613
timestamp 1624857261
transform 1 0 90304 0 1 121589
box 0 0 1 1
use contact_33  contact_33_1107
timestamp 1624857261
transform 1 0 79832 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1095
timestamp 1624857261
transform 1 0 82552 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1085
timestamp 1624857261
transform 1 0 85000 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1071
timestamp 1624857261
transform 1 0 87312 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1061
timestamp 1624857261
transform 1 0 89896 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1108
timestamp 1624857261
transform 1 0 79832 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1111
timestamp 1624857261
transform 1 0 79696 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3735
timestamp 1624857261
transform 1 0 79832 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3765
timestamp 1624857261
transform 1 0 79560 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3707
timestamp 1624857261
transform 1 0 82280 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3733
timestamp 1624857261
transform 1 0 82008 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1096
timestamp 1624857261
transform 1 0 82552 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1101
timestamp 1624857261
transform 1 0 82416 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1086
timestamp 1624857261
transform 1 0 85000 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1089
timestamp 1624857261
transform 1 0 84864 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3675
timestamp 1624857261
transform 1 0 84592 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3705
timestamp 1624857261
transform 1 0 84456 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1072
timestamp 1624857261
transform 1 0 87312 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1075
timestamp 1624857261
transform 1 0 87176 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3643
timestamp 1624857261
transform 1 0 87856 0 1 126349
box 0 0 1 1
use contact_33  contact_33_3645
timestamp 1624857261
transform 1 0 87312 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1062
timestamp 1624857261
transform 1 0 89896 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1063
timestamp 1624857261
transform 1 0 89760 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3619
timestamp 1624857261
transform 1 0 89624 0 1 126485
box 0 0 1 1
use contact_7  contact_7_339
timestamp 1624857261
transform 1 0 79477 0 1 127542
box 0 0 1 1
use contact_19  contact_19_945
timestamp 1624857261
transform 1 0 79478 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1112
timestamp 1624857261
transform 1 0 79832 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3734
timestamp 1624857261
transform 1 0 79832 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3764
timestamp 1624857261
transform 1 0 79560 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5429
timestamp 1624857261
transform 1 0 79424 0 1 127573
box 0 0 1 1
use contact_7  contact_7_338
timestamp 1624857261
transform 1 0 81973 0 1 127542
box 0 0 1 1
use contact_19  contact_19_944
timestamp 1624857261
transform 1 0 81974 0 1 127547
box 0 0 1 1
use contact_33  contact_33_3706
timestamp 1624857261
transform 1 0 82280 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3732
timestamp 1624857261
transform 1 0 82008 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5428
timestamp 1624857261
transform 1 0 82008 0 1 127573
box 0 0 1 1
use contact_33  contact_33_1102
timestamp 1624857261
transform 1 0 82416 0 1 127437
box 0 0 1 1
use contact_7  contact_7_337
timestamp 1624857261
transform 1 0 84469 0 1 127542
box 0 0 1 1
use contact_19  contact_19_943
timestamp 1624857261
transform 1 0 84470 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1090
timestamp 1624857261
transform 1 0 84864 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3674
timestamp 1624857261
transform 1 0 84592 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3704
timestamp 1624857261
transform 1 0 84456 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5427
timestamp 1624857261
transform 1 0 84456 0 1 127573
box 0 0 1 1
use contact_7  contact_7_336
timestamp 1624857261
transform 1 0 86965 0 1 127542
box 0 0 1 1
use contact_19  contact_19_942
timestamp 1624857261
transform 1 0 86966 0 1 127547
box 0 0 1 1
use contact_33  contact_33_5426
timestamp 1624857261
transform 1 0 87040 0 1 127573
box 0 0 1 1
use contact_33  contact_33_1076
timestamp 1624857261
transform 1 0 87312 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3644
timestamp 1624857261
transform 1 0 87312 0 1 127165
box 0 0 1 1
use contact_7  contact_7_335
timestamp 1624857261
transform 1 0 89461 0 1 127542
box 0 0 1 1
use contact_19  contact_19_941
timestamp 1624857261
transform 1 0 89462 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1064
timestamp 1624857261
transform 1 0 89760 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3618
timestamp 1624857261
transform 1 0 89624 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5425
timestamp 1624857261
transform 1 0 89488 0 1 127573
box 0 0 1 1
use contact_33  contact_33_3603
timestamp 1624857261
transform 1 0 91528 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3608
timestamp 1624857261
transform 1 0 90848 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3582
timestamp 1624857261
transform 1 0 93296 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3589
timestamp 1624857261
transform 1 0 92752 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3560
timestamp 1624857261
transform 1 0 95472 0 1 121453
box 0 0 1 1
use contact_33  contact_33_3576
timestamp 1624857261
transform 1 0 94248 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3550
timestamp 1624857261
transform 1 0 97104 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3527
timestamp 1624857261
transform 1 0 99008 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3530
timestamp 1624857261
transform 1 0 98328 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3539
timestamp 1624857261
transform 1 0 97784 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3506
timestamp 1624857261
transform 1 0 100776 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3524
timestamp 1624857261
transform 1 0 99552 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3496
timestamp 1624857261
transform 1 0 102000 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3499
timestamp 1624857261
transform 1 0 101592 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3602
timestamp 1624857261
transform 1 0 91528 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3609
timestamp 1624857261
transform 1 0 90848 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3583
timestamp 1624857261
transform 1 0 93296 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3588
timestamp 1624857261
transform 1 0 92752 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3561
timestamp 1624857261
transform 1 0 95472 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3577
timestamp 1624857261
transform 1 0 94248 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3551
timestamp 1624857261
transform 1 0 97104 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3526
timestamp 1624857261
transform 1 0 99008 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3531
timestamp 1624857261
transform 1 0 98328 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3538
timestamp 1624857261
transform 1 0 97784 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3507
timestamp 1624857261
transform 1 0 100776 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3525
timestamp 1624857261
transform 1 0 99552 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3497
timestamp 1624857261
transform 1 0 102000 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3498
timestamp 1624857261
transform 1 0 101592 0 1 121997
box 0 0 1 1
use contact_33  contact_33_1049
timestamp 1624857261
transform 1 0 92480 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1037
timestamp 1624857261
transform 1 0 94928 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1025
timestamp 1624857261
transform 1 0 97512 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1013
timestamp 1624857261
transform 1 0 99960 0 1 123765
box 0 0 1 1
use contact_33  contact_33_1053
timestamp 1624857261
transform 1 0 92344 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3593
timestamp 1624857261
transform 1 0 92208 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1050
timestamp 1624857261
transform 1 0 92480 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1038
timestamp 1624857261
transform 1 0 94928 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1039
timestamp 1624857261
transform 1 0 94792 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3565
timestamp 1624857261
transform 1 0 94656 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1026
timestamp 1624857261
transform 1 0 97512 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1027
timestamp 1624857261
transform 1 0 97376 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3543
timestamp 1624857261
transform 1 0 97240 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1014
timestamp 1624857261
transform 1 0 99960 0 1 125669
box 0 0 1 1
use contact_33  contact_33_1015
timestamp 1624857261
transform 1 0 99824 0 1 125669
box 0 0 1 1
use contact_33  contact_33_3511
timestamp 1624857261
transform 1 0 99688 0 1 126485
box 0 0 1 1
use contact_33  contact_33_3541
timestamp 1624857261
transform 1 0 99416 0 1 126485
box 0 0 1 1
use contact_33  contact_33_1005
timestamp 1624857261
transform 1 0 102136 0 1 125669
box 0 0 1 1
use contact_7  contact_7_334
timestamp 1624857261
transform 1 0 91957 0 1 127542
box 0 0 1 1
use contact_19  contact_19_940
timestamp 1624857261
transform 1 0 91958 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1054
timestamp 1624857261
transform 1 0 92344 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3592
timestamp 1624857261
transform 1 0 92208 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5424
timestamp 1624857261
transform 1 0 91936 0 1 127573
box 0 0 1 1
use contact_7  contact_7_333
timestamp 1624857261
transform 1 0 94453 0 1 127542
box 0 0 1 1
use contact_19  contact_19_939
timestamp 1624857261
transform 1 0 94454 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1040
timestamp 1624857261
transform 1 0 94792 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3564
timestamp 1624857261
transform 1 0 94656 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5423
timestamp 1624857261
transform 1 0 94384 0 1 127573
box 0 0 1 1
use contact_7  contact_7_332
timestamp 1624857261
transform 1 0 96949 0 1 127542
box 0 0 1 1
use contact_19  contact_19_938
timestamp 1624857261
transform 1 0 96950 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1028
timestamp 1624857261
transform 1 0 97376 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3542
timestamp 1624857261
transform 1 0 97240 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5422
timestamp 1624857261
transform 1 0 96832 0 1 127573
box 0 0 1 1
use contact_7  contact_7_331
timestamp 1624857261
transform 1 0 99445 0 1 127542
box 0 0 1 1
use contact_19  contact_19_937
timestamp 1624857261
transform 1 0 99446 0 1 127547
box 0 0 1 1
use contact_33  contact_33_1016
timestamp 1624857261
transform 1 0 99824 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3510
timestamp 1624857261
transform 1 0 99688 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3540
timestamp 1624857261
transform 1 0 99416 0 1 127165
box 0 0 1 1
use contact_33  contact_33_5421
timestamp 1624857261
transform 1 0 99416 0 1 127573
box 0 0 1 1
use contact_7  contact_7_330
timestamp 1624857261
transform 1 0 101941 0 1 127542
box 0 0 1 1
use contact_19  contact_19_936
timestamp 1624857261
transform 1 0 101942 0 1 127547
box 0 0 1 1
use contact_33  contact_33_5420
timestamp 1624857261
transform 1 0 102000 0 1 127573
box 0 0 1 1
use contact_33  contact_33_911
timestamp 1624857261
transform 1 0 110296 0 1 112069
box 0 0 1 1
use contact_33  contact_33_912
timestamp 1624857261
transform 1 0 110296 0 1 112341
box 0 0 1 1
use contact_33  contact_33_833
timestamp 1624857261
transform 1 0 110432 0 1 113565
box 0 0 1 1
use contact_33  contact_33_834
timestamp 1624857261
transform 1 0 110432 0 1 113293
box 0 0 1 1
use contact_33  contact_33_851
timestamp 1624857261
transform 1 0 110296 0 1 114517
box 0 0 1 1
use contact_33  contact_33_852
timestamp 1624857261
transform 1 0 110296 0 1 114789
box 0 0 1 1
use contact_33  contact_33_847
timestamp 1624857261
transform 1 0 110160 0 1 117237
box 0 0 1 1
use contact_33  contact_33_848
timestamp 1624857261
transform 1 0 110160 0 1 117509
box 0 0 1 1
use contact_33  contact_33_849
timestamp 1624857261
transform 1 0 110432 0 1 117917
box 0 0 1 1
use contact_33  contact_33_850
timestamp 1624857261
transform 1 0 110432 0 1 117645
box 0 0 1 1
use contact_33  contact_33_883
timestamp 1624857261
transform 1 0 110296 0 1 118189
box 0 0 1 1
use contact_33  contact_33_884
timestamp 1624857261
transform 1 0 110296 0 1 117917
box 0 0 1 1
use contact_33  contact_33_901
timestamp 1624857261
transform 1 0 110296 0 1 118461
box 0 0 1 1
use contact_33  contact_33_902
timestamp 1624857261
transform 1 0 110296 0 1 118733
box 0 0 1 1
use contact_33  contact_33_3472
timestamp 1624857261
transform 1 0 104040 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3473
timestamp 1624857261
transform 1 0 104040 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3476
timestamp 1624857261
transform 1 0 103904 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3477
timestamp 1624857261
transform 1 0 103904 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3478
timestamp 1624857261
transform 1 0 103360 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3479
timestamp 1624857261
transform 1 0 103360 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3450
timestamp 1624857261
transform 1 0 105808 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3451
timestamp 1624857261
transform 1 0 105808 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3468
timestamp 1624857261
transform 1 0 104584 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3469
timestamp 1624857261
transform 1 0 104584 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3440
timestamp 1624857261
transform 1 0 107032 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3441
timestamp 1624857261
transform 1 0 107032 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3418
timestamp 1624857261
transform 1 0 109480 0 1 121589
box 0 0 1 1
use contact_33  contact_33_3419
timestamp 1624857261
transform 1 0 109480 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3428
timestamp 1624857261
transform 1 0 108120 0 1 121997
box 0 0 1 1
use contact_33  contact_33_3429
timestamp 1624857261
transform 1 0 108120 0 1 121589
box 0 0 1 1
use contact_33  contact_33_969
timestamp 1624857261
transform 1 0 110160 0 1 121045
box 0 0 1 1
use contact_33  contact_33_3416
timestamp 1624857261
transform 1 0 111656 0 1 121181
box 0 0 1 1
use contact_33  contact_33_3417
timestamp 1624857261
transform 1 0 111656 0 1 121453
box 0 0 1 1
use contact_33  contact_33_1001
timestamp 1624857261
transform 1 0 102408 0 1 123765
box 0 0 1 1
use contact_33  contact_33_989
timestamp 1624857261
transform 1 0 104992 0 1 123765
box 0 0 1 1
use contact_33  contact_33_975
timestamp 1624857261
transform 1 0 107440 0 1 123765
box 0 0 1 1
use contact_7  contact_7_479
timestamp 1624857261
transform 1 0 111124 0 1 123964
box 0 0 1 1
use contact_33  contact_33_970
timestamp 1624857261
transform 1 0 110160 0 1 123493
box 0 0 1 1
use contact_33  contact_33_1002
timestamp 1624857261
transform 1 0 102408 0 1 125669
box 0 0 1 1
use contact_33  contact_33_990
timestamp 1624857261
transform 1 0 104992 0 1 125669
box 0 0 1 1
use contact_33  contact_33_991
timestamp 1624857261
transform 1 0 104856 0 1 125669
box 0 0 1 1
use contact_33  contact_33_976
timestamp 1624857261
transform 1 0 107440 0 1 125669
box 0 0 1 1
use contact_33  contact_33_979
timestamp 1624857261
transform 1 0 107304 0 1 125669
box 0 0 1 1
use contact_7  contact_7_481
timestamp 1624857261
transform 1 0 111000 0 1 125378
box 0 0 1 1
use contact_33  contact_33_1006
timestamp 1624857261
transform 1 0 102272 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3486
timestamp 1624857261
transform 1 0 102272 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3487
timestamp 1624857261
transform 1 0 102272 0 1 126485
box 0 0 1 1
use contact_7  contact_7_329
timestamp 1624857261
transform 1 0 104437 0 1 127542
box 0 0 1 1
use contact_19  contact_19_935
timestamp 1624857261
transform 1 0 104438 0 1 127547
box 0 0 1 1
use contact_33  contact_33_992
timestamp 1624857261
transform 1 0 104856 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3456
timestamp 1624857261
transform 1 0 104720 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3457
timestamp 1624857261
transform 1 0 104720 0 1 126485
box 0 0 1 1
use contact_33  contact_33_5419
timestamp 1624857261
transform 1 0 104448 0 1 127573
box 0 0 1 1
use contact_7  contact_7_328
timestamp 1624857261
transform 1 0 106933 0 1 127542
box 0 0 1 1
use contact_19  contact_19_934
timestamp 1624857261
transform 1 0 106934 0 1 127547
box 0 0 1 1
use contact_33  contact_33_980
timestamp 1624857261
transform 1 0 107304 0 1 127437
box 0 0 1 1
use contact_33  contact_33_3430
timestamp 1624857261
transform 1 0 107168 0 1 127165
box 0 0 1 1
use contact_33  contact_33_3431
timestamp 1624857261
transform 1 0 107168 0 1 126485
box 0 0 1 1
use contact_33  contact_33_5418
timestamp 1624857261
transform 1 0 107032 0 1 127573
box 0 0 1 1
use contact_33  contact_33_3283
timestamp 1624857261
transform 1 0 115328 0 1 111525
box 0 0 1 1
use contact_33  contact_33_3282
timestamp 1624857261
transform 1 0 115328 0 1 111797
box 0 0 1 1
use contact_33  contact_33_3281
timestamp 1624857261
transform 1 0 115328 0 1 111389
box 0 0 1 1
use contact_33  contact_33_3167
timestamp 1624857261
transform 1 0 115192 0 1 111933
box 0 0 1 1
use contact_33  contact_33_3009
timestamp 1624857261
transform 1 0 116008 0 1 111525
box 0 0 1 1
use contact_33  contact_33_3008
timestamp 1624857261
transform 1 0 116008 0 1 111797
box 0 0 1 1
use contact_33  contact_33_2845
timestamp 1624857261
transform 1 0 116008 0 1 111933
box 0 0 1 1
use contact_33  contact_33_777
timestamp 1624857261
transform 1 0 115736 0 1 111933
box 0 0 1 1
use contact_33  contact_33_526
timestamp 1624857261
transform 1 0 115600 0 1 111797
box 0 0 1 1
use contact_33  contact_33_525
timestamp 1624857261
transform 1 0 115600 0 1 111525
box 0 0 1 1
use contact_33  contact_33_480
timestamp 1624857261
transform 1 0 115736 0 1 111389
box 0 0 1 1
use contact_33  contact_33_2612
timestamp 1624857261
transform 1 0 116416 0 1 111933
box 0 0 1 1
use contact_33  contact_33_2599
timestamp 1624857261
transform 1 0 116416 0 1 111389
box 0 0 1 1
use contact_33  contact_33_231
timestamp 1624857261
transform 1 0 116824 0 1 111933
box 0 0 1 1
use contact_33  contact_33_138
timestamp 1624857261
transform 1 0 116960 0 1 111797
box 0 0 1 1
use contact_33  contact_33_137
timestamp 1624857261
transform 1 0 116960 0 1 111525
box 0 0 1 1
use contact_33  contact_33_113
timestamp 1624857261
transform 1 0 116824 0 1 111389
box 0 0 1 1
use contact_33  contact_33_3393
timestamp 1624857261
transform 1 0 115192 0 1 112749
box 0 0 1 1
use contact_33  contact_33_3391
timestamp 1624857261
transform 1 0 115192 0 1 112613
box 0 0 1 1
use contact_33  contact_33_3390
timestamp 1624857261
transform 1 0 115192 0 1 112341
box 0 0 1 1
use contact_33  contact_33_3166
timestamp 1624857261
transform 1 0 115192 0 1 112205
box 0 0 1 1
use contact_33  contact_33_2844
timestamp 1624857261
transform 1 0 116008 0 1 112205
box 0 0 1 1
use contact_33  contact_33_2809
timestamp 1624857261
transform 1 0 116144 0 1 112341
box 0 0 1 1
use contact_33  contact_33_2808
timestamp 1624857261
transform 1 0 116144 0 1 112613
box 0 0 1 1
use contact_33  contact_33_780
timestamp 1624857261
transform 1 0 115736 0 1 112341
box 0 0 1 1
use contact_33  contact_33_779
timestamp 1624857261
transform 1 0 115736 0 1 112613
box 0 0 1 1
use contact_33  contact_33_778
timestamp 1624857261
transform 1 0 115736 0 1 112205
box 0 0 1 1
use contact_33  contact_33_618
timestamp 1624857261
transform 1 0 115600 0 1 112749
box 0 0 1 1
use contact_33  contact_33_2613
timestamp 1624857261
transform 1 0 116416 0 1 112205
box 0 0 1 1
use contact_33  contact_33_232
timestamp 1624857261
transform 1 0 116824 0 1 112205
box 0 0 1 1
use contact_33  contact_33_230
timestamp 1624857261
transform 1 0 116824 0 1 112341
box 0 0 1 1
use contact_33  contact_33_229
timestamp 1624857261
transform 1 0 116824 0 1 112613
box 0 0 1 1
use contact_33  contact_33_107
timestamp 1624857261
transform 1 0 116960 0 1 112749
box 0 0 1 1
use contact_33  contact_33_3392
timestamp 1624857261
transform 1 0 115192 0 1 113021
box 0 0 1 1
use contact_33  contact_33_617
timestamp 1624857261
transform 1 0 115600 0 1 113021
box 0 0 1 1
use contact_33  contact_33_286
timestamp 1624857261
transform 1 0 116824 0 1 113429
box 0 0 1 1
use contact_33  contact_33_285
timestamp 1624857261
transform 1 0 116824 0 1 113157
box 0 0 1 1
use contact_33  contact_33_284
timestamp 1624857261
transform 1 0 116824 0 1 113565
box 0 0 1 1
use contact_33  contact_33_108
timestamp 1624857261
transform 1 0 116960 0 1 113021
box 0 0 1 1
use contact_33  contact_33_3345
timestamp 1624857261
transform 1 0 115192 0 1 113837
box 0 0 1 1
use contact_33  contact_33_3344
timestamp 1624857261
transform 1 0 115192 0 1 114109
box 0 0 1 1
use contact_33  contact_33_3195
timestamp 1624857261
transform 1 0 115192 0 1 114245
box 0 0 1 1
use contact_33  contact_33_3194
timestamp 1624857261
transform 1 0 115192 0 1 114517
box 0 0 1 1
use contact_33  contact_33_716
timestamp 1624857261
transform 1 0 115736 0 1 114517
box 0 0 1 1
use contact_33  contact_33_715
timestamp 1624857261
transform 1 0 115736 0 1 114245
box 0 0 1 1
use contact_33  contact_33_696
timestamp 1624857261
transform 1 0 115600 0 1 113837
box 0 0 1 1
use contact_33  contact_33_695
timestamp 1624857261
transform 1 0 115600 0 1 114109
box 0 0 1 1
use contact_33  contact_33_2631
timestamp 1624857261
transform 1 0 116416 0 1 114109
box 0 0 1 1
use contact_33  contact_33_2630
timestamp 1624857261
transform 1 0 116416 0 1 113837
box 0 0 1 1
use contact_33  contact_33_283
timestamp 1624857261
transform 1 0 116824 0 1 113837
box 0 0 1 1
use contact_33  contact_33_3383
timestamp 1624857261
transform 1 0 115328 0 1 115469
box 0 0 1 1
use contact_33  contact_33_3381
timestamp 1624857261
transform 1 0 115328 0 1 115333
box 0 0 1 1
use contact_33  contact_33_3380
timestamp 1624857261
transform 1 0 115328 0 1 115061
box 0 0 1 1
use contact_33  contact_33_3155
timestamp 1624857261
transform 1 0 115328 0 1 114653
box 0 0 1 1
use contact_33  contact_33_3154
timestamp 1624857261
transform 1 0 115328 0 1 114925
box 0 0 1 1
use contact_33  contact_33_2783
timestamp 1624857261
transform 1 0 116144 0 1 114925
box 0 0 1 1
use contact_33  contact_33_2782
timestamp 1624857261
transform 1 0 116144 0 1 114653
box 0 0 1 1
use contact_33  contact_33_714
timestamp 1624857261
transform 1 0 115736 0 1 114653
box 0 0 1 1
use contact_33  contact_33_713
timestamp 1624857261
transform 1 0 115736 0 1 114925
box 0 0 1 1
use contact_33  contact_33_685
timestamp 1624857261
transform 1 0 115736 0 1 115469
box 0 0 1 1
use contact_33  contact_33_468
timestamp 1624857261
transform 1 0 115600 0 1 115061
box 0 0 1 1
use contact_33  contact_33_467
timestamp 1624857261
transform 1 0 115600 0 1 115333
box 0 0 1 1
use contact_33  contact_33_2643
timestamp 1624857261
transform 1 0 116552 0 1 115333
box 0 0 1 1
use contact_33  contact_33_2642
timestamp 1624857261
transform 1 0 116552 0 1 115061
box 0 0 1 1
use contact_33  contact_33_247
timestamp 1624857261
transform 1 0 116824 0 1 115469
box 0 0 1 1
use contact_33  contact_33_88
timestamp 1624857261
transform 1 0 116960 0 1 115333
box 0 0 1 1
use contact_33  contact_33_87
timestamp 1624857261
transform 1 0 116960 0 1 115061
box 0 0 1 1
use contact_33  contact_33_3382
timestamp 1624857261
transform 1 0 115328 0 1 115741
box 0 0 1 1
use contact_33  contact_33_3139
timestamp 1624857261
transform 1 0 115192 0 1 116285
box 0 0 1 1
use contact_33  contact_33_3137
timestamp 1624857261
transform 1 0 115192 0 1 116149
box 0 0 1 1
use contact_33  contact_33_3136
timestamp 1624857261
transform 1 0 115192 0 1 115877
box 0 0 1 1
use contact_33  contact_33_2985
timestamp 1624857261
transform 1 0 116008 0 1 115877
box 0 0 1 1
use contact_33  contact_33_2984
timestamp 1624857261
transform 1 0 116008 0 1 116149
box 0 0 1 1
use contact_33  contact_33_2943
timestamp 1624857261
transform 1 0 116280 0 1 116149
box 0 0 1 1
use contact_33  contact_33_2942
timestamp 1624857261
transform 1 0 116280 0 1 115877
box 0 0 1 1
use contact_33  contact_33_686
timestamp 1624857261
transform 1 0 115736 0 1 115741
box 0 0 1 1
use contact_33  contact_33_684
timestamp 1624857261
transform 1 0 115736 0 1 115877
box 0 0 1 1
use contact_33  contact_33_683
timestamp 1624857261
transform 1 0 115736 0 1 116149
box 0 0 1 1
use contact_33  contact_33_485
timestamp 1624857261
transform 1 0 115736 0 1 116285
box 0 0 1 1
use contact_33  contact_33_2605
timestamp 1624857261
transform 1 0 116552 0 1 116285
box 0 0 1 1
use contact_33  contact_33_282
timestamp 1624857261
transform 1 0 116960 0 1 116285
box 0 0 1 1
use contact_33  contact_33_280
timestamp 1624857261
transform 1 0 116960 0 1 116149
box 0 0 1 1
use contact_33  contact_33_279
timestamp 1624857261
transform 1 0 116960 0 1 115877
box 0 0 1 1
use contact_33  contact_33_248
timestamp 1624857261
transform 1 0 116824 0 1 115741
box 0 0 1 1
use contact_33  contact_33_3138
timestamp 1624857261
transform 1 0 115192 0 1 116557
box 0 0 1 1
use contact_33  contact_33_3053
timestamp 1624857261
transform 1 0 115328 0 1 116693
box 0 0 1 1
use contact_33  contact_33_3052
timestamp 1624857261
transform 1 0 115328 0 1 116965
box 0 0 1 1
use contact_33  contact_33_488
timestamp 1624857261
transform 1 0 115736 0 1 116693
box 0 0 1 1
use contact_33  contact_33_487
timestamp 1624857261
transform 1 0 115736 0 1 116965
box 0 0 1 1
use contact_33  contact_33_486
timestamp 1624857261
transform 1 0 115736 0 1 116557
box 0 0 1 1
use contact_33  contact_33_2679
timestamp 1624857261
transform 1 0 116552 0 1 117101
box 0 0 1 1
use contact_33  contact_33_2604
timestamp 1624857261
transform 1 0 116552 0 1 116557
box 0 0 1 1
use contact_33  contact_33_281
timestamp 1624857261
transform 1 0 116960 0 1 116557
box 0 0 1 1
use contact_33  contact_33_262
timestamp 1624857261
transform 1 0 116824 0 1 116693
box 0 0 1 1
use contact_33  contact_33_261
timestamp 1624857261
transform 1 0 116824 0 1 116965
box 0 0 1 1
use contact_33  contact_33_98
timestamp 1624857261
transform 1 0 116960 0 1 117101
box 0 0 1 1
use contact_33  contact_33_2759
timestamp 1624857261
transform 1 0 116280 0 1 118053
box 0 0 1 1
use contact_33  contact_33_2758
timestamp 1624857261
transform 1 0 116280 0 1 117781
box 0 0 1 1
use contact_33  contact_33_2678
timestamp 1624857261
transform 1 0 116552 0 1 117373
box 0 0 1 1
use contact_33  contact_33_264
timestamp 1624857261
transform 1 0 116824 0 1 117781
box 0 0 1 1
use contact_33  contact_33_263
timestamp 1624857261
transform 1 0 116824 0 1 117509
box 0 0 1 1
use contact_33  contact_33_97
timestamp 1624857261
transform 1 0 116960 0 1 117373
box 0 0 1 1
use contact_33  contact_33_3287
timestamp 1624857261
transform 1 0 115192 0 1 118597
box 0 0 1 1
use contact_33  contact_33_3286
timestamp 1624857261
transform 1 0 115192 0 1 118869
box 0 0 1 1
use contact_33  contact_33_3285
timestamp 1624857261
transform 1 0 115192 0 1 118461
box 0 0 1 1
use contact_33  contact_33_3284
timestamp 1624857261
transform 1 0 115192 0 1 118189
box 0 0 1 1
use contact_33  contact_33_3279
timestamp 1624857261
transform 1 0 115328 0 1 119005
box 0 0 1 1
use contact_33  contact_33_2881
timestamp 1624857261
transform 1 0 116008 0 1 119005
box 0 0 1 1
use contact_33  contact_33_2840
timestamp 1624857261
transform 1 0 116280 0 1 119005
box 0 0 1 1
use contact_33  contact_33_2815
timestamp 1624857261
transform 1 0 116280 0 1 118597
box 0 0 1 1
use contact_33  contact_33_2814
timestamp 1624857261
transform 1 0 116280 0 1 118869
box 0 0 1 1
use contact_33  contact_33_706
timestamp 1624857261
transform 1 0 115600 0 1 118189
box 0 0 1 1
use contact_33  contact_33_705
timestamp 1624857261
transform 1 0 115600 0 1 118461
box 0 0 1 1
use contact_33  contact_33_586
timestamp 1624857261
transform 1 0 115600 0 1 118597
box 0 0 1 1
use contact_33  contact_33_585
timestamp 1624857261
transform 1 0 115600 0 1 118869
box 0 0 1 1
use contact_33  contact_33_578
timestamp 1624857261
transform 1 0 115736 0 1 119005
box 0 0 1 1
use contact_33  contact_33_395
timestamp 1624857261
transform 1 0 116960 0 1 119005
box 0 0 1 1
use contact_33  contact_33_3278
timestamp 1624857261
transform 1 0 115328 0 1 119277
box 0 0 1 1
use contact_33  contact_33_3153
timestamp 1624857261
transform 1 0 115192 0 1 119685
box 0 0 1 1
use contact_33  contact_33_3152
timestamp 1624857261
transform 1 0 115192 0 1 119413
box 0 0 1 1
use contact_33  contact_33_3151
timestamp 1624857261
transform 1 0 115328 0 1 119821
box 0 0 1 1
use contact_33  contact_33_2880
timestamp 1624857261
transform 1 0 116008 0 1 119277
box 0 0 1 1
use contact_33  contact_33_2841
timestamp 1624857261
transform 1 0 116280 0 1 119277
box 0 0 1 1
use contact_33  contact_33_577
timestamp 1624857261
transform 1 0 115736 0 1 119277
box 0 0 1 1
use contact_33  contact_33_507
timestamp 1624857261
transform 1 0 115736 0 1 119821
box 0 0 1 1
use contact_33  contact_33_458
timestamp 1624857261
transform 1 0 115600 0 1 119685
box 0 0 1 1
use contact_33  contact_33_457
timestamp 1624857261
transform 1 0 115600 0 1 119413
box 0 0 1 1
use contact_33  contact_33_2645
timestamp 1624857261
transform 1 0 116552 0 1 119685
box 0 0 1 1
use contact_33  contact_33_2644
timestamp 1624857261
transform 1 0 116552 0 1 119413
box 0 0 1 1
use contact_33  contact_33_408
timestamp 1624857261
transform 1 0 116960 0 1 119685
box 0 0 1 1
use contact_33  contact_33_407
timestamp 1624857261
transform 1 0 116960 0 1 119413
box 0 0 1 1
use contact_33  contact_33_406
timestamp 1624857261
transform 1 0 116824 0 1 119821
box 0 0 1 1
use contact_33  contact_33_396
timestamp 1624857261
transform 1 0 116960 0 1 119277
box 0 0 1 1
use contact_33  contact_33_3164
timestamp 1624857261
transform 1 0 115192 0 1 120229
box 0 0 1 1
use contact_33  contact_33_3150
timestamp 1624857261
transform 1 0 115328 0 1 120093
box 0 0 1 1
use contact_33  contact_33_2755
timestamp 1624857261
transform 1 0 116008 0 1 120229
box 0 0 1 1
use contact_33  contact_33_510
timestamp 1624857261
transform 1 0 115736 0 1 120229
box 0 0 1 1
use contact_33  contact_33_508
timestamp 1624857261
transform 1 0 115736 0 1 120093
box 0 0 1 1
use contact_33  contact_33_405
timestamp 1624857261
transform 1 0 116824 0 1 120093
box 0 0 1 1
use contact_33  contact_33_347
timestamp 1624857261
transform 1 0 116960 0 1 120229
box 0 0 1 1
use contact_33  contact_33_3399
timestamp 1624857261
transform 1 0 115328 0 1 121045
box 0 0 1 1
use contact_33  contact_33_3398
timestamp 1624857261
transform 1 0 115328 0 1 120637
box 0 0 1 1
use contact_33  contact_33_3165
timestamp 1624857261
transform 1 0 115192 0 1 120501
box 0 0 1 1
use contact_33  contact_33_3397
timestamp 1624857261
transform 1 0 116280 0 1 121181
box 0 0 1 1
use contact_33  contact_33_2754
timestamp 1624857261
transform 1 0 116008 0 1 120501
box 0 0 1 1
use contact_33  contact_33_509
timestamp 1624857261
transform 1 0 115736 0 1 120501
box 0 0 1 1
use contact_33  contact_33_348
timestamp 1624857261
transform 1 0 116960 0 1 120501
box 0 0 1 1
use contact_33  contact_33_346
timestamp 1624857261
transform 1 0 117368 0 1 120637
box 0 0 1 1
use contact_33  contact_33_24
timestamp 1624857261
transform 1 0 123624 0 1 121861
box 0 0 1 1
use contact_7  contact_7_477
timestamp 1624857261
transform 1 0 114985 0 1 122550
box 0 0 1 1
use contact_33  contact_33_447
timestamp 1624857261
transform 1 0 117368 0 1 123629
box 0 0 1 1
use contact_33  contact_33_345
timestamp 1624857261
transform 1 0 117368 0 1 123357
box 0 0 1 1
use contact_33  contact_33_2479
timestamp 1624857261
transform 1 0 123760 0 1 123357
box 0 0 1 1
use contact_7  contact_7_480
timestamp 1624857261
transform 1 0 123611 0 1 123964
box 0 0 1 1
use contact_7  contact_7_478
timestamp 1624857261
transform 1 0 123611 0 1 122550
box 0 0 1 1
use contact_33  contact_33_3396
timestamp 1624857261
transform 1 0 116280 0 1 124853
box 0 0 1 1
use contact_33  contact_33_2535
timestamp 1624857261
transform 1 0 117368 0 1 124989
box 0 0 1 1
use contact_33  contact_33_23
timestamp 1624857261
transform 1 0 123624 0 1 124581
box 0 0 1 1
use contact_33  contact_33_22
timestamp 1624857261
transform 1 0 123896 0 1 124717
box 0 0 1 1
use contact_7  contact_7_482
timestamp 1624857261
transform 1 0 123611 0 1 125378
box 0 0 1 1
use contact_33  contact_33_448
timestamp 1624857261
transform 1 0 117232 0 1 126213
box 0 0 1 1
use contact_33  contact_33_63
timestamp 1624857261
transform 1 0 117504 0 1 126349
box 0 0 1 1
use contact_33  contact_33_2478
timestamp 1624857261
transform 1 0 123760 0 1 126077
box 0 0 1 1
use contact_33  contact_33_2476
timestamp 1624857261
transform 1 0 123624 0 1 126213
box 0 0 1 1
use contact_33  contact_33_21
timestamp 1624857261
transform 1 0 123896 0 1 127437
box 0 0 1 1
use contact_33  contact_33_20
timestamp 1624857261
transform 1 0 123760 0 1 127573
box 0 0 1 1
use contact_33  contact_33_2534
timestamp 1624857261
transform 1 0 117368 0 1 127709
box 0 0 1 1
use contact_33  contact_33_64
timestamp 1624857261
transform 1 0 117504 0 1 129069
box 0 0 1 1
use contact_33  contact_33_2533
timestamp 1624857261
transform 1 0 119408 0 1 127845
box 0 0 1 1
use contact_33  contact_33_62
timestamp 1624857261
transform 1 0 119544 0 1 129205
box 0 0 1 1
use contact_33  contact_33_2490
timestamp 1624857261
transform 1 0 123624 0 1 128933
box 0 0 1 1
use contact_33  contact_33_2477
timestamp 1624857261
transform 1 0 123624 0 1 128797
box 0 0 1 1
use control_logic_r  control_logic_r_0
timestamp 1624857261
transform -1 0 136182 0 -1 130364
box -75 -49 11458 18431
use contact_33  contact_33_8
timestamp 1624857261
transform 1 0 134640 0 1 123221
box 0 0 1 1
use contact_33  contact_33_7
timestamp 1624857261
transform 1 0 134640 0 1 120501
box 0 0 1 1
use contact_33  contact_33_4
timestamp 1624857261
transform 1 0 134640 0 1 117645
box 0 0 1 1
use contact_33  contact_33_3
timestamp 1624857261
transform 1 0 134640 0 1 120365
box 0 0 1 1
use contact_33  contact_33_3885
timestamp 1624857261
transform 1 0 67728 0 1 132061
box 0 0 1 1
use contact_13  contact_13_977
timestamp 1624857261
transform 1 0 67657 0 1 131992
box 0 0 1 1
use contact_13  contact_13_976
timestamp 1624857261
transform 1 0 67993 0 1 131992
box 0 0 1 1
use contact_19  contact_19_813
timestamp 1624857261
transform 1 0 67650 0 1 132001
box 0 0 1 1
use contact_14  contact_14_977
timestamp 1624857261
transform 1 0 67653 0 1 132000
box 0 0 1 1
use contact_14  contact_14_976
timestamp 1624857261
transform 1 0 67989 0 1 132000
box 0 0 1 1
use contact_7  contact_7_197
timestamp 1624857261
transform 1 0 67649 0 1 131996
box 0 0 1 1
use contact_13  contact_13_975
timestamp 1624857261
transform 1 0 68329 0 1 131992
box 0 0 1 1
use contact_14  contact_14_975
timestamp 1624857261
transform 1 0 68325 0 1 132000
box 0 0 1 1
use contact_13  contact_13_974
timestamp 1624857261
transform 1 0 68665 0 1 131992
box 0 0 1 1
use contact_14  contact_14_974
timestamp 1624857261
transform 1 0 68661 0 1 132000
box 0 0 1 1
use contact_13  contact_13_973
timestamp 1624857261
transform 1 0 69001 0 1 131992
box 0 0 1 1
use contact_14  contact_14_973
timestamp 1624857261
transform 1 0 68997 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3884
timestamp 1624857261
transform 1 0 67728 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3867
timestamp 1624857261
transform 1 0 69224 0 1 132061
box 0 0 1 1
use contact_13  contact_13_972
timestamp 1624857261
transform 1 0 69337 0 1 131992
box 0 0 1 1
use contact_19  contact_19_812
timestamp 1624857261
transform 1 0 69330 0 1 132001
box 0 0 1 1
use contact_14  contact_14_972
timestamp 1624857261
transform 1 0 69333 0 1 132000
box 0 0 1 1
use contact_7  contact_7_196
timestamp 1624857261
transform 1 0 69329 0 1 131996
box 0 0 1 1
use contact_13  contact_13_971
timestamp 1624857261
transform 1 0 69673 0 1 131992
box 0 0 1 1
use contact_14  contact_14_971
timestamp 1624857261
transform 1 0 69669 0 1 132000
box 0 0 1 1
use contact_13  contact_13_970
timestamp 1624857261
transform 1 0 70009 0 1 131992
box 0 0 1 1
use contact_13  contact_13_969
timestamp 1624857261
transform 1 0 70345 0 1 131992
box 0 0 1 1
use contact_14  contact_14_970
timestamp 1624857261
transform 1 0 70005 0 1 132000
box 0 0 1 1
use contact_14  contact_14_969
timestamp 1624857261
transform 1 0 70341 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3866
timestamp 1624857261
transform 1 0 69224 0 1 132469
box 0 0 1 1
use contact_13  contact_13_968
timestamp 1624857261
transform 1 0 70681 0 1 131992
box 0 0 1 1
use contact_14  contact_14_968
timestamp 1624857261
transform 1 0 70677 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3845
timestamp 1624857261
transform 1 0 71128 0 1 132061
box 0 0 1 1
use contact_13  contact_13_967
timestamp 1624857261
transform 1 0 71017 0 1 131992
box 0 0 1 1
use contact_19  contact_19_811
timestamp 1624857261
transform 1 0 71010 0 1 132001
box 0 0 1 1
use contact_14  contact_14_967
timestamp 1624857261
transform 1 0 71013 0 1 132000
box 0 0 1 1
use contact_7  contact_7_195
timestamp 1624857261
transform 1 0 71009 0 1 131996
box 0 0 1 1
use contact_13  contact_13_966
timestamp 1624857261
transform 1 0 71353 0 1 131992
box 0 0 1 1
use contact_13  contact_13_965
timestamp 1624857261
transform 1 0 71689 0 1 131992
box 0 0 1 1
use contact_14  contact_14_966
timestamp 1624857261
transform 1 0 71349 0 1 132000
box 0 0 1 1
use contact_14  contact_14_965
timestamp 1624857261
transform 1 0 71685 0 1 132000
box 0 0 1 1
use contact_13  contact_13_964
timestamp 1624857261
transform 1 0 72025 0 1 131992
box 0 0 1 1
use contact_14  contact_14_964
timestamp 1624857261
transform 1 0 72021 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3844
timestamp 1624857261
transform 1 0 71128 0 1 132469
box 0 0 1 1
use contact_13  contact_13_963
timestamp 1624857261
transform 1 0 72361 0 1 131992
box 0 0 1 1
use contact_14  contact_14_963
timestamp 1624857261
transform 1 0 72357 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3823
timestamp 1624857261
transform 1 0 72624 0 1 132061
box 0 0 1 1
use contact_13  contact_13_962
timestamp 1624857261
transform 1 0 72697 0 1 131992
box 0 0 1 1
use contact_19  contact_19_810
timestamp 1624857261
transform 1 0 72690 0 1 132001
box 0 0 1 1
use contact_14  contact_14_962
timestamp 1624857261
transform 1 0 72693 0 1 132000
box 0 0 1 1
use contact_7  contact_7_194
timestamp 1624857261
transform 1 0 72689 0 1 131996
box 0 0 1 1
use contact_13  contact_13_961
timestamp 1624857261
transform 1 0 73033 0 1 131992
box 0 0 1 1
use contact_14  contact_14_961
timestamp 1624857261
transform 1 0 73029 0 1 132000
box 0 0 1 1
use contact_13  contact_13_960
timestamp 1624857261
transform 1 0 73369 0 1 131992
box 0 0 1 1
use contact_14  contact_14_960
timestamp 1624857261
transform 1 0 73365 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3822
timestamp 1624857261
transform 1 0 72624 0 1 132469
box 0 0 1 1
use contact_13  contact_13_959
timestamp 1624857261
transform 1 0 73705 0 1 131992
box 0 0 1 1
use contact_14  contact_14_959
timestamp 1624857261
transform 1 0 73701 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3813
timestamp 1624857261
transform 1 0 74256 0 1 132061
box 0 0 1 1
use contact_13  contact_13_958
timestamp 1624857261
transform 1 0 74041 0 1 131992
box 0 0 1 1
use contact_14  contact_14_958
timestamp 1624857261
transform 1 0 74037 0 1 132000
box 0 0 1 1
use contact_13  contact_13_957
timestamp 1624857261
transform 1 0 74377 0 1 131992
box 0 0 1 1
use contact_13  contact_13_956
timestamp 1624857261
transform 1 0 74713 0 1 131992
box 0 0 1 1
use contact_19  contact_19_809
timestamp 1624857261
transform 1 0 74370 0 1 132001
box 0 0 1 1
use contact_14  contact_14_957
timestamp 1624857261
transform 1 0 74373 0 1 132000
box 0 0 1 1
use contact_14  contact_14_956
timestamp 1624857261
transform 1 0 74709 0 1 132000
box 0 0 1 1
use contact_7  contact_7_193
timestamp 1624857261
transform 1 0 74369 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3812
timestamp 1624857261
transform 1 0 74256 0 1 132469
box 0 0 1 1
use contact_13  contact_13_955
timestamp 1624857261
transform 1 0 75049 0 1 131992
box 0 0 1 1
use contact_14  contact_14_955
timestamp 1624857261
transform 1 0 75045 0 1 132000
box 0 0 1 1
use contact_13  contact_13_954
timestamp 1624857261
transform 1 0 75385 0 1 131992
box 0 0 1 1
use contact_13  contact_13_953
timestamp 1624857261
transform 1 0 75721 0 1 131992
box 0 0 1 1
use contact_14  contact_14_954
timestamp 1624857261
transform 1 0 75381 0 1 132000
box 0 0 1 1
use contact_14  contact_14_953
timestamp 1624857261
transform 1 0 75717 0 1 132000
box 0 0 1 1
use contact_13  contact_13_952
timestamp 1624857261
transform 1 0 76057 0 1 131992
box 0 0 1 1
use contact_19  contact_19_808
timestamp 1624857261
transform 1 0 76050 0 1 132001
box 0 0 1 1
use contact_14  contact_14_952
timestamp 1624857261
transform 1 0 76053 0 1 132000
box 0 0 1 1
use contact_7  contact_7_192
timestamp 1624857261
transform 1 0 76049 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3785
timestamp 1624857261
transform 1 0 76160 0 1 132061
box 0 0 1 1
use contact_13  contact_13_951
timestamp 1624857261
transform 1 0 76393 0 1 131992
box 0 0 1 1
use contact_14  contact_14_951
timestamp 1624857261
transform 1 0 76389 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3784
timestamp 1624857261
transform 1 0 76160 0 1 132469
box 0 0 1 1
use contact_13  contact_13_950
timestamp 1624857261
transform 1 0 76729 0 1 131992
box 0 0 1 1
use contact_14  contact_14_950
timestamp 1624857261
transform 1 0 76725 0 1 132000
box 0 0 1 1
use contact_13  contact_13_949
timestamp 1624857261
transform 1 0 77065 0 1 131992
box 0 0 1 1
use contact_14  contact_14_949
timestamp 1624857261
transform 1 0 77061 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3759
timestamp 1624857261
transform 1 0 77656 0 1 132061
box 0 0 1 1
use contact_13  contact_13_948
timestamp 1624857261
transform 1 0 77401 0 1 131992
box 0 0 1 1
use contact_14  contact_14_948
timestamp 1624857261
transform 1 0 77397 0 1 132000
box 0 0 1 1
use contact_13  contact_13_947
timestamp 1624857261
transform 1 0 77737 0 1 131992
box 0 0 1 1
use contact_19  contact_19_807
timestamp 1624857261
transform 1 0 77730 0 1 132001
box 0 0 1 1
use contact_14  contact_14_947
timestamp 1624857261
transform 1 0 77733 0 1 132000
box 0 0 1 1
use contact_7  contact_7_191
timestamp 1624857261
transform 1 0 77729 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3758
timestamp 1624857261
transform 1 0 77656 0 1 132469
box 0 0 1 1
use contact_14  contact_14_943
timestamp 1624857261
transform 1 0 79077 0 1 132000
box 0 0 1 1
use contact_14  contact_14_944
timestamp 1624857261
transform 1 0 78741 0 1 132000
box 0 0 1 1
use contact_14  contact_14_945
timestamp 1624857261
transform 1 0 78405 0 1 132000
box 0 0 1 1
use contact_14  contact_14_946
timestamp 1624857261
transform 1 0 78069 0 1 132000
box 0 0 1 1
use contact_13  contact_13_943
timestamp 1624857261
transform 1 0 79081 0 1 131992
box 0 0 1 1
use contact_13  contact_13_944
timestamp 1624857261
transform 1 0 78745 0 1 131992
box 0 0 1 1
use contact_13  contact_13_945
timestamp 1624857261
transform 1 0 78409 0 1 131992
box 0 0 1 1
use contact_13  contact_13_946
timestamp 1624857261
transform 1 0 78073 0 1 131992
box 0 0 1 1
use contact_13  contact_13_942
timestamp 1624857261
transform 1 0 79417 0 1 131992
box 0 0 1 1
use contact_13  contact_13_941
timestamp 1624857261
transform 1 0 79753 0 1 131992
box 0 0 1 1
use contact_13  contact_13_940
timestamp 1624857261
transform 1 0 80089 0 1 131992
box 0 0 1 1
use contact_13  contact_13_939
timestamp 1624857261
transform 1 0 80425 0 1 131992
box 0 0 1 1
use contact_33  contact_33_3747
timestamp 1624857261
transform 1 0 79288 0 1 132061
box 0 0 1 1
use contact_19  contact_19_806
timestamp 1624857261
transform 1 0 79410 0 1 132001
box 0 0 1 1
use contact_14  contact_14_942
timestamp 1624857261
transform 1 0 79413 0 1 132000
box 0 0 1 1
use contact_7  contact_7_190
timestamp 1624857261
transform 1 0 79409 0 1 131996
box 0 0 1 1
use contact_14  contact_14_941
timestamp 1624857261
transform 1 0 79749 0 1 132000
box 0 0 1 1
use contact_14  contact_14_940
timestamp 1624857261
transform 1 0 80085 0 1 132000
box 0 0 1 1
use contact_14  contact_14_939
timestamp 1624857261
transform 1 0 80421 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3746
timestamp 1624857261
transform 1 0 79288 0 1 132469
box 0 0 1 1
use contact_13  contact_13_938
timestamp 1624857261
transform 1 0 80761 0 1 131992
box 0 0 1 1
use contact_14  contact_14_938
timestamp 1624857261
transform 1 0 80757 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3723
timestamp 1624857261
transform 1 0 81192 0 1 132061
box 0 0 1 1
use contact_13  contact_13_937
timestamp 1624857261
transform 1 0 81097 0 1 131992
box 0 0 1 1
use contact_19  contact_19_805
timestamp 1624857261
transform 1 0 81090 0 1 132001
box 0 0 1 1
use contact_14  contact_14_937
timestamp 1624857261
transform 1 0 81093 0 1 132000
box 0 0 1 1
use contact_7  contact_7_189
timestamp 1624857261
transform 1 0 81089 0 1 131996
box 0 0 1 1
use contact_13  contact_13_936
timestamp 1624857261
transform 1 0 81433 0 1 131992
box 0 0 1 1
use contact_13  contact_13_935
timestamp 1624857261
transform 1 0 81769 0 1 131992
box 0 0 1 1
use contact_14  contact_14_936
timestamp 1624857261
transform 1 0 81429 0 1 132000
box 0 0 1 1
use contact_14  contact_14_935
timestamp 1624857261
transform 1 0 81765 0 1 132000
box 0 0 1 1
use contact_13  contact_13_934
timestamp 1624857261
transform 1 0 82105 0 1 131992
box 0 0 1 1
use contact_14  contact_14_934
timestamp 1624857261
transform 1 0 82101 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3722
timestamp 1624857261
transform 1 0 81192 0 1 132469
box 0 0 1 1
use contact_13  contact_13_933
timestamp 1624857261
transform 1 0 82441 0 1 131992
box 0 0 1 1
use contact_13  contact_13_932
timestamp 1624857261
transform 1 0 82777 0 1 131992
box 0 0 1 1
use contact_13  contact_13_931
timestamp 1624857261
transform 1 0 83113 0 1 131992
box 0 0 1 1
use contact_13  contact_13_930
timestamp 1624857261
transform 1 0 83449 0 1 131992
box 0 0 1 1
use contact_14  contact_14_933
timestamp 1624857261
transform 1 0 82437 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3703
timestamp 1624857261
transform 1 0 82688 0 1 132061
box 0 0 1 1
use contact_19  contact_19_804
timestamp 1624857261
transform 1 0 82770 0 1 132001
box 0 0 1 1
use contact_14  contact_14_932
timestamp 1624857261
transform 1 0 82773 0 1 132000
box 0 0 1 1
use contact_7  contact_7_188
timestamp 1624857261
transform 1 0 82769 0 1 131996
box 0 0 1 1
use contact_14  contact_14_931
timestamp 1624857261
transform 1 0 83109 0 1 132000
box 0 0 1 1
use contact_14  contact_14_930
timestamp 1624857261
transform 1 0 83445 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3702
timestamp 1624857261
transform 1 0 82688 0 1 132469
box 0 0 1 1
use contact_13  contact_13_929
timestamp 1624857261
transform 1 0 83785 0 1 131992
box 0 0 1 1
use contact_13  contact_13_928
timestamp 1624857261
transform 1 0 84121 0 1 131992
box 0 0 1 1
use contact_13  contact_13_927
timestamp 1624857261
transform 1 0 84457 0 1 131992
box 0 0 1 1
use contact_13  contact_13_926
timestamp 1624857261
transform 1 0 84793 0 1 131992
box 0 0 1 1
use contact_14  contact_14_929
timestamp 1624857261
transform 1 0 83781 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3685
timestamp 1624857261
transform 1 0 84320 0 1 132061
box 0 0 1 1
use contact_19  contact_19_803
timestamp 1624857261
transform 1 0 84450 0 1 132001
box 0 0 1 1
use contact_14  contact_14_928
timestamp 1624857261
transform 1 0 84117 0 1 132000
box 0 0 1 1
use contact_14  contact_14_927
timestamp 1624857261
transform 1 0 84453 0 1 132000
box 0 0 1 1
use contact_7  contact_7_187
timestamp 1624857261
transform 1 0 84449 0 1 131996
box 0 0 1 1
use contact_14  contact_14_926
timestamp 1624857261
transform 1 0 84789 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3684
timestamp 1624857261
transform 1 0 84320 0 1 132469
box 0 0 1 1
use contact_13  contact_13_925
timestamp 1624857261
transform 1 0 85129 0 1 131992
box 0 0 1 1
use contact_13  contact_13_924
timestamp 1624857261
transform 1 0 85465 0 1 131992
box 0 0 1 1
use contact_14  contact_14_925
timestamp 1624857261
transform 1 0 85125 0 1 132000
box 0 0 1 1
use contact_14  contact_14_924
timestamp 1624857261
transform 1 0 85461 0 1 132000
box 0 0 1 1
use contact_13  contact_13_923
timestamp 1624857261
transform 1 0 85801 0 1 131992
box 0 0 1 1
use contact_14  contact_14_923
timestamp 1624857261
transform 1 0 85797 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3661
timestamp 1624857261
transform 1 0 86088 0 1 132061
box 0 0 1 1
use contact_13  contact_13_922
timestamp 1624857261
transform 1 0 86137 0 1 131992
box 0 0 1 1
use contact_19  contact_19_802
timestamp 1624857261
transform 1 0 86130 0 1 132001
box 0 0 1 1
use contact_14  contact_14_922
timestamp 1624857261
transform 1 0 86133 0 1 132000
box 0 0 1 1
use contact_7  contact_7_186
timestamp 1624857261
transform 1 0 86129 0 1 131996
box 0 0 1 1
use contact_13  contact_13_921
timestamp 1624857261
transform 1 0 86473 0 1 131992
box 0 0 1 1
use contact_14  contact_14_921
timestamp 1624857261
transform 1 0 86469 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3660
timestamp 1624857261
transform 1 0 86088 0 1 132469
box 0 0 1 1
use contact_13  contact_13_920
timestamp 1624857261
transform 1 0 86809 0 1 131992
box 0 0 1 1
use contact_13  contact_13_919
timestamp 1624857261
transform 1 0 87145 0 1 131992
box 0 0 1 1
use contact_13  contact_13_918
timestamp 1624857261
transform 1 0 87481 0 1 131992
box 0 0 1 1
use contact_13  contact_13_917
timestamp 1624857261
transform 1 0 87817 0 1 131992
box 0 0 1 1
use contact_14  contact_14_920
timestamp 1624857261
transform 1 0 86805 0 1 132000
box 0 0 1 1
use contact_14  contact_14_919
timestamp 1624857261
transform 1 0 87141 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3637
timestamp 1624857261
transform 1 0 87720 0 1 132061
box 0 0 1 1
use contact_19  contact_19_801
timestamp 1624857261
transform 1 0 87810 0 1 132001
box 0 0 1 1
use contact_14  contact_14_918
timestamp 1624857261
transform 1 0 87477 0 1 132000
box 0 0 1 1
use contact_14  contact_14_917
timestamp 1624857261
transform 1 0 87813 0 1 132000
box 0 0 1 1
use contact_7  contact_7_185
timestamp 1624857261
transform 1 0 87809 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3636
timestamp 1624857261
transform 1 0 87720 0 1 132469
box 0 0 1 1
use contact_13  contact_13_916
timestamp 1624857261
transform 1 0 88153 0 1 131992
box 0 0 1 1
use contact_13  contact_13_915
timestamp 1624857261
transform 1 0 88489 0 1 131992
box 0 0 1 1
use contact_13  contact_13_914
timestamp 1624857261
transform 1 0 88825 0 1 131992
box 0 0 1 1
use contact_13  contact_13_913
timestamp 1624857261
transform 1 0 89161 0 1 131992
box 0 0 1 1
use contact_13  contact_13_912
timestamp 1624857261
transform 1 0 89497 0 1 131992
box 0 0 1 1
use contact_14  contact_14_916
timestamp 1624857261
transform 1 0 88149 0 1 132000
box 0 0 1 1
use contact_14  contact_14_915
timestamp 1624857261
transform 1 0 88485 0 1 132000
box 0 0 1 1
use contact_14  contact_14_914
timestamp 1624857261
transform 1 0 88821 0 1 132000
box 0 0 1 1
use contact_14  contact_14_913
timestamp 1624857261
transform 1 0 89157 0 1 132000
box 0 0 1 1
use contact_19  contact_19_800
timestamp 1624857261
transform 1 0 89490 0 1 132001
box 0 0 1 1
use contact_14  contact_14_912
timestamp 1624857261
transform 1 0 89493 0 1 132000
box 0 0 1 1
use contact_7  contact_7_184
timestamp 1624857261
transform 1 0 89489 0 1 131996
box 0 0 1 1
use contact_14  contact_14_909
timestamp 1624857261
transform 1 0 90501 0 1 132000
box 0 0 1 1
use contact_14  contact_14_910
timestamp 1624857261
transform 1 0 90165 0 1 132000
box 0 0 1 1
use contact_14  contact_14_911
timestamp 1624857261
transform 1 0 89829 0 1 132000
box 0 0 1 1
use contact_13  contact_13_909
timestamp 1624857261
transform 1 0 90505 0 1 131992
box 0 0 1 1
use contact_13  contact_13_910
timestamp 1624857261
transform 1 0 90169 0 1 131992
box 0 0 1 1
use contact_13  contact_13_911
timestamp 1624857261
transform 1 0 89833 0 1 131992
box 0 0 1 1
use contact_33  contact_33_3626
timestamp 1624857261
transform 1 0 89760 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3627
timestamp 1624857261
transform 1 0 89760 0 1 132061
box 0 0 1 1
use contact_13  contact_13_908
timestamp 1624857261
transform 1 0 90841 0 1 131992
box 0 0 1 1
use contact_13  contact_13_907
timestamp 1624857261
transform 1 0 91177 0 1 131992
box 0 0 1 1
use contact_13  contact_13_906
timestamp 1624857261
transform 1 0 91513 0 1 131992
box 0 0 1 1
use contact_13  contact_13_905
timestamp 1624857261
transform 1 0 91849 0 1 131992
box 0 0 1 1
use contact_14  contact_14_908
timestamp 1624857261
transform 1 0 90837 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3605
timestamp 1624857261
transform 1 0 91120 0 1 132061
box 0 0 1 1
use contact_19  contact_19_799
timestamp 1624857261
transform 1 0 91170 0 1 132001
box 0 0 1 1
use contact_14  contact_14_907
timestamp 1624857261
transform 1 0 91173 0 1 132000
box 0 0 1 1
use contact_14  contact_14_906
timestamp 1624857261
transform 1 0 91509 0 1 132000
box 0 0 1 1
use contact_7  contact_7_183
timestamp 1624857261
transform 1 0 91169 0 1 131996
box 0 0 1 1
use contact_14  contact_14_905
timestamp 1624857261
transform 1 0 91845 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3604
timestamp 1624857261
transform 1 0 91120 0 1 132469
box 0 0 1 1
use contact_13  contact_13_904
timestamp 1624857261
transform 1 0 92185 0 1 131992
box 0 0 1 1
use contact_13  contact_13_903
timestamp 1624857261
transform 1 0 92521 0 1 131992
box 0 0 1 1
use contact_14  contact_14_904
timestamp 1624857261
transform 1 0 92181 0 1 132000
box 0 0 1 1
use contact_14  contact_14_903
timestamp 1624857261
transform 1 0 92517 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3587
timestamp 1624857261
transform 1 0 92888 0 1 132061
box 0 0 1 1
use contact_13  contact_13_902
timestamp 1624857261
transform 1 0 92857 0 1 131992
box 0 0 1 1
use contact_19  contact_19_798
timestamp 1624857261
transform 1 0 92850 0 1 132001
box 0 0 1 1
use contact_14  contact_14_902
timestamp 1624857261
transform 1 0 92853 0 1 132000
box 0 0 1 1
use contact_7  contact_7_182
timestamp 1624857261
transform 1 0 92849 0 1 131996
box 0 0 1 1
use contact_13  contact_13_901
timestamp 1624857261
transform 1 0 93193 0 1 131992
box 0 0 1 1
use contact_14  contact_14_901
timestamp 1624857261
transform 1 0 93189 0 1 132000
box 0 0 1 1
use contact_13  contact_13_900
timestamp 1624857261
transform 1 0 93529 0 1 131992
box 0 0 1 1
use contact_14  contact_14_900
timestamp 1624857261
transform 1 0 93525 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3586
timestamp 1624857261
transform 1 0 92888 0 1 132469
box 0 0 1 1
use contact_13  contact_13_899
timestamp 1624857261
transform 1 0 93865 0 1 131992
box 0 0 1 1
use contact_13  contact_13_898
timestamp 1624857261
transform 1 0 94201 0 1 131992
box 0 0 1 1
use contact_13  contact_13_897
timestamp 1624857261
transform 1 0 94537 0 1 131992
box 0 0 1 1
use contact_13  contact_13_896
timestamp 1624857261
transform 1 0 94873 0 1 131992
box 0 0 1 1
use contact_14  contact_14_899
timestamp 1624857261
transform 1 0 93861 0 1 132000
box 0 0 1 1
use contact_14  contact_14_898
timestamp 1624857261
transform 1 0 94197 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3573
timestamp 1624857261
transform 1 0 94656 0 1 132061
box 0 0 1 1
use contact_19  contact_19_797
timestamp 1624857261
transform 1 0 94530 0 1 132001
box 0 0 1 1
use contact_14  contact_14_897
timestamp 1624857261
transform 1 0 94533 0 1 132000
box 0 0 1 1
use contact_14  contact_14_896
timestamp 1624857261
transform 1 0 94869 0 1 132000
box 0 0 1 1
use contact_7  contact_7_181
timestamp 1624857261
transform 1 0 94529 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3572
timestamp 1624857261
transform 1 0 94656 0 1 132469
box 0 0 1 1
use contact_13  contact_13_895
timestamp 1624857261
transform 1 0 95209 0 1 131992
box 0 0 1 1
use contact_14  contact_14_895
timestamp 1624857261
transform 1 0 95205 0 1 132000
box 0 0 1 1
use contact_14  contact_14_894
timestamp 1624857261
transform 1 0 95541 0 1 132000
box 0 0 1 1
use contact_13  contact_13_894
timestamp 1624857261
transform 1 0 95545 0 1 131992
box 0 0 1 1
use contact_13  contact_13_893
timestamp 1624857261
transform 1 0 95881 0 1 131992
box 0 0 1 1
use contact_14  contact_14_893
timestamp 1624857261
transform 1 0 95877 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3557
timestamp 1624857261
transform 1 0 96152 0 1 132061
box 0 0 1 1
use contact_13  contact_13_892
timestamp 1624857261
transform 1 0 96217 0 1 131992
box 0 0 1 1
use contact_19  contact_19_796
timestamp 1624857261
transform 1 0 96210 0 1 132001
box 0 0 1 1
use contact_14  contact_14_892
timestamp 1624857261
transform 1 0 96213 0 1 132000
box 0 0 1 1
use contact_7  contact_7_180
timestamp 1624857261
transform 1 0 96209 0 1 131996
box 0 0 1 1
use contact_13  contact_13_891
timestamp 1624857261
transform 1 0 96553 0 1 131992
box 0 0 1 1
use contact_14  contact_14_891
timestamp 1624857261
transform 1 0 96549 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3556
timestamp 1624857261
transform 1 0 96152 0 1 132469
box 0 0 1 1
use contact_13  contact_13_890
timestamp 1624857261
transform 1 0 96889 0 1 131992
box 0 0 1 1
use contact_13  contact_13_889
timestamp 1624857261
transform 1 0 97225 0 1 131992
box 0 0 1 1
use contact_13  contact_13_888
timestamp 1624857261
transform 1 0 97561 0 1 131992
box 0 0 1 1
use contact_13  contact_13_887
timestamp 1624857261
transform 1 0 97897 0 1 131992
box 0 0 1 1
use contact_14  contact_14_890
timestamp 1624857261
transform 1 0 96885 0 1 132000
box 0 0 1 1
use contact_14  contact_14_889
timestamp 1624857261
transform 1 0 97221 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3535
timestamp 1624857261
transform 1 0 97920 0 1 132061
box 0 0 1 1
use contact_19  contact_19_795
timestamp 1624857261
transform 1 0 97890 0 1 132001
box 0 0 1 1
use contact_14  contact_14_888
timestamp 1624857261
transform 1 0 97557 0 1 132000
box 0 0 1 1
use contact_14  contact_14_887
timestamp 1624857261
transform 1 0 97893 0 1 132000
box 0 0 1 1
use contact_7  contact_7_179
timestamp 1624857261
transform 1 0 97889 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3534
timestamp 1624857261
transform 1 0 97920 0 1 132469
box 0 0 1 1
use contact_13  contact_13_886
timestamp 1624857261
transform 1 0 98233 0 1 131992
box 0 0 1 1
use contact_13  contact_13_885
timestamp 1624857261
transform 1 0 98569 0 1 131992
box 0 0 1 1
use contact_13  contact_13_884
timestamp 1624857261
transform 1 0 98905 0 1 131992
box 0 0 1 1
use contact_13  contact_13_883
timestamp 1624857261
transform 1 0 99241 0 1 131992
box 0 0 1 1
use contact_13  contact_13_882
timestamp 1624857261
transform 1 0 99577 0 1 131992
box 0 0 1 1
use contact_14  contact_14_886
timestamp 1624857261
transform 1 0 98229 0 1 132000
box 0 0 1 1
use contact_14  contact_14_885
timestamp 1624857261
transform 1 0 98565 0 1 132000
box 0 0 1 1
use contact_14  contact_14_884
timestamp 1624857261
transform 1 0 98901 0 1 132000
box 0 0 1 1
use contact_14  contact_14_883
timestamp 1624857261
transform 1 0 99237 0 1 132000
box 0 0 1 1
use contact_19  contact_19_794
timestamp 1624857261
transform 1 0 99570 0 1 132001
box 0 0 1 1
use contact_14  contact_14_882
timestamp 1624857261
transform 1 0 99573 0 1 132000
box 0 0 1 1
use contact_7  contact_7_178
timestamp 1624857261
transform 1 0 99569 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3521
timestamp 1624857261
transform 1 0 99688 0 1 132061
box 0 0 1 1
use contact_13  contact_13_881
timestamp 1624857261
transform 1 0 99913 0 1 131992
box 0 0 1 1
use contact_14  contact_14_881
timestamp 1624857261
transform 1 0 99909 0 1 132000
box 0 0 1 1
use contact_13  contact_13_880
timestamp 1624857261
transform 1 0 100249 0 1 131992
box 0 0 1 1
use contact_14  contact_14_880
timestamp 1624857261
transform 1 0 100245 0 1 132000
box 0 0 1 1
use contact_13  contact_13_879
timestamp 1624857261
transform 1 0 100585 0 1 131992
box 0 0 1 1
use contact_13  contact_13_878
timestamp 1624857261
transform 1 0 100921 0 1 131992
box 0 0 1 1
use contact_14  contact_14_879
timestamp 1624857261
transform 1 0 100581 0 1 132000
box 0 0 1 1
use contact_14  contact_14_878
timestamp 1624857261
transform 1 0 100917 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3520
timestamp 1624857261
transform 1 0 99688 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3505
timestamp 1624857261
transform 1 0 101184 0 1 132061
box 0 0 1 1
use contact_13  contact_13_877
timestamp 1624857261
transform 1 0 101257 0 1 131992
box 0 0 1 1
use contact_19  contact_19_793
timestamp 1624857261
transform 1 0 101250 0 1 132001
box 0 0 1 1
use contact_14  contact_14_877
timestamp 1624857261
transform 1 0 101253 0 1 132000
box 0 0 1 1
use contact_7  contact_7_177
timestamp 1624857261
transform 1 0 101249 0 1 131996
box 0 0 1 1
use contact_13  contact_13_876
timestamp 1624857261
transform 1 0 101593 0 1 131992
box 0 0 1 1
use contact_13  contact_13_875
timestamp 1624857261
transform 1 0 101929 0 1 131992
box 0 0 1 1
use contact_14  contact_14_876
timestamp 1624857261
transform 1 0 101589 0 1 132000
box 0 0 1 1
use contact_14  contact_14_875
timestamp 1624857261
transform 1 0 101925 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3504
timestamp 1624857261
transform 1 0 101184 0 1 132469
box 0 0 1 1
use contact_13  contact_13_874
timestamp 1624857261
transform 1 0 102265 0 1 131992
box 0 0 1 1
use contact_13  contact_13_873
timestamp 1624857261
transform 1 0 102601 0 1 131992
box 0 0 1 1
use contact_14  contact_14_874
timestamp 1624857261
transform 1 0 102261 0 1 132000
box 0 0 1 1
use contact_14  contact_14_873
timestamp 1624857261
transform 1 0 102597 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3481
timestamp 1624857261
transform 1 0 102952 0 1 132061
box 0 0 1 1
use contact_13  contact_13_872
timestamp 1624857261
transform 1 0 102937 0 1 131992
box 0 0 1 1
use contact_19  contact_19_792
timestamp 1624857261
transform 1 0 102930 0 1 132001
box 0 0 1 1
use contact_14  contact_14_872
timestamp 1624857261
transform 1 0 102933 0 1 132000
box 0 0 1 1
use contact_7  contact_7_176
timestamp 1624857261
transform 1 0 102929 0 1 131996
box 0 0 1 1
use contact_13  contact_13_871
timestamp 1624857261
transform 1 0 103273 0 1 131992
box 0 0 1 1
use contact_14  contact_14_871
timestamp 1624857261
transform 1 0 103269 0 1 132000
box 0 0 1 1
use contact_13  contact_13_870
timestamp 1624857261
transform 1 0 103609 0 1 131992
box 0 0 1 1
use contact_14  contact_14_870
timestamp 1624857261
transform 1 0 103605 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3480
timestamp 1624857261
transform 1 0 102952 0 1 132469
box 0 0 1 1
use contact_13  contact_13_869
timestamp 1624857261
transform 1 0 103945 0 1 131992
box 0 0 1 1
use contact_14  contact_14_869
timestamp 1624857261
transform 1 0 103941 0 1 132000
box 0 0 1 1
use contact_13  contact_13_868
timestamp 1624857261
transform 1 0 104281 0 1 131992
box 0 0 1 1
use contact_14  contact_14_868
timestamp 1624857261
transform 1 0 104277 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3463
timestamp 1624857261
transform 1 0 104720 0 1 132061
box 0 0 1 1
use contact_13  contact_13_867
timestamp 1624857261
transform 1 0 104617 0 1 131992
box 0 0 1 1
use contact_13  contact_13_866
timestamp 1624857261
transform 1 0 104953 0 1 131992
box 0 0 1 1
use contact_19  contact_19_791
timestamp 1624857261
transform 1 0 104610 0 1 132001
box 0 0 1 1
use contact_14  contact_14_867
timestamp 1624857261
transform 1 0 104613 0 1 132000
box 0 0 1 1
use contact_14  contact_14_866
timestamp 1624857261
transform 1 0 104949 0 1 132000
box 0 0 1 1
use contact_7  contact_7_175
timestamp 1624857261
transform 1 0 104609 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3462
timestamp 1624857261
transform 1 0 104720 0 1 132469
box 0 0 1 1
use contact_13  contact_13_865
timestamp 1624857261
transform 1 0 105289 0 1 131992
box 0 0 1 1
use contact_14  contact_14_865
timestamp 1624857261
transform 1 0 105285 0 1 132000
box 0 0 1 1
use contact_13  contact_13_864
timestamp 1624857261
transform 1 0 105625 0 1 131992
box 0 0 1 1
use contact_13  contact_13_863
timestamp 1624857261
transform 1 0 105961 0 1 131992
box 0 0 1 1
use contact_14  contact_14_864
timestamp 1624857261
transform 1 0 105621 0 1 132000
box 0 0 1 1
use contact_14  contact_14_863
timestamp 1624857261
transform 1 0 105957 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3447
timestamp 1624857261
transform 1 0 106216 0 1 132061
box 0 0 1 1
use contact_13  contact_13_862
timestamp 1624857261
transform 1 0 106297 0 1 131992
box 0 0 1 1
use contact_19  contact_19_790
timestamp 1624857261
transform 1 0 106290 0 1 132001
box 0 0 1 1
use contact_14  contact_14_862
timestamp 1624857261
transform 1 0 106293 0 1 132000
box 0 0 1 1
use contact_7  contact_7_174
timestamp 1624857261
transform 1 0 106289 0 1 131996
box 0 0 1 1
use contact_14  contact_14_861
timestamp 1624857261
transform 1 0 106629 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3446
timestamp 1624857261
transform 1 0 106216 0 1 132469
box 0 0 1 1
use contact_13  contact_13_861
timestamp 1624857261
transform 1 0 106633 0 1 131992
box 0 0 1 1
use contact_13  contact_13_860
timestamp 1624857261
transform 1 0 106969 0 1 131992
box 0 0 1 1
use contact_14  contact_14_860
timestamp 1624857261
transform 1 0 106965 0 1 132000
box 0 0 1 1
use contact_13  contact_13_859
timestamp 1624857261
transform 1 0 107305 0 1 131992
box 0 0 1 1
use contact_14  contact_14_859
timestamp 1624857261
transform 1 0 107301 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3427
timestamp 1624857261
transform 1 0 107848 0 1 132061
box 0 0 1 1
use contact_13  contact_13_858
timestamp 1624857261
transform 1 0 107641 0 1 131992
box 0 0 1 1
use contact_14  contact_14_858
timestamp 1624857261
transform 1 0 107637 0 1 132000
box 0 0 1 1
use contact_13  contact_13_857
timestamp 1624857261
transform 1 0 107977 0 1 131992
box 0 0 1 1
use contact_19  contact_19_789
timestamp 1624857261
transform 1 0 107970 0 1 132001
box 0 0 1 1
use contact_14  contact_14_857
timestamp 1624857261
transform 1 0 107973 0 1 132000
box 0 0 1 1
use contact_7  contact_7_173
timestamp 1624857261
transform 1 0 107969 0 1 131996
box 0 0 1 1
use contact_33  contact_33_3426
timestamp 1624857261
transform 1 0 107848 0 1 132469
box 0 0 1 1
use contact_14  contact_14_853
timestamp 1624857261
transform 1 0 109317 0 1 132000
box 0 0 1 1
use contact_14  contact_14_854
timestamp 1624857261
transform 1 0 108981 0 1 132000
box 0 0 1 1
use contact_14  contact_14_855
timestamp 1624857261
transform 1 0 108645 0 1 132000
box 0 0 1 1
use contact_14  contact_14_856
timestamp 1624857261
transform 1 0 108309 0 1 132000
box 0 0 1 1
use contact_13  contact_13_853
timestamp 1624857261
transform 1 0 109321 0 1 131992
box 0 0 1 1
use contact_13  contact_13_854
timestamp 1624857261
transform 1 0 108985 0 1 131992
box 0 0 1 1
use contact_13  contact_13_855
timestamp 1624857261
transform 1 0 108649 0 1 131992
box 0 0 1 1
use contact_13  contact_13_856
timestamp 1624857261
transform 1 0 108313 0 1 131992
box 0 0 1 1
use contact_33  contact_33_3413
timestamp 1624857261
transform 1 0 109616 0 1 132061
box 0 0 1 1
use contact_13  contact_13_852
timestamp 1624857261
transform 1 0 109657 0 1 131992
box 0 0 1 1
use contact_19  contact_19_788
timestamp 1624857261
transform 1 0 109650 0 1 132001
box 0 0 1 1
use contact_14  contact_14_852
timestamp 1624857261
transform 1 0 109653 0 1 132000
box 0 0 1 1
use contact_7  contact_7_172
timestamp 1624857261
transform 1 0 109649 0 1 131996
box 0 0 1 1
use contact_13  contact_13_851
timestamp 1624857261
transform 1 0 109993 0 1 131992
box 0 0 1 1
use contact_13  contact_13_850
timestamp 1624857261
transform 1 0 110329 0 1 131992
box 0 0 1 1
use contact_14  contact_14_851
timestamp 1624857261
transform 1 0 109989 0 1 132000
box 0 0 1 1
use contact_14  contact_14_850
timestamp 1624857261
transform 1 0 110325 0 1 132000
box 0 0 1 1
use contact_13  contact_13_849
timestamp 1624857261
transform 1 0 110665 0 1 131992
box 0 0 1 1
use contact_14  contact_14_849
timestamp 1624857261
transform 1 0 110661 0 1 132000
box 0 0 1 1
use contact_13  contact_13_848
timestamp 1624857261
transform 1 0 111001 0 1 131992
box 0 0 1 1
use contact_14  contact_14_848
timestamp 1624857261
transform 1 0 110997 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3412
timestamp 1624857261
transform 1 0 109616 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3409
timestamp 1624857261
transform 1 0 111384 0 1 132061
box 0 0 1 1
use contact_13  contact_13_847
timestamp 1624857261
transform 1 0 111337 0 1 131992
box 0 0 1 1
use contact_19  contact_19_787
timestamp 1624857261
transform 1 0 111330 0 1 132001
box 0 0 1 1
use contact_14  contact_14_847
timestamp 1624857261
transform 1 0 111333 0 1 132000
box 0 0 1 1
use contact_7  contact_7_171
timestamp 1624857261
transform 1 0 111329 0 1 131996
box 0 0 1 1
use contact_13  contact_13_846
timestamp 1624857261
transform 1 0 111673 0 1 131992
box 0 0 1 1
use contact_14  contact_14_846
timestamp 1624857261
transform 1 0 111669 0 1 132000
box 0 0 1 1
use contact_13  contact_13_845
timestamp 1624857261
transform 1 0 112009 0 1 131992
box 0 0 1 1
use contact_14  contact_14_845
timestamp 1624857261
transform 1 0 112005 0 1 132000
box 0 0 1 1
use contact_13  contact_13_844
timestamp 1624857261
transform 1 0 112345 0 1 131992
box 0 0 1 1
use contact_14  contact_14_844
timestamp 1624857261
transform 1 0 112341 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3408
timestamp 1624857261
transform 1 0 111384 0 1 132469
box 0 0 1 1
use contact_33  contact_33_3405
timestamp 1624857261
transform 1 0 112880 0 1 132061
box 0 0 1 1
use contact_13  contact_13_843
timestamp 1624857261
transform 1 0 112681 0 1 131992
box 0 0 1 1
use contact_14  contact_14_843
timestamp 1624857261
transform 1 0 112677 0 1 132000
box 0 0 1 1
use contact_13  contact_13_842
timestamp 1624857261
transform 1 0 113017 0 1 131992
box 0 0 1 1
use contact_13  contact_13_841
timestamp 1624857261
transform 1 0 113353 0 1 131992
box 0 0 1 1
use contact_19  contact_19_786
timestamp 1624857261
transform 1 0 113010 0 1 132001
box 0 0 1 1
use contact_14  contact_14_842
timestamp 1624857261
transform 1 0 113013 0 1 132000
box 0 0 1 1
use contact_14  contact_14_841
timestamp 1624857261
transform 1 0 113349 0 1 132000
box 0 0 1 1
use contact_7  contact_7_170
timestamp 1624857261
transform 1 0 113009 0 1 131996
box 0 0 1 1
use contact_13  contact_13_840
timestamp 1624857261
transform 1 0 113689 0 1 131992
box 0 0 1 1
use contact_14  contact_14_840
timestamp 1624857261
transform 1 0 113685 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3404
timestamp 1624857261
transform 1 0 112880 0 1 132469
box 0 0 1 1
use contact_33  contact_33_2532
timestamp 1624857261
transform 1 0 119408 0 1 129885
box 0 0 1 1
use contact_7  contact_7_326
timestamp 1624857261
transform 1 0 119937 0 1 130760
box 0 0 1 1
use contact_33  contact_33_2513
timestamp 1624857261
transform 1 0 119680 0 1 130021
box 0 0 1 1
use contact_33  contact_33_5489
timestamp 1624857261
transform 1 0 119952 0 1 130837
box 0 0 1 1
use col_addr_dff  col_addr_dff_0
timestamp 1624857261
transform -1 0 121308 0 -1 131361
box -36 -49 1204 1467
use contact_7  contact_7_327
timestamp 1624857261
transform 1 0 121105 0 1 130760
box 0 0 1 1
use contact_33  contact_33_5490
timestamp 1624857261
transform 1 0 121176 0 1 130837
box 0 0 1 1
use contact_32  contact_32_0
timestamp 1624857261
transform 1 0 123527 0 1 131016
box 0 0 1 1
use contact_33  contact_33_18
timestamp 1624857261
transform 1 0 123624 0 1 130429
box 0 0 1 1
use contact_33  contact_33_19
timestamp 1624857261
transform 1 0 123760 0 1 130293
box 0 0 1 1
use contact_33  contact_33_2491
timestamp 1624857261
transform 1 0 123624 0 1 129885
box 0 0 1 1
use contact_13  contact_13_839
timestamp 1624857261
transform 1 0 114025 0 1 131992
box 0 0 1 1
use contact_14  contact_14_839
timestamp 1624857261
transform 1 0 114021 0 1 132000
box 0 0 1 1
use contact_13  contact_13_838
timestamp 1624857261
transform 1 0 114361 0 1 131992
box 0 0 1 1
use contact_14  contact_14_838
timestamp 1624857261
transform 1 0 114357 0 1 132000
box 0 0 1 1
use contact_13  contact_13_837
timestamp 1624857261
transform 1 0 114697 0 1 131992
box 0 0 1 1
use contact_19  contact_19_785
timestamp 1624857261
transform 1 0 114690 0 1 132001
box 0 0 1 1
use contact_14  contact_14_837
timestamp 1624857261
transform 1 0 114693 0 1 132000
box 0 0 1 1
use contact_7  contact_7_169
timestamp 1624857261
transform 1 0 114689 0 1 131996
box 0 0 1 1
use contact_13  contact_13_836
timestamp 1624857261
transform 1 0 115033 0 1 131992
box 0 0 1 1
use contact_14  contact_14_836
timestamp 1624857261
transform 1 0 115029 0 1 132000
box 0 0 1 1
use contact_33  contact_33_3401
timestamp 1624857261
transform 1 0 114648 0 1 132061
box 0 0 1 1
use contact_33  contact_33_3400
timestamp 1624857261
transform 1 0 114648 0 1 132469
box 0 0 1 1
use contact_13  contact_13_835
timestamp 1624857261
transform 1 0 115369 0 1 131992
box 0 0 1 1
use contact_14  contact_14_835
timestamp 1624857261
transform 1 0 115365 0 1 132000
box 0 0 1 1
use contact_13  contact_13_834
timestamp 1624857261
transform 1 0 115705 0 1 131992
box 0 0 1 1
use contact_14  contact_14_834
timestamp 1624857261
transform 1 0 115701 0 1 132000
box 0 0 1 1
use contact_13  contact_13_833
timestamp 1624857261
transform 1 0 116041 0 1 131992
box 0 0 1 1
use contact_13  contact_13_832
timestamp 1624857261
transform 1 0 116377 0 1 131992
box 0 0 1 1
use contact_19  contact_19_784
timestamp 1624857261
transform 1 0 116370 0 1 132001
box 0 0 1 1
use contact_14  contact_14_833
timestamp 1624857261
transform 1 0 116037 0 1 132000
box 0 0 1 1
use contact_14  contact_14_832
timestamp 1624857261
transform 1 0 116373 0 1 132000
box 0 0 1 1
use contact_7  contact_7_168
timestamp 1624857261
transform 1 0 116369 0 1 131996
box 0 0 1 1
use contact_33  contact_33_2693
timestamp 1624857261
transform 1 0 116416 0 1 132061
box 0 0 1 1
use contact_33  contact_33_2692
timestamp 1624857261
transform 1 0 116416 0 1 132469
box 0 0 1 1
use contact_13  contact_13_831
timestamp 1624857261
transform 1 0 116713 0 1 131992
box 0 0 1 1
use contact_14  contact_14_831
timestamp 1624857261
transform 1 0 116709 0 1 132000
box 0 0 1 1
use contact_13  contact_13_830
timestamp 1624857261
transform 1 0 117049 0 1 131992
box 0 0 1 1
use contact_13  contact_13_829
timestamp 1624857261
transform 1 0 117385 0 1 131992
box 0 0 1 1
use contact_14  contact_14_830
timestamp 1624857261
transform 1 0 117045 0 1 132000
box 0 0 1 1
use contact_14  contact_14_829
timestamp 1624857261
transform 1 0 117381 0 1 132000
box 0 0 1 1
use contact_13  contact_13_828
timestamp 1624857261
transform 1 0 117721 0 1 131992
box 0 0 1 1
use contact_14  contact_14_828
timestamp 1624857261
transform 1 0 117717 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2531
timestamp 1624857261
transform 1 0 117912 0 1 132061
box 0 0 1 1
use contact_13  contact_13_827
timestamp 1624857261
transform 1 0 118057 0 1 131992
box 0 0 1 1
use contact_19  contact_19_783
timestamp 1624857261
transform 1 0 118050 0 1 132001
box 0 0 1 1
use contact_14  contact_14_827
timestamp 1624857261
transform 1 0 118053 0 1 132000
box 0 0 1 1
use contact_7  contact_7_167
timestamp 1624857261
transform 1 0 118049 0 1 131996
box 0 0 1 1
use contact_33  contact_33_2530
timestamp 1624857261
transform 1 0 117912 0 1 132469
box 0 0 1 1
use contact_14  contact_14_823
timestamp 1624857261
transform 1 0 119397 0 1 132000
box 0 0 1 1
use contact_14  contact_14_824
timestamp 1624857261
transform 1 0 119061 0 1 132000
box 0 0 1 1
use contact_14  contact_14_825
timestamp 1624857261
transform 1 0 118725 0 1 132000
box 0 0 1 1
use contact_14  contact_14_826
timestamp 1624857261
transform 1 0 118389 0 1 132000
box 0 0 1 1
use contact_13  contact_13_823
timestamp 1624857261
transform 1 0 119401 0 1 131992
box 0 0 1 1
use contact_13  contact_13_824
timestamp 1624857261
transform 1 0 119065 0 1 131992
box 0 0 1 1
use contact_13  contact_13_825
timestamp 1624857261
transform 1 0 118729 0 1 131992
box 0 0 1 1
use contact_13  contact_13_826
timestamp 1624857261
transform 1 0 118393 0 1 131992
box 0 0 1 1
use contact_33  contact_33_61
timestamp 1624857261
transform 1 0 119544 0 1 131245
box 0 0 1 1
use contact_33  contact_33_28
timestamp 1624857261
transform 1 0 120632 0 1 131381
box 0 0 1 1
use contact_33  contact_33_2512
timestamp 1624857261
transform 1 0 119680 0 1 131925
box 0 0 1 1
use contact_33  contact_33_2511
timestamp 1624857261
transform 1 0 119680 0 1 132061
box 0 0 1 1
use contact_13  contact_13_822
timestamp 1624857261
transform 1 0 119737 0 1 131992
box 0 0 1 1
use contact_19  contact_19_782
timestamp 1624857261
transform 1 0 119730 0 1 132001
box 0 0 1 1
use contact_14  contact_14_822
timestamp 1624857261
transform 1 0 119733 0 1 132000
box 0 0 1 1
use contact_7  contact_7_166
timestamp 1624857261
transform 1 0 119729 0 1 131996
box 0 0 1 1
use contact_13  contact_13_821
timestamp 1624857261
transform 1 0 120073 0 1 131992
box 0 0 1 1
use contact_14  contact_14_821
timestamp 1624857261
transform 1 0 120069 0 1 132000
box 0 0 1 1
use contact_13  contact_13_820
timestamp 1624857261
transform 1 0 120409 0 1 131992
box 0 0 1 1
use contact_14  contact_14_820
timestamp 1624857261
transform 1 0 120405 0 1 132000
box 0 0 1 1
use contact_13  contact_13_819
timestamp 1624857261
transform 1 0 120745 0 1 131992
box 0 0 1 1
use contact_14  contact_14_819
timestamp 1624857261
transform 1 0 120741 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2510
timestamp 1624857261
transform 1 0 119680 0 1 132469
box 0 0 1 1
use contact_13  contact_13_818
timestamp 1624857261
transform 1 0 121081 0 1 131992
box 0 0 1 1
use contact_14  contact_14_818
timestamp 1624857261
transform 1 0 121077 0 1 132000
box 0 0 1 1
use contact_13  contact_13_817
timestamp 1624857261
transform 1 0 121417 0 1 131992
box 0 0 1 1
use contact_13  contact_13_816
timestamp 1624857261
transform 1 0 121753 0 1 131992
box 0 0 1 1
use contact_19  contact_19_781
timestamp 1624857261
transform 1 0 121410 0 1 132001
box 0 0 1 1
use contact_14  contact_14_817
timestamp 1624857261
transform 1 0 121413 0 1 132000
box 0 0 1 1
use contact_14  contact_14_816
timestamp 1624857261
transform 1 0 121749 0 1 132000
box 0 0 1 1
use contact_7  contact_7_165
timestamp 1624857261
transform 1 0 121409 0 1 131996
box 0 0 1 1
use contact_13  contact_13_815
timestamp 1624857261
transform 1 0 122089 0 1 131992
box 0 0 1 1
use contact_14  contact_14_815
timestamp 1624857261
transform 1 0 122085 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2485
timestamp 1624857261
transform 1 0 121448 0 1 132061
box 0 0 1 1
use contact_33  contact_33_2484
timestamp 1624857261
transform 1 0 121448 0 1 132469
box 0 0 1 1
use contact_13  contact_13_814
timestamp 1624857261
transform 1 0 122425 0 1 131992
box 0 0 1 1
use contact_13  contact_13_813
timestamp 1624857261
transform 1 0 122761 0 1 131992
box 0 0 1 1
use contact_14  contact_14_814
timestamp 1624857261
transform 1 0 122421 0 1 132000
box 0 0 1 1
use contact_14  contact_14_813
timestamp 1624857261
transform 1 0 122757 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2483
timestamp 1624857261
transform 1 0 123080 0 1 132061
box 0 0 1 1
use contact_13  contact_13_812
timestamp 1624857261
transform 1 0 123097 0 1 131992
box 0 0 1 1
use contact_19  contact_19_780
timestamp 1624857261
transform 1 0 123090 0 1 132001
box 0 0 1 1
use contact_14  contact_14_812
timestamp 1624857261
transform 1 0 123093 0 1 132000
box 0 0 1 1
use contact_7  contact_7_164
timestamp 1624857261
transform 1 0 123089 0 1 131996
box 0 0 1 1
use contact_13  contact_13_811
timestamp 1624857261
transform 1 0 123433 0 1 131992
box 0 0 1 1
use contact_14  contact_14_811
timestamp 1624857261
transform 1 0 123429 0 1 132000
box 0 0 1 1
use contact_13  contact_13_810
timestamp 1624857261
transform 1 0 123769 0 1 131992
box 0 0 1 1
use contact_14  contact_14_810
timestamp 1624857261
transform 1 0 123765 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2482
timestamp 1624857261
transform 1 0 123080 0 1 132469
box 0 0 1 1
use contact_13  contact_13_809
timestamp 1624857261
transform 1 0 124105 0 1 131992
box 0 0 1 1
use contact_14  contact_14_809
timestamp 1624857261
transform 1 0 124101 0 1 132000
box 0 0 1 1
use contact_13  contact_13_808
timestamp 1624857261
transform 1 0 124441 0 1 131992
box 0 0 1 1
use contact_14  contact_14_808
timestamp 1624857261
transform 1 0 124437 0 1 132000
box 0 0 1 1
use contact_13  contact_13_807
timestamp 1624857261
transform 1 0 124777 0 1 131992
box 0 0 1 1
use contact_19  contact_19_779
timestamp 1624857261
transform 1 0 124770 0 1 132001
box 0 0 1 1
use contact_14  contact_14_807
timestamp 1624857261
transform 1 0 124773 0 1 132000
box 0 0 1 1
use contact_7  contact_7_163
timestamp 1624857261
transform 1 0 124769 0 1 131996
box 0 0 1 1
use contact_13  contact_13_806
timestamp 1624857261
transform 1 0 125113 0 1 131992
box 0 0 1 1
use contact_14  contact_14_806
timestamp 1624857261
transform 1 0 125109 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2467
timestamp 1624857261
transform 1 0 124712 0 1 132061
box 0 0 1 1
use contact_33  contact_33_2466
timestamp 1624857261
transform 1 0 124712 0 1 132469
box 0 0 1 1
use contact_33  contact_33_27
timestamp 1624857261
transform 1 0 120632 0 1 133149
box 0 0 1 1
use contact_33  contact_33_17
timestamp 1624857261
transform 1 0 123624 0 1 133149
box 0 0 1 1
use contact_7  contact_7_360
timestamp 1624857261
transform 1 0 132842 0 1 129658
box 0 0 1 1
use contact_33  contact_33_5450
timestamp 1624857261
transform 1 0 132736 0 1 129749
box 0 0 1 1
use contact_13  contact_13_805
timestamp 1624857261
transform 1 0 125449 0 1 131992
box 0 0 1 1
use contact_14  contact_14_805
timestamp 1624857261
transform 1 0 125445 0 1 132000
box 0 0 1 1
use contact_13  contact_13_804
timestamp 1624857261
transform 1 0 125785 0 1 131992
box 0 0 1 1
use contact_13  contact_13_803
timestamp 1624857261
transform 1 0 126121 0 1 131992
box 0 0 1 1
use contact_14  contact_14_804
timestamp 1624857261
transform 1 0 125781 0 1 132000
box 0 0 1 1
use contact_14  contact_14_803
timestamp 1624857261
transform 1 0 126117 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2465
timestamp 1624857261
transform 1 0 126344 0 1 132061
box 0 0 1 1
use contact_13  contact_13_802
timestamp 1624857261
transform 1 0 126457 0 1 131992
box 0 0 1 1
use contact_19  contact_19_778
timestamp 1624857261
transform 1 0 126450 0 1 132001
box 0 0 1 1
use contact_14  contact_14_802
timestamp 1624857261
transform 1 0 126453 0 1 132000
box 0 0 1 1
use contact_7  contact_7_162
timestamp 1624857261
transform 1 0 126449 0 1 131996
box 0 0 1 1
use contact_13  contact_13_801
timestamp 1624857261
transform 1 0 126793 0 1 131992
box 0 0 1 1
use contact_14  contact_14_801
timestamp 1624857261
transform 1 0 126789 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2464
timestamp 1624857261
transform 1 0 126344 0 1 132469
box 0 0 1 1
use contact_13  contact_13_800
timestamp 1624857261
transform 1 0 127129 0 1 131992
box 0 0 1 1
use contact_14  contact_14_800
timestamp 1624857261
transform 1 0 127125 0 1 132000
box 0 0 1 1
use contact_13  contact_13_799
timestamp 1624857261
transform 1 0 127465 0 1 131992
box 0 0 1 1
use contact_14  contact_14_799
timestamp 1624857261
transform 1 0 127461 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2461
timestamp 1624857261
transform 1 0 128112 0 1 132061
box 0 0 1 1
use contact_13  contact_13_798
timestamp 1624857261
transform 1 0 127801 0 1 131992
box 0 0 1 1
use contact_13  contact_13_797
timestamp 1624857261
transform 1 0 128137 0 1 131992
box 0 0 1 1
use contact_19  contact_19_777
timestamp 1624857261
transform 1 0 128130 0 1 132001
box 0 0 1 1
use contact_14  contact_14_798
timestamp 1624857261
transform 1 0 127797 0 1 132000
box 0 0 1 1
use contact_14  contact_14_797
timestamp 1624857261
transform 1 0 128133 0 1 132000
box 0 0 1 1
use contact_7  contact_7_161
timestamp 1624857261
transform 1 0 128129 0 1 131996
box 0 0 1 1
use contact_33  contact_33_2460
timestamp 1624857261
transform 1 0 128112 0 1 132469
box 0 0 1 1
use contact_13  contact_13_796
timestamp 1624857261
transform 1 0 128473 0 1 131992
box 0 0 1 1
use contact_13  contact_13_795
timestamp 1624857261
transform 1 0 128809 0 1 131992
box 0 0 1 1
use contact_14  contact_14_796
timestamp 1624857261
transform 1 0 128469 0 1 132000
box 0 0 1 1
use contact_14  contact_14_795
timestamp 1624857261
transform 1 0 128805 0 1 132000
box 0 0 1 1
use contact_13  contact_13_794
timestamp 1624857261
transform 1 0 129145 0 1 131992
box 0 0 1 1
use contact_14  contact_14_794
timestamp 1624857261
transform 1 0 129141 0 1 132000
box 0 0 1 1
use contact_13  contact_13_793
timestamp 1624857261
transform 1 0 129481 0 1 131992
box 0 0 1 1
use contact_14  contact_14_793
timestamp 1624857261
transform 1 0 129477 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2457
timestamp 1624857261
transform 1 0 129880 0 1 132061
box 0 0 1 1
use contact_13  contact_13_792
timestamp 1624857261
transform 1 0 129817 0 1 131992
box 0 0 1 1
use contact_19  contact_19_776
timestamp 1624857261
transform 1 0 129810 0 1 132001
box 0 0 1 1
use contact_14  contact_14_792
timestamp 1624857261
transform 1 0 129813 0 1 132000
box 0 0 1 1
use contact_7  contact_7_160
timestamp 1624857261
transform 1 0 129809 0 1 131996
box 0 0 1 1
use contact_33  contact_33_2456
timestamp 1624857261
transform 1 0 129880 0 1 132469
box 0 0 1 1
use contact_13  contact_13_791
timestamp 1624857261
transform 1 0 130153 0 1 131992
box 0 0 1 1
use contact_14  contact_14_791
timestamp 1624857261
transform 1 0 130149 0 1 132000
box 0 0 1 1
use contact_13  contact_13_790
timestamp 1624857261
transform 1 0 130489 0 1 131992
box 0 0 1 1
use contact_13  contact_13_789
timestamp 1624857261
transform 1 0 130825 0 1 131992
box 0 0 1 1
use contact_14  contact_14_790
timestamp 1624857261
transform 1 0 130485 0 1 132000
box 0 0 1 1
use contact_14  contact_14_789
timestamp 1624857261
transform 1 0 130821 0 1 132000
box 0 0 1 1
use contact_13  contact_13_788
timestamp 1624857261
transform 1 0 131161 0 1 131992
box 0 0 1 1
use contact_14  contact_14_788
timestamp 1624857261
transform 1 0 131157 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2451
timestamp 1624857261
transform 1 0 131376 0 1 132061
box 0 0 1 1
use contact_13  contact_13_787
timestamp 1624857261
transform 1 0 131497 0 1 131992
box 0 0 1 1
use contact_19  contact_19_775
timestamp 1624857261
transform 1 0 131490 0 1 132001
box 0 0 1 1
use contact_14  contact_14_787
timestamp 1624857261
transform 1 0 131493 0 1 132000
box 0 0 1 1
use contact_7  contact_7_159
timestamp 1624857261
transform 1 0 131489 0 1 131996
box 0 0 1 1
use contact_33  contact_33_2450
timestamp 1624857261
transform 1 0 131376 0 1 132469
box 0 0 1 1
use contact_13  contact_13_786
timestamp 1624857261
transform 1 0 131833 0 1 131992
box 0 0 1 1
use contact_14  contact_14_786
timestamp 1624857261
transform 1 0 131829 0 1 132000
box 0 0 1 1
use contact_13  contact_13_785
timestamp 1624857261
transform 1 0 132169 0 1 131992
box 0 0 1 1
use contact_14  contact_14_785
timestamp 1624857261
transform 1 0 132165 0 1 132000
box 0 0 1 1
use contact_13  contact_13_784
timestamp 1624857261
transform 1 0 132505 0 1 131992
box 0 0 1 1
use contact_13  contact_13_783
timestamp 1624857261
transform 1 0 132841 0 1 131992
box 0 0 1 1
use contact_14  contact_14_784
timestamp 1624857261
transform 1 0 132501 0 1 132000
box 0 0 1 1
use contact_14  contact_14_783
timestamp 1624857261
transform 1 0 132837 0 1 132000
box 0 0 1 1
use contact_33  contact_33_2449
timestamp 1624857261
transform 1 0 133144 0 1 132061
box 0 0 1 1
use contact_13  contact_13_782
timestamp 1624857261
transform 1 0 133177 0 1 131992
box 0 0 1 1
use contact_19  contact_19_774
timestamp 1624857261
transform 1 0 133170 0 1 132001
box 0 0 1 1
use contact_14  contact_14_782
timestamp 1624857261
transform 1 0 133173 0 1 132000
box 0 0 1 1
use contact_7  contact_7_158
timestamp 1624857261
transform 1 0 133169 0 1 131996
box 0 0 1 1
use contact_33  contact_33_2448
timestamp 1624857261
transform 1 0 133144 0 1 132469
box 0 0 1 1
use contact_14  contact_14_778
timestamp 1624857261
transform 1 0 134517 0 1 132000
box 0 0 1 1
use contact_14  contact_14_779
timestamp 1624857261
transform 1 0 134181 0 1 132000
box 0 0 1 1
use contact_14  contact_14_780
timestamp 1624857261
transform 1 0 133845 0 1 132000
box 0 0 1 1
use contact_14  contact_14_781
timestamp 1624857261
transform 1 0 133509 0 1 132000
box 0 0 1 1
use contact_13  contact_13_778
timestamp 1624857261
transform 1 0 134521 0 1 131992
box 0 0 1 1
use contact_13  contact_13_779
timestamp 1624857261
transform 1 0 134185 0 1 131992
box 0 0 1 1
use contact_13  contact_13_780
timestamp 1624857261
transform 1 0 133849 0 1 131992
box 0 0 1 1
use contact_13  contact_13_781
timestamp 1624857261
transform 1 0 133513 0 1 131992
box 0 0 1 1
use contact_7  contact_7_157
timestamp 1624857261
transform 1 0 134849 0 1 131996
box 0 0 1 1
use contact_14  contact_14_777
timestamp 1624857261
transform 1 0 134853 0 1 132000
box 0 0 1 1
use contact_19  contact_19_773
timestamp 1624857261
transform 1 0 134850 0 1 132001
box 0 0 1 1
use contact_13  contact_13_777
timestamp 1624857261
transform 1 0 134857 0 1 131992
box 0 0 1 1
use contact_33  contact_33_2444
timestamp 1624857261
transform 1 0 134912 0 1 132469
box 0 0 1 1
use contact_33  contact_33_2445
timestamp 1624857261
transform 1 0 134912 0 1 132061
box 0 0 1 1
use contact_33  contact_33_2432
timestamp 1624857261
transform 1 0 136544 0 1 1229
box 0 0 1 1
use contact_14  contact_14_1177
timestamp 1624857261
transform 1 0 135189 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1177
timestamp 1624857261
transform 1 0 135193 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1175
timestamp 1624857261
transform 1 0 135861 0 1 1691
box 0 0 1 1
use contact_14  contact_14_1176
timestamp 1624857261
transform 1 0 135525 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1175
timestamp 1624857261
transform 1 0 135865 0 1 1683
box 0 0 1 1
use contact_13  contact_13_1176
timestamp 1624857261
transform 1 0 135529 0 1 1683
box 0 0 1 1
use contact_14  contact_14_1174
timestamp 1624857261
transform 1 0 136197 0 1 1691
box 0 0 1 1
use contact_13  contact_13_1174
timestamp 1624857261
transform 1 0 136201 0 1 1683
box 0 0 1 1
use contact_38  contact_38_2
timestamp 1624857261
transform 1 0 136876 0 1 1628
box 0 0 192 192
use contact_7  contact_7_237
timestamp 1624857261
transform 1 0 136529 0 1 1687
box 0 0 1 1
use contact_14  contact_14_1173
timestamp 1624857261
transform 1 0 136533 0 1 1691
box 0 0 1 1
use contact_19  contact_19_853
timestamp 1624857261
transform 1 0 136530 0 1 1692
box 0 0 1 1
use contact_13  contact_13_1173
timestamp 1624857261
transform 1 0 136537 0 1 1683
box 0 0 1 1
use contact_33  contact_33_2433
timestamp 1624857261
transform 1 0 136544 0 1 1637
box 0 0 1 1
use contact_7  contact_7_77
timestamp 1624857261
transform 1 0 136939 0 1 2023
box 0 0 1 1
use contact_14  contact_14_385
timestamp 1624857261
transform 1 0 136943 0 1 2027
box 0 0 1 1
use contact_19  contact_19_385
timestamp 1624857261
transform 1 0 136940 0 1 2028
box 0 0 1 1
use contact_13  contact_13_385
timestamp 1624857261
transform 1 0 136947 0 1 2019
box 0 0 1 1
use contact_14  contact_14_383
timestamp 1624857261
transform 1 0 136943 0 1 2699
box 0 0 1 1
use contact_14  contact_14_384
timestamp 1624857261
transform 1 0 136943 0 1 2363
box 0 0 1 1
use contact_19  contact_19_383
timestamp 1624857261
transform 1 0 136940 0 1 2700
box 0 0 1 1
use contact_19  contact_19_384
timestamp 1624857261
transform 1 0 136940 0 1 2364
box 0 0 1 1
use contact_13  contact_13_383
timestamp 1624857261
transform 1 0 136947 0 1 2691
box 0 0 1 1
use contact_13  contact_13_384
timestamp 1624857261
transform 1 0 136947 0 1 2355
box 0 0 1 1
use contact_39  contact_39_2
timestamp 1624857261
transform 1 0 138448 0 1 277
box 0 0 192 192
use contact_39  contact_39_3
timestamp 1624857261
transform 1 0 138176 0 1 413
box 0 0 192 192
use contact_39  contact_39_6
timestamp 1624857261
transform 1 0 138176 0 1 277
box 0 0 192 192
use contact_39  contact_39_8
timestamp 1624857261
transform 1 0 138312 0 1 549
box 0 0 192 192
use contact_39  contact_39_10
timestamp 1624857261
transform 1 0 138448 0 1 413
box 0 0 192 192
use contact_39  contact_39_19
timestamp 1624857261
transform 1 0 138176 0 1 549
box 0 0 192 192
use contact_39  contact_39_21
timestamp 1624857261
transform 1 0 138312 0 1 413
box 0 0 192 192
use contact_39  contact_39_24
timestamp 1624857261
transform 1 0 138448 0 1 549
box 0 0 192 192
use contact_39  contact_39_27
timestamp 1624857261
transform 1 0 138312 0 1 277
box 0 0 192 192
use contact_39  contact_39_40
timestamp 1624857261
transform 1 0 137768 0 1 1093
box 0 0 192 192
use contact_39  contact_39_44
timestamp 1624857261
transform 1 0 137496 0 1 1093
box 0 0 192 192
use contact_39  contact_39_47
timestamp 1624857261
transform 1 0 137496 0 1 1229
box 0 0 192 192
use contact_39  contact_39_49
timestamp 1624857261
transform 1 0 137632 0 1 1229
box 0 0 192 192
use contact_39  contact_39_50
timestamp 1624857261
transform 1 0 137632 0 1 1093
box 0 0 192 192
use contact_39  contact_39_52
timestamp 1624857261
transform 1 0 137768 0 1 1229
box 0 0 192 192
use contact_39  contact_39_59
timestamp 1624857261
transform 1 0 137768 0 1 957
box 0 0 192 192
use contact_39  contact_39_61
timestamp 1624857261
transform 1 0 137496 0 1 957
box 0 0 192 192
use contact_39  contact_39_71
timestamp 1624857261
transform 1 0 137632 0 1 957
box 0 0 192 192
use contact_14  contact_14_382
timestamp 1624857261
transform 1 0 136943 0 1 3035
box 0 0 1 1
use contact_19  contact_19_382
timestamp 1624857261
transform 1 0 136940 0 1 3036
box 0 0 1 1
use contact_13  contact_13_382
timestamp 1624857261
transform 1 0 136947 0 1 3027
box 0 0 1 1
use contact_7  contact_7_76
timestamp 1624857261
transform 1 0 136939 0 1 3703
box 0 0 1 1
use contact_14  contact_14_380
timestamp 1624857261
transform 1 0 136943 0 1 3707
box 0 0 1 1
use contact_14  contact_14_381
timestamp 1624857261
transform 1 0 136943 0 1 3371
box 0 0 1 1
use contact_19  contact_19_380
timestamp 1624857261
transform 1 0 136940 0 1 3708
box 0 0 1 1
use contact_19  contact_19_381
timestamp 1624857261
transform 1 0 136940 0 1 3372
box 0 0 1 1
use contact_13  contact_13_380
timestamp 1624857261
transform 1 0 136947 0 1 3699
box 0 0 1 1
use contact_13  contact_13_381
timestamp 1624857261
transform 1 0 136947 0 1 3363
box 0 0 1 1
use contact_14  contact_14_378
timestamp 1624857261
transform 1 0 136943 0 1 4379
box 0 0 1 1
use contact_14  contact_14_379
timestamp 1624857261
transform 1 0 136943 0 1 4043
box 0 0 1 1
use contact_19  contact_19_378
timestamp 1624857261
transform 1 0 136940 0 1 4380
box 0 0 1 1
use contact_19  contact_19_379
timestamp 1624857261
transform 1 0 136940 0 1 4044
box 0 0 1 1
use contact_13  contact_13_378
timestamp 1624857261
transform 1 0 136947 0 1 4371
box 0 0 1 1
use contact_13  contact_13_379
timestamp 1624857261
transform 1 0 136947 0 1 4035
box 0 0 1 1
use contact_14  contact_14_377
timestamp 1624857261
transform 1 0 136943 0 1 4715
box 0 0 1 1
use contact_19  contact_19_377
timestamp 1624857261
transform 1 0 136940 0 1 4716
box 0 0 1 1
use contact_13  contact_13_377
timestamp 1624857261
transform 1 0 136947 0 1 4707
box 0 0 1 1
use contact_14  contact_14_376
timestamp 1624857261
transform 1 0 136943 0 1 5051
box 0 0 1 1
use contact_19  contact_19_376
timestamp 1624857261
transform 1 0 136940 0 1 5052
box 0 0 1 1
use contact_13  contact_13_376
timestamp 1624857261
transform 1 0 136947 0 1 5043
box 0 0 1 1
use contact_33  contact_33_2377
timestamp 1624857261
transform 1 0 137496 0 1 3813
box 0 0 1 1
use contact_7  contact_7_75
timestamp 1624857261
transform 1 0 136939 0 1 5383
box 0 0 1 1
use contact_14  contact_14_374
timestamp 1624857261
transform 1 0 136943 0 1 5723
box 0 0 1 1
use contact_14  contact_14_375
timestamp 1624857261
transform 1 0 136943 0 1 5387
box 0 0 1 1
use contact_19  contact_19_374
timestamp 1624857261
transform 1 0 136940 0 1 5724
box 0 0 1 1
use contact_19  contact_19_375
timestamp 1624857261
transform 1 0 136940 0 1 5388
box 0 0 1 1
use contact_13  contact_13_374
timestamp 1624857261
transform 1 0 136947 0 1 5715
box 0 0 1 1
use contact_13  contact_13_375
timestamp 1624857261
transform 1 0 136947 0 1 5379
box 0 0 1 1
use contact_14  contact_14_373
timestamp 1624857261
transform 1 0 136943 0 1 6059
box 0 0 1 1
use contact_19  contact_19_373
timestamp 1624857261
transform 1 0 136940 0 1 6060
box 0 0 1 1
use contact_13  contact_13_373
timestamp 1624857261
transform 1 0 136947 0 1 6051
box 0 0 1 1
use contact_14  contact_14_371
timestamp 1624857261
transform 1 0 136943 0 1 6731
box 0 0 1 1
use contact_14  contact_14_372
timestamp 1624857261
transform 1 0 136943 0 1 6395
box 0 0 1 1
use contact_19  contact_19_371
timestamp 1624857261
transform 1 0 136940 0 1 6732
box 0 0 1 1
use contact_19  contact_19_372
timestamp 1624857261
transform 1 0 136940 0 1 6396
box 0 0 1 1
use contact_13  contact_13_371
timestamp 1624857261
transform 1 0 136947 0 1 6723
box 0 0 1 1
use contact_13  contact_13_372
timestamp 1624857261
transform 1 0 136947 0 1 6387
box 0 0 1 1
use contact_7  contact_7_74
timestamp 1624857261
transform 1 0 136939 0 1 7063
box 0 0 1 1
use contact_14  contact_14_370
timestamp 1624857261
transform 1 0 136943 0 1 7067
box 0 0 1 1
use contact_19  contact_19_370
timestamp 1624857261
transform 1 0 136940 0 1 7068
box 0 0 1 1
use contact_13  contact_13_370
timestamp 1624857261
transform 1 0 136947 0 1 7059
box 0 0 1 1
use contact_14  contact_14_368
timestamp 1624857261
transform 1 0 136943 0 1 7739
box 0 0 1 1
use contact_14  contact_14_369
timestamp 1624857261
transform 1 0 136943 0 1 7403
box 0 0 1 1
use contact_19  contact_19_368
timestamp 1624857261
transform 1 0 136940 0 1 7740
box 0 0 1 1
use contact_19  contact_19_369
timestamp 1624857261
transform 1 0 136940 0 1 7404
box 0 0 1 1
use contact_13  contact_13_368
timestamp 1624857261
transform 1 0 136947 0 1 7731
box 0 0 1 1
use contact_13  contact_13_369
timestamp 1624857261
transform 1 0 136947 0 1 7395
box 0 0 1 1
use contact_33  contact_33_2427
timestamp 1624857261
transform 1 0 137496 0 1 5445
box 0 0 1 1
use contact_33  contact_33_2383
timestamp 1624857261
transform 1 0 137496 0 1 7077
box 0 0 1 1
use contact_14  contact_14_366
timestamp 1624857261
transform 1 0 136943 0 1 8411
box 0 0 1 1
use contact_14  contact_14_367
timestamp 1624857261
transform 1 0 136943 0 1 8075
box 0 0 1 1
use contact_19  contact_19_366
timestamp 1624857261
transform 1 0 136940 0 1 8412
box 0 0 1 1
use contact_19  contact_19_367
timestamp 1624857261
transform 1 0 136940 0 1 8076
box 0 0 1 1
use contact_13  contact_13_366
timestamp 1624857261
transform 1 0 136947 0 1 8403
box 0 0 1 1
use contact_13  contact_13_367
timestamp 1624857261
transform 1 0 136947 0 1 8067
box 0 0 1 1
use contact_7  contact_7_73
timestamp 1624857261
transform 1 0 136939 0 1 8743
box 0 0 1 1
use contact_14  contact_14_365
timestamp 1624857261
transform 1 0 136943 0 1 8747
box 0 0 1 1
use contact_19  contact_19_365
timestamp 1624857261
transform 1 0 136940 0 1 8748
box 0 0 1 1
use contact_13  contact_13_365
timestamp 1624857261
transform 1 0 136947 0 1 8739
box 0 0 1 1
use contact_14  contact_14_363
timestamp 1624857261
transform 1 0 136943 0 1 9419
box 0 0 1 1
use contact_14  contact_14_364
timestamp 1624857261
transform 1 0 136943 0 1 9083
box 0 0 1 1
use contact_19  contact_19_363
timestamp 1624857261
transform 1 0 136940 0 1 9420
box 0 0 1 1
use contact_19  contact_19_364
timestamp 1624857261
transform 1 0 136940 0 1 9084
box 0 0 1 1
use contact_13  contact_13_363
timestamp 1624857261
transform 1 0 136947 0 1 9411
box 0 0 1 1
use contact_13  contact_13_364
timestamp 1624857261
transform 1 0 136947 0 1 9075
box 0 0 1 1
use contact_14  contact_14_362
timestamp 1624857261
transform 1 0 136943 0 1 9755
box 0 0 1 1
use contact_19  contact_19_362
timestamp 1624857261
transform 1 0 136940 0 1 9756
box 0 0 1 1
use contact_13  contact_13_362
timestamp 1624857261
transform 1 0 136947 0 1 9747
box 0 0 1 1
use contact_14  contact_14_361
timestamp 1624857261
transform 1 0 136943 0 1 10091
box 0 0 1 1
use contact_19  contact_19_361
timestamp 1624857261
transform 1 0 136940 0 1 10092
box 0 0 1 1
use contact_13  contact_13_361
timestamp 1624857261
transform 1 0 136947 0 1 10083
box 0 0 1 1
use contact_33  contact_33_2367
timestamp 1624857261
transform 1 0 137496 0 1 8709
box 0 0 1 1
use contact_7  contact_7_72
timestamp 1624857261
transform 1 0 136939 0 1 10423
box 0 0 1 1
use contact_14  contact_14_359
timestamp 1624857261
transform 1 0 136943 0 1 10763
box 0 0 1 1
use contact_14  contact_14_360
timestamp 1624857261
transform 1 0 136943 0 1 10427
box 0 0 1 1
use contact_19  contact_19_359
timestamp 1624857261
transform 1 0 136940 0 1 10764
box 0 0 1 1
use contact_19  contact_19_360
timestamp 1624857261
transform 1 0 136940 0 1 10428
box 0 0 1 1
use contact_13  contact_13_359
timestamp 1624857261
transform 1 0 136947 0 1 10755
box 0 0 1 1
use contact_13  contact_13_360
timestamp 1624857261
transform 1 0 136947 0 1 10419
box 0 0 1 1
use contact_14  contact_14_358
timestamp 1624857261
transform 1 0 136943 0 1 11099
box 0 0 1 1
use contact_19  contact_19_358
timestamp 1624857261
transform 1 0 136940 0 1 11100
box 0 0 1 1
use contact_13  contact_13_358
timestamp 1624857261
transform 1 0 136947 0 1 11091
box 0 0 1 1
use contact_14  contact_14_356
timestamp 1624857261
transform 1 0 136943 0 1 11771
box 0 0 1 1
use contact_14  contact_14_357
timestamp 1624857261
transform 1 0 136943 0 1 11435
box 0 0 1 1
use contact_19  contact_19_356
timestamp 1624857261
transform 1 0 136940 0 1 11772
box 0 0 1 1
use contact_19  contact_19_357
timestamp 1624857261
transform 1 0 136940 0 1 11436
box 0 0 1 1
use contact_13  contact_13_356
timestamp 1624857261
transform 1 0 136947 0 1 11763
box 0 0 1 1
use contact_13  contact_13_357
timestamp 1624857261
transform 1 0 136947 0 1 11427
box 0 0 1 1
use contact_7  contact_7_71
timestamp 1624857261
transform 1 0 136939 0 1 12103
box 0 0 1 1
use contact_14  contact_14_355
timestamp 1624857261
transform 1 0 136943 0 1 12107
box 0 0 1 1
use contact_19  contact_19_355
timestamp 1624857261
transform 1 0 136940 0 1 12108
box 0 0 1 1
use contact_13  contact_13_355
timestamp 1624857261
transform 1 0 136947 0 1 12099
box 0 0 1 1
use contact_14  contact_14_353
timestamp 1624857261
transform 1 0 136943 0 1 12779
box 0 0 1 1
use contact_14  contact_14_354
timestamp 1624857261
transform 1 0 136943 0 1 12443
box 0 0 1 1
use contact_19  contact_19_353
timestamp 1624857261
transform 1 0 136940 0 1 12780
box 0 0 1 1
use contact_19  contact_19_354
timestamp 1624857261
transform 1 0 136940 0 1 12444
box 0 0 1 1
use contact_13  contact_13_353
timestamp 1624857261
transform 1 0 136947 0 1 12771
box 0 0 1 1
use contact_13  contact_13_354
timestamp 1624857261
transform 1 0 136947 0 1 12435
box 0 0 1 1
use contact_33  contact_33_2411
timestamp 1624857261
transform 1 0 137496 0 1 11973
box 0 0 1 1
use contact_33  contact_33_2389
timestamp 1624857261
transform 1 0 137496 0 1 10477
box 0 0 1 1
use contact_14  contact_14_352
timestamp 1624857261
transform 1 0 136943 0 1 13115
box 0 0 1 1
use contact_19  contact_19_352
timestamp 1624857261
transform 1 0 136940 0 1 13116
box 0 0 1 1
use contact_13  contact_13_351
timestamp 1624857261
transform 1 0 136947 0 1 13443
box 0 0 1 1
use contact_13  contact_13_352
timestamp 1624857261
transform 1 0 136947 0 1 13107
box 0 0 1 1
use contact_7  contact_7_70
timestamp 1624857261
transform 1 0 136939 0 1 13783
box 0 0 1 1
use contact_14  contact_14_350
timestamp 1624857261
transform 1 0 136943 0 1 13787
box 0 0 1 1
use contact_14  contact_14_351
timestamp 1624857261
transform 1 0 136943 0 1 13451
box 0 0 1 1
use contact_19  contact_19_350
timestamp 1624857261
transform 1 0 136940 0 1 13788
box 0 0 1 1
use contact_19  contact_19_351
timestamp 1624857261
transform 1 0 136940 0 1 13452
box 0 0 1 1
use contact_13  contact_13_350
timestamp 1624857261
transform 1 0 136947 0 1 13779
box 0 0 1 1
use contact_14  contact_14_349
timestamp 1624857261
transform 1 0 136943 0 1 14123
box 0 0 1 1
use contact_19  contact_19_349
timestamp 1624857261
transform 1 0 136940 0 1 14124
box 0 0 1 1
use contact_13  contact_13_349
timestamp 1624857261
transform 1 0 136947 0 1 14115
box 0 0 1 1
use contact_14  contact_14_347
timestamp 1624857261
transform 1 0 136943 0 1 14795
box 0 0 1 1
use contact_14  contact_14_348
timestamp 1624857261
transform 1 0 136943 0 1 14459
box 0 0 1 1
use contact_19  contact_19_347
timestamp 1624857261
transform 1 0 136940 0 1 14796
box 0 0 1 1
use contact_19  contact_19_348
timestamp 1624857261
transform 1 0 136940 0 1 14460
box 0 0 1 1
use contact_13  contact_13_347
timestamp 1624857261
transform 1 0 136947 0 1 14787
box 0 0 1 1
use contact_13  contact_13_348
timestamp 1624857261
transform 1 0 136947 0 1 14451
box 0 0 1 1
use contact_14  contact_14_346
timestamp 1624857261
transform 1 0 136943 0 1 15131
box 0 0 1 1
use contact_19  contact_19_346
timestamp 1624857261
transform 1 0 136940 0 1 15132
box 0 0 1 1
use contact_13  contact_13_346
timestamp 1624857261
transform 1 0 136947 0 1 15123
box 0 0 1 1
use contact_7  contact_7_69
timestamp 1624857261
transform 1 0 136939 0 1 15463
box 0 0 1 1
use contact_14  contact_14_345
timestamp 1624857261
transform 1 0 136943 0 1 15467
box 0 0 1 1
use contact_19  contact_19_345
timestamp 1624857261
transform 1 0 136940 0 1 15468
box 0 0 1 1
use contact_13  contact_13_345
timestamp 1624857261
transform 1 0 136947 0 1 15459
box 0 0 1 1
use contact_33  contact_33_2392
timestamp 1624857261
transform 1 0 137496 0 1 13877
box 0 0 1 1
use contact_14  contact_14_344
timestamp 1624857261
transform 1 0 136943 0 1 15803
box 0 0 1 1
use contact_19  contact_19_344
timestamp 1624857261
transform 1 0 136940 0 1 15804
box 0 0 1 1
use contact_13  contact_13_344
timestamp 1624857261
transform 1 0 136947 0 1 15795
box 0 0 1 1
use contact_14  contact_14_342
timestamp 1624857261
transform 1 0 136943 0 1 16475
box 0 0 1 1
use contact_14  contact_14_343
timestamp 1624857261
transform 1 0 136943 0 1 16139
box 0 0 1 1
use contact_19  contact_19_342
timestamp 1624857261
transform 1 0 136940 0 1 16476
box 0 0 1 1
use contact_19  contact_19_343
timestamp 1624857261
transform 1 0 136940 0 1 16140
box 0 0 1 1
use contact_13  contact_13_342
timestamp 1624857261
transform 1 0 136947 0 1 16467
box 0 0 1 1
use contact_13  contact_13_343
timestamp 1624857261
transform 1 0 136947 0 1 16131
box 0 0 1 1
use contact_14  contact_14_341
timestamp 1624857261
transform 1 0 136943 0 1 16811
box 0 0 1 1
use contact_19  contact_19_341
timestamp 1624857261
transform 1 0 136940 0 1 16812
box 0 0 1 1
use contact_13  contact_13_341
timestamp 1624857261
transform 1 0 136947 0 1 16803
box 0 0 1 1
use contact_7  contact_7_68
timestamp 1624857261
transform 1 0 136939 0 1 17143
box 0 0 1 1
use contact_14  contact_14_339
timestamp 1624857261
transform 1 0 136943 0 1 17483
box 0 0 1 1
use contact_14  contact_14_340
timestamp 1624857261
transform 1 0 136943 0 1 17147
box 0 0 1 1
use contact_19  contact_19_339
timestamp 1624857261
transform 1 0 136940 0 1 17484
box 0 0 1 1
use contact_19  contact_19_340
timestamp 1624857261
transform 1 0 136940 0 1 17148
box 0 0 1 1
use contact_13  contact_13_339
timestamp 1624857261
transform 1 0 136947 0 1 17475
box 0 0 1 1
use contact_13  contact_13_340
timestamp 1624857261
transform 1 0 136947 0 1 17139
box 0 0 1 1
use contact_14  contact_14_338
timestamp 1624857261
transform 1 0 136943 0 1 17819
box 0 0 1 1
use contact_19  contact_19_338
timestamp 1624857261
transform 1 0 136940 0 1 17820
box 0 0 1 1
use contact_13  contact_13_338
timestamp 1624857261
transform 1 0 136947 0 1 17811
box 0 0 1 1
use contact_33  contact_33_2413
timestamp 1624857261
transform 1 0 137496 0 1 17005
box 0 0 1 1
use contact_33  contact_33_2398
timestamp 1624857261
transform 1 0 137496 0 1 15509
box 0 0 1 1
use contact_14  contact_14_336
timestamp 1624857261
transform 1 0 136943 0 1 18491
box 0 0 1 1
use contact_14  contact_14_337
timestamp 1624857261
transform 1 0 136943 0 1 18155
box 0 0 1 1
use contact_19  contact_19_336
timestamp 1624857261
transform 1 0 136940 0 1 18492
box 0 0 1 1
use contact_19  contact_19_337
timestamp 1624857261
transform 1 0 136940 0 1 18156
box 0 0 1 1
use contact_13  contact_13_336
timestamp 1624857261
transform 1 0 136947 0 1 18483
box 0 0 1 1
use contact_13  contact_13_337
timestamp 1624857261
transform 1 0 136947 0 1 18147
box 0 0 1 1
use contact_7  contact_7_67
timestamp 1624857261
transform 1 0 136939 0 1 18823
box 0 0 1 1
use contact_14  contact_14_335
timestamp 1624857261
transform 1 0 136943 0 1 18827
box 0 0 1 1
use contact_19  contact_19_335
timestamp 1624857261
transform 1 0 136940 0 1 18828
box 0 0 1 1
use contact_13  contact_13_335
timestamp 1624857261
transform 1 0 136947 0 1 18819
box 0 0 1 1
use contact_14  contact_14_333
timestamp 1624857261
transform 1 0 136943 0 1 19499
box 0 0 1 1
use contact_14  contact_14_334
timestamp 1624857261
transform 1 0 136943 0 1 19163
box 0 0 1 1
use contact_19  contact_19_333
timestamp 1624857261
transform 1 0 136940 0 1 19500
box 0 0 1 1
use contact_19  contact_19_334
timestamp 1624857261
transform 1 0 136940 0 1 19164
box 0 0 1 1
use contact_13  contact_13_333
timestamp 1624857261
transform 1 0 136947 0 1 19491
box 0 0 1 1
use contact_13  contact_13_334
timestamp 1624857261
transform 1 0 136947 0 1 19155
box 0 0 1 1
use contact_14  contact_14_332
timestamp 1624857261
transform 1 0 136943 0 1 19835
box 0 0 1 1
use contact_19  contact_19_332
timestamp 1624857261
transform 1 0 136940 0 1 19836
box 0 0 1 1
use contact_13  contact_13_332
timestamp 1624857261
transform 1 0 136947 0 1 19827
box 0 0 1 1
use contact_7  contact_7_66
timestamp 1624857261
transform 1 0 136939 0 1 20503
box 0 0 1 1
use contact_14  contact_14_331
timestamp 1624857261
transform 1 0 136943 0 1 20171
box 0 0 1 1
use contact_19  contact_19_331
timestamp 1624857261
transform 1 0 136940 0 1 20172
box 0 0 1 1
use contact_13  contact_13_330
timestamp 1624857261
transform 1 0 136947 0 1 20499
box 0 0 1 1
use contact_13  contact_13_331
timestamp 1624857261
transform 1 0 136947 0 1 20163
box 0 0 1 1
use contact_14  contact_14_330
timestamp 1624857261
transform 1 0 136943 0 1 20507
box 0 0 1 1
use contact_19  contact_19_330
timestamp 1624857261
transform 1 0 136940 0 1 20508
box 0 0 1 1
use contact_33  contact_33_2420
timestamp 1624857261
transform 1 0 137496 0 1 18773
box 0 0 1 1
use contact_33  contact_33_2356
timestamp 1624857261
transform 1 0 137496 0 1 20405
box 0 0 1 1
use contact_14  contact_14_329
timestamp 1624857261
transform 1 0 136943 0 1 20843
box 0 0 1 1
use contact_19  contact_19_329
timestamp 1624857261
transform 1 0 136940 0 1 20844
box 0 0 1 1
use contact_13  contact_13_329
timestamp 1624857261
transform 1 0 136947 0 1 20835
box 0 0 1 1
use contact_14  contact_14_327
timestamp 1624857261
transform 1 0 136943 0 1 21515
box 0 0 1 1
use contact_14  contact_14_328
timestamp 1624857261
transform 1 0 136943 0 1 21179
box 0 0 1 1
use contact_19  contact_19_327
timestamp 1624857261
transform 1 0 136940 0 1 21516
box 0 0 1 1
use contact_19  contact_19_328
timestamp 1624857261
transform 1 0 136940 0 1 21180
box 0 0 1 1
use contact_13  contact_13_327
timestamp 1624857261
transform 1 0 136947 0 1 21507
box 0 0 1 1
use contact_13  contact_13_328
timestamp 1624857261
transform 1 0 136947 0 1 21171
box 0 0 1 1
use contact_14  contact_14_326
timestamp 1624857261
transform 1 0 136943 0 1 21851
box 0 0 1 1
use contact_19  contact_19_326
timestamp 1624857261
transform 1 0 136940 0 1 21852
box 0 0 1 1
use contact_13  contact_13_326
timestamp 1624857261
transform 1 0 136947 0 1 21843
box 0 0 1 1
use contact_7  contact_7_65
timestamp 1624857261
transform 1 0 136939 0 1 22183
box 0 0 1 1
use contact_14  contact_14_324
timestamp 1624857261
transform 1 0 136943 0 1 22523
box 0 0 1 1
use contact_14  contact_14_325
timestamp 1624857261
transform 1 0 136943 0 1 22187
box 0 0 1 1
use contact_19  contact_19_324
timestamp 1624857261
transform 1 0 136940 0 1 22524
box 0 0 1 1
use contact_19  contact_19_325
timestamp 1624857261
transform 1 0 136940 0 1 22188
box 0 0 1 1
use contact_13  contact_13_324
timestamp 1624857261
transform 1 0 136947 0 1 22515
box 0 0 1 1
use contact_13  contact_13_325
timestamp 1624857261
transform 1 0 136947 0 1 22179
box 0 0 1 1
use contact_14  contact_14_323
timestamp 1624857261
transform 1 0 136943 0 1 22859
box 0 0 1 1
use contact_19  contact_19_323
timestamp 1624857261
transform 1 0 136940 0 1 22860
box 0 0 1 1
use contact_13  contact_13_323
timestamp 1624857261
transform 1 0 136947 0 1 22851
box 0 0 1 1
use contact_33  contact_33_2380
timestamp 1624857261
transform 1 0 137496 0 1 22309
box 0 0 1 1
use contact_14  contact_14_321
timestamp 1624857261
transform 1 0 136943 0 1 23531
box 0 0 1 1
use contact_14  contact_14_322
timestamp 1624857261
transform 1 0 136943 0 1 23195
box 0 0 1 1
use contact_19  contact_19_321
timestamp 1624857261
transform 1 0 136940 0 1 23532
box 0 0 1 1
use contact_19  contact_19_322
timestamp 1624857261
transform 1 0 136940 0 1 23196
box 0 0 1 1
use contact_13  contact_13_321
timestamp 1624857261
transform 1 0 136947 0 1 23523
box 0 0 1 1
use contact_13  contact_13_322
timestamp 1624857261
transform 1 0 136947 0 1 23187
box 0 0 1 1
use contact_7  contact_7_64
timestamp 1624857261
transform 1 0 136939 0 1 23863
box 0 0 1 1
use contact_14  contact_14_320
timestamp 1624857261
transform 1 0 136943 0 1 23867
box 0 0 1 1
use contact_19  contact_19_320
timestamp 1624857261
transform 1 0 136940 0 1 23868
box 0 0 1 1
use contact_13  contact_13_320
timestamp 1624857261
transform 1 0 136947 0 1 23859
box 0 0 1 1
use contact_14  contact_14_318
timestamp 1624857261
transform 1 0 136943 0 1 24539
box 0 0 1 1
use contact_14  contact_14_319
timestamp 1624857261
transform 1 0 136943 0 1 24203
box 0 0 1 1
use contact_19  contact_19_318
timestamp 1624857261
transform 1 0 136940 0 1 24540
box 0 0 1 1
use contact_19  contact_19_319
timestamp 1624857261
transform 1 0 136940 0 1 24204
box 0 0 1 1
use contact_13  contact_13_318
timestamp 1624857261
transform 1 0 136947 0 1 24531
box 0 0 1 1
use contact_13  contact_13_319
timestamp 1624857261
transform 1 0 136947 0 1 24195
box 0 0 1 1
use contact_14  contact_14_317
timestamp 1624857261
transform 1 0 136943 0 1 24875
box 0 0 1 1
use contact_19  contact_19_317
timestamp 1624857261
transform 1 0 136940 0 1 24876
box 0 0 1 1
use contact_13  contact_13_317
timestamp 1624857261
transform 1 0 136947 0 1 24867
box 0 0 1 1
use contact_7  contact_7_63
timestamp 1624857261
transform 1 0 136939 0 1 25543
box 0 0 1 1
use contact_14  contact_14_315
timestamp 1624857261
transform 1 0 136943 0 1 25547
box 0 0 1 1
use contact_14  contact_14_316
timestamp 1624857261
transform 1 0 136943 0 1 25211
box 0 0 1 1
use contact_19  contact_19_315
timestamp 1624857261
transform 1 0 136940 0 1 25548
box 0 0 1 1
use contact_19  contact_19_316
timestamp 1624857261
transform 1 0 136940 0 1 25212
box 0 0 1 1
use contact_13  contact_13_315
timestamp 1624857261
transform 1 0 136947 0 1 25539
box 0 0 1 1
use contact_13  contact_13_316
timestamp 1624857261
transform 1 0 136947 0 1 25203
box 0 0 1 1
use contact_33  contact_33_2402
timestamp 1624857261
transform 1 0 137496 0 1 25573
box 0 0 1 1
use contact_33  contact_33_2355
timestamp 1624857261
transform 1 0 137496 0 1 23941
box 0 0 1 1
use contact_14  contact_14_314
timestamp 1624857261
transform 1 0 136943 0 1 25883
box 0 0 1 1
use contact_19  contact_19_314
timestamp 1624857261
transform 1 0 136940 0 1 25884
box 0 0 1 1
use contact_13  contact_13_314
timestamp 1624857261
transform 1 0 136947 0 1 25875
box 0 0 1 1
use contact_14  contact_14_312
timestamp 1624857261
transform 1 0 136943 0 1 26555
box 0 0 1 1
use contact_14  contact_14_313
timestamp 1624857261
transform 1 0 136943 0 1 26219
box 0 0 1 1
use contact_19  contact_19_312
timestamp 1624857261
transform 1 0 136940 0 1 26556
box 0 0 1 1
use contact_19  contact_19_313
timestamp 1624857261
transform 1 0 136940 0 1 26220
box 0 0 1 1
use contact_13  contact_13_312
timestamp 1624857261
transform 1 0 136947 0 1 26547
box 0 0 1 1
use contact_13  contact_13_313
timestamp 1624857261
transform 1 0 136947 0 1 26211
box 0 0 1 1
use contact_7  contact_7_62
timestamp 1624857261
transform 1 0 136939 0 1 27223
box 0 0 1 1
use contact_14  contact_14_310
timestamp 1624857261
transform 1 0 136943 0 1 27227
box 0 0 1 1
use contact_14  contact_14_311
timestamp 1624857261
transform 1 0 136943 0 1 26891
box 0 0 1 1
use contact_19  contact_19_310
timestamp 1624857261
transform 1 0 136940 0 1 27228
box 0 0 1 1
use contact_19  contact_19_311
timestamp 1624857261
transform 1 0 136940 0 1 26892
box 0 0 1 1
use contact_13  contact_13_310
timestamp 1624857261
transform 1 0 136947 0 1 27219
box 0 0 1 1
use contact_13  contact_13_311
timestamp 1624857261
transform 1 0 136947 0 1 26883
box 0 0 1 1
use contact_14  contact_14_309
timestamp 1624857261
transform 1 0 136943 0 1 27563
box 0 0 1 1
use contact_19  contact_19_309
timestamp 1624857261
transform 1 0 136940 0 1 27564
box 0 0 1 1
use contact_13  contact_13_309
timestamp 1624857261
transform 1 0 136947 0 1 27555
box 0 0 1 1
use contact_14  contact_14_308
timestamp 1624857261
transform 1 0 136943 0 1 27899
box 0 0 1 1
use contact_19  contact_19_308
timestamp 1624857261
transform 1 0 136940 0 1 27900
box 0 0 1 1
use contact_13  contact_13_308
timestamp 1624857261
transform 1 0 136947 0 1 27891
box 0 0 1 1
use contact_33  contact_33_2368
timestamp 1624857261
transform 1 0 137496 0 1 27205
box 0 0 1 1
use contact_14  contact_14_306
timestamp 1624857261
transform 1 0 136943 0 1 28571
box 0 0 1 1
use contact_14  contact_14_307
timestamp 1624857261
transform 1 0 136943 0 1 28235
box 0 0 1 1
use contact_19  contact_19_306
timestamp 1624857261
transform 1 0 136940 0 1 28572
box 0 0 1 1
use contact_19  contact_19_307
timestamp 1624857261
transform 1 0 136940 0 1 28236
box 0 0 1 1
use contact_13  contact_13_306
timestamp 1624857261
transform 1 0 136947 0 1 28563
box 0 0 1 1
use contact_13  contact_13_307
timestamp 1624857261
transform 1 0 136947 0 1 28227
box 0 0 1 1
use contact_7  contact_7_61
timestamp 1624857261
transform 1 0 136939 0 1 28903
box 0 0 1 1
use contact_14  contact_14_305
timestamp 1624857261
transform 1 0 136943 0 1 28907
box 0 0 1 1
use contact_19  contact_19_305
timestamp 1624857261
transform 1 0 136940 0 1 28908
box 0 0 1 1
use contact_13  contact_13_305
timestamp 1624857261
transform 1 0 136947 0 1 28899
box 0 0 1 1
use contact_14  contact_14_303
timestamp 1624857261
transform 1 0 136943 0 1 29579
box 0 0 1 1
use contact_14  contact_14_304
timestamp 1624857261
transform 1 0 136943 0 1 29243
box 0 0 1 1
use contact_19  contact_19_303
timestamp 1624857261
transform 1 0 136940 0 1 29580
box 0 0 1 1
use contact_19  contact_19_304
timestamp 1624857261
transform 1 0 136940 0 1 29244
box 0 0 1 1
use contact_13  contact_13_303
timestamp 1624857261
transform 1 0 136947 0 1 29571
box 0 0 1 1
use contact_13  contact_13_304
timestamp 1624857261
transform 1 0 136947 0 1 29235
box 0 0 1 1
use contact_14  contact_14_302
timestamp 1624857261
transform 1 0 136943 0 1 29915
box 0 0 1 1
use contact_19  contact_19_302
timestamp 1624857261
transform 1 0 136940 0 1 29916
box 0 0 1 1
use contact_13  contact_13_302
timestamp 1624857261
transform 1 0 136947 0 1 29907
box 0 0 1 1
use contact_7  contact_7_60
timestamp 1624857261
transform 1 0 136939 0 1 30583
box 0 0 1 1
use contact_14  contact_14_300
timestamp 1624857261
transform 1 0 136943 0 1 30587
box 0 0 1 1
use contact_14  contact_14_301
timestamp 1624857261
transform 1 0 136943 0 1 30251
box 0 0 1 1
use contact_19  contact_19_300
timestamp 1624857261
transform 1 0 136940 0 1 30588
box 0 0 1 1
use contact_19  contact_19_301
timestamp 1624857261
transform 1 0 136940 0 1 30252
box 0 0 1 1
use contact_13  contact_13_300
timestamp 1624857261
transform 1 0 136947 0 1 30579
box 0 0 1 1
use contact_13  contact_13_301
timestamp 1624857261
transform 1 0 136947 0 1 30243
box 0 0 1 1
use contact_33  contact_33_2421
timestamp 1624857261
transform 1 0 137496 0 1 28973
box 0 0 1 1
use contact_33  contact_33_2408
timestamp 1624857261
transform 1 0 137496 0 1 30469
box 0 0 1 1
use contact_14  contact_14_299
timestamp 1624857261
transform 1 0 136943 0 1 30923
box 0 0 1 1
use contact_19  contact_19_299
timestamp 1624857261
transform 1 0 136940 0 1 30924
box 0 0 1 1
use contact_13  contact_13_299
timestamp 1624857261
transform 1 0 136947 0 1 30915
box 0 0 1 1
use contact_14  contact_14_297
timestamp 1624857261
transform 1 0 136943 0 1 31595
box 0 0 1 1
use contact_14  contact_14_298
timestamp 1624857261
transform 1 0 136943 0 1 31259
box 0 0 1 1
use contact_19  contact_19_297
timestamp 1624857261
transform 1 0 136940 0 1 31596
box 0 0 1 1
use contact_19  contact_19_298
timestamp 1624857261
transform 1 0 136940 0 1 31260
box 0 0 1 1
use contact_13  contact_13_297
timestamp 1624857261
transform 1 0 136947 0 1 31587
box 0 0 1 1
use contact_13  contact_13_298
timestamp 1624857261
transform 1 0 136947 0 1 31251
box 0 0 1 1
use contact_7  contact_7_59
timestamp 1624857261
transform 1 0 136939 0 1 32263
box 0 0 1 1
use contact_14  contact_14_295
timestamp 1624857261
transform 1 0 136943 0 1 32267
box 0 0 1 1
use contact_14  contact_14_296
timestamp 1624857261
transform 1 0 136943 0 1 31931
box 0 0 1 1
use contact_19  contact_19_295
timestamp 1624857261
transform 1 0 136940 0 1 32268
box 0 0 1 1
use contact_19  contact_19_296
timestamp 1624857261
transform 1 0 136940 0 1 31932
box 0 0 1 1
use contact_13  contact_13_295
timestamp 1624857261
transform 1 0 136947 0 1 32259
box 0 0 1 1
use contact_13  contact_13_296
timestamp 1624857261
transform 1 0 136947 0 1 31923
box 0 0 1 1
use contact_14  contact_14_294
timestamp 1624857261
transform 1 0 136943 0 1 32603
box 0 0 1 1
use contact_19  contact_19_294
timestamp 1624857261
transform 1 0 136940 0 1 32604
box 0 0 1 1
use contact_13  contact_13_294
timestamp 1624857261
transform 1 0 136947 0 1 32595
box 0 0 1 1
use contact_14  contact_14_293
timestamp 1624857261
transform 1 0 136943 0 1 32939
box 0 0 1 1
use contact_19  contact_19_293
timestamp 1624857261
transform 1 0 136940 0 1 32940
box 0 0 1 1
use contact_13  contact_13_293
timestamp 1624857261
transform 1 0 136947 0 1 32931
box 0 0 1 1
use contact_33  contact_33_2409
timestamp 1624857261
transform 1 0 137496 0 1 32373
box 0 0 1 1
use contact_14  contact_14_291
timestamp 1624857261
transform 1 0 136943 0 1 33611
box 0 0 1 1
use contact_14  contact_14_292
timestamp 1624857261
transform 1 0 136943 0 1 33275
box 0 0 1 1
use contact_19  contact_19_291
timestamp 1624857261
transform 1 0 136940 0 1 33612
box 0 0 1 1
use contact_19  contact_19_292
timestamp 1624857261
transform 1 0 136940 0 1 33276
box 0 0 1 1
use contact_13  contact_13_291
timestamp 1624857261
transform 1 0 136947 0 1 33603
box 0 0 1 1
use contact_13  contact_13_292
timestamp 1624857261
transform 1 0 136947 0 1 33267
box 0 0 1 1
use contact_7  contact_7_58
timestamp 1624857261
transform 1 0 136939 0 1 33943
box 0 0 1 1
use contact_14  contact_14_290
timestamp 1624857261
transform 1 0 136943 0 1 33947
box 0 0 1 1
use contact_19  contact_19_290
timestamp 1624857261
transform 1 0 136940 0 1 33948
box 0 0 1 1
use contact_13  contact_13_290
timestamp 1624857261
transform 1 0 136947 0 1 33939
box 0 0 1 1
use contact_14  contact_14_288
timestamp 1624857261
transform 1 0 136943 0 1 34619
box 0 0 1 1
use contact_14  contact_14_289
timestamp 1624857261
transform 1 0 136943 0 1 34283
box 0 0 1 1
use contact_19  contact_19_288
timestamp 1624857261
transform 1 0 136940 0 1 34620
box 0 0 1 1
use contact_19  contact_19_289
timestamp 1624857261
transform 1 0 136940 0 1 34284
box 0 0 1 1
use contact_13  contact_13_288
timestamp 1624857261
transform 1 0 136947 0 1 34611
box 0 0 1 1
use contact_13  contact_13_289
timestamp 1624857261
transform 1 0 136947 0 1 34275
box 0 0 1 1
use contact_14  contact_14_287
timestamp 1624857261
transform 1 0 136943 0 1 34955
box 0 0 1 1
use contact_19  contact_19_287
timestamp 1624857261
transform 1 0 136940 0 1 34956
box 0 0 1 1
use contact_13  contact_13_287
timestamp 1624857261
transform 1 0 136947 0 1 34947
box 0 0 1 1
use contact_7  contact_7_57
timestamp 1624857261
transform 1 0 136939 0 1 35623
box 0 0 1 1
use contact_14  contact_14_285
timestamp 1624857261
transform 1 0 136943 0 1 35627
box 0 0 1 1
use contact_14  contact_14_286
timestamp 1624857261
transform 1 0 136943 0 1 35291
box 0 0 1 1
use contact_19  contact_19_285
timestamp 1624857261
transform 1 0 136940 0 1 35628
box 0 0 1 1
use contact_19  contact_19_286
timestamp 1624857261
transform 1 0 136940 0 1 35292
box 0 0 1 1
use contact_13  contact_13_285
timestamp 1624857261
transform 1 0 136947 0 1 35619
box 0 0 1 1
use contact_13  contact_13_286
timestamp 1624857261
transform 1 0 136947 0 1 35283
box 0 0 1 1
use contact_33  contact_33_2388
timestamp 1624857261
transform 1 0 137496 0 1 35637
box 0 0 1 1
use contact_33  contact_33_2373
timestamp 1624857261
transform 1 0 137496 0 1 34005
box 0 0 1 1
use contact_14  contact_14_283
timestamp 1624857261
transform 1 0 136943 0 1 36299
box 0 0 1 1
use contact_14  contact_14_284
timestamp 1624857261
transform 1 0 136943 0 1 35963
box 0 0 1 1
use contact_19  contact_19_283
timestamp 1624857261
transform 1 0 136940 0 1 36300
box 0 0 1 1
use contact_19  contact_19_284
timestamp 1624857261
transform 1 0 136940 0 1 35964
box 0 0 1 1
use contact_13  contact_13_283
timestamp 1624857261
transform 1 0 136947 0 1 36291
box 0 0 1 1
use contact_13  contact_13_284
timestamp 1624857261
transform 1 0 136947 0 1 35955
box 0 0 1 1
use contact_14  contact_14_282
timestamp 1624857261
transform 1 0 136943 0 1 36635
box 0 0 1 1
use contact_19  contact_19_282
timestamp 1624857261
transform 1 0 136940 0 1 36636
box 0 0 1 1
use contact_13  contact_13_282
timestamp 1624857261
transform 1 0 136947 0 1 36627
box 0 0 1 1
use contact_7  contact_7_56
timestamp 1624857261
transform 1 0 136939 0 1 37303
box 0 0 1 1
use contact_14  contact_14_280
timestamp 1624857261
transform 1 0 136943 0 1 37307
box 0 0 1 1
use contact_14  contact_14_281
timestamp 1624857261
transform 1 0 136943 0 1 36971
box 0 0 1 1
use contact_19  contact_19_280
timestamp 1624857261
transform 1 0 136940 0 1 37308
box 0 0 1 1
use contact_19  contact_19_281
timestamp 1624857261
transform 1 0 136940 0 1 36972
box 0 0 1 1
use contact_13  contact_13_280
timestamp 1624857261
transform 1 0 136947 0 1 37299
box 0 0 1 1
use contact_13  contact_13_281
timestamp 1624857261
transform 1 0 136947 0 1 36963
box 0 0 1 1
use contact_14  contact_14_279
timestamp 1624857261
transform 1 0 136943 0 1 37643
box 0 0 1 1
use contact_19  contact_19_279
timestamp 1624857261
transform 1 0 136940 0 1 37644
box 0 0 1 1
use contact_13  contact_13_279
timestamp 1624857261
transform 1 0 136947 0 1 37635
box 0 0 1 1
use contact_14  contact_14_278
timestamp 1624857261
transform 1 0 136943 0 1 37979
box 0 0 1 1
use contact_19  contact_19_278
timestamp 1624857261
transform 1 0 136940 0 1 37980
box 0 0 1 1
use contact_13  contact_13_278
timestamp 1624857261
transform 1 0 136947 0 1 37971
box 0 0 1 1
use contact_33  contact_33_2422
timestamp 1624857261
transform 1 0 137496 0 1 37269
box 0 0 1 1
use contact_14  contact_14_276
timestamp 1624857261
transform 1 0 136943 0 1 38651
box 0 0 1 1
use contact_14  contact_14_277
timestamp 1624857261
transform 1 0 136943 0 1 38315
box 0 0 1 1
use contact_19  contact_19_276
timestamp 1624857261
transform 1 0 136940 0 1 38652
box 0 0 1 1
use contact_19  contact_19_277
timestamp 1624857261
transform 1 0 136940 0 1 38316
box 0 0 1 1
use contact_13  contact_13_276
timestamp 1624857261
transform 1 0 136947 0 1 38643
box 0 0 1 1
use contact_13  contact_13_277
timestamp 1624857261
transform 1 0 136947 0 1 38307
box 0 0 1 1
use contact_7  contact_7_55
timestamp 1624857261
transform 1 0 136939 0 1 38983
box 0 0 1 1
use contact_14  contact_14_275
timestamp 1624857261
transform 1 0 136943 0 1 38987
box 0 0 1 1
use contact_19  contact_19_275
timestamp 1624857261
transform 1 0 136940 0 1 38988
box 0 0 1 1
use contact_13  contact_13_275
timestamp 1624857261
transform 1 0 136947 0 1 38979
box 0 0 1 1
use contact_14  contact_14_273
timestamp 1624857261
transform 1 0 136943 0 1 39659
box 0 0 1 1
use contact_14  contact_14_274
timestamp 1624857261
transform 1 0 136943 0 1 39323
box 0 0 1 1
use contact_19  contact_19_273
timestamp 1624857261
transform 1 0 136940 0 1 39660
box 0 0 1 1
use contact_19  contact_19_274
timestamp 1624857261
transform 1 0 136940 0 1 39324
box 0 0 1 1
use contact_13  contact_13_273
timestamp 1624857261
transform 1 0 136947 0 1 39651
box 0 0 1 1
use contact_13  contact_13_274
timestamp 1624857261
transform 1 0 136947 0 1 39315
box 0 0 1 1
use contact_14  contact_14_272
timestamp 1624857261
transform 1 0 136943 0 1 39995
box 0 0 1 1
use contact_19  contact_19_272
timestamp 1624857261
transform 1 0 136940 0 1 39996
box 0 0 1 1
use contact_13  contact_13_272
timestamp 1624857261
transform 1 0 136947 0 1 39987
box 0 0 1 1
use contact_7  contact_7_54
timestamp 1624857261
transform 1 0 136939 0 1 40663
box 0 0 1 1
use contact_14  contact_14_270
timestamp 1624857261
transform 1 0 136943 0 1 40667
box 0 0 1 1
use contact_14  contact_14_271
timestamp 1624857261
transform 1 0 136943 0 1 40331
box 0 0 1 1
use contact_19  contact_19_270
timestamp 1624857261
transform 1 0 136940 0 1 40668
box 0 0 1 1
use contact_19  contact_19_271
timestamp 1624857261
transform 1 0 136940 0 1 40332
box 0 0 1 1
use contact_13  contact_13_270
timestamp 1624857261
transform 1 0 136947 0 1 40659
box 0 0 1 1
use contact_13  contact_13_271
timestamp 1624857261
transform 1 0 136947 0 1 40323
box 0 0 1 1
use contact_33  contact_33_2363
timestamp 1624857261
transform 1 0 137496 0 1 40669
box 0 0 1 1
use contact_33  contact_33_2357
timestamp 1624857261
transform 1 0 137496 0 1 38901
box 0 0 1 1
use contact_14  contact_14_268
timestamp 1624857261
transform 1 0 136943 0 1 41339
box 0 0 1 1
use contact_14  contact_14_269
timestamp 1624857261
transform 1 0 136943 0 1 41003
box 0 0 1 1
use contact_19  contact_19_268
timestamp 1624857261
transform 1 0 136940 0 1 41340
box 0 0 1 1
use contact_19  contact_19_269
timestamp 1624857261
transform 1 0 136940 0 1 41004
box 0 0 1 1
use contact_13  contact_13_268
timestamp 1624857261
transform 1 0 136947 0 1 41331
box 0 0 1 1
use contact_13  contact_13_269
timestamp 1624857261
transform 1 0 136947 0 1 40995
box 0 0 1 1
use contact_14  contact_14_267
timestamp 1624857261
transform 1 0 136943 0 1 41675
box 0 0 1 1
use contact_19  contact_19_267
timestamp 1624857261
transform 1 0 136940 0 1 41676
box 0 0 1 1
use contact_13  contact_13_267
timestamp 1624857261
transform 1 0 136947 0 1 41667
box 0 0 1 1
use contact_7  contact_7_53
timestamp 1624857261
transform 1 0 136939 0 1 42343
box 0 0 1 1
use contact_14  contact_14_265
timestamp 1624857261
transform 1 0 136943 0 1 42347
box 0 0 1 1
use contact_14  contact_14_266
timestamp 1624857261
transform 1 0 136943 0 1 42011
box 0 0 1 1
use contact_19  contact_19_265
timestamp 1624857261
transform 1 0 136940 0 1 42348
box 0 0 1 1
use contact_19  contact_19_266
timestamp 1624857261
transform 1 0 136940 0 1 42012
box 0 0 1 1
use contact_13  contact_13_265
timestamp 1624857261
transform 1 0 136947 0 1 42339
box 0 0 1 1
use contact_13  contact_13_266
timestamp 1624857261
transform 1 0 136947 0 1 42003
box 0 0 1 1
use contact_14  contact_14_264
timestamp 1624857261
transform 1 0 136943 0 1 42683
box 0 0 1 1
use contact_19  contact_19_264
timestamp 1624857261
transform 1 0 136940 0 1 42684
box 0 0 1 1
use contact_13  contact_13_264
timestamp 1624857261
transform 1 0 136947 0 1 42675
box 0 0 1 1
use contact_14  contact_14_262
timestamp 1624857261
transform 1 0 136943 0 1 43355
box 0 0 1 1
use contact_14  contact_14_263
timestamp 1624857261
transform 1 0 136943 0 1 43019
box 0 0 1 1
use contact_19  contact_19_262
timestamp 1624857261
transform 1 0 136940 0 1 43356
box 0 0 1 1
use contact_19  contact_19_263
timestamp 1624857261
transform 1 0 136940 0 1 43020
box 0 0 1 1
use contact_13  contact_13_262
timestamp 1624857261
transform 1 0 136947 0 1 43347
box 0 0 1 1
use contact_13  contact_13_263
timestamp 1624857261
transform 1 0 136947 0 1 43011
box 0 0 1 1
use contact_33  contact_33_2366
timestamp 1624857261
transform 1 0 137496 0 1 42437
box 0 0 1 1
use contact_14  contact_14_261
timestamp 1624857261
transform 1 0 136943 0 1 43691
box 0 0 1 1
use contact_19  contact_19_261
timestamp 1624857261
transform 1 0 136940 0 1 43692
box 0 0 1 1
use contact_13  contact_13_261
timestamp 1624857261
transform 1 0 136947 0 1 43683
box 0 0 1 1
use contact_7  contact_7_52
timestamp 1624857261
transform 1 0 136939 0 1 44023
box 0 0 1 1
use contact_14  contact_14_259
timestamp 1624857261
transform 1 0 136943 0 1 44363
box 0 0 1 1
use contact_14  contact_14_260
timestamp 1624857261
transform 1 0 136943 0 1 44027
box 0 0 1 1
use contact_19  contact_19_259
timestamp 1624857261
transform 1 0 136940 0 1 44364
box 0 0 1 1
use contact_19  contact_19_260
timestamp 1624857261
transform 1 0 136940 0 1 44028
box 0 0 1 1
use contact_13  contact_13_259
timestamp 1624857261
transform 1 0 136947 0 1 44355
box 0 0 1 1
use contact_13  contact_13_260
timestamp 1624857261
transform 1 0 136947 0 1 44019
box 0 0 1 1
use contact_14  contact_14_258
timestamp 1624857261
transform 1 0 136943 0 1 44699
box 0 0 1 1
use contact_19  contact_19_258
timestamp 1624857261
transform 1 0 136940 0 1 44700
box 0 0 1 1
use contact_13  contact_13_258
timestamp 1624857261
transform 1 0 136947 0 1 44691
box 0 0 1 1
use contact_14  contact_14_256
timestamp 1624857261
transform 1 0 136943 0 1 45371
box 0 0 1 1
use contact_14  contact_14_257
timestamp 1624857261
transform 1 0 136943 0 1 45035
box 0 0 1 1
use contact_19  contact_19_256
timestamp 1624857261
transform 1 0 136940 0 1 45372
box 0 0 1 1
use contact_19  contact_19_257
timestamp 1624857261
transform 1 0 136940 0 1 45036
box 0 0 1 1
use contact_13  contact_13_256
timestamp 1624857261
transform 1 0 136947 0 1 45363
box 0 0 1 1
use contact_13  contact_13_257
timestamp 1624857261
transform 1 0 136947 0 1 45027
box 0 0 1 1
use contact_7  contact_7_51
timestamp 1624857261
transform 1 0 136939 0 1 45703
box 0 0 1 1
use contact_14  contact_14_255
timestamp 1624857261
transform 1 0 136943 0 1 45707
box 0 0 1 1
use contact_19  contact_19_255
timestamp 1624857261
transform 1 0 136940 0 1 45708
box 0 0 1 1
use contact_13  contact_13_255
timestamp 1624857261
transform 1 0 136947 0 1 45699
box 0 0 1 1
use contact_33  contact_33_2424
timestamp 1624857261
transform 1 0 137496 0 1 44069
box 0 0 1 1
use contact_33  contact_33_2365
timestamp 1624857261
transform 1 0 137496 0 1 45565
box 0 0 1 1
use contact_14  contact_14_253
timestamp 1624857261
transform 1 0 136943 0 1 46379
box 0 0 1 1
use contact_14  contact_14_254
timestamp 1624857261
transform 1 0 136943 0 1 46043
box 0 0 1 1
use contact_19  contact_19_253
timestamp 1624857261
transform 1 0 136940 0 1 46380
box 0 0 1 1
use contact_19  contact_19_254
timestamp 1624857261
transform 1 0 136940 0 1 46044
box 0 0 1 1
use contact_13  contact_13_253
timestamp 1624857261
transform 1 0 136947 0 1 46371
box 0 0 1 1
use contact_13  contact_13_254
timestamp 1624857261
transform 1 0 136947 0 1 46035
box 0 0 1 1
use contact_14  contact_14_252
timestamp 1624857261
transform 1 0 136943 0 1 46715
box 0 0 1 1
use contact_19  contact_19_252
timestamp 1624857261
transform 1 0 136940 0 1 46716
box 0 0 1 1
use contact_13  contact_13_252
timestamp 1624857261
transform 1 0 136947 0 1 46707
box 0 0 1 1
use contact_7  contact_7_50
timestamp 1624857261
transform 1 0 136939 0 1 47383
box 0 0 1 1
use contact_14  contact_14_250
timestamp 1624857261
transform 1 0 136943 0 1 47387
box 0 0 1 1
use contact_14  contact_14_251
timestamp 1624857261
transform 1 0 136943 0 1 47051
box 0 0 1 1
use contact_19  contact_19_250
timestamp 1624857261
transform 1 0 136940 0 1 47388
box 0 0 1 1
use contact_19  contact_19_251
timestamp 1624857261
transform 1 0 136940 0 1 47052
box 0 0 1 1
use contact_13  contact_13_250
timestamp 1624857261
transform 1 0 136947 0 1 47379
box 0 0 1 1
use contact_13  contact_13_251
timestamp 1624857261
transform 1 0 136947 0 1 47043
box 0 0 1 1
use contact_14  contact_14_249
timestamp 1624857261
transform 1 0 136943 0 1 47723
box 0 0 1 1
use contact_19  contact_19_249
timestamp 1624857261
transform 1 0 136940 0 1 47724
box 0 0 1 1
use contact_13  contact_13_249
timestamp 1624857261
transform 1 0 136947 0 1 47715
box 0 0 1 1
use contact_14  contact_14_247
timestamp 1624857261
transform 1 0 136943 0 1 48395
box 0 0 1 1
use contact_14  contact_14_248
timestamp 1624857261
transform 1 0 136943 0 1 48059
box 0 0 1 1
use contact_19  contact_19_247
timestamp 1624857261
transform 1 0 136940 0 1 48396
box 0 0 1 1
use contact_19  contact_19_248
timestamp 1624857261
transform 1 0 136940 0 1 48060
box 0 0 1 1
use contact_13  contact_13_247
timestamp 1624857261
transform 1 0 136947 0 1 48387
box 0 0 1 1
use contact_13  contact_13_248
timestamp 1624857261
transform 1 0 136947 0 1 48051
box 0 0 1 1
use contact_33  contact_33_2376
timestamp 1624857261
transform 1 0 137496 0 1 47469
box 0 0 1 1
use contact_14  contact_14_246
timestamp 1624857261
transform 1 0 136943 0 1 48731
box 0 0 1 1
use contact_19  contact_19_246
timestamp 1624857261
transform 1 0 136940 0 1 48732
box 0 0 1 1
use contact_13  contact_13_246
timestamp 1624857261
transform 1 0 136947 0 1 48723
box 0 0 1 1
use contact_7  contact_7_49
timestamp 1624857261
transform 1 0 136939 0 1 49063
box 0 0 1 1
use contact_14  contact_14_244
timestamp 1624857261
transform 1 0 136943 0 1 49403
box 0 0 1 1
use contact_14  contact_14_245
timestamp 1624857261
transform 1 0 136943 0 1 49067
box 0 0 1 1
use contact_19  contact_19_244
timestamp 1624857261
transform 1 0 136940 0 1 49404
box 0 0 1 1
use contact_19  contact_19_245
timestamp 1624857261
transform 1 0 136940 0 1 49068
box 0 0 1 1
use contact_13  contact_13_244
timestamp 1624857261
transform 1 0 136947 0 1 49395
box 0 0 1 1
use contact_13  contact_13_245
timestamp 1624857261
transform 1 0 136947 0 1 49059
box 0 0 1 1
use contact_14  contact_14_243
timestamp 1624857261
transform 1 0 136943 0 1 49739
box 0 0 1 1
use contact_19  contact_19_243
timestamp 1624857261
transform 1 0 136940 0 1 49740
box 0 0 1 1
use contact_13  contact_13_243
timestamp 1624857261
transform 1 0 136947 0 1 49731
box 0 0 1 1
use contact_14  contact_14_241
timestamp 1624857261
transform 1 0 136943 0 1 50411
box 0 0 1 1
use contact_14  contact_14_242
timestamp 1624857261
transform 1 0 136943 0 1 50075
box 0 0 1 1
use contact_19  contact_19_241
timestamp 1624857261
transform 1 0 136940 0 1 50412
box 0 0 1 1
use contact_19  contact_19_242
timestamp 1624857261
transform 1 0 136940 0 1 50076
box 0 0 1 1
use contact_13  contact_13_241
timestamp 1624857261
transform 1 0 136947 0 1 50403
box 0 0 1 1
use contact_13  contact_13_242
timestamp 1624857261
transform 1 0 136947 0 1 50067
box 0 0 1 1
use contact_7  contact_7_48
timestamp 1624857261
transform 1 0 136939 0 1 50743
box 0 0 1 1
use contact_14  contact_14_240
timestamp 1624857261
transform 1 0 136943 0 1 50747
box 0 0 1 1
use contact_19  contact_19_240
timestamp 1624857261
transform 1 0 136940 0 1 50748
box 0 0 1 1
use contact_13  contact_13_240
timestamp 1624857261
transform 1 0 136947 0 1 50739
box 0 0 1 1
use contact_33  contact_33_2404
timestamp 1624857261
transform 1 0 137496 0 1 50869
box 0 0 1 1
use contact_33  contact_33_2354
timestamp 1624857261
transform 1 0 137496 0 1 48965
box 0 0 1 1
use contact_14  contact_14_238
timestamp 1624857261
transform 1 0 136943 0 1 51419
box 0 0 1 1
use contact_14  contact_14_239
timestamp 1624857261
transform 1 0 136943 0 1 51083
box 0 0 1 1
use contact_19  contact_19_238
timestamp 1624857261
transform 1 0 136940 0 1 51420
box 0 0 1 1
use contact_19  contact_19_239
timestamp 1624857261
transform 1 0 136940 0 1 51084
box 0 0 1 1
use contact_13  contact_13_238
timestamp 1624857261
transform 1 0 136947 0 1 51411
box 0 0 1 1
use contact_13  contact_13_239
timestamp 1624857261
transform 1 0 136947 0 1 51075
box 0 0 1 1
use contact_14  contact_14_237
timestamp 1624857261
transform 1 0 136943 0 1 51755
box 0 0 1 1
use contact_19  contact_19_237
timestamp 1624857261
transform 1 0 136940 0 1 51756
box 0 0 1 1
use contact_13  contact_13_237
timestamp 1624857261
transform 1 0 136947 0 1 51747
box 0 0 1 1
use contact_7  contact_7_47
timestamp 1624857261
transform 1 0 136939 0 1 52423
box 0 0 1 1
use contact_14  contact_14_235
timestamp 1624857261
transform 1 0 136943 0 1 52427
box 0 0 1 1
use contact_14  contact_14_236
timestamp 1624857261
transform 1 0 136943 0 1 52091
box 0 0 1 1
use contact_19  contact_19_235
timestamp 1624857261
transform 1 0 136940 0 1 52428
box 0 0 1 1
use contact_19  contact_19_236
timestamp 1624857261
transform 1 0 136940 0 1 52092
box 0 0 1 1
use contact_13  contact_13_235
timestamp 1624857261
transform 1 0 136947 0 1 52419
box 0 0 1 1
use contact_13  contact_13_236
timestamp 1624857261
transform 1 0 136947 0 1 52083
box 0 0 1 1
use contact_14  contact_14_234
timestamp 1624857261
transform 1 0 136943 0 1 52763
box 0 0 1 1
use contact_19  contact_19_234
timestamp 1624857261
transform 1 0 136940 0 1 52764
box 0 0 1 1
use contact_13  contact_13_234
timestamp 1624857261
transform 1 0 136947 0 1 52755
box 0 0 1 1
use contact_14  contact_14_232
timestamp 1624857261
transform 1 0 136943 0 1 53435
box 0 0 1 1
use contact_14  contact_14_233
timestamp 1624857261
transform 1 0 136943 0 1 53099
box 0 0 1 1
use contact_19  contact_19_232
timestamp 1624857261
transform 1 0 136940 0 1 53436
box 0 0 1 1
use contact_19  contact_19_233
timestamp 1624857261
transform 1 0 136940 0 1 53100
box 0 0 1 1
use contact_13  contact_13_232
timestamp 1624857261
transform 1 0 136947 0 1 53427
box 0 0 1 1
use contact_13  contact_13_233
timestamp 1624857261
transform 1 0 136947 0 1 53091
box 0 0 1 1
use contact_33  contact_33_2405
timestamp 1624857261
transform 1 0 137496 0 1 52501
box 0 0 1 1
use contact_14  contact_14_231
timestamp 1624857261
transform 1 0 136943 0 1 53771
box 0 0 1 1
use contact_19  contact_19_231
timestamp 1624857261
transform 1 0 136940 0 1 53772
box 0 0 1 1
use contact_13  contact_13_231
timestamp 1624857261
transform 1 0 136947 0 1 53763
box 0 0 1 1
use contact_7  contact_7_46
timestamp 1624857261
transform 1 0 136939 0 1 54103
box 0 0 1 1
use contact_14  contact_14_229
timestamp 1624857261
transform 1 0 136943 0 1 54443
box 0 0 1 1
use contact_14  contact_14_230
timestamp 1624857261
transform 1 0 136943 0 1 54107
box 0 0 1 1
use contact_19  contact_19_229
timestamp 1624857261
transform 1 0 136940 0 1 54444
box 0 0 1 1
use contact_19  contact_19_230
timestamp 1624857261
transform 1 0 136940 0 1 54108
box 0 0 1 1
use contact_13  contact_13_229
timestamp 1624857261
transform 1 0 136947 0 1 54435
box 0 0 1 1
use contact_13  contact_13_230
timestamp 1624857261
transform 1 0 136947 0 1 54099
box 0 0 1 1
use contact_14  contact_14_228
timestamp 1624857261
transform 1 0 136943 0 1 54779
box 0 0 1 1
use contact_19  contact_19_228
timestamp 1624857261
transform 1 0 136940 0 1 54780
box 0 0 1 1
use contact_13  contact_13_228
timestamp 1624857261
transform 1 0 136947 0 1 54771
box 0 0 1 1
use contact_14  contact_14_226
timestamp 1624857261
transform 1 0 136943 0 1 55451
box 0 0 1 1
use contact_14  contact_14_227
timestamp 1624857261
transform 1 0 136943 0 1 55115
box 0 0 1 1
use contact_19  contact_19_226
timestamp 1624857261
transform 1 0 136940 0 1 55452
box 0 0 1 1
use contact_19  contact_19_227
timestamp 1624857261
transform 1 0 136940 0 1 55116
box 0 0 1 1
use contact_13  contact_13_226
timestamp 1624857261
transform 1 0 136947 0 1 55443
box 0 0 1 1
use contact_13  contact_13_227
timestamp 1624857261
transform 1 0 136947 0 1 55107
box 0 0 1 1
use contact_7  contact_7_45
timestamp 1624857261
transform 1 0 136939 0 1 55783
box 0 0 1 1
use contact_14  contact_14_225
timestamp 1624857261
transform 1 0 136943 0 1 55787
box 0 0 1 1
use contact_19  contact_19_225
timestamp 1624857261
transform 1 0 136940 0 1 55788
box 0 0 1 1
use contact_13  contact_13_225
timestamp 1624857261
transform 1 0 136947 0 1 55779
box 0 0 1 1
use contact_33  contact_33_2387
timestamp 1624857261
transform 1 0 137496 0 1 55765
box 0 0 1 1
use contact_33  contact_33_2375
timestamp 1624857261
transform 1 0 137496 0 1 54133
box 0 0 1 1
use contact_14  contact_14_223
timestamp 1624857261
transform 1 0 136943 0 1 56459
box 0 0 1 1
use contact_14  contact_14_224
timestamp 1624857261
transform 1 0 136943 0 1 56123
box 0 0 1 1
use contact_19  contact_19_223
timestamp 1624857261
transform 1 0 136940 0 1 56460
box 0 0 1 1
use contact_19  contact_19_224
timestamp 1624857261
transform 1 0 136940 0 1 56124
box 0 0 1 1
use contact_13  contact_13_223
timestamp 1624857261
transform 1 0 136947 0 1 56451
box 0 0 1 1
use contact_13  contact_13_224
timestamp 1624857261
transform 1 0 136947 0 1 56115
box 0 0 1 1
use contact_14  contact_14_222
timestamp 1624857261
transform 1 0 136943 0 1 56795
box 0 0 1 1
use contact_19  contact_19_222
timestamp 1624857261
transform 1 0 136940 0 1 56796
box 0 0 1 1
use contact_13  contact_13_222
timestamp 1624857261
transform 1 0 136947 0 1 56787
box 0 0 1 1
use contact_7  contact_7_44
timestamp 1624857261
transform 1 0 136939 0 1 57463
box 0 0 1 1
use contact_14  contact_14_220
timestamp 1624857261
transform 1 0 136943 0 1 57467
box 0 0 1 1
use contact_14  contact_14_221
timestamp 1624857261
transform 1 0 136943 0 1 57131
box 0 0 1 1
use contact_19  contact_19_220
timestamp 1624857261
transform 1 0 136940 0 1 57468
box 0 0 1 1
use contact_19  contact_19_221
timestamp 1624857261
transform 1 0 136940 0 1 57132
box 0 0 1 1
use contact_13  contact_13_220
timestamp 1624857261
transform 1 0 136947 0 1 57459
box 0 0 1 1
use contact_13  contact_13_221
timestamp 1624857261
transform 1 0 136947 0 1 57123
box 0 0 1 1
use contact_14  contact_14_219
timestamp 1624857261
transform 1 0 136943 0 1 57803
box 0 0 1 1
use contact_19  contact_19_219
timestamp 1624857261
transform 1 0 136940 0 1 57804
box 0 0 1 1
use contact_13  contact_13_219
timestamp 1624857261
transform 1 0 136947 0 1 57795
box 0 0 1 1
use contact_14  contact_14_217
timestamp 1624857261
transform 1 0 136943 0 1 58475
box 0 0 1 1
use contact_14  contact_14_218
timestamp 1624857261
transform 1 0 136943 0 1 58139
box 0 0 1 1
use contact_19  contact_19_217
timestamp 1624857261
transform 1 0 136940 0 1 58476
box 0 0 1 1
use contact_19  contact_19_218
timestamp 1624857261
transform 1 0 136940 0 1 58140
box 0 0 1 1
use contact_13  contact_13_217
timestamp 1624857261
transform 1 0 136947 0 1 58467
box 0 0 1 1
use contact_13  contact_13_218
timestamp 1624857261
transform 1 0 136947 0 1 58131
box 0 0 1 1
use contact_33  contact_33_2364
timestamp 1624857261
transform 1 0 137496 0 1 57397
box 0 0 1 1
use contact_14  contact_14_216
timestamp 1624857261
transform 1 0 136943 0 1 58811
box 0 0 1 1
use contact_19  contact_19_216
timestamp 1624857261
transform 1 0 136940 0 1 58812
box 0 0 1 1
use contact_13  contact_13_216
timestamp 1624857261
transform 1 0 136947 0 1 58803
box 0 0 1 1
use contact_7  contact_7_43
timestamp 1624857261
transform 1 0 136939 0 1 59143
box 0 0 1 1
use contact_14  contact_14_214
timestamp 1624857261
transform 1 0 136943 0 1 59483
box 0 0 1 1
use contact_14  contact_14_215
timestamp 1624857261
transform 1 0 136943 0 1 59147
box 0 0 1 1
use contact_19  contact_19_214
timestamp 1624857261
transform 1 0 136940 0 1 59484
box 0 0 1 1
use contact_19  contact_19_215
timestamp 1624857261
transform 1 0 136940 0 1 59148
box 0 0 1 1
use contact_13  contact_13_214
timestamp 1624857261
transform 1 0 136947 0 1 59475
box 0 0 1 1
use contact_13  contact_13_215
timestamp 1624857261
transform 1 0 136947 0 1 59139
box 0 0 1 1
use contact_14  contact_14_212
timestamp 1624857261
transform 1 0 136943 0 1 60155
box 0 0 1 1
use contact_14  contact_14_213
timestamp 1624857261
transform 1 0 136943 0 1 59819
box 0 0 1 1
use contact_19  contact_19_212
timestamp 1624857261
transform 1 0 136940 0 1 60156
box 0 0 1 1
use contact_19  contact_19_213
timestamp 1624857261
transform 1 0 136940 0 1 59820
box 0 0 1 1
use contact_13  contact_13_212
timestamp 1624857261
transform 1 0 136947 0 1 60147
box 0 0 1 1
use contact_13  contact_13_213
timestamp 1624857261
transform 1 0 136947 0 1 59811
box 0 0 1 1
use contact_14  contact_14_211
timestamp 1624857261
transform 1 0 136943 0 1 60491
box 0 0 1 1
use contact_19  contact_19_211
timestamp 1624857261
transform 1 0 136940 0 1 60492
box 0 0 1 1
use contact_13  contact_13_211
timestamp 1624857261
transform 1 0 136947 0 1 60483
box 0 0 1 1
use contact_7  contact_7_42
timestamp 1624857261
transform 1 0 136939 0 1 60823
box 0 0 1 1
use contact_14  contact_14_210
timestamp 1624857261
transform 1 0 136943 0 1 60827
box 0 0 1 1
use contact_19  contact_19_210
timestamp 1624857261
transform 1 0 136940 0 1 60828
box 0 0 1 1
use contact_13  contact_13_210
timestamp 1624857261
transform 1 0 136947 0 1 60819
box 0 0 1 1
use contact_33  contact_33_2399
timestamp 1624857261
transform 1 0 137496 0 1 60933
box 0 0 1 1
use contact_33  contact_33_2394
timestamp 1624857261
transform 1 0 137496 0 1 59029
box 0 0 1 1
use contact_14  contact_14_208
timestamp 1624857261
transform 1 0 136943 0 1 61499
box 0 0 1 1
use contact_14  contact_14_209
timestamp 1624857261
transform 1 0 136943 0 1 61163
box 0 0 1 1
use contact_19  contact_19_208
timestamp 1624857261
transform 1 0 136940 0 1 61500
box 0 0 1 1
use contact_19  contact_19_209
timestamp 1624857261
transform 1 0 136940 0 1 61164
box 0 0 1 1
use contact_13  contact_13_208
timestamp 1624857261
transform 1 0 136947 0 1 61491
box 0 0 1 1
use contact_13  contact_13_209
timestamp 1624857261
transform 1 0 136947 0 1 61155
box 0 0 1 1
use contact_14  contact_14_207
timestamp 1624857261
transform 1 0 136943 0 1 61835
box 0 0 1 1
use contact_19  contact_19_207
timestamp 1624857261
transform 1 0 136940 0 1 61836
box 0 0 1 1
use contact_13  contact_13_207
timestamp 1624857261
transform 1 0 136947 0 1 61827
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1624857261
transform 1 0 136939 0 1 62503
box 0 0 1 1
use contact_14  contact_14_205
timestamp 1624857261
transform 1 0 136943 0 1 62507
box 0 0 1 1
use contact_14  contact_14_206
timestamp 1624857261
transform 1 0 136943 0 1 62171
box 0 0 1 1
use contact_19  contact_19_205
timestamp 1624857261
transform 1 0 136940 0 1 62508
box 0 0 1 1
use contact_19  contact_19_206
timestamp 1624857261
transform 1 0 136940 0 1 62172
box 0 0 1 1
use contact_13  contact_13_205
timestamp 1624857261
transform 1 0 136947 0 1 62499
box 0 0 1 1
use contact_13  contact_13_206
timestamp 1624857261
transform 1 0 136947 0 1 62163
box 0 0 1 1
use contact_14  contact_14_204
timestamp 1624857261
transform 1 0 136943 0 1 62843
box 0 0 1 1
use contact_19  contact_19_204
timestamp 1624857261
transform 1 0 136940 0 1 62844
box 0 0 1 1
use contact_13  contact_13_204
timestamp 1624857261
transform 1 0 136947 0 1 62835
box 0 0 1 1
use contact_14  contact_14_202
timestamp 1624857261
transform 1 0 136943 0 1 63515
box 0 0 1 1
use contact_14  contact_14_203
timestamp 1624857261
transform 1 0 136943 0 1 63179
box 0 0 1 1
use contact_19  contact_19_202
timestamp 1624857261
transform 1 0 136940 0 1 63516
box 0 0 1 1
use contact_19  contact_19_203
timestamp 1624857261
transform 1 0 136940 0 1 63180
box 0 0 1 1
use contact_13  contact_13_202
timestamp 1624857261
transform 1 0 136947 0 1 63507
box 0 0 1 1
use contact_13  contact_13_203
timestamp 1624857261
transform 1 0 136947 0 1 63171
box 0 0 1 1
use contact_33  contact_33_2374
timestamp 1624857261
transform 1 0 137496 0 1 62565
box 0 0 1 1
use contact_14  contact_14_201
timestamp 1624857261
transform 1 0 136943 0 1 63851
box 0 0 1 1
use contact_19  contact_19_201
timestamp 1624857261
transform 1 0 136940 0 1 63852
box 0 0 1 1
use contact_13  contact_13_200
timestamp 1624857261
transform 1 0 136947 0 1 64179
box 0 0 1 1
use contact_13  contact_13_201
timestamp 1624857261
transform 1 0 136947 0 1 63843
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1624857261
transform 1 0 136939 0 1 64183
box 0 0 1 1
use contact_14  contact_14_199
timestamp 1624857261
transform 1 0 136943 0 1 64523
box 0 0 1 1
use contact_14  contact_14_200
timestamp 1624857261
transform 1 0 136943 0 1 64187
box 0 0 1 1
use contact_19  contact_19_199
timestamp 1624857261
transform 1 0 136940 0 1 64524
box 0 0 1 1
use contact_19  contact_19_200
timestamp 1624857261
transform 1 0 136940 0 1 64188
box 0 0 1 1
use contact_13  contact_13_199
timestamp 1624857261
transform 1 0 136947 0 1 64515
box 0 0 1 1
use contact_14  contact_14_197
timestamp 1624857261
transform 1 0 136943 0 1 65195
box 0 0 1 1
use contact_14  contact_14_198
timestamp 1624857261
transform 1 0 136943 0 1 64859
box 0 0 1 1
use contact_19  contact_19_197
timestamp 1624857261
transform 1 0 136940 0 1 65196
box 0 0 1 1
use contact_19  contact_19_198
timestamp 1624857261
transform 1 0 136940 0 1 64860
box 0 0 1 1
use contact_13  contact_13_197
timestamp 1624857261
transform 1 0 136947 0 1 65187
box 0 0 1 1
use contact_13  contact_13_198
timestamp 1624857261
transform 1 0 136947 0 1 64851
box 0 0 1 1
use contact_14  contact_14_196
timestamp 1624857261
transform 1 0 136943 0 1 65531
box 0 0 1 1
use contact_19  contact_19_196
timestamp 1624857261
transform 1 0 136940 0 1 65532
box 0 0 1 1
use contact_13  contact_13_196
timestamp 1624857261
transform 1 0 136947 0 1 65523
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1624857261
transform 1 0 136939 0 1 65863
box 0 0 1 1
use contact_14  contact_14_195
timestamp 1624857261
transform 1 0 136943 0 1 65867
box 0 0 1 1
use contact_19  contact_19_195
timestamp 1624857261
transform 1 0 136940 0 1 65868
box 0 0 1 1
use contact_13  contact_13_195
timestamp 1624857261
transform 1 0 136947 0 1 65859
box 0 0 1 1
use contact_33  contact_33_2401
timestamp 1624857261
transform 1 0 137496 0 1 65965
box 0 0 1 1
use contact_33  contact_33_2362
timestamp 1624857261
transform 1 0 137496 0 1 64197
box 0 0 1 1
use contact_14  contact_14_193
timestamp 1624857261
transform 1 0 136943 0 1 66539
box 0 0 1 1
use contact_14  contact_14_194
timestamp 1624857261
transform 1 0 136943 0 1 66203
box 0 0 1 1
use contact_19  contact_19_193
timestamp 1624857261
transform 1 0 136940 0 1 66540
box 0 0 1 1
use contact_19  contact_19_194
timestamp 1624857261
transform 1 0 136940 0 1 66204
box 0 0 1 1
use contact_13  contact_13_193
timestamp 1624857261
transform 1 0 136947 0 1 66531
box 0 0 1 1
use contact_13  contact_13_194
timestamp 1624857261
transform 1 0 136947 0 1 66195
box 0 0 1 1
use contact_14  contact_14_192
timestamp 1624857261
transform 1 0 136943 0 1 66875
box 0 0 1 1
use contact_19  contact_19_192
timestamp 1624857261
transform 1 0 136940 0 1 66876
box 0 0 1 1
use contact_13  contact_13_192
timestamp 1624857261
transform 1 0 136947 0 1 66867
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1624857261
transform 1 0 136939 0 1 67543
box 0 0 1 1
use contact_14  contact_14_190
timestamp 1624857261
transform 1 0 136943 0 1 67547
box 0 0 1 1
use contact_14  contact_14_191
timestamp 1624857261
transform 1 0 136943 0 1 67211
box 0 0 1 1
use contact_19  contact_19_190
timestamp 1624857261
transform 1 0 136940 0 1 67548
box 0 0 1 1
use contact_19  contact_19_191
timestamp 1624857261
transform 1 0 136940 0 1 67212
box 0 0 1 1
use contact_13  contact_13_190
timestamp 1624857261
transform 1 0 136947 0 1 67539
box 0 0 1 1
use contact_13  contact_13_191
timestamp 1624857261
transform 1 0 136947 0 1 67203
box 0 0 1 1
use contact_14  contact_14_189
timestamp 1624857261
transform 1 0 136943 0 1 67883
box 0 0 1 1
use contact_19  contact_19_189
timestamp 1624857261
transform 1 0 136940 0 1 67884
box 0 0 1 1
use contact_13  contact_13_188
timestamp 1624857261
transform 1 0 136947 0 1 68211
box 0 0 1 1
use contact_13  contact_13_189
timestamp 1624857261
transform 1 0 136947 0 1 67875
box 0 0 1 1
use contact_14  contact_14_187
timestamp 1624857261
transform 1 0 136943 0 1 68555
box 0 0 1 1
use contact_14  contact_14_188
timestamp 1624857261
transform 1 0 136943 0 1 68219
box 0 0 1 1
use contact_19  contact_19_187
timestamp 1624857261
transform 1 0 136940 0 1 68556
box 0 0 1 1
use contact_19  contact_19_188
timestamp 1624857261
transform 1 0 136940 0 1 68220
box 0 0 1 1
use contact_13  contact_13_187
timestamp 1624857261
transform 1 0 136947 0 1 68547
box 0 0 1 1
use contact_33  contact_33_2390
timestamp 1624857261
transform 1 0 137496 0 1 67461
box 0 0 1 1
use contact_14  contact_14_186
timestamp 1624857261
transform 1 0 136943 0 1 68891
box 0 0 1 1
use contact_19  contact_19_186
timestamp 1624857261
transform 1 0 136940 0 1 68892
box 0 0 1 1
use contact_13  contact_13_186
timestamp 1624857261
transform 1 0 136947 0 1 68883
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1624857261
transform 1 0 136939 0 1 69223
box 0 0 1 1
use contact_14  contact_14_184
timestamp 1624857261
transform 1 0 136943 0 1 69563
box 0 0 1 1
use contact_14  contact_14_185
timestamp 1624857261
transform 1 0 136943 0 1 69227
box 0 0 1 1
use contact_19  contact_19_184
timestamp 1624857261
transform 1 0 136940 0 1 69564
box 0 0 1 1
use contact_19  contact_19_185
timestamp 1624857261
transform 1 0 136940 0 1 69228
box 0 0 1 1
use contact_13  contact_13_184
timestamp 1624857261
transform 1 0 136947 0 1 69555
box 0 0 1 1
use contact_13  contact_13_185
timestamp 1624857261
transform 1 0 136947 0 1 69219
box 0 0 1 1
use contact_14  contact_14_183
timestamp 1624857261
transform 1 0 136943 0 1 69899
box 0 0 1 1
use contact_19  contact_19_183
timestamp 1624857261
transform 1 0 136940 0 1 69900
box 0 0 1 1
use contact_13  contact_13_183
timestamp 1624857261
transform 1 0 136947 0 1 69891
box 0 0 1 1
use contact_14  contact_14_181
timestamp 1624857261
transform 1 0 136943 0 1 70571
box 0 0 1 1
use contact_14  contact_14_182
timestamp 1624857261
transform 1 0 136943 0 1 70235
box 0 0 1 1
use contact_19  contact_19_181
timestamp 1624857261
transform 1 0 136940 0 1 70572
box 0 0 1 1
use contact_19  contact_19_182
timestamp 1624857261
transform 1 0 136940 0 1 70236
box 0 0 1 1
use contact_13  contact_13_181
timestamp 1624857261
transform 1 0 136947 0 1 70563
box 0 0 1 1
use contact_13  contact_13_182
timestamp 1624857261
transform 1 0 136947 0 1 70227
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1624857261
transform 1 0 136939 0 1 70903
box 0 0 1 1
use contact_14  contact_14_180
timestamp 1624857261
transform 1 0 136943 0 1 70907
box 0 0 1 1
use contact_19  contact_19_180
timestamp 1624857261
transform 1 0 136940 0 1 70908
box 0 0 1 1
use contact_13  contact_13_180
timestamp 1624857261
transform 1 0 136947 0 1 70899
box 0 0 1 1
use contact_14  contact_14_179
timestamp 1624857261
transform 1 0 136943 0 1 71243
box 0 0 1 1
use contact_19  contact_19_179
timestamp 1624857261
transform 1 0 136940 0 1 71244
box 0 0 1 1
use contact_13  contact_13_179
timestamp 1624857261
transform 1 0 136947 0 1 71235
box 0 0 1 1
use contact_33  contact_33_2371
timestamp 1624857261
transform 1 0 137496 0 1 70997
box 0 0 1 1
use contact_33  contact_33_2361
timestamp 1624857261
transform 1 0 137496 0 1 69229
box 0 0 1 1
use contact_14  contact_14_178
timestamp 1624857261
transform 1 0 136943 0 1 71579
box 0 0 1 1
use contact_19  contact_19_178
timestamp 1624857261
transform 1 0 136940 0 1 71580
box 0 0 1 1
use contact_13  contact_13_178
timestamp 1624857261
transform 1 0 136947 0 1 71571
box 0 0 1 1
use contact_14  contact_14_176
timestamp 1624857261
transform 1 0 136943 0 1 72251
box 0 0 1 1
use contact_14  contact_14_177
timestamp 1624857261
transform 1 0 136943 0 1 71915
box 0 0 1 1
use contact_19  contact_19_176
timestamp 1624857261
transform 1 0 136940 0 1 72252
box 0 0 1 1
use contact_19  contact_19_177
timestamp 1624857261
transform 1 0 136940 0 1 71916
box 0 0 1 1
use contact_13  contact_13_176
timestamp 1624857261
transform 1 0 136947 0 1 72243
box 0 0 1 1
use contact_13  contact_13_177
timestamp 1624857261
transform 1 0 136947 0 1 71907
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1624857261
transform 1 0 136939 0 1 72583
box 0 0 1 1
use contact_14  contact_14_175
timestamp 1624857261
transform 1 0 136943 0 1 72587
box 0 0 1 1
use contact_19  contact_19_175
timestamp 1624857261
transform 1 0 136940 0 1 72588
box 0 0 1 1
use contact_13  contact_13_175
timestamp 1624857261
transform 1 0 136947 0 1 72579
box 0 0 1 1
use contact_14  contact_14_173
timestamp 1624857261
transform 1 0 136943 0 1 73259
box 0 0 1 1
use contact_14  contact_14_174
timestamp 1624857261
transform 1 0 136943 0 1 72923
box 0 0 1 1
use contact_19  contact_19_173
timestamp 1624857261
transform 1 0 136940 0 1 73260
box 0 0 1 1
use contact_19  contact_19_174
timestamp 1624857261
transform 1 0 136940 0 1 72924
box 0 0 1 1
use contact_13  contact_13_173
timestamp 1624857261
transform 1 0 136947 0 1 73251
box 0 0 1 1
use contact_13  contact_13_174
timestamp 1624857261
transform 1 0 136947 0 1 72915
box 0 0 1 1
use contact_14  contact_14_172
timestamp 1624857261
transform 1 0 136943 0 1 73595
box 0 0 1 1
use contact_19  contact_19_172
timestamp 1624857261
transform 1 0 136940 0 1 73596
box 0 0 1 1
use contact_13  contact_13_172
timestamp 1624857261
transform 1 0 136947 0 1 73587
box 0 0 1 1
use contact_33  contact_33_2391
timestamp 1624857261
transform 1 0 137496 0 1 72629
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1624857261
transform 1 0 136939 0 1 74263
box 0 0 1 1
use contact_14  contact_14_170
timestamp 1624857261
transform 1 0 136943 0 1 74267
box 0 0 1 1
use contact_14  contact_14_171
timestamp 1624857261
transform 1 0 136943 0 1 73931
box 0 0 1 1
use contact_19  contact_19_170
timestamp 1624857261
transform 1 0 136940 0 1 74268
box 0 0 1 1
use contact_19  contact_19_171
timestamp 1624857261
transform 1 0 136940 0 1 73932
box 0 0 1 1
use contact_13  contact_13_170
timestamp 1624857261
transform 1 0 136947 0 1 74259
box 0 0 1 1
use contact_13  contact_13_171
timestamp 1624857261
transform 1 0 136947 0 1 73923
box 0 0 1 1
use contact_14  contact_14_169
timestamp 1624857261
transform 1 0 136943 0 1 74603
box 0 0 1 1
use contact_19  contact_19_169
timestamp 1624857261
transform 1 0 136940 0 1 74604
box 0 0 1 1
use contact_13  contact_13_169
timestamp 1624857261
transform 1 0 136947 0 1 74595
box 0 0 1 1
use contact_14  contact_14_167
timestamp 1624857261
transform 1 0 136943 0 1 75275
box 0 0 1 1
use contact_14  contact_14_168
timestamp 1624857261
transform 1 0 136943 0 1 74939
box 0 0 1 1
use contact_19  contact_19_167
timestamp 1624857261
transform 1 0 136940 0 1 75276
box 0 0 1 1
use contact_19  contact_19_168
timestamp 1624857261
transform 1 0 136940 0 1 74940
box 0 0 1 1
use contact_13  contact_13_167
timestamp 1624857261
transform 1 0 136947 0 1 75267
box 0 0 1 1
use contact_13  contact_13_168
timestamp 1624857261
transform 1 0 136947 0 1 74931
box 0 0 1 1
use contact_14  contact_14_166
timestamp 1624857261
transform 1 0 136943 0 1 75611
box 0 0 1 1
use contact_19  contact_19_166
timestamp 1624857261
transform 1 0 136940 0 1 75612
box 0 0 1 1
use contact_13  contact_13_166
timestamp 1624857261
transform 1 0 136947 0 1 75603
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1624857261
transform 1 0 136939 0 1 75943
box 0 0 1 1
use contact_14  contact_14_165
timestamp 1624857261
transform 1 0 136943 0 1 75947
box 0 0 1 1
use contact_19  contact_19_165
timestamp 1624857261
transform 1 0 136940 0 1 75948
box 0 0 1 1
use contact_13  contact_13_164
timestamp 1624857261
transform 1 0 136947 0 1 76275
box 0 0 1 1
use contact_13  contact_13_165
timestamp 1624857261
transform 1 0 136947 0 1 75939
box 0 0 1 1
use contact_14  contact_14_164
timestamp 1624857261
transform 1 0 136943 0 1 76283
box 0 0 1 1
use contact_19  contact_19_164
timestamp 1624857261
transform 1 0 136940 0 1 76284
box 0 0 1 1
use contact_33  contact_33_2384
timestamp 1624857261
transform 1 0 137496 0 1 74261
box 0 0 1 1
use contact_33  contact_33_2353
timestamp 1624857261
transform 1 0 137496 0 1 75893
box 0 0 1 1
use contact_14  contact_14_163
timestamp 1624857261
transform 1 0 136943 0 1 76619
box 0 0 1 1
use contact_19  contact_19_163
timestamp 1624857261
transform 1 0 136940 0 1 76620
box 0 0 1 1
use contact_13  contact_13_163
timestamp 1624857261
transform 1 0 136947 0 1 76611
box 0 0 1 1
use contact_14  contact_14_161
timestamp 1624857261
transform 1 0 136943 0 1 77291
box 0 0 1 1
use contact_14  contact_14_162
timestamp 1624857261
transform 1 0 136943 0 1 76955
box 0 0 1 1
use contact_19  contact_19_161
timestamp 1624857261
transform 1 0 136940 0 1 77292
box 0 0 1 1
use contact_19  contact_19_162
timestamp 1624857261
transform 1 0 136940 0 1 76956
box 0 0 1 1
use contact_13  contact_13_161
timestamp 1624857261
transform 1 0 136947 0 1 77283
box 0 0 1 1
use contact_13  contact_13_162
timestamp 1624857261
transform 1 0 136947 0 1 76947
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1624857261
transform 1 0 136939 0 1 77623
box 0 0 1 1
use contact_14  contact_14_160
timestamp 1624857261
transform 1 0 136943 0 1 77627
box 0 0 1 1
use contact_19  contact_19_160
timestamp 1624857261
transform 1 0 136940 0 1 77628
box 0 0 1 1
use contact_13  contact_13_160
timestamp 1624857261
transform 1 0 136947 0 1 77619
box 0 0 1 1
use contact_14  contact_14_158
timestamp 1624857261
transform 1 0 136943 0 1 78299
box 0 0 1 1
use contact_14  contact_14_159
timestamp 1624857261
transform 1 0 136943 0 1 77963
box 0 0 1 1
use contact_19  contact_19_158
timestamp 1624857261
transform 1 0 136940 0 1 78300
box 0 0 1 1
use contact_19  contact_19_159
timestamp 1624857261
transform 1 0 136940 0 1 77964
box 0 0 1 1
use contact_13  contact_13_158
timestamp 1624857261
transform 1 0 136947 0 1 78291
box 0 0 1 1
use contact_13  contact_13_159
timestamp 1624857261
transform 1 0 136947 0 1 77955
box 0 0 1 1
use contact_14  contact_14_157
timestamp 1624857261
transform 1 0 136943 0 1 78635
box 0 0 1 1
use contact_19  contact_19_157
timestamp 1624857261
transform 1 0 136940 0 1 78636
box 0 0 1 1
use contact_13  contact_13_157
timestamp 1624857261
transform 1 0 136947 0 1 78627
box 0 0 1 1
use contact_33  contact_33_2378
timestamp 1624857261
transform 1 0 137496 0 1 77525
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1624857261
transform 1 0 136939 0 1 79303
box 0 0 1 1
use contact_14  contact_14_155
timestamp 1624857261
transform 1 0 136943 0 1 79307
box 0 0 1 1
use contact_14  contact_14_156
timestamp 1624857261
transform 1 0 136943 0 1 78971
box 0 0 1 1
use contact_19  contact_19_155
timestamp 1624857261
transform 1 0 136940 0 1 79308
box 0 0 1 1
use contact_19  contact_19_156
timestamp 1624857261
transform 1 0 136940 0 1 78972
box 0 0 1 1
use contact_13  contact_13_155
timestamp 1624857261
transform 1 0 136947 0 1 79299
box 0 0 1 1
use contact_13  contact_13_156
timestamp 1624857261
transform 1 0 136947 0 1 78963
box 0 0 1 1
use contact_14  contact_14_154
timestamp 1624857261
transform 1 0 136943 0 1 79643
box 0 0 1 1
use contact_19  contact_19_154
timestamp 1624857261
transform 1 0 136940 0 1 79644
box 0 0 1 1
use contact_13  contact_13_154
timestamp 1624857261
transform 1 0 136947 0 1 79635
box 0 0 1 1
use contact_14  contact_14_152
timestamp 1624857261
transform 1 0 136943 0 1 80315
box 0 0 1 1
use contact_14  contact_14_153
timestamp 1624857261
transform 1 0 136943 0 1 79979
box 0 0 1 1
use contact_19  contact_19_152
timestamp 1624857261
transform 1 0 136940 0 1 80316
box 0 0 1 1
use contact_19  contact_19_153
timestamp 1624857261
transform 1 0 136940 0 1 79980
box 0 0 1 1
use contact_13  contact_13_152
timestamp 1624857261
transform 1 0 136947 0 1 80307
box 0 0 1 1
use contact_13  contact_13_153
timestamp 1624857261
transform 1 0 136947 0 1 79971
box 0 0 1 1
use contact_14  contact_14_151
timestamp 1624857261
transform 1 0 136943 0 1 80651
box 0 0 1 1
use contact_19  contact_19_151
timestamp 1624857261
transform 1 0 136940 0 1 80652
box 0 0 1 1
use contact_13  contact_13_151
timestamp 1624857261
transform 1 0 136947 0 1 80643
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1624857261
transform 1 0 136939 0 1 80983
box 0 0 1 1
use contact_14  contact_14_149
timestamp 1624857261
transform 1 0 136943 0 1 81323
box 0 0 1 1
use contact_14  contact_14_150
timestamp 1624857261
transform 1 0 136943 0 1 80987
box 0 0 1 1
use contact_19  contact_19_149
timestamp 1624857261
transform 1 0 136940 0 1 81324
box 0 0 1 1
use contact_19  contact_19_150
timestamp 1624857261
transform 1 0 136940 0 1 80988
box 0 0 1 1
use contact_13  contact_13_149
timestamp 1624857261
transform 1 0 136947 0 1 81315
box 0 0 1 1
use contact_13  contact_13_150
timestamp 1624857261
transform 1 0 136947 0 1 80979
box 0 0 1 1
use contact_33  contact_33_2418
timestamp 1624857261
transform 1 0 137496 0 1 79429
box 0 0 1 1
use contact_33  contact_33_2359
timestamp 1624857261
transform 1 0 137496 0 1 81061
box 0 0 1 1
use contact_14  contact_14_148
timestamp 1624857261
transform 1 0 136943 0 1 81659
box 0 0 1 1
use contact_19  contact_19_148
timestamp 1624857261
transform 1 0 136940 0 1 81660
box 0 0 1 1
use contact_13  contact_13_148
timestamp 1624857261
transform 1 0 136947 0 1 81651
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1624857261
transform 1 0 136943 0 1 82331
box 0 0 1 1
use contact_14  contact_14_147
timestamp 1624857261
transform 1 0 136943 0 1 81995
box 0 0 1 1
use contact_19  contact_19_146
timestamp 1624857261
transform 1 0 136940 0 1 82332
box 0 0 1 1
use contact_19  contact_19_147
timestamp 1624857261
transform 1 0 136940 0 1 81996
box 0 0 1 1
use contact_13  contact_13_146
timestamp 1624857261
transform 1 0 136947 0 1 82323
box 0 0 1 1
use contact_13  contact_13_147
timestamp 1624857261
transform 1 0 136947 0 1 81987
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1624857261
transform 1 0 136939 0 1 82663
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1624857261
transform 1 0 136943 0 1 83003
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1624857261
transform 1 0 136943 0 1 82667
box 0 0 1 1
use contact_19  contact_19_144
timestamp 1624857261
transform 1 0 136940 0 1 83004
box 0 0 1 1
use contact_19  contact_19_145
timestamp 1624857261
transform 1 0 136940 0 1 82668
box 0 0 1 1
use contact_13  contact_13_144
timestamp 1624857261
transform 1 0 136947 0 1 82995
box 0 0 1 1
use contact_13  contact_13_145
timestamp 1624857261
transform 1 0 136947 0 1 82659
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1624857261
transform 1 0 136943 0 1 83339
box 0 0 1 1
use contact_19  contact_19_143
timestamp 1624857261
transform 1 0 136940 0 1 83340
box 0 0 1 1
use contact_13  contact_13_143
timestamp 1624857261
transform 1 0 136947 0 1 83331
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1624857261
transform 1 0 136943 0 1 83675
box 0 0 1 1
use contact_19  contact_19_142
timestamp 1624857261
transform 1 0 136940 0 1 83676
box 0 0 1 1
use contact_13  contact_13_142
timestamp 1624857261
transform 1 0 136947 0 1 83667
box 0 0 1 1
use contact_33  contact_33_2395
timestamp 1624857261
transform 1 0 137496 0 1 82693
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1624857261
transform 1 0 136939 0 1 84343
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1624857261
transform 1 0 136943 0 1 84347
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1624857261
transform 1 0 136943 0 1 84011
box 0 0 1 1
use contact_19  contact_19_140
timestamp 1624857261
transform 1 0 136940 0 1 84348
box 0 0 1 1
use contact_19  contact_19_141
timestamp 1624857261
transform 1 0 136940 0 1 84012
box 0 0 1 1
use contact_13  contact_13_140
timestamp 1624857261
transform 1 0 136947 0 1 84339
box 0 0 1 1
use contact_13  contact_13_141
timestamp 1624857261
transform 1 0 136947 0 1 84003
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1624857261
transform 1 0 136943 0 1 84683
box 0 0 1 1
use contact_19  contact_19_139
timestamp 1624857261
transform 1 0 136940 0 1 84684
box 0 0 1 1
use contact_13  contact_13_139
timestamp 1624857261
transform 1 0 136947 0 1 84675
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1624857261
transform 1 0 136943 0 1 85355
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1624857261
transform 1 0 136943 0 1 85019
box 0 0 1 1
use contact_19  contact_19_137
timestamp 1624857261
transform 1 0 136940 0 1 85356
box 0 0 1 1
use contact_19  contact_19_138
timestamp 1624857261
transform 1 0 136940 0 1 85020
box 0 0 1 1
use contact_13  contact_13_137
timestamp 1624857261
transform 1 0 136947 0 1 85347
box 0 0 1 1
use contact_13  contact_13_138
timestamp 1624857261
transform 1 0 136947 0 1 85011
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1624857261
transform 1 0 136943 0 1 85691
box 0 0 1 1
use contact_19  contact_19_136
timestamp 1624857261
transform 1 0 136940 0 1 85692
box 0 0 1 1
use contact_13  contact_13_136
timestamp 1624857261
transform 1 0 136947 0 1 85683
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1624857261
transform 1 0 136939 0 1 86023
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1624857261
transform 1 0 136943 0 1 86363
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1624857261
transform 1 0 136943 0 1 86027
box 0 0 1 1
use contact_19  contact_19_134
timestamp 1624857261
transform 1 0 136940 0 1 86364
box 0 0 1 1
use contact_19  contact_19_135
timestamp 1624857261
transform 1 0 136940 0 1 86028
box 0 0 1 1
use contact_13  contact_13_134
timestamp 1624857261
transform 1 0 136947 0 1 86355
box 0 0 1 1
use contact_13  contact_13_135
timestamp 1624857261
transform 1 0 136947 0 1 86019
box 0 0 1 1
use contact_33  contact_33_2381
timestamp 1624857261
transform 1 0 137496 0 1 85957
box 0 0 1 1
use contact_33  contact_33_2370
timestamp 1624857261
transform 1 0 137496 0 1 84461
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1624857261
transform 1 0 136943 0 1 86699
box 0 0 1 1
use contact_19  contact_19_133
timestamp 1624857261
transform 1 0 136940 0 1 86700
box 0 0 1 1
use contact_13  contact_13_133
timestamp 1624857261
transform 1 0 136947 0 1 86691
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1624857261
transform 1 0 136943 0 1 87371
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1624857261
transform 1 0 136943 0 1 87035
box 0 0 1 1
use contact_19  contact_19_131
timestamp 1624857261
transform 1 0 136940 0 1 87372
box 0 0 1 1
use contact_19  contact_19_132
timestamp 1624857261
transform 1 0 136940 0 1 87036
box 0 0 1 1
use contact_13  contact_13_131
timestamp 1624857261
transform 1 0 136947 0 1 87363
box 0 0 1 1
use contact_13  contact_13_132
timestamp 1624857261
transform 1 0 136947 0 1 87027
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1624857261
transform 1 0 136939 0 1 87703
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1624857261
transform 1 0 136943 0 1 88043
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1624857261
transform 1 0 136943 0 1 87707
box 0 0 1 1
use contact_19  contact_19_129
timestamp 1624857261
transform 1 0 136940 0 1 88044
box 0 0 1 1
use contact_19  contact_19_130
timestamp 1624857261
transform 1 0 136940 0 1 87708
box 0 0 1 1
use contact_13  contact_13_129
timestamp 1624857261
transform 1 0 136947 0 1 88035
box 0 0 1 1
use contact_13  contact_13_130
timestamp 1624857261
transform 1 0 136947 0 1 87699
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1624857261
transform 1 0 136943 0 1 88379
box 0 0 1 1
use contact_19  contact_19_128
timestamp 1624857261
transform 1 0 136940 0 1 88380
box 0 0 1 1
use contact_13  contact_13_128
timestamp 1624857261
transform 1 0 136947 0 1 88371
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1624857261
transform 1 0 136943 0 1 88715
box 0 0 1 1
use contact_19  contact_19_127
timestamp 1624857261
transform 1 0 136940 0 1 88716
box 0 0 1 1
use contact_13  contact_13_127
timestamp 1624857261
transform 1 0 136947 0 1 88707
box 0 0 1 1
use contact_33  contact_33_2360
timestamp 1624857261
transform 1 0 137496 0 1 87725
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1624857261
transform 1 0 136939 0 1 89383
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1624857261
transform 1 0 136943 0 1 89387
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1624857261
transform 1 0 136943 0 1 89051
box 0 0 1 1
use contact_19  contact_19_125
timestamp 1624857261
transform 1 0 136940 0 1 89388
box 0 0 1 1
use contact_19  contact_19_126
timestamp 1624857261
transform 1 0 136940 0 1 89052
box 0 0 1 1
use contact_13  contact_13_125
timestamp 1624857261
transform 1 0 136947 0 1 89379
box 0 0 1 1
use contact_13  contact_13_126
timestamp 1624857261
transform 1 0 136947 0 1 89043
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1624857261
transform 1 0 136943 0 1 89723
box 0 0 1 1
use contact_19  contact_19_124
timestamp 1624857261
transform 1 0 136940 0 1 89724
box 0 0 1 1
use contact_13  contact_13_124
timestamp 1624857261
transform 1 0 136947 0 1 89715
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1624857261
transform 1 0 136943 0 1 90395
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1624857261
transform 1 0 136943 0 1 90059
box 0 0 1 1
use contact_19  contact_19_122
timestamp 1624857261
transform 1 0 136940 0 1 90396
box 0 0 1 1
use contact_19  contact_19_123
timestamp 1624857261
transform 1 0 136940 0 1 90060
box 0 0 1 1
use contact_13  contact_13_122
timestamp 1624857261
transform 1 0 136947 0 1 90387
box 0 0 1 1
use contact_13  contact_13_123
timestamp 1624857261
transform 1 0 136947 0 1 90051
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1624857261
transform 1 0 136943 0 1 90731
box 0 0 1 1
use contact_19  contact_19_121
timestamp 1624857261
transform 1 0 136940 0 1 90732
box 0 0 1 1
use contact_13  contact_13_121
timestamp 1624857261
transform 1 0 136947 0 1 90723
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1624857261
transform 1 0 136939 0 1 91063
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1624857261
transform 1 0 136943 0 1 91403
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1624857261
transform 1 0 136943 0 1 91067
box 0 0 1 1
use contact_19  contact_19_119
timestamp 1624857261
transform 1 0 136940 0 1 91404
box 0 0 1 1
use contact_19  contact_19_120
timestamp 1624857261
transform 1 0 136940 0 1 91068
box 0 0 1 1
use contact_13  contact_13_119
timestamp 1624857261
transform 1 0 136947 0 1 91395
box 0 0 1 1
use contact_13  contact_13_120
timestamp 1624857261
transform 1 0 136947 0 1 91059
box 0 0 1 1
use contact_33  contact_33_2423
timestamp 1624857261
transform 1 0 137496 0 1 89493
box 0 0 1 1
use contact_33  contact_33_2416
timestamp 1624857261
transform 1 0 137496 0 1 91125
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1624857261
transform 1 0 136943 0 1 92075
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1624857261
transform 1 0 136943 0 1 91739
box 0 0 1 1
use contact_19  contact_19_117
timestamp 1624857261
transform 1 0 136940 0 1 92076
box 0 0 1 1
use contact_19  contact_19_118
timestamp 1624857261
transform 1 0 136940 0 1 91740
box 0 0 1 1
use contact_13  contact_13_117
timestamp 1624857261
transform 1 0 136947 0 1 92067
box 0 0 1 1
use contact_13  contact_13_118
timestamp 1624857261
transform 1 0 136947 0 1 91731
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1624857261
transform 1 0 136943 0 1 92411
box 0 0 1 1
use contact_19  contact_19_116
timestamp 1624857261
transform 1 0 136940 0 1 92412
box 0 0 1 1
use contact_13  contact_13_116
timestamp 1624857261
transform 1 0 136947 0 1 92403
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1624857261
transform 1 0 136939 0 1 92743
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1624857261
transform 1 0 136943 0 1 93083
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1624857261
transform 1 0 136943 0 1 92747
box 0 0 1 1
use contact_19  contact_19_114
timestamp 1624857261
transform 1 0 136940 0 1 93084
box 0 0 1 1
use contact_19  contact_19_115
timestamp 1624857261
transform 1 0 136940 0 1 92748
box 0 0 1 1
use contact_13  contact_13_114
timestamp 1624857261
transform 1 0 136947 0 1 93075
box 0 0 1 1
use contact_13  contact_13_115
timestamp 1624857261
transform 1 0 136947 0 1 92739
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1624857261
transform 1 0 136943 0 1 93419
box 0 0 1 1
use contact_19  contact_19_113
timestamp 1624857261
transform 1 0 136940 0 1 93420
box 0 0 1 1
use contact_13  contact_13_113
timestamp 1624857261
transform 1 0 136947 0 1 93411
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1624857261
transform 1 0 136943 0 1 93755
box 0 0 1 1
use contact_19  contact_19_112
timestamp 1624857261
transform 1 0 136940 0 1 93756
box 0 0 1 1
use contact_13  contact_13_112
timestamp 1624857261
transform 1 0 136947 0 1 93747
box 0 0 1 1
use contact_33  contact_33_2410
timestamp 1624857261
transform 1 0 137496 0 1 92893
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1624857261
transform 1 0 136939 0 1 94423
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1624857261
transform 1 0 136943 0 1 94427
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1624857261
transform 1 0 136943 0 1 94091
box 0 0 1 1
use contact_19  contact_19_110
timestamp 1624857261
transform 1 0 136940 0 1 94428
box 0 0 1 1
use contact_19  contact_19_111
timestamp 1624857261
transform 1 0 136940 0 1 94092
box 0 0 1 1
use contact_13  contact_13_110
timestamp 1624857261
transform 1 0 136947 0 1 94419
box 0 0 1 1
use contact_13  contact_13_111
timestamp 1624857261
transform 1 0 136947 0 1 94083
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1624857261
transform 1 0 136943 0 1 94763
box 0 0 1 1
use contact_19  contact_19_109
timestamp 1624857261
transform 1 0 136940 0 1 94764
box 0 0 1 1
use contact_13  contact_13_109
timestamp 1624857261
transform 1 0 136947 0 1 94755
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1624857261
transform 1 0 136943 0 1 95435
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1624857261
transform 1 0 136943 0 1 95099
box 0 0 1 1
use contact_19  contact_19_107
timestamp 1624857261
transform 1 0 136940 0 1 95436
box 0 0 1 1
use contact_19  contact_19_108
timestamp 1624857261
transform 1 0 136940 0 1 95100
box 0 0 1 1
use contact_13  contact_13_107
timestamp 1624857261
transform 1 0 136947 0 1 95427
box 0 0 1 1
use contact_13  contact_13_108
timestamp 1624857261
transform 1 0 136947 0 1 95091
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1624857261
transform 1 0 136943 0 1 95771
box 0 0 1 1
use contact_19  contact_19_106
timestamp 1624857261
transform 1 0 136940 0 1 95772
box 0 0 1 1
use contact_13  contact_13_106
timestamp 1624857261
transform 1 0 136947 0 1 95763
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1624857261
transform 1 0 136939 0 1 96103
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1624857261
transform 1 0 136943 0 1 96443
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1624857261
transform 1 0 136943 0 1 96107
box 0 0 1 1
use contact_19  contact_19_104
timestamp 1624857261
transform 1 0 136940 0 1 96444
box 0 0 1 1
use contact_19  contact_19_105
timestamp 1624857261
transform 1 0 136940 0 1 96108
box 0 0 1 1
use contact_13  contact_13_104
timestamp 1624857261
transform 1 0 136947 0 1 96435
box 0 0 1 1
use contact_13  contact_13_105
timestamp 1624857261
transform 1 0 136947 0 1 96099
box 0 0 1 1
use contact_33  contact_33_2425
timestamp 1624857261
transform 1 0 137496 0 1 94389
box 0 0 1 1
use contact_33  contact_33_2397
timestamp 1624857261
transform 1 0 137496 0 1 96021
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1624857261
transform 1 0 136943 0 1 96779
box 0 0 1 1
use contact_19  contact_19_103
timestamp 1624857261
transform 1 0 136940 0 1 96780
box 0 0 1 1
use contact_13  contact_13_102
timestamp 1624857261
transform 1 0 136947 0 1 97107
box 0 0 1 1
use contact_13  contact_13_103
timestamp 1624857261
transform 1 0 136947 0 1 96771
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1624857261
transform 1 0 136943 0 1 97451
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1624857261
transform 1 0 136943 0 1 97115
box 0 0 1 1
use contact_19  contact_19_101
timestamp 1624857261
transform 1 0 136940 0 1 97452
box 0 0 1 1
use contact_19  contact_19_102
timestamp 1624857261
transform 1 0 136940 0 1 97116
box 0 0 1 1
use contact_13  contact_13_101
timestamp 1624857261
transform 1 0 136947 0 1 97443
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1624857261
transform 1 0 136939 0 1 97783
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1624857261
transform 1 0 136943 0 1 98123
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1624857261
transform 1 0 136943 0 1 97787
box 0 0 1 1
use contact_19  contact_19_99
timestamp 1624857261
transform 1 0 136940 0 1 98124
box 0 0 1 1
use contact_19  contact_19_100
timestamp 1624857261
transform 1 0 136940 0 1 97788
box 0 0 1 1
use contact_13  contact_13_99
timestamp 1624857261
transform 1 0 136947 0 1 98115
box 0 0 1 1
use contact_13  contact_13_100
timestamp 1624857261
transform 1 0 136947 0 1 97779
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1624857261
transform 1 0 136943 0 1 98459
box 0 0 1 1
use contact_19  contact_19_98
timestamp 1624857261
transform 1 0 136940 0 1 98460
box 0 0 1 1
use contact_13  contact_13_98
timestamp 1624857261
transform 1 0 136947 0 1 98451
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1624857261
transform 1 0 136943 0 1 99131
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1624857261
transform 1 0 136943 0 1 98795
box 0 0 1 1
use contact_19  contact_19_96
timestamp 1624857261
transform 1 0 136940 0 1 99132
box 0 0 1 1
use contact_19  contact_19_97
timestamp 1624857261
transform 1 0 136940 0 1 98796
box 0 0 1 1
use contact_13  contact_13_96
timestamp 1624857261
transform 1 0 136947 0 1 99123
box 0 0 1 1
use contact_13  contact_13_97
timestamp 1624857261
transform 1 0 136947 0 1 98787
box 0 0 1 1
use contact_33  contact_33_2426
timestamp 1624857261
transform 1 0 137496 0 1 97789
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1624857261
transform 1 0 136939 0 1 99463
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1624857261
transform 1 0 136943 0 1 99467
box 0 0 1 1
use contact_19  contact_19_95
timestamp 1624857261
transform 1 0 136940 0 1 99468
box 0 0 1 1
use contact_13  contact_13_95
timestamp 1624857261
transform 1 0 136947 0 1 99459
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1624857261
transform 1 0 136943 0 1 100139
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1624857261
transform 1 0 136943 0 1 99803
box 0 0 1 1
use contact_19  contact_19_93
timestamp 1624857261
transform 1 0 136940 0 1 100140
box 0 0 1 1
use contact_19  contact_19_94
timestamp 1624857261
transform 1 0 136940 0 1 99804
box 0 0 1 1
use contact_13  contact_13_93
timestamp 1624857261
transform 1 0 136947 0 1 100131
box 0 0 1 1
use contact_13  contact_13_94
timestamp 1624857261
transform 1 0 136947 0 1 99795
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1624857261
transform 1 0 136943 0 1 100475
box 0 0 1 1
use contact_19  contact_19_92
timestamp 1624857261
transform 1 0 136940 0 1 100476
box 0 0 1 1
use contact_13  contact_13_92
timestamp 1624857261
transform 1 0 136947 0 1 100467
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1624857261
transform 1 0 136939 0 1 101143
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1624857261
transform 1 0 136943 0 1 101147
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1624857261
transform 1 0 136943 0 1 100811
box 0 0 1 1
use contact_19  contact_19_90
timestamp 1624857261
transform 1 0 136940 0 1 101148
box 0 0 1 1
use contact_19  contact_19_91
timestamp 1624857261
transform 1 0 136940 0 1 100812
box 0 0 1 1
use contact_13  contact_13_90
timestamp 1624857261
transform 1 0 136947 0 1 101139
box 0 0 1 1
use contact_13  contact_13_91
timestamp 1624857261
transform 1 0 136947 0 1 100803
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1624857261
transform 1 0 136943 0 1 101483
box 0 0 1 1
use contact_19  contact_19_89
timestamp 1624857261
transform 1 0 136940 0 1 101484
box 0 0 1 1
use contact_13  contact_13_89
timestamp 1624857261
transform 1 0 136947 0 1 101475
box 0 0 1 1
use contact_33  contact_33_2415
timestamp 1624857261
transform 1 0 137496 0 1 101189
box 0 0 1 1
use contact_33  contact_33_2412
timestamp 1624857261
transform 1 0 137496 0 1 99557
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1624857261
transform 1 0 136943 0 1 102155
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1624857261
transform 1 0 136943 0 1 101819
box 0 0 1 1
use contact_19  contact_19_87
timestamp 1624857261
transform 1 0 136940 0 1 102156
box 0 0 1 1
use contact_19  contact_19_88
timestamp 1624857261
transform 1 0 136940 0 1 101820
box 0 0 1 1
use contact_13  contact_13_87
timestamp 1624857261
transform 1 0 136947 0 1 102147
box 0 0 1 1
use contact_13  contact_13_88
timestamp 1624857261
transform 1 0 136947 0 1 101811
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1624857261
transform 1 0 136943 0 1 102491
box 0 0 1 1
use contact_19  contact_19_86
timestamp 1624857261
transform 1 0 136940 0 1 102492
box 0 0 1 1
use contact_13  contact_13_86
timestamp 1624857261
transform 1 0 136947 0 1 102483
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1624857261
transform 1 0 136939 0 1 102823
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1624857261
transform 1 0 136943 0 1 103163
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1624857261
transform 1 0 136943 0 1 102827
box 0 0 1 1
use contact_19  contact_19_84
timestamp 1624857261
transform 1 0 136940 0 1 103164
box 0 0 1 1
use contact_19  contact_19_85
timestamp 1624857261
transform 1 0 136940 0 1 102828
box 0 0 1 1
use contact_13  contact_13_84
timestamp 1624857261
transform 1 0 136947 0 1 103155
box 0 0 1 1
use contact_13  contact_13_85
timestamp 1624857261
transform 1 0 136947 0 1 102819
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1624857261
transform 1 0 136943 0 1 103499
box 0 0 1 1
use contact_19  contact_19_83
timestamp 1624857261
transform 1 0 136940 0 1 103500
box 0 0 1 1
use contact_13  contact_13_83
timestamp 1624857261
transform 1 0 136947 0 1 103491
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1624857261
transform 1 0 136943 0 1 104171
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1624857261
transform 1 0 136943 0 1 103835
box 0 0 1 1
use contact_19  contact_19_81
timestamp 1624857261
transform 1 0 136940 0 1 104172
box 0 0 1 1
use contact_19  contact_19_82
timestamp 1624857261
transform 1 0 136940 0 1 103836
box 0 0 1 1
use contact_13  contact_13_81
timestamp 1624857261
transform 1 0 136947 0 1 104163
box 0 0 1 1
use contact_13  contact_13_82
timestamp 1624857261
transform 1 0 136947 0 1 103827
box 0 0 1 1
use contact_33  contact_33_2414
timestamp 1624857261
transform 1 0 137496 0 1 102821
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1624857261
transform 1 0 136939 0 1 104503
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1624857261
transform 1 0 136943 0 1 104507
box 0 0 1 1
use contact_19  contact_19_80
timestamp 1624857261
transform 1 0 136940 0 1 104508
box 0 0 1 1
use contact_13  contact_13_80
timestamp 1624857261
transform 1 0 136947 0 1 104499
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1624857261
transform 1 0 136943 0 1 105179
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1624857261
transform 1 0 136943 0 1 104843
box 0 0 1 1
use contact_19  contact_19_78
timestamp 1624857261
transform 1 0 136940 0 1 105180
box 0 0 1 1
use contact_19  contact_19_79
timestamp 1624857261
transform 1 0 136940 0 1 104844
box 0 0 1 1
use contact_13  contact_13_78
timestamp 1624857261
transform 1 0 136947 0 1 105171
box 0 0 1 1
use contact_13  contact_13_79
timestamp 1624857261
transform 1 0 136947 0 1 104835
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1624857261
transform 1 0 136943 0 1 105515
box 0 0 1 1
use contact_19  contact_19_77
timestamp 1624857261
transform 1 0 136940 0 1 105516
box 0 0 1 1
use contact_13  contact_13_77
timestamp 1624857261
transform 1 0 136947 0 1 105507
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1624857261
transform 1 0 136939 0 1 106183
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1624857261
transform 1 0 136943 0 1 106187
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1624857261
transform 1 0 136943 0 1 105851
box 0 0 1 1
use contact_19  contact_19_75
timestamp 1624857261
transform 1 0 136940 0 1 106188
box 0 0 1 1
use contact_19  contact_19_76
timestamp 1624857261
transform 1 0 136940 0 1 105852
box 0 0 1 1
use contact_13  contact_13_75
timestamp 1624857261
transform 1 0 136947 0 1 106179
box 0 0 1 1
use contact_13  contact_13_76
timestamp 1624857261
transform 1 0 136947 0 1 105843
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1624857261
transform 1 0 136943 0 1 106523
box 0 0 1 1
use contact_19  contact_19_74
timestamp 1624857261
transform 1 0 136940 0 1 106524
box 0 0 1 1
use contact_13  contact_13_74
timestamp 1624857261
transform 1 0 136947 0 1 106515
box 0 0 1 1
use contact_33  contact_33_2407
timestamp 1624857261
transform 1 0 137496 0 1 104453
box 0 0 1 1
use contact_33  contact_33_2358
timestamp 1624857261
transform 1 0 137496 0 1 106221
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1624857261
transform 1 0 136943 0 1 107195
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1624857261
transform 1 0 136943 0 1 106859
box 0 0 1 1
use contact_19  contact_19_72
timestamp 1624857261
transform 1 0 136940 0 1 107196
box 0 0 1 1
use contact_19  contact_19_73
timestamp 1624857261
transform 1 0 136940 0 1 106860
box 0 0 1 1
use contact_13  contact_13_72
timestamp 1624857261
transform 1 0 136947 0 1 107187
box 0 0 1 1
use contact_13  contact_13_73
timestamp 1624857261
transform 1 0 136947 0 1 106851
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1624857261
transform 1 0 136943 0 1 107531
box 0 0 1 1
use contact_19  contact_19_71
timestamp 1624857261
transform 1 0 136940 0 1 107532
box 0 0 1 1
use contact_13  contact_13_71
timestamp 1624857261
transform 1 0 136947 0 1 107523
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1624857261
transform 1 0 136939 0 1 107863
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1624857261
transform 1 0 136943 0 1 108203
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1624857261
transform 1 0 136943 0 1 107867
box 0 0 1 1
use contact_19  contact_19_69
timestamp 1624857261
transform 1 0 136940 0 1 108204
box 0 0 1 1
use contact_19  contact_19_70
timestamp 1624857261
transform 1 0 136940 0 1 107868
box 0 0 1 1
use contact_13  contact_13_69
timestamp 1624857261
transform 1 0 136947 0 1 108195
box 0 0 1 1
use contact_13  contact_13_70
timestamp 1624857261
transform 1 0 136947 0 1 107859
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1624857261
transform 1 0 136943 0 1 108539
box 0 0 1 1
use contact_19  contact_19_68
timestamp 1624857261
transform 1 0 136940 0 1 108540
box 0 0 1 1
use contact_13  contact_13_68
timestamp 1624857261
transform 1 0 136947 0 1 108531
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1624857261
transform 1 0 136943 0 1 109211
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1624857261
transform 1 0 136943 0 1 108875
box 0 0 1 1
use contact_19  contact_19_66
timestamp 1624857261
transform 1 0 136940 0 1 109212
box 0 0 1 1
use contact_19  contact_19_67
timestamp 1624857261
transform 1 0 136940 0 1 108876
box 0 0 1 1
use contact_13  contact_13_66
timestamp 1624857261
transform 1 0 136947 0 1 109203
box 0 0 1 1
use contact_13  contact_13_67
timestamp 1624857261
transform 1 0 136947 0 1 108867
box 0 0 1 1
use contact_33  contact_33_2400
timestamp 1624857261
transform 1 0 137496 0 1 107989
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1624857261
transform 1 0 136939 0 1 109543
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1624857261
transform 1 0 136943 0 1 109547
box 0 0 1 1
use contact_19  contact_19_65
timestamp 1624857261
transform 1 0 136940 0 1 109548
box 0 0 1 1
use contact_13  contact_13_65
timestamp 1624857261
transform 1 0 136947 0 1 109539
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1624857261
transform 1 0 136943 0 1 110219
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1624857261
transform 1 0 136943 0 1 109883
box 0 0 1 1
use contact_19  contact_19_63
timestamp 1624857261
transform 1 0 136940 0 1 110220
box 0 0 1 1
use contact_19  contact_19_64
timestamp 1624857261
transform 1 0 136940 0 1 109884
box 0 0 1 1
use contact_13  contact_13_63
timestamp 1624857261
transform 1 0 136947 0 1 110211
box 0 0 1 1
use contact_13  contact_13_64
timestamp 1624857261
transform 1 0 136947 0 1 109875
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1624857261
transform 1 0 136943 0 1 110555
box 0 0 1 1
use contact_19  contact_19_62
timestamp 1624857261
transform 1 0 136940 0 1 110556
box 0 0 1 1
use contact_13  contact_13_62
timestamp 1624857261
transform 1 0 136947 0 1 110547
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1624857261
transform 1 0 136939 0 1 111223
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1624857261
transform 1 0 136943 0 1 111227
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1624857261
transform 1 0 136943 0 1 110891
box 0 0 1 1
use contact_19  contact_19_60
timestamp 1624857261
transform 1 0 136940 0 1 111228
box 0 0 1 1
use contact_19  contact_19_61
timestamp 1624857261
transform 1 0 136940 0 1 110892
box 0 0 1 1
use contact_13  contact_13_60
timestamp 1624857261
transform 1 0 136947 0 1 111219
box 0 0 1 1
use contact_13  contact_13_61
timestamp 1624857261
transform 1 0 136947 0 1 110883
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1624857261
transform 1 0 136943 0 1 111563
box 0 0 1 1
use contact_19  contact_19_59
timestamp 1624857261
transform 1 0 136940 0 1 111564
box 0 0 1 1
use contact_13  contact_13_59
timestamp 1624857261
transform 1 0 136947 0 1 111555
box 0 0 1 1
use contact_33  contact_33_2382
timestamp 1624857261
transform 1 0 137496 0 1 111253
box 0 0 1 1
use contact_33  contact_33_2379
timestamp 1624857261
transform 1 0 137496 0 1 109621
box 0 0 1 1
use contact_33  contact_33_6
timestamp 1624857261
transform 1 0 135320 0 1 112069
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1624857261
transform 1 0 136943 0 1 112235
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1624857261
transform 1 0 136943 0 1 111899
box 0 0 1 1
use contact_19  contact_19_57
timestamp 1624857261
transform 1 0 136940 0 1 112236
box 0 0 1 1
use contact_19  contact_19_58
timestamp 1624857261
transform 1 0 136940 0 1 111900
box 0 0 1 1
use contact_13  contact_13_57
timestamp 1624857261
transform 1 0 136947 0 1 112227
box 0 0 1 1
use contact_13  contact_13_58
timestamp 1624857261
transform 1 0 136947 0 1 111891
box 0 0 1 1
use contact_7  contact_7_475
timestamp 1624857261
transform 1 0 136192 0 1 112614
box 0 0 1 1
use contact_33  contact_33_5491
timestamp 1624857261
transform 1 0 136187 0 1 112618
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1624857261
transform 1 0 136943 0 1 112571
box 0 0 1 1
use contact_19  contact_19_56
timestamp 1624857261
transform 1 0 136940 0 1 112572
box 0 0 1 1
use contact_13  contact_13_56
timestamp 1624857261
transform 1 0 136947 0 1 112563
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1624857261
transform 1 0 136939 0 1 112903
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1624857261
transform 1 0 136943 0 1 112907
box 0 0 1 1
use contact_19  contact_19_55
timestamp 1624857261
transform 1 0 136940 0 1 112908
box 0 0 1 1
use contact_13  contact_13_55
timestamp 1624857261
transform 1 0 136947 0 1 112899
box 0 0 1 1
use contact_33  contact_33_2440
timestamp 1624857261
transform 1 0 136816 0 1 113021
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1624857261
transform 1 0 136943 0 1 113579
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1624857261
transform 1 0 136943 0 1 113243
box 0 0 1 1
use contact_19  contact_19_53
timestamp 1624857261
transform 1 0 136940 0 1 113580
box 0 0 1 1
use contact_19  contact_19_54
timestamp 1624857261
transform 1 0 136940 0 1 113244
box 0 0 1 1
use contact_13  contact_13_53
timestamp 1624857261
transform 1 0 136947 0 1 113571
box 0 0 1 1
use contact_13  contact_13_54
timestamp 1624857261
transform 1 0 136947 0 1 113235
box 0 0 1 1
use contact_33  contact_33_2441
timestamp 1624857261
transform 1 0 136816 0 1 113293
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1624857261
transform 1 0 136943 0 1 113915
box 0 0 1 1
use contact_19  contact_19_52
timestamp 1624857261
transform 1 0 136940 0 1 113916
box 0 0 1 1
use contact_13  contact_13_52
timestamp 1624857261
transform 1 0 136947 0 1 113907
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1624857261
transform 1 0 136943 0 1 114251
box 0 0 1 1
use contact_19  contact_19_51
timestamp 1624857261
transform 1 0 136940 0 1 114252
box 0 0 1 1
use contact_13  contact_13_51
timestamp 1624857261
transform 1 0 136947 0 1 114243
box 0 0 1 1
use contact_33  contact_33_2393
timestamp 1624857261
transform 1 0 137496 0 1 112885
box 0 0 1 1
use contact_33  contact_33_5
timestamp 1624857261
transform 1 0 135320 0 1 114653
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1624857261
transform 1 0 136939 0 1 114583
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1624857261
transform 1 0 136943 0 1 114587
box 0 0 1 1
use contact_19  contact_19_50
timestamp 1624857261
transform 1 0 136940 0 1 114588
box 0 0 1 1
use contact_13  contact_13_50
timestamp 1624857261
transform 1 0 136947 0 1 114579
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1624857261
transform 1 0 136943 0 1 115259
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1624857261
transform 1 0 136943 0 1 114923
box 0 0 1 1
use contact_19  contact_19_48
timestamp 1624857261
transform 1 0 136940 0 1 115260
box 0 0 1 1
use contact_19  contact_19_49
timestamp 1624857261
transform 1 0 136940 0 1 114924
box 0 0 1 1
use contact_13  contact_13_48
timestamp 1624857261
transform 1 0 136947 0 1 115251
box 0 0 1 1
use contact_13  contact_13_49
timestamp 1624857261
transform 1 0 136947 0 1 114915
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1624857261
transform 1 0 136943 0 1 115595
box 0 0 1 1
use contact_19  contact_19_47
timestamp 1624857261
transform 1 0 136940 0 1 115596
box 0 0 1 1
use contact_13  contact_13_47
timestamp 1624857261
transform 1 0 136947 0 1 115587
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1624857261
transform 1 0 136939 0 1 116263
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1624857261
transform 1 0 136943 0 1 116267
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1624857261
transform 1 0 136943 0 1 115931
box 0 0 1 1
use contact_19  contact_19_45
timestamp 1624857261
transform 1 0 136940 0 1 116268
box 0 0 1 1
use contact_19  contact_19_46
timestamp 1624857261
transform 1 0 136940 0 1 115932
box 0 0 1 1
use contact_13  contact_13_45
timestamp 1624857261
transform 1 0 136947 0 1 116259
box 0 0 1 1
use contact_13  contact_13_46
timestamp 1624857261
transform 1 0 136947 0 1 115923
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1624857261
transform 1 0 136943 0 1 116603
box 0 0 1 1
use contact_19  contact_19_44
timestamp 1624857261
transform 1 0 136940 0 1 116604
box 0 0 1 1
use contact_13  contact_13_44
timestamp 1624857261
transform 1 0 136947 0 1 116595
box 0 0 1 1
use contact_33  contact_33_2386
timestamp 1624857261
transform 1 0 137496 0 1 114517
box 0 0 1 1
use contact_33  contact_33_2369
timestamp 1624857261
transform 1 0 137496 0 1 116149
box 0 0 1 1
use contact_33  contact_33_2
timestamp 1624857261
transform 1 0 138176 0 1 114789
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1624857261
transform 1 0 136943 0 1 117275
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1624857261
transform 1 0 136943 0 1 116939
box 0 0 1 1
use contact_19  contact_19_42
timestamp 1624857261
transform 1 0 136940 0 1 117276
box 0 0 1 1
use contact_19  contact_19_43
timestamp 1624857261
transform 1 0 136940 0 1 116940
box 0 0 1 1
use contact_13  contact_13_42
timestamp 1624857261
transform 1 0 136947 0 1 117267
box 0 0 1 1
use contact_13  contact_13_43
timestamp 1624857261
transform 1 0 136947 0 1 116931
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1624857261
transform 1 0 136943 0 1 117611
box 0 0 1 1
use contact_19  contact_19_41
timestamp 1624857261
transform 1 0 136940 0 1 117612
box 0 0 1 1
use contact_13  contact_13_41
timestamp 1624857261
transform 1 0 136947 0 1 117603
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1624857261
transform 1 0 136939 0 1 117943
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1624857261
transform 1 0 136943 0 1 118283
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1624857261
transform 1 0 136943 0 1 117947
box 0 0 1 1
use contact_19  contact_19_39
timestamp 1624857261
transform 1 0 136940 0 1 118284
box 0 0 1 1
use contact_19  contact_19_40
timestamp 1624857261
transform 1 0 136940 0 1 117948
box 0 0 1 1
use contact_13  contact_13_39
timestamp 1624857261
transform 1 0 136947 0 1 118275
box 0 0 1 1
use contact_13  contact_13_40
timestamp 1624857261
transform 1 0 136947 0 1 117939
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1624857261
transform 1 0 136943 0 1 118619
box 0 0 1 1
use contact_19  contact_19_38
timestamp 1624857261
transform 1 0 136940 0 1 118620
box 0 0 1 1
use contact_13  contact_13_38
timestamp 1624857261
transform 1 0 136947 0 1 118611
box 0 0 1 1
use contact_33  contact_33_2437
timestamp 1624857261
transform 1 0 136816 0 1 119141
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1624857261
transform 1 0 136943 0 1 119291
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1624857261
transform 1 0 136943 0 1 118955
box 0 0 1 1
use contact_19  contact_19_36
timestamp 1624857261
transform 1 0 136940 0 1 119292
box 0 0 1 1
use contact_19  contact_19_37
timestamp 1624857261
transform 1 0 136940 0 1 118956
box 0 0 1 1
use contact_13  contact_13_36
timestamp 1624857261
transform 1 0 136947 0 1 119283
box 0 0 1 1
use contact_13  contact_13_37
timestamp 1624857261
transform 1 0 136947 0 1 118947
box 0 0 1 1
use contact_33  contact_33_2372
timestamp 1624857261
transform 1 0 137496 0 1 118053
box 0 0 1 1
use contact_33  contact_33_2436
timestamp 1624857261
transform 1 0 136816 0 1 119549
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1624857261
transform 1 0 136939 0 1 119623
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1624857261
transform 1 0 136943 0 1 119627
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1624857261
transform 1 0 136940 0 1 119628
box 0 0 1 1
use contact_13  contact_13_35
timestamp 1624857261
transform 1 0 136947 0 1 119619
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1624857261
transform 1 0 136943 0 1 120299
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1624857261
transform 1 0 136943 0 1 119963
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1624857261
transform 1 0 136940 0 1 120300
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1624857261
transform 1 0 136940 0 1 119964
box 0 0 1 1
use contact_13  contact_13_33
timestamp 1624857261
transform 1 0 136947 0 1 120291
box 0 0 1 1
use contact_13  contact_13_34
timestamp 1624857261
transform 1 0 136947 0 1 119955
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1624857261
transform 1 0 136943 0 1 120635
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1624857261
transform 1 0 136940 0 1 120636
box 0 0 1 1
use contact_13  contact_13_32
timestamp 1624857261
transform 1 0 136947 0 1 120627
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1624857261
transform 1 0 136939 0 1 121303
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1624857261
transform 1 0 136943 0 1 121307
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1624857261
transform 1 0 136943 0 1 120971
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1624857261
transform 1 0 136940 0 1 121308
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1624857261
transform 1 0 136940 0 1 120972
box 0 0 1 1
use contact_13  contact_13_30
timestamp 1624857261
transform 1 0 136947 0 1 121299
box 0 0 1 1
use contact_13  contact_13_31
timestamp 1624857261
transform 1 0 136947 0 1 120963
box 0 0 1 1
use contact_33  contact_33_2438
timestamp 1624857261
transform 1 0 136816 0 1 121453
box 0 0 1 1
use contact_33  contact_33_2439
timestamp 1624857261
transform 1 0 136816 0 1 121725
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1624857261
transform 1 0 136943 0 1 121643
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1624857261
transform 1 0 136940 0 1 121644
box 0 0 1 1
use contact_13  contact_13_29
timestamp 1624857261
transform 1 0 136947 0 1 121635
box 0 0 1 1
use contact_33  contact_33_2419
timestamp 1624857261
transform 1 0 137496 0 1 121453
box 0 0 1 1
use contact_33  contact_33_2396
timestamp 1624857261
transform 1 0 137496 0 1 119685
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1624857261
transform 1 0 136943 0 1 122315
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1624857261
transform 1 0 136943 0 1 121979
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1624857261
transform 1 0 136940 0 1 122316
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1624857261
transform 1 0 136940 0 1 121980
box 0 0 1 1
use contact_13  contact_13_27
timestamp 1624857261
transform 1 0 136947 0 1 122307
box 0 0 1 1
use contact_13  contact_13_28
timestamp 1624857261
transform 1 0 136947 0 1 121971
box 0 0 1 1
use contact_33  contact_33_5492
timestamp 1624857261
transform 1 0 136187 0 1 122853
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1624857261
transform 1 0 136943 0 1 122651
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1624857261
transform 1 0 136940 0 1 122652
box 0 0 1 1
use contact_13  contact_13_26
timestamp 1624857261
transform 1 0 136947 0 1 122643
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1624857261
transform 1 0 136939 0 1 122983
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1624857261
transform 1 0 136943 0 1 123323
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1624857261
transform 1 0 136943 0 1 122987
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1624857261
transform 1 0 136940 0 1 123324
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1624857261
transform 1 0 136940 0 1 122988
box 0 0 1 1
use contact_13  contact_13_24
timestamp 1624857261
transform 1 0 136947 0 1 123315
box 0 0 1 1
use contact_13  contact_13_25
timestamp 1624857261
transform 1 0 136947 0 1 122979
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1624857261
transform 1 0 136943 0 1 123659
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1624857261
transform 1 0 136940 0 1 123660
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1624857261
transform 1 0 136947 0 1 123651
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1624857261
transform 1 0 136943 0 1 124331
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1624857261
transform 1 0 136943 0 1 123995
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1624857261
transform 1 0 136940 0 1 124332
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1624857261
transform 1 0 136940 0 1 123996
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1624857261
transform 1 0 136947 0 1 124323
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1624857261
transform 1 0 136947 0 1 123987
box 0 0 1 1
use contact_33  contact_33_2403
timestamp 1624857261
transform 1 0 137496 0 1 122949
box 0 0 1 1
use contact_33  contact_33_1
timestamp 1624857261
transform 1 0 138176 0 1 123357
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1624857261
transform 1 0 136939 0 1 124663
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1624857261
transform 1 0 136943 0 1 124667
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1624857261
transform 1 0 136940 0 1 124668
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1624857261
transform 1 0 136947 0 1 124659
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1624857261
transform 1 0 136943 0 1 125339
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1624857261
transform 1 0 136943 0 1 125003
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1624857261
transform 1 0 136940 0 1 125340
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1624857261
transform 1 0 136940 0 1 125004
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1624857261
transform 1 0 136947 0 1 125331
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1624857261
transform 1 0 136947 0 1 124995
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1624857261
transform 1 0 136943 0 1 125675
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1624857261
transform 1 0 136940 0 1 125676
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1624857261
transform 1 0 136947 0 1 125667
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1624857261
transform 1 0 136939 0 1 126343
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1624857261
transform 1 0 136943 0 1 126347
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1624857261
transform 1 0 136943 0 1 126011
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1624857261
transform 1 0 136940 0 1 126348
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1624857261
transform 1 0 136940 0 1 126012
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1624857261
transform 1 0 136947 0 1 126339
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1624857261
transform 1 0 136947 0 1 126003
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1624857261
transform 1 0 136943 0 1 126683
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1624857261
transform 1 0 136940 0 1 126684
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1624857261
transform 1 0 136947 0 1 126675
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1624857261
transform 1 0 136943 0 1 127019
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1624857261
transform 1 0 136940 0 1 127020
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1624857261
transform 1 0 136947 0 1 127011
box 0 0 1 1
use contact_33  contact_33_2417
timestamp 1624857261
transform 1 0 137496 0 1 124717
box 0 0 1 1
use contact_33  contact_33_2406
timestamp 1624857261
transform 1 0 137496 0 1 126485
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1624857261
transform 1 0 136943 0 1 127355
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1624857261
transform 1 0 136940 0 1 127356
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1624857261
transform 1 0 136947 0 1 127347
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1624857261
transform 1 0 136939 0 1 128023
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1624857261
transform 1 0 136943 0 1 128027
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1624857261
transform 1 0 136943 0 1 127691
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1624857261
transform 1 0 136940 0 1 128028
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1624857261
transform 1 0 136940 0 1 127692
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1624857261
transform 1 0 136947 0 1 128019
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1624857261
transform 1 0 136947 0 1 127683
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1624857261
transform 1 0 136943 0 1 128363
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1624857261
transform 1 0 136940 0 1 128364
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1624857261
transform 1 0 136947 0 1 128355
box 0 0 1 1
use contact_33  contact_33_2434
timestamp 1624857261
transform 1 0 136816 0 1 128117
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1624857261
transform 1 0 136943 0 1 129035
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1624857261
transform 1 0 136943 0 1 128699
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1624857261
transform 1 0 136940 0 1 129036
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1624857261
transform 1 0 136940 0 1 128700
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1624857261
transform 1 0 136947 0 1 129027
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1624857261
transform 1 0 136947 0 1 128691
box 0 0 1 1
use contact_33  contact_33_2435
timestamp 1624857261
transform 1 0 136816 0 1 128797
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1624857261
transform 1 0 136943 0 1 129371
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1624857261
transform 1 0 136940 0 1 129372
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1624857261
transform 1 0 136947 0 1 129363
box 0 0 1 1
use contact_33  contact_33_2385
timestamp 1624857261
transform 1 0 137496 0 1 128117
box 0 0 1 1
use contact_7  contact_7_361
timestamp 1624857261
transform 1 0 135979 0 1 129763
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1624857261
transform 1 0 136939 0 1 129703
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1624857261
transform 1 0 136943 0 1 129707
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1624857261
transform 1 0 136940 0 1 129708
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1624857261
transform 1 0 136947 0 1 129699
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1624857261
transform 1 0 136943 0 1 130379
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1624857261
transform 1 0 136943 0 1 130043
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1624857261
transform 1 0 136940 0 1 130380
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1624857261
transform 1 0 136940 0 1 130044
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1624857261
transform 1 0 136947 0 1 130371
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1624857261
transform 1 0 136947 0 1 130035
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1624857261
transform 1 0 136943 0 1 130715
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1624857261
transform 1 0 136940 0 1 130716
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1624857261
transform 1 0 136947 0 1 130707
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1624857261
transform 1 0 136943 0 1 131051
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1624857261
transform 1 0 136940 0 1 131052
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1624857261
transform 1 0 136947 0 1 131043
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1624857261
transform 1 0 136939 0 1 131383
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1624857261
transform 1 0 136943 0 1 131387
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1624857261
transform 1 0 136940 0 1 131388
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1624857261
transform 1 0 136947 0 1 131379
box 0 0 1 1
use contact_33  contact_33_2430
timestamp 1624857261
transform 1 0 136816 0 1 131517
box 0 0 1 1
use contact_14  contact_14_776
timestamp 1624857261
transform 1 0 135189 0 1 132000
box 0 0 1 1
use contact_13  contact_13_776
timestamp 1624857261
transform 1 0 135193 0 1 131992
box 0 0 1 1
use contact_14  contact_14_775
timestamp 1624857261
transform 1 0 135525 0 1 132000
box 0 0 1 1
use contact_13  contact_13_775
timestamp 1624857261
transform 1 0 135529 0 1 131992
box 0 0 1 1
use contact_14  contact_14_774
timestamp 1624857261
transform 1 0 135861 0 1 132000
box 0 0 1 1
use contact_13  contact_13_774
timestamp 1624857261
transform 1 0 135865 0 1 131992
box 0 0 1 1
use contact_7  contact_7_156
timestamp 1624857261
transform 1 0 136529 0 1 131996
box 0 0 1 1
use contact_14  contact_14_772
timestamp 1624857261
transform 1 0 136533 0 1 132000
box 0 0 1 1
use contact_14  contact_14_773
timestamp 1624857261
transform 1 0 136197 0 1 132000
box 0 0 1 1
use contact_19  contact_19_772
timestamp 1624857261
transform 1 0 136530 0 1 132001
box 0 0 1 1
use contact_13  contact_13_772
timestamp 1624857261
transform 1 0 136537 0 1 131992
box 0 0 1 1
use contact_13  contact_13_773
timestamp 1624857261
transform 1 0 136201 0 1 131992
box 0 0 1 1
use contact_38  contact_38_1
timestamp 1624857261
transform 1 0 136876 0 1 131937
box 0 0 192 192
use contact_33  contact_33_2431
timestamp 1624857261
transform 1 0 136816 0 1 131925
box 0 0 1 1
use contact_33  contact_33_2429
timestamp 1624857261
transform 1 0 136408 0 1 132061
box 0 0 1 1
use contact_33  contact_33_2352
timestamp 1624857261
transform 1 0 137496 0 1 129749
box 0 0 1 1
use contact_33  contact_33_0
timestamp 1624857261
transform 1 0 138176 0 1 130429
box 0 0 1 1
use contact_33  contact_33_2428
timestamp 1624857261
transform 1 0 136408 0 1 132469
box 0 0 1 1
use contact_39  contact_39_36
timestamp 1624857261
transform 1 0 137632 0 1 132605
box 0 0 192 192
use contact_39  contact_39_37
timestamp 1624857261
transform 1 0 137632 0 1 132469
box 0 0 192 192
use contact_39  contact_39_56
timestamp 1624857261
transform 1 0 137496 0 1 132469
box 0 0 192 192
use contact_39  contact_39_58
timestamp 1624857261
transform 1 0 137496 0 1 132605
box 0 0 192 192
use contact_39  contact_39_62
timestamp 1624857261
transform 1 0 137768 0 1 132605
box 0 0 192 192
use contact_39  contact_39_69
timestamp 1624857261
transform 1 0 137768 0 1 132469
box 0 0 192 192
use contact_39  contact_39_39
timestamp 1624857261
transform 1 0 137496 0 1 132741
box 0 0 192 192
use contact_39  contact_39_45
timestamp 1624857261
transform 1 0 137768 0 1 132741
box 0 0 192 192
use contact_39  contact_39_51
timestamp 1624857261
transform 1 0 137632 0 1 132741
box 0 0 192 192
use contact_39  contact_39_0
timestamp 1624857261
transform 1 0 138312 0 1 133285
box 0 0 192 192
use contact_39  contact_39_7
timestamp 1624857261
transform 1 0 138448 0 1 133149
box 0 0 192 192
use contact_39  contact_39_16
timestamp 1624857261
transform 1 0 138176 0 1 133149
box 0 0 192 192
use contact_39  contact_39_17
timestamp 1624857261
transform 1 0 138312 0 1 133149
box 0 0 192 192
use contact_39  contact_39_20
timestamp 1624857261
transform 1 0 138448 0 1 133285
box 0 0 192 192
use contact_39  contact_39_34
timestamp 1624857261
transform 1 0 138176 0 1 133285
box 0 0 192 192
use contact_39  contact_39_11
timestamp 1624857261
transform 1 0 138176 0 1 133421
box 0 0 192 192
use contact_39  contact_39_22
timestamp 1624857261
transform 1 0 138312 0 1 133421
box 0 0 192 192
use contact_39  contact_39_32
timestamp 1624857261
transform 1 0 138448 0 1 133421
box 0 0 192 192
<< labels >>
rlabel metal3 s 0 8024 212 8100 4 csb0
port 53 nsew default input
rlabel metal3 s 0 9792 212 9868 4 web0
port 55 nsew default input
rlabel metal3 s 0 8296 212 8372 4 clk0
port 56 nsew default input
rlabel metal4 s 23664 0 23740 212 4 din0[0]
port 1 nsew default input
rlabel metal4 s 24752 0 24828 212 4 din0[1]
port 2 nsew default input
rlabel metal4 s 25976 0 26052 212 4 din0[2]
port 3 nsew default input
rlabel metal4 s 27064 0 27140 212 4 din0[3]
port 4 nsew default input
rlabel metal4 s 28152 0 28228 212 4 din0[4]
port 5 nsew default input
rlabel metal4 s 29240 0 29316 212 4 din0[5]
port 6 nsew default input
rlabel metal4 s 30600 0 30676 212 4 din0[6]
port 7 nsew default input
rlabel metal4 s 31824 0 31900 212 4 din0[7]
port 8 nsew default input
rlabel metal4 s 32912 0 32988 212 4 din0[8]
port 9 nsew default input
rlabel metal4 s 34000 0 34076 212 4 din0[9]
port 10 nsew default input
rlabel metal4 s 35088 0 35164 212 4 din0[10]
port 11 nsew default input
rlabel metal4 s 36448 0 36524 212 4 din0[11]
port 12 nsew default input
rlabel metal4 s 37536 0 37612 212 4 din0[12]
port 13 nsew default input
rlabel metal4 s 38624 0 38700 212 4 din0[13]
port 14 nsew default input
rlabel metal4 s 39984 0 40060 212 4 din0[14]
port 15 nsew default input
rlabel metal4 s 41208 0 41284 212 4 din0[15]
port 16 nsew default input
rlabel metal4 s 42296 0 42372 212 4 din0[16]
port 17 nsew default input
rlabel metal4 s 43384 0 43460 212 4 din0[17]
port 18 nsew default input
rlabel metal4 s 44472 0 44548 212 4 din0[18]
port 19 nsew default input
rlabel metal4 s 45832 0 45908 212 4 din0[19]
port 20 nsew default input
rlabel metal4 s 46920 0 46996 212 4 din0[20]
port 21 nsew default input
rlabel metal4 s 48144 0 48220 212 4 din0[21]
port 22 nsew default input
rlabel metal4 s 49232 0 49308 212 4 din0[22]
port 23 nsew default input
rlabel metal4 s 50320 0 50396 212 4 din0[23]
port 24 nsew default input
rlabel metal4 s 51680 0 51756 212 4 din0[24]
port 25 nsew default input
rlabel metal4 s 52768 0 52844 212 4 din0[25]
port 26 nsew default input
rlabel metal4 s 53856 0 53932 212 4 din0[26]
port 27 nsew default input
rlabel metal4 s 54944 0 55020 212 4 din0[27]
port 28 nsew default input
rlabel metal4 s 56304 0 56380 212 4 din0[28]
port 29 nsew default input
rlabel metal4 s 57528 0 57604 212 4 din0[29]
port 30 nsew default input
rlabel metal4 s 58616 0 58692 212 4 din0[30]
port 31 nsew default input
rlabel metal4 s 59704 0 59780 212 4 din0[31]
port 32 nsew default input
rlabel metal4 s 28968 0 29044 212 4 dout0[0]
port 62 nsew default output
rlabel metal4 s 31960 0 32036 212 4 dout0[1]
port 63 nsew default output
rlabel metal4 s 34408 0 34484 212 4 dout0[2]
port 64 nsew default output
rlabel metal4 s 36992 0 37068 212 4 dout0[3]
port 65 nsew default output
rlabel metal4 s 39440 0 39516 212 4 dout0[4]
port 66 nsew default output
rlabel metal4 s 41752 0 41828 212 4 dout0[5]
port 67 nsew default output
rlabel metal4 s 44200 0 44276 212 4 dout0[6]
port 68 nsew default output
rlabel metal4 s 46512 0 46588 212 4 dout0[7]
port 69 nsew default output
rlabel metal4 s 49912 0 49988 212 4 dout0[8]
port 70 nsew default output
rlabel metal4 s 51952 0 52028 212 4 dout0[9]
port 71 nsew default output
rlabel metal4 s 54536 0 54612 212 4 dout0[10]
port 72 nsew default output
rlabel metal4 s 56984 0 57060 212 4 dout0[11]
port 73 nsew default output
rlabel metal4 s 59296 0 59372 212 4 dout0[12]
port 74 nsew default output
rlabel metal4 s 61880 0 61956 212 4 dout0[13]
port 75 nsew default output
rlabel metal4 s 64464 0 64540 212 4 dout0[14]
port 76 nsew default output
rlabel metal4 s 66912 0 66988 212 4 dout0[15]
port 77 nsew default output
rlabel metal4 s 69496 0 69572 212 4 dout0[16]
port 78 nsew default output
rlabel metal4 s 71944 0 72020 212 4 dout0[17]
port 79 nsew default output
rlabel metal4 s 74392 0 74468 212 4 dout0[18]
port 80 nsew default output
rlabel metal4 s 76840 0 76916 212 4 dout0[19]
port 81 nsew default output
rlabel metal4 s 79424 0 79500 212 4 dout0[20]
port 82 nsew default output
rlabel metal4 s 81872 0 81948 212 4 dout0[21]
port 83 nsew default output
rlabel metal4 s 84320 0 84396 212 4 dout0[22]
port 84 nsew default output
rlabel metal4 s 86904 0 86980 212 4 dout0[23]
port 85 nsew default output
rlabel metal4 s 89080 0 89156 212 4 dout0[24]
port 86 nsew default output
rlabel metal4 s 91936 0 92012 212 4 dout0[25]
port 87 nsew default output
rlabel metal4 s 94384 0 94460 212 4 dout0[26]
port 88 nsew default output
rlabel metal4 s 96832 0 96908 212 4 dout0[27]
port 89 nsew default output
rlabel metal4 s 99416 0 99492 212 4 dout0[28]
port 90 nsew default output
rlabel metal4 s 101864 0 101940 212 4 dout0[29]
port 91 nsew default output
rlabel metal4 s 104312 0 104388 212 4 dout0[30]
port 92 nsew default output
rlabel metal4 s 106896 0 106972 212 4 dout0[31]
port 93 nsew default output
rlabel metal4 s 16592 0 16668 212 4 addr0[0]
port 33 nsew default input
rlabel metal4 s 17680 0 17756 212 4 addr0[1]
port 34 nsew default input
rlabel metal3 s 0 29784 212 29860 4 addr0[2]
port 35 nsew default input
rlabel metal3 s 0 31416 212 31492 4 addr0[3]
port 36 nsew default input
rlabel metal3 s 0 32776 212 32852 4 addr0[4]
port 37 nsew default input
rlabel metal3 s 0 34272 212 34348 4 addr0[5]
port 38 nsew default input
rlabel metal3 s 0 35360 212 35436 4 addr0[6]
port 39 nsew default input
rlabel metal3 s 0 37128 212 37204 4 addr0[7]
port 40 nsew default input
rlabel metal3 s 0 38216 212 38292 4 addr0[8]
port 41 nsew default input
rlabel metal3 s 0 40120 212 40196 4 addr0[9]
port 42 nsew default input
rlabel metal4 s 18768 0 18844 212 4 wmask0[0]
port 58 nsew default input
rlabel metal4 s 20128 0 20204 212 4 wmask0[1]
port 59 nsew default input
rlabel metal4 s 21080 0 21156 212 4 wmask0[2]
port 60 nsew default input
rlabel metal4 s 22304 0 22380 212 4 wmask0[3]
port 61 nsew default input
rlabel metal3 s 138584 129880 138796 129956 4 csb1
port 54 nsew default input
rlabel metal4 s 132736 133552 132812 133764 4 clk1
port 57 nsew default input
rlabel metal4 s 29648 133552 29724 133764 4 dout1[0]
port 94 nsew default output
rlabel metal4 s 31960 133552 32036 133764 4 dout1[1]
port 95 nsew default output
rlabel metal4 s 34544 133552 34620 133764 4 dout1[2]
port 96 nsew default output
rlabel metal4 s 36992 133552 37068 133764 4 dout1[3]
port 97 nsew default output
rlabel metal4 s 39576 133552 39652 133764 4 dout1[4]
port 98 nsew default output
rlabel metal4 s 42024 133552 42100 133764 4 dout1[5]
port 99 nsew default output
rlabel metal4 s 44608 133552 44684 133764 4 dout1[6]
port 100 nsew default output
rlabel metal4 s 47056 133552 47132 133764 4 dout1[7]
port 101 nsew default output
rlabel metal4 s 49504 133552 49580 133764 4 dout1[8]
port 102 nsew default output
rlabel metal4 s 51952 133552 52028 133764 4 dout1[9]
port 103 nsew default output
rlabel metal4 s 54400 133552 54476 133764 4 dout1[10]
port 104 nsew default output
rlabel metal4 s 56984 133552 57060 133764 4 dout1[11]
port 105 nsew default output
rlabel metal4 s 59568 133552 59644 133764 4 dout1[12]
port 106 nsew default output
rlabel metal4 s 62016 133552 62092 133764 4 dout1[13]
port 107 nsew default output
rlabel metal4 s 64600 133552 64676 133764 4 dout1[14]
port 108 nsew default output
rlabel metal4 s 67048 133552 67124 133764 4 dout1[15]
port 109 nsew default output
rlabel metal4 s 69360 133552 69436 133764 4 dout1[16]
port 110 nsew default output
rlabel metal4 s 72080 133552 72156 133764 4 dout1[17]
port 111 nsew default output
rlabel metal4 s 74392 133552 74468 133764 4 dout1[18]
port 112 nsew default output
rlabel metal4 s 76976 133552 77052 133764 4 dout1[19]
port 113 nsew default output
rlabel metal4 s 79424 133552 79500 133764 4 dout1[20]
port 114 nsew default output
rlabel metal4 s 82008 133552 82084 133764 4 dout1[21]
port 115 nsew default output
rlabel metal4 s 84456 133552 84532 133764 4 dout1[22]
port 116 nsew default output
rlabel metal4 s 87040 133552 87116 133764 4 dout1[23]
port 117 nsew default output
rlabel metal4 s 89488 133552 89564 133764 4 dout1[24]
port 118 nsew default output
rlabel metal4 s 91936 133552 92012 133764 4 dout1[25]
port 119 nsew default output
rlabel metal4 s 94384 133552 94460 133764 4 dout1[26]
port 120 nsew default output
rlabel metal4 s 96832 133552 96908 133764 4 dout1[27]
port 121 nsew default output
rlabel metal4 s 99416 133552 99492 133764 4 dout1[28]
port 122 nsew default output
rlabel metal4 s 102000 133552 102076 133764 4 dout1[29]
port 123 nsew default output
rlabel metal4 s 104448 133552 104524 133764 4 dout1[30]
port 124 nsew default output
rlabel metal4 s 107032 133552 107108 133764 4 dout1[31]
port 125 nsew default output
rlabel metal4 s 121176 133552 121252 133764 4 addr1[0]
port 43 nsew default input
rlabel metal4 s 119952 133552 120028 133764 4 addr1[1]
port 44 nsew default input
rlabel metal3 s 138584 19312 138796 19388 4 addr1[2]
port 45 nsew default input
rlabel metal3 s 138584 17408 138796 17484 4 addr1[3]
port 46 nsew default input
rlabel metal3 s 138584 16456 138796 16532 4 addr1[4]
port 47 nsew default input
rlabel metal3 s 138584 14688 138796 14764 4 addr1[5]
port 48 nsew default input
rlabel metal4 s 124848 0 124924 212 4 addr1[6]
port 49 nsew default input
rlabel metal4 s 124440 0 124516 212 4 addr1[7]
port 50 nsew default input
rlabel metal4 s 124576 0 124652 212 4 addr1[8]
port 51 nsew default input
rlabel metal4 s 124712 0 124788 212 4 addr1[9]
port 52 nsew default input
rlabel metal4 s 952 952 1300 132812 4 vccd1
port 126 nsew power bidirectional abutment
rlabel metal3 s 952 952 137844 1300 4 vccd1
port 126 nsew power bidirectional abutment
rlabel metal4 s 137496 952 137844 132812 4 vccd1
port 126 nsew power bidirectional abutment
rlabel metal3 s 952 132464 137844 132812 4 vccd1
port 126 nsew power bidirectional abutment
rlabel metal4 s 272 272 620 133492 4 vssd1
port 127 nsew ground bidirectional abutment
rlabel metal3 s 272 133144 138524 133492 4 vssd1
port 127 nsew ground bidirectional abutment
rlabel metal3 s 272 272 138524 620 4 vssd1
port 127 nsew ground bidirectional abutment
rlabel metal4 s 138176 272 138524 133492 4 vssd1
port 127 nsew ground bidirectional abutment
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 138796 133764
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_4kbyte_1rw1r_32x1024_8.gds
string LEFsymmetry X Y R90
string GDS_END 2602142
string GDS_START 134
<< end >>
