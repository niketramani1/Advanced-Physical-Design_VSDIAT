magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1294 19147 16306 34747
<< metal4 >>
tri 979 33194 1272 33487 se
rect 1272 33485 13740 33487
tri 13740 33485 13742 33487 sw
rect 1272 33463 13742 33485
tri 13742 33463 13764 33485 sw
rect 1272 33227 1355 33463
rect 1591 33227 1675 33463
rect 1911 33227 1995 33463
rect 2231 33227 2315 33463
rect 2551 33227 2635 33463
rect 2871 33227 2955 33463
rect 3191 33227 3275 33463
rect 3511 33227 3595 33463
rect 3831 33227 3915 33463
rect 4151 33227 4235 33463
rect 4471 33227 4555 33463
rect 4791 33227 4875 33463
rect 5111 33227 5195 33463
rect 5431 33227 5515 33463
rect 5751 33227 5835 33463
rect 6071 33227 6155 33463
rect 6391 33227 6475 33463
rect 6711 33227 6795 33463
rect 7031 33227 7115 33463
rect 7351 33227 7435 33463
rect 7671 33227 7755 33463
rect 7991 33227 8075 33463
rect 8311 33227 8395 33463
rect 8631 33227 8715 33463
rect 8951 33227 9035 33463
rect 9271 33227 9355 33463
rect 9591 33227 9675 33463
rect 9911 33227 9995 33463
rect 10231 33227 10315 33463
rect 10551 33227 10635 33463
rect 10871 33227 10955 33463
rect 11191 33227 11275 33463
rect 11511 33227 11595 33463
rect 11831 33227 11915 33463
rect 12151 33227 12235 33463
rect 12471 33227 12555 33463
rect 12791 33227 12875 33463
rect 13111 33227 13195 33463
rect 13431 33227 13515 33463
rect 13751 33227 13764 33463
rect 1272 33194 13764 33227
tri 732 32947 979 33194 se
rect 979 32958 992 33194
rect 1228 33140 13764 33194
tri 13764 33140 14087 33463 sw
rect 1228 32958 13838 33140
rect 979 32947 13838 32958
tri 659 32874 732 32947 se
rect 732 32874 1270 32947
tri 506 32721 659 32874 se
rect 659 32721 672 32874
tri 339 32554 506 32721 se
rect 506 32638 672 32721
rect 908 32721 1270 32874
tri 1270 32721 1496 32947 nw
tri 13516 32723 13740 32947 ne
rect 13740 32904 13838 32947
rect 14074 32947 14087 33140
tri 14087 32947 14280 33140 sw
rect 14074 32904 14280 32947
rect 13740 32820 14280 32904
tri 14280 32820 14407 32947 sw
rect 13740 32723 14158 32820
tri 13740 32721 13742 32723 ne
rect 13742 32721 14158 32723
rect 908 32638 1187 32721
tri 1187 32638 1270 32721 nw
rect 506 32554 732 32638
tri -23 32192 339 32554 se
rect 339 32318 352 32554
rect 588 32318 732 32554
rect 339 32192 732 32318
tri -34 32181 -23 32192 se
rect -23 32181 -10 32192
rect -34 31956 -10 32181
rect 226 32183 732 32192
tri 732 32183 1187 32638 nw
tri 13742 32584 13879 32721 ne
rect 13879 32584 14158 32721
rect 14394 32721 14407 32820
tri 14407 32721 14506 32820 sw
rect 14394 32584 14506 32721
tri 13879 32183 14280 32584 ne
rect 14280 32500 14506 32584
tri 14506 32500 14727 32721 sw
rect 14280 32264 14478 32500
rect 14714 32264 14727 32500
rect 14280 32183 14727 32264
rect 226 31956 506 32183
tri 506 31957 732 32183 nw
tri 14280 31957 14506 32183 ne
rect 14506 32181 14727 32183
tri 14727 32181 15046 32500 sw
rect 14506 32178 15046 32181
rect -34 31872 506 31956
rect -34 31636 -10 31872
rect 226 31636 506 31872
rect -34 31552 506 31636
rect -34 31316 -10 31552
rect 226 31316 506 31552
rect -34 31232 506 31316
rect -34 30996 -10 31232
rect 226 30996 506 31232
rect -34 30912 506 30996
rect -34 30676 -10 30912
rect 226 30676 506 30912
rect -34 30592 506 30676
rect -34 30356 -10 30592
rect 226 30356 506 30592
rect -34 30272 506 30356
rect -34 30036 -10 30272
rect 226 30036 506 30272
rect -34 29952 506 30036
rect -34 29716 -10 29952
rect 226 29716 506 29952
rect -34 29632 506 29716
rect -34 29396 -10 29632
rect 226 29396 506 29632
rect -34 29312 506 29396
rect -34 29076 -10 29312
rect 226 29076 506 29312
rect -34 28992 506 29076
rect -34 28756 -10 28992
rect 226 28756 506 28992
rect -34 28672 506 28756
rect -34 28436 -10 28672
rect 226 28436 506 28672
rect -34 28352 506 28436
rect -34 28116 -10 28352
rect 226 28116 506 28352
rect -34 28032 506 28116
rect -34 27796 -10 28032
rect 226 27796 506 28032
rect -34 27712 506 27796
rect -34 27476 -10 27712
rect 226 27476 506 27712
rect -34 27392 506 27476
rect -34 27156 -10 27392
rect 226 27156 506 27392
rect -34 27072 506 27156
rect -34 26836 -10 27072
rect 226 26836 506 27072
rect -34 26752 506 26836
rect -34 26516 -10 26752
rect 226 26516 506 26752
rect -34 26432 506 26516
rect -34 26196 -10 26432
rect 226 26196 506 26432
rect -34 26112 506 26196
rect -34 25876 -10 26112
rect 226 25876 506 26112
rect -34 25792 506 25876
rect -34 25556 -10 25792
rect 226 25556 506 25792
rect -34 25472 506 25556
rect -34 25236 -10 25472
rect 226 25236 506 25472
rect -34 25152 506 25236
rect -34 24916 -10 25152
rect 226 24916 506 25152
rect -34 24832 506 24916
rect -34 24596 -10 24832
rect 226 24596 506 24832
rect -34 24512 506 24596
rect -34 24276 -10 24512
rect 226 24276 506 24512
rect -34 24192 506 24276
rect -34 23956 -10 24192
rect 226 23956 506 24192
rect -34 23872 506 23956
rect -34 23636 -10 23872
rect 226 23636 506 23872
rect -34 23552 506 23636
rect -34 23316 -10 23552
rect 226 23316 506 23552
rect -34 23232 506 23316
rect -34 22996 -10 23232
rect 226 22996 506 23232
rect -34 22912 506 22996
rect -34 22676 -10 22912
rect 226 22676 506 22912
rect -34 22592 506 22676
rect -34 22356 -10 22592
rect 226 22356 506 22592
rect -34 22272 506 22356
rect -34 22036 -10 22272
rect 226 22036 506 22272
rect -34 21952 506 22036
rect -34 21716 -10 21952
rect 226 21716 506 21952
rect 14506 31942 14786 32178
rect 15022 31942 15046 32178
rect 14506 31858 15046 31942
rect 14506 31622 14786 31858
rect 15022 31622 15046 31858
rect 14506 31538 15046 31622
rect 14506 31302 14786 31538
rect 15022 31302 15046 31538
rect 14506 31218 15046 31302
rect 14506 30982 14786 31218
rect 15022 30982 15046 31218
rect 14506 30898 15046 30982
rect 14506 30662 14786 30898
rect 15022 30662 15046 30898
rect 14506 30578 15046 30662
rect 14506 30342 14786 30578
rect 15022 30342 15046 30578
rect 14506 30258 15046 30342
rect 14506 30022 14786 30258
rect 15022 30022 15046 30258
rect 14506 29938 15046 30022
rect 14506 29702 14786 29938
rect 15022 29702 15046 29938
rect 14506 29618 15046 29702
rect 14506 29382 14786 29618
rect 15022 29382 15046 29618
rect 14506 29298 15046 29382
rect 14506 29062 14786 29298
rect 15022 29062 15046 29298
rect 14506 28978 15046 29062
rect 14506 28742 14786 28978
rect 15022 28742 15046 28978
rect 14506 28658 15046 28742
rect 14506 28422 14786 28658
rect 15022 28422 15046 28658
rect 14506 28338 15046 28422
rect 14506 28102 14786 28338
rect 15022 28102 15046 28338
rect 14506 28018 15046 28102
rect 14506 27782 14786 28018
rect 15022 27782 15046 28018
rect 14506 27698 15046 27782
rect 14506 27462 14786 27698
rect 15022 27462 15046 27698
rect 14506 27378 15046 27462
rect 14506 27142 14786 27378
rect 15022 27142 15046 27378
rect 14506 27058 15046 27142
rect 14506 26822 14786 27058
rect 15022 26822 15046 27058
rect 14506 26738 15046 26822
rect 14506 26502 14786 26738
rect 15022 26502 15046 26738
rect 14506 26418 15046 26502
rect 14506 26182 14786 26418
rect 15022 26182 15046 26418
rect 14506 26098 15046 26182
rect 14506 25862 14786 26098
rect 15022 25862 15046 26098
rect 14506 25778 15046 25862
rect 14506 25542 14786 25778
rect 15022 25542 15046 25778
rect 14506 25458 15046 25542
rect 14506 25222 14786 25458
rect 15022 25222 15046 25458
rect 14506 25138 15046 25222
rect 14506 24902 14786 25138
rect 15022 24902 15046 25138
rect 14506 24818 15046 24902
rect 14506 24582 14786 24818
rect 15022 24582 15046 24818
rect 14506 24498 15046 24582
rect 14506 24262 14786 24498
rect 15022 24262 15046 24498
rect 14506 24178 15046 24262
rect 14506 23942 14786 24178
rect 15022 23942 15046 24178
rect 14506 23858 15046 23942
rect 14506 23622 14786 23858
rect 15022 23622 15046 23858
rect 14506 23538 15046 23622
rect 14506 23302 14786 23538
rect 15022 23302 15046 23538
rect 14506 23218 15046 23302
rect 14506 22982 14786 23218
rect 15022 22982 15046 23218
rect 14506 22898 15046 22982
rect 14506 22662 14786 22898
rect 15022 22662 15046 22898
rect 14506 22578 15046 22662
rect 14506 22342 14786 22578
rect 15022 22342 15046 22578
rect 14506 22258 15046 22342
rect 14506 22022 14786 22258
rect 15022 22022 15046 22258
rect 14506 21938 15046 22022
rect -34 21713 506 21716
tri -34 21630 49 21713 ne
rect 49 21630 506 21713
tri 506 21630 813 21937 sw
tri 14280 21711 14506 21937 se
rect 14506 21711 14786 21938
tri 49 21394 285 21630 ne
rect 285 21394 298 21630
rect 534 21394 813 21630
tri 285 21173 506 21394 ne
rect 506 21310 813 21394
tri 813 21310 1133 21630 sw
rect 506 21173 618 21310
tri 506 21074 605 21173 ne
rect 605 21074 618 21173
rect 854 21173 1133 21310
tri 1133 21173 1270 21310 sw
tri 13825 21256 14280 21711 se
rect 14280 21702 14786 21711
rect 15022 21713 15046 21938
rect 15022 21702 15035 21713
tri 15035 21702 15046 21713 nw
rect 14280 21576 14909 21702
tri 14909 21576 15035 21702 nw
rect 14280 21340 14424 21576
rect 14660 21340 14673 21576
tri 14673 21340 14909 21576 nw
rect 14280 21256 14506 21340
tri 13742 21173 13825 21256 se
rect 13825 21173 14104 21256
rect 854 21074 1270 21173
tri 605 20947 732 21074 ne
rect 732 20990 1270 21074
rect 732 20947 938 20990
tri 732 20754 925 20947 ne
rect 925 20754 938 20947
rect 1174 20947 1270 20990
tri 1270 20947 1496 21173 sw
tri 13740 21171 13742 21173 se
rect 13742 21171 14104 21173
tri 13516 20947 13740 21171 se
rect 13740 21020 14104 21171
rect 14340 21173 14506 21256
tri 14506 21173 14673 21340 nw
rect 14340 21020 14353 21173
tri 14353 21020 14506 21173 nw
rect 13740 20947 14280 21020
tri 14280 20947 14353 21020 nw
rect 1174 20936 14269 20947
tri 14269 20936 14280 20947 nw
rect 1174 20754 13784 20936
tri 925 20667 1012 20754 ne
rect 1012 20700 13784 20754
rect 14020 20700 14033 20936
tri 14033 20700 14269 20936 nw
rect 1012 20667 13740 20700
tri 1012 20431 1248 20667 ne
rect 1248 20431 1261 20667
rect 1497 20431 1581 20667
rect 1817 20431 1901 20667
rect 2137 20431 2221 20667
rect 2457 20431 2541 20667
rect 2777 20431 2861 20667
rect 3097 20431 3181 20667
rect 3417 20431 3501 20667
rect 3737 20431 3821 20667
rect 4057 20431 4141 20667
rect 4377 20431 4461 20667
rect 4697 20431 4781 20667
rect 5017 20431 5101 20667
rect 5337 20431 5421 20667
rect 5657 20431 5741 20667
rect 5977 20431 6061 20667
rect 6297 20431 6381 20667
rect 6617 20431 6701 20667
rect 6937 20431 7021 20667
rect 7257 20431 7341 20667
rect 7577 20431 7661 20667
rect 7897 20431 7981 20667
rect 8217 20431 8301 20667
rect 8537 20431 8621 20667
rect 8857 20431 8941 20667
rect 9177 20431 9261 20667
rect 9497 20431 9581 20667
rect 9817 20431 9901 20667
rect 10137 20431 10221 20667
rect 10457 20431 10541 20667
rect 10777 20431 10861 20667
rect 11097 20431 11181 20667
rect 11417 20431 11501 20667
rect 11737 20431 11821 20667
rect 12057 20431 12141 20667
rect 12377 20431 12461 20667
rect 12697 20431 12781 20667
rect 13017 20431 13101 20667
rect 13337 20431 13421 20667
rect 13657 20431 13740 20667
tri 1248 20409 1270 20431 ne
rect 1270 20409 13740 20431
tri 1270 20407 1272 20409 ne
rect 1272 20407 13740 20409
tri 13740 20407 14033 20700 nw
<< via4 >>
rect 1355 33227 1591 33463
rect 1675 33227 1911 33463
rect 1995 33227 2231 33463
rect 2315 33227 2551 33463
rect 2635 33227 2871 33463
rect 2955 33227 3191 33463
rect 3275 33227 3511 33463
rect 3595 33227 3831 33463
rect 3915 33227 4151 33463
rect 4235 33227 4471 33463
rect 4555 33227 4791 33463
rect 4875 33227 5111 33463
rect 5195 33227 5431 33463
rect 5515 33227 5751 33463
rect 5835 33227 6071 33463
rect 6155 33227 6391 33463
rect 6475 33227 6711 33463
rect 6795 33227 7031 33463
rect 7115 33227 7351 33463
rect 7435 33227 7671 33463
rect 7755 33227 7991 33463
rect 8075 33227 8311 33463
rect 8395 33227 8631 33463
rect 8715 33227 8951 33463
rect 9035 33227 9271 33463
rect 9355 33227 9591 33463
rect 9675 33227 9911 33463
rect 9995 33227 10231 33463
rect 10315 33227 10551 33463
rect 10635 33227 10871 33463
rect 10955 33227 11191 33463
rect 11275 33227 11511 33463
rect 11595 33227 11831 33463
rect 11915 33227 12151 33463
rect 12235 33227 12471 33463
rect 12555 33227 12791 33463
rect 12875 33227 13111 33463
rect 13195 33227 13431 33463
rect 13515 33227 13751 33463
rect 992 32958 1228 33194
rect 672 32638 908 32874
rect 13838 32904 14074 33140
rect 352 32318 588 32554
rect -10 31956 226 32192
rect 14158 32584 14394 32820
rect 14478 32264 14714 32500
rect -10 31636 226 31872
rect -10 31316 226 31552
rect -10 30996 226 31232
rect -10 30676 226 30912
rect -10 30356 226 30592
rect -10 30036 226 30272
rect -10 29716 226 29952
rect -10 29396 226 29632
rect -10 29076 226 29312
rect -10 28756 226 28992
rect -10 28436 226 28672
rect -10 28116 226 28352
rect -10 27796 226 28032
rect -10 27476 226 27712
rect -10 27156 226 27392
rect -10 26836 226 27072
rect -10 26516 226 26752
rect -10 26196 226 26432
rect -10 25876 226 26112
rect -10 25556 226 25792
rect -10 25236 226 25472
rect -10 24916 226 25152
rect -10 24596 226 24832
rect -10 24276 226 24512
rect -10 23956 226 24192
rect -10 23636 226 23872
rect -10 23316 226 23552
rect -10 22996 226 23232
rect -10 22676 226 22912
rect -10 22356 226 22592
rect -10 22036 226 22272
rect -10 21716 226 21952
rect 14786 31942 15022 32178
rect 14786 31622 15022 31858
rect 14786 31302 15022 31538
rect 14786 30982 15022 31218
rect 14786 30662 15022 30898
rect 14786 30342 15022 30578
rect 14786 30022 15022 30258
rect 14786 29702 15022 29938
rect 14786 29382 15022 29618
rect 14786 29062 15022 29298
rect 14786 28742 15022 28978
rect 14786 28422 15022 28658
rect 14786 28102 15022 28338
rect 14786 27782 15022 28018
rect 14786 27462 15022 27698
rect 14786 27142 15022 27378
rect 14786 26822 15022 27058
rect 14786 26502 15022 26738
rect 14786 26182 15022 26418
rect 14786 25862 15022 26098
rect 14786 25542 15022 25778
rect 14786 25222 15022 25458
rect 14786 24902 15022 25138
rect 14786 24582 15022 24818
rect 14786 24262 15022 24498
rect 14786 23942 15022 24178
rect 14786 23622 15022 23858
rect 14786 23302 15022 23538
rect 14786 22982 15022 23218
rect 14786 22662 15022 22898
rect 14786 22342 15022 22578
rect 14786 22022 15022 22258
rect 298 21394 534 21630
rect 618 21074 854 21310
rect 14786 21702 15022 21938
rect 14424 21340 14660 21576
rect 938 20754 1174 20990
rect 14104 21020 14340 21256
rect 13784 20700 14020 20936
rect 1261 20431 1497 20667
rect 1581 20431 1817 20667
rect 1901 20431 2137 20667
rect 2221 20431 2457 20667
rect 2541 20431 2777 20667
rect 2861 20431 3097 20667
rect 3181 20431 3417 20667
rect 3501 20431 3737 20667
rect 3821 20431 4057 20667
rect 4141 20431 4377 20667
rect 4461 20431 4697 20667
rect 4781 20431 5017 20667
rect 5101 20431 5337 20667
rect 5421 20431 5657 20667
rect 5741 20431 5977 20667
rect 6061 20431 6297 20667
rect 6381 20431 6617 20667
rect 6701 20431 6937 20667
rect 7021 20431 7257 20667
rect 7341 20431 7577 20667
rect 7661 20431 7897 20667
rect 7981 20431 8217 20667
rect 8301 20431 8537 20667
rect 8621 20431 8857 20667
rect 8941 20431 9177 20667
rect 9261 20431 9497 20667
rect 9581 20431 9817 20667
rect 9901 20431 10137 20667
rect 10221 20431 10457 20667
rect 10541 20431 10777 20667
rect 10861 20431 11097 20667
rect 11181 20431 11417 20667
rect 11501 20431 11737 20667
rect 11821 20431 12057 20667
rect 12141 20431 12377 20667
rect 12461 20431 12697 20667
rect 12781 20431 13017 20667
rect 13101 20431 13337 20667
rect 13421 20431 13657 20667
<< metal5 >>
tri 979 33194 1272 33487 se
rect 1272 33463 13740 33487
tri 13740 33463 13764 33487 sw
rect 1272 33227 1355 33463
rect 1591 33227 1675 33463
rect 1911 33227 1995 33463
rect 2231 33227 2315 33463
rect 2551 33227 2635 33463
rect 2871 33227 2955 33463
rect 3191 33227 3275 33463
rect 3511 33227 3595 33463
rect 3831 33227 3915 33463
rect 4151 33227 4235 33463
rect 4471 33227 4555 33463
rect 4791 33227 4875 33463
rect 5111 33227 5195 33463
rect 5431 33227 5515 33463
rect 5751 33227 5835 33463
rect 6071 33227 6155 33463
rect 6391 33227 6475 33463
rect 6711 33227 6795 33463
rect 7031 33227 7115 33463
rect 7351 33227 7435 33463
rect 7671 33227 7755 33463
rect 7991 33227 8075 33463
rect 8311 33227 8395 33463
rect 8631 33227 8715 33463
rect 8951 33227 9035 33463
rect 9271 33227 9355 33463
rect 9591 33227 9675 33463
rect 9911 33227 9995 33463
rect 10231 33227 10315 33463
rect 10551 33227 10635 33463
rect 10871 33227 10955 33463
rect 11191 33227 11275 33463
rect 11511 33227 11595 33463
rect 11831 33227 11915 33463
rect 12151 33227 12235 33463
rect 12471 33227 12555 33463
rect 12791 33227 12875 33463
rect 13111 33227 13195 33463
rect 13431 33227 13515 33463
rect 13751 33227 13764 33463
rect 1272 33194 13764 33227
tri 659 32874 979 33194 se
rect 979 32958 992 33194
rect 1228 33140 13764 33194
tri 13764 33140 14087 33463 sw
rect 1228 32958 13838 33140
rect 979 32904 13838 32958
rect 14074 32904 14087 33140
rect 979 32874 14087 32904
tri 339 32554 659 32874 se
rect 659 32638 672 32874
rect 908 32820 14087 32874
tri 14087 32820 14407 33140 sw
rect 908 32638 14158 32820
rect 659 32584 14158 32638
rect 14394 32584 14407 32820
rect 659 32554 14407 32584
tri -23 32192 339 32554 se
rect 339 32318 352 32554
rect 588 32500 14407 32554
tri 14407 32500 14727 32820 sw
rect 588 32318 14478 32500
rect 339 32264 14478 32318
rect 14714 32264 14727 32500
rect 339 32192 14727 32264
tri -34 32181 -23 32192 se
rect -23 32181 -10 32192
rect -34 31956 -10 32181
rect 226 32181 14727 32192
tri 14727 32181 15046 32500 sw
rect 226 32178 15046 32181
rect 226 31956 14786 32178
rect -34 31942 14786 31956
rect 15022 31942 15046 32178
rect -34 31872 15046 31942
rect -34 31636 -10 31872
rect 226 31858 15046 31872
rect 226 31636 14786 31858
rect -34 31622 14786 31636
rect 15022 31622 15046 31858
rect -34 31552 15046 31622
rect -34 31316 -10 31552
rect 226 31538 15046 31552
rect 226 31316 14786 31538
rect -34 31302 14786 31316
rect 15022 31302 15046 31538
rect -34 31232 15046 31302
rect -34 30996 -10 31232
rect 226 31218 15046 31232
rect 226 30996 14786 31218
rect -34 30982 14786 30996
rect 15022 30982 15046 31218
rect -34 30912 15046 30982
rect -34 30676 -10 30912
rect 226 30898 15046 30912
rect 226 30676 14786 30898
rect -34 30662 14786 30676
rect 15022 30662 15046 30898
rect -34 30592 15046 30662
rect -34 30356 -10 30592
rect 226 30578 15046 30592
rect 226 30356 14786 30578
rect -34 30342 14786 30356
rect 15022 30342 15046 30578
rect -34 30272 15046 30342
rect -34 30036 -10 30272
rect 226 30258 15046 30272
rect 226 30036 14786 30258
rect -34 30022 14786 30036
rect 15022 30022 15046 30258
rect -34 29952 15046 30022
rect -34 29716 -10 29952
rect 226 29938 15046 29952
rect 226 29716 14786 29938
rect -34 29702 14786 29716
rect 15022 29702 15046 29938
rect -34 29632 15046 29702
rect -34 29396 -10 29632
rect 226 29618 15046 29632
rect 226 29396 14786 29618
rect -34 29382 14786 29396
rect 15022 29382 15046 29618
rect -34 29312 15046 29382
rect -34 29076 -10 29312
rect 226 29298 15046 29312
rect 226 29076 14786 29298
rect -34 29062 14786 29076
rect 15022 29062 15046 29298
rect -34 28992 15046 29062
rect -34 28756 -10 28992
rect 226 28978 15046 28992
rect 226 28756 14786 28978
rect -34 28742 14786 28756
rect 15022 28742 15046 28978
rect -34 28672 15046 28742
rect -34 28436 -10 28672
rect 226 28658 15046 28672
rect 226 28436 14786 28658
rect -34 28422 14786 28436
rect 15022 28422 15046 28658
rect -34 28352 15046 28422
rect -34 28116 -10 28352
rect 226 28338 15046 28352
rect 226 28116 14786 28338
rect -34 28102 14786 28116
rect 15022 28102 15046 28338
rect -34 28032 15046 28102
rect -34 27796 -10 28032
rect 226 28018 15046 28032
rect 226 27796 14786 28018
rect -34 27782 14786 27796
rect 15022 27782 15046 28018
rect -34 27712 15046 27782
rect -34 27476 -10 27712
rect 226 27698 15046 27712
rect 226 27476 14786 27698
rect -34 27462 14786 27476
rect 15022 27462 15046 27698
rect -34 27392 15046 27462
rect -34 27156 -10 27392
rect 226 27378 15046 27392
rect 226 27156 14786 27378
rect -34 27142 14786 27156
rect 15022 27142 15046 27378
rect -34 27072 15046 27142
rect -34 26836 -10 27072
rect 226 27058 15046 27072
rect 226 26836 14786 27058
rect -34 26822 14786 26836
rect 15022 26822 15046 27058
rect -34 26752 15046 26822
rect -34 26516 -10 26752
rect 226 26738 15046 26752
rect 226 26516 14786 26738
rect -34 26502 14786 26516
rect 15022 26502 15046 26738
rect -34 26432 15046 26502
rect -34 26196 -10 26432
rect 226 26418 15046 26432
rect 226 26196 14786 26418
rect -34 26182 14786 26196
rect 15022 26182 15046 26418
rect -34 26112 15046 26182
rect -34 25876 -10 26112
rect 226 26098 15046 26112
rect 226 25876 14786 26098
rect -34 25862 14786 25876
rect 15022 25862 15046 26098
rect -34 25792 15046 25862
rect -34 25556 -10 25792
rect 226 25778 15046 25792
rect 226 25556 14786 25778
rect -34 25542 14786 25556
rect 15022 25542 15046 25778
rect -34 25472 15046 25542
rect -34 25236 -10 25472
rect 226 25458 15046 25472
rect 226 25236 14786 25458
rect -34 25222 14786 25236
rect 15022 25222 15046 25458
rect -34 25152 15046 25222
rect -34 24916 -10 25152
rect 226 25138 15046 25152
rect 226 24916 14786 25138
rect -34 24902 14786 24916
rect 15022 24902 15046 25138
rect -34 24832 15046 24902
rect -34 24596 -10 24832
rect 226 24818 15046 24832
rect 226 24596 14786 24818
rect -34 24582 14786 24596
rect 15022 24582 15046 24818
rect -34 24512 15046 24582
rect -34 24276 -10 24512
rect 226 24498 15046 24512
rect 226 24276 14786 24498
rect -34 24262 14786 24276
rect 15022 24262 15046 24498
rect -34 24192 15046 24262
rect -34 23956 -10 24192
rect 226 24178 15046 24192
rect 226 23956 14786 24178
rect -34 23942 14786 23956
rect 15022 23942 15046 24178
rect -34 23872 15046 23942
rect -34 23636 -10 23872
rect 226 23858 15046 23872
rect 226 23636 14786 23858
rect -34 23622 14786 23636
rect 15022 23622 15046 23858
rect -34 23552 15046 23622
rect -34 23316 -10 23552
rect 226 23538 15046 23552
rect 226 23316 14786 23538
rect -34 23302 14786 23316
rect 15022 23302 15046 23538
rect -34 23232 15046 23302
rect -34 22996 -10 23232
rect 226 23218 15046 23232
rect 226 22996 14786 23218
rect -34 22982 14786 22996
rect 15022 22982 15046 23218
rect -34 22912 15046 22982
rect -34 22676 -10 22912
rect 226 22898 15046 22912
rect 226 22676 14786 22898
rect -34 22662 14786 22676
rect 15022 22662 15046 22898
rect -34 22592 15046 22662
rect -34 22356 -10 22592
rect 226 22578 15046 22592
rect 226 22356 14786 22578
rect -34 22342 14786 22356
rect 15022 22342 15046 22578
rect -34 22272 15046 22342
rect -34 22036 -10 22272
rect 226 22258 15046 22272
rect 226 22036 14786 22258
rect -34 22022 14786 22036
rect 15022 22022 15046 22258
rect -34 21952 15046 22022
rect -34 21716 -10 21952
rect 226 21938 15046 21952
rect 226 21716 14786 21938
rect -34 21713 14786 21716
tri -34 21630 49 21713 ne
rect 49 21702 14786 21713
rect 15022 21713 15046 21938
rect 15022 21702 15035 21713
tri 15035 21702 15046 21713 nw
rect 49 21630 14909 21702
tri 49 21394 285 21630 ne
rect 285 21394 298 21630
rect 534 21576 14909 21630
tri 14909 21576 15035 21702 nw
rect 534 21394 14424 21576
tri 285 21310 369 21394 ne
rect 369 21340 14424 21394
rect 14660 21340 14673 21576
tri 14673 21340 14909 21576 nw
rect 369 21310 14589 21340
tri 369 21074 605 21310 ne
rect 605 21074 618 21310
rect 854 21256 14589 21310
tri 14589 21256 14673 21340 nw
rect 854 21074 14104 21256
tri 605 20990 689 21074 ne
rect 689 21020 14104 21074
rect 14340 21020 14353 21256
tri 14353 21020 14589 21256 nw
rect 689 20990 14269 21020
tri 689 20754 925 20990 ne
rect 925 20754 938 20990
rect 1174 20936 14269 20990
tri 14269 20936 14353 21020 nw
rect 1174 20754 13784 20936
tri 925 20667 1012 20754 ne
rect 1012 20700 13784 20754
rect 14020 20700 14033 20936
tri 14033 20700 14269 20936 nw
rect 1012 20667 13740 20700
tri 1012 20431 1248 20667 ne
rect 1248 20431 1261 20667
rect 1497 20431 1581 20667
rect 1817 20431 1901 20667
rect 2137 20431 2221 20667
rect 2457 20431 2541 20667
rect 2777 20431 2861 20667
rect 3097 20431 3181 20667
rect 3417 20431 3501 20667
rect 3737 20431 3821 20667
rect 4057 20431 4141 20667
rect 4377 20431 4461 20667
rect 4697 20431 4781 20667
rect 5017 20431 5101 20667
rect 5337 20431 5421 20667
rect 5657 20431 5741 20667
rect 5977 20431 6061 20667
rect 6297 20431 6381 20667
rect 6617 20431 6701 20667
rect 6937 20431 7021 20667
rect 7257 20431 7341 20667
rect 7577 20431 7661 20667
rect 7897 20431 7981 20667
rect 8217 20431 8301 20667
rect 8537 20431 8621 20667
rect 8857 20431 8941 20667
rect 9177 20431 9261 20667
rect 9497 20431 9581 20667
rect 9817 20431 9901 20667
rect 10137 20431 10221 20667
rect 10457 20431 10541 20667
rect 10777 20431 10861 20667
rect 11097 20431 11181 20667
rect 11417 20431 11501 20667
rect 11737 20431 11821 20667
rect 12057 20431 12141 20667
rect 12377 20431 12461 20667
rect 12697 20431 12781 20667
rect 13017 20431 13101 20667
rect 13337 20431 13421 20667
rect 13657 20431 13740 20667
tri 1248 20407 1272 20431 ne
rect 1272 20407 13740 20431
tri 13740 20407 14033 20700 nw
<< glass >>
tri 506 31957 1496 32947 se
rect 1496 31957 13516 32947
tri 13516 31957 14506 32947 sw
rect 506 21937 14506 31957
tri 506 20947 1496 21937 ne
rect 1496 20947 13516 21937
tri 13516 20947 14506 21937 nw
use sky130_fd_pr__padplhp__example_559591418080  sky130_fd_pr__padplhp__example_559591418080_0
timestamp 1624855509
transform 0 -1 14506 1 0 20947
box -478 -478 6000 7000
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 49858642
string GDS_START 49858552
<< end >>
