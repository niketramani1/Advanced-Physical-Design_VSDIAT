magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1114 -1260 4421 5060
<< nwell >>
rect 737 168 905 890
rect 1971 168 2139 890
rect 737 0 2139 168
<< pwell >>
rect 804 890 838 956
rect 2038 890 2072 956
rect 1005 756 1871 790
rect 1005 302 1039 756
rect 1837 302 1871 756
rect 1005 268 1871 302
<< mvnmos >>
rect 1163 429 1763 629
<< mvndiff >>
rect 1163 674 1763 682
rect 1163 640 1241 674
rect 1275 640 1309 674
rect 1343 640 1377 674
rect 1411 640 1445 674
rect 1479 640 1513 674
rect 1547 640 1581 674
rect 1615 640 1649 674
rect 1683 640 1717 674
rect 1751 640 1763 674
rect 1163 629 1763 640
rect 1163 418 1763 429
rect 1163 384 1241 418
rect 1275 384 1309 418
rect 1343 384 1377 418
rect 1411 384 1445 418
rect 1479 384 1513 418
rect 1547 384 1581 418
rect 1615 384 1649 418
rect 1683 384 1717 418
rect 1751 384 1763 418
rect 1163 376 1763 384
<< mvndiffc >>
rect 1241 640 1275 674
rect 1309 640 1343 674
rect 1377 640 1411 674
rect 1445 640 1479 674
rect 1513 640 1547 674
rect 1581 640 1615 674
rect 1649 640 1683 674
rect 1717 640 1751 674
rect 1241 384 1275 418
rect 1309 384 1343 418
rect 1377 384 1411 418
rect 1445 384 1479 418
rect 1513 384 1547 418
rect 1581 384 1615 418
rect 1649 384 1683 418
rect 1717 384 1751 418
<< mvpsubdiff >>
rect 1005 756 1107 790
rect 1141 756 1175 790
rect 1209 756 1243 790
rect 1277 756 1311 790
rect 1345 756 1379 790
rect 1413 756 1447 790
rect 1481 756 1515 790
rect 1549 756 1583 790
rect 1617 756 1651 790
rect 1685 756 1803 790
rect 1005 688 1039 722
rect 1005 620 1039 654
rect 1837 676 1871 790
rect 1005 552 1039 586
rect 1005 484 1039 518
rect 1005 416 1039 450
rect 1837 608 1871 642
rect 1837 540 1871 574
rect 1837 472 1871 506
rect 1005 268 1039 382
rect 1837 404 1871 438
rect 1837 336 1871 370
rect 1073 268 1107 302
rect 1141 268 1175 302
rect 1209 268 1243 302
rect 1277 268 1311 302
rect 1345 268 1379 302
rect 1413 268 1447 302
rect 1481 268 1515 302
rect 1549 268 1583 302
rect 1617 268 1651 302
rect 1685 268 1719 302
rect 1753 268 1871 302
<< mvnsubdiff >>
rect 804 789 838 890
rect 804 721 838 755
rect 804 653 838 687
rect 804 585 838 619
rect 804 517 838 551
rect 804 449 838 483
rect 804 381 838 415
rect 804 313 838 347
rect 804 245 838 279
rect 2038 781 2072 890
rect 2038 713 2072 747
rect 2038 645 2072 679
rect 2038 577 2072 611
rect 2038 509 2072 543
rect 2038 441 2072 475
rect 2038 373 2072 407
rect 2038 305 2072 339
rect 804 177 838 211
rect 804 101 838 143
rect 2038 237 2072 271
rect 2038 169 2072 203
rect 2038 101 2072 135
rect 804 67 872 101
rect 906 67 940 101
rect 974 67 1008 101
rect 1042 67 1076 101
rect 1110 67 1144 101
rect 1178 67 1212 101
rect 1246 67 1280 101
rect 1314 67 1348 101
rect 1382 67 1416 101
rect 1450 67 1484 101
rect 1518 67 1552 101
rect 1586 67 1620 101
rect 1654 67 1688 101
rect 1722 67 1756 101
rect 1790 67 1824 101
rect 1858 67 1892 101
rect 1926 67 1960 101
rect 1994 67 2072 101
<< mvpsubdiffcont >>
rect 1107 756 1141 790
rect 1175 756 1209 790
rect 1243 756 1277 790
rect 1311 756 1345 790
rect 1379 756 1413 790
rect 1447 756 1481 790
rect 1515 756 1549 790
rect 1583 756 1617 790
rect 1651 756 1685 790
rect 1803 756 1837 790
rect 1005 722 1039 756
rect 1005 654 1039 688
rect 1837 642 1871 676
rect 1005 586 1039 620
rect 1005 518 1039 552
rect 1005 450 1039 484
rect 1837 574 1871 608
rect 1837 506 1871 540
rect 1837 438 1871 472
rect 1005 382 1039 416
rect 1837 370 1871 404
rect 1837 302 1871 336
rect 1039 268 1073 302
rect 1107 268 1141 302
rect 1175 268 1209 302
rect 1243 268 1277 302
rect 1311 268 1345 302
rect 1379 268 1413 302
rect 1447 268 1481 302
rect 1515 268 1549 302
rect 1583 268 1617 302
rect 1651 268 1685 302
rect 1719 268 1753 302
<< mvnsubdiffcont >>
rect 804 755 838 789
rect 804 687 838 721
rect 804 619 838 653
rect 804 551 838 585
rect 804 483 838 517
rect 804 415 838 449
rect 804 347 838 381
rect 804 279 838 313
rect 2038 747 2072 781
rect 2038 679 2072 713
rect 2038 611 2072 645
rect 2038 543 2072 577
rect 2038 475 2072 509
rect 2038 407 2072 441
rect 2038 339 2072 373
rect 2038 271 2072 305
rect 804 211 838 245
rect 804 143 838 177
rect 2038 203 2072 237
rect 2038 135 2072 169
rect 872 67 906 101
rect 940 67 974 101
rect 1008 67 1042 101
rect 1076 67 1110 101
rect 1144 67 1178 101
rect 1212 67 1246 101
rect 1280 67 1314 101
rect 1348 67 1382 101
rect 1416 67 1450 101
rect 1484 67 1518 101
rect 1552 67 1586 101
rect 1620 67 1654 101
rect 1688 67 1722 101
rect 1756 67 1790 101
rect 1824 67 1858 101
rect 1892 67 1926 101
rect 1960 67 1994 101
<< poly >>
rect 1071 613 1163 629
rect 1071 579 1087 613
rect 1121 579 1163 613
rect 1071 545 1163 579
rect 1071 511 1087 545
rect 1121 511 1163 545
rect 1071 477 1163 511
rect 1071 443 1087 477
rect 1121 443 1163 477
rect 1071 429 1163 443
rect 1763 429 1789 629
rect 1071 427 1137 429
<< polycont >>
rect 1087 579 1121 613
rect 1087 511 1121 545
rect 1087 443 1121 477
<< locali >>
rect 804 789 838 956
rect 2038 823 2072 972
rect 804 754 838 755
rect 804 681 838 687
rect 804 608 838 619
rect 804 535 838 551
rect 804 462 838 483
rect 804 389 838 415
rect 804 317 838 347
rect 804 245 838 279
rect 999 790 1877 796
rect 999 756 1097 790
rect 1141 756 1175 790
rect 1224 756 1243 790
rect 1277 756 1283 790
rect 1345 756 1379 790
rect 1415 756 1447 790
rect 1491 756 1515 790
rect 1567 756 1583 790
rect 1643 756 1651 790
rect 1719 756 1761 790
rect 1795 756 1803 790
rect 1837 756 1877 790
rect 999 722 1005 756
rect 1039 750 1877 756
rect 1039 722 1045 750
rect 999 718 1045 722
rect 999 654 1005 718
rect 1039 654 1045 718
rect 1831 712 1877 750
rect 1831 678 1837 712
rect 1871 678 1877 712
rect 1831 676 1877 678
rect 999 634 1045 654
rect 1225 640 1226 674
rect 1275 640 1298 674
rect 1343 640 1370 674
rect 1411 640 1442 674
rect 1479 640 1513 674
rect 1548 640 1581 674
rect 1620 640 1649 674
rect 1692 640 1717 674
rect 1764 640 1767 674
rect 1831 642 1837 676
rect 1871 642 1877 676
rect 999 586 1005 634
rect 1039 586 1045 634
rect 999 552 1045 586
rect 999 517 1005 552
rect 1039 517 1045 552
rect 999 484 1045 517
rect 999 434 1005 484
rect 1039 434 1045 484
rect 999 416 1045 434
rect 1087 613 1121 629
rect 1087 545 1121 552
rect 1087 477 1121 480
rect 1087 427 1121 443
rect 1831 608 1877 642
rect 1831 573 1837 608
rect 1871 573 1877 608
rect 1831 540 1877 573
rect 1831 496 1837 540
rect 1871 496 1877 540
rect 1831 472 1877 496
rect 1831 418 1837 472
rect 1871 418 1877 472
rect 999 351 1005 416
rect 1039 351 1045 416
rect 1275 384 1307 418
rect 1343 384 1377 418
rect 1422 384 1445 418
rect 1503 384 1513 418
rect 1547 384 1550 418
rect 1615 384 1631 418
rect 1683 384 1712 418
rect 1751 384 1767 418
rect 1831 404 1877 418
rect 999 308 1045 351
rect 1831 340 1837 404
rect 1871 340 1877 404
rect 1831 336 1877 340
rect 1831 308 1837 336
rect 999 302 1837 308
rect 1871 302 1877 336
rect 999 268 1039 302
rect 1073 268 1077 302
rect 1141 268 1153 302
rect 1209 268 1229 302
rect 1277 268 1305 302
rect 1345 268 1379 302
rect 1415 268 1447 302
rect 1491 268 1515 302
rect 1567 268 1583 302
rect 1643 268 1651 302
rect 1753 268 1761 302
rect 1795 268 1877 302
rect 999 262 1877 268
rect 2038 781 2072 789
rect 2038 713 2072 717
rect 2038 607 2072 611
rect 2038 535 2072 543
rect 2038 463 2072 475
rect 2038 391 2072 407
rect 2038 319 2072 339
rect 804 177 838 211
rect 804 101 838 139
rect 2038 246 2072 271
rect 2038 173 2072 203
rect 2038 101 2072 135
rect 804 67 872 101
rect 910 67 940 101
rect 983 67 1008 101
rect 1056 67 1076 101
rect 1129 67 1144 101
rect 1202 67 1212 101
rect 1275 67 1280 101
rect 1382 67 1387 101
rect 1450 67 1460 101
rect 1518 67 1533 101
rect 1586 67 1606 101
rect 1654 67 1678 101
rect 1722 67 1750 101
rect 1790 67 1822 101
rect 1858 67 1892 101
rect 1928 67 1960 101
rect 2000 67 2072 101
<< viali >>
rect 804 721 838 754
rect 804 720 838 721
rect 804 653 838 681
rect 804 647 838 653
rect 804 585 838 608
rect 804 574 838 585
rect 804 517 838 535
rect 804 501 838 517
rect 804 449 838 462
rect 804 428 838 449
rect 804 381 838 389
rect 804 355 838 381
rect 804 313 838 317
rect 804 283 838 313
rect 1097 756 1107 790
rect 1107 756 1131 790
rect 1190 756 1209 790
rect 1209 756 1224 790
rect 1283 756 1311 790
rect 1311 756 1317 790
rect 1381 756 1413 790
rect 1413 756 1415 790
rect 1457 756 1481 790
rect 1481 756 1491 790
rect 1533 756 1549 790
rect 1549 756 1567 790
rect 1609 756 1617 790
rect 1617 756 1643 790
rect 1685 756 1719 790
rect 1761 756 1795 790
rect 1005 688 1039 718
rect 1005 684 1039 688
rect 1837 678 1871 712
rect 1226 640 1241 674
rect 1241 640 1260 674
rect 1298 640 1309 674
rect 1309 640 1332 674
rect 1370 640 1377 674
rect 1377 640 1404 674
rect 1442 640 1445 674
rect 1445 640 1476 674
rect 1514 640 1547 674
rect 1547 640 1548 674
rect 1586 640 1615 674
rect 1615 640 1620 674
rect 1658 640 1683 674
rect 1683 640 1692 674
rect 1730 640 1751 674
rect 1751 640 1764 674
rect 1005 620 1039 634
rect 1005 600 1039 620
rect 1005 518 1039 551
rect 1005 517 1039 518
rect 1005 450 1039 468
rect 1005 434 1039 450
rect 1087 579 1121 586
rect 1087 552 1121 579
rect 1087 511 1121 514
rect 1087 480 1121 511
rect 1837 574 1871 607
rect 1837 573 1871 574
rect 1837 506 1871 530
rect 1837 496 1871 506
rect 1837 438 1871 452
rect 1837 418 1871 438
rect 1005 382 1039 385
rect 1005 351 1039 382
rect 1225 384 1241 418
rect 1241 384 1259 418
rect 1307 384 1309 418
rect 1309 384 1341 418
rect 1388 384 1411 418
rect 1411 384 1422 418
rect 1469 384 1479 418
rect 1479 384 1503 418
rect 1550 384 1581 418
rect 1581 384 1584 418
rect 1631 384 1649 418
rect 1649 384 1665 418
rect 1712 384 1717 418
rect 1717 384 1746 418
rect 1837 370 1871 374
rect 1837 340 1871 370
rect 1077 268 1107 302
rect 1107 268 1111 302
rect 1153 268 1175 302
rect 1175 268 1187 302
rect 1229 268 1243 302
rect 1243 268 1263 302
rect 1305 268 1311 302
rect 1311 268 1339 302
rect 1381 268 1413 302
rect 1413 268 1415 302
rect 1457 268 1481 302
rect 1481 268 1491 302
rect 1533 268 1549 302
rect 1549 268 1567 302
rect 1609 268 1617 302
rect 1617 268 1643 302
rect 1685 268 1719 302
rect 1761 268 1795 302
rect 2038 789 2072 823
rect 2038 747 2072 751
rect 2038 717 2072 747
rect 2038 645 2072 679
rect 2038 577 2072 607
rect 2038 573 2072 577
rect 2038 509 2072 535
rect 2038 501 2072 509
rect 2038 441 2072 463
rect 2038 429 2072 441
rect 2038 373 2072 391
rect 2038 357 2072 373
rect 2038 305 2072 319
rect 2038 285 2072 305
rect 804 211 838 245
rect 804 143 838 173
rect 804 139 838 143
rect 2038 237 2072 246
rect 2038 212 2072 237
rect 2038 169 2072 173
rect 2038 139 2072 169
rect 876 67 906 101
rect 906 67 910 101
rect 949 67 974 101
rect 974 67 983 101
rect 1022 67 1042 101
rect 1042 67 1056 101
rect 1095 67 1110 101
rect 1110 67 1129 101
rect 1168 67 1178 101
rect 1178 67 1202 101
rect 1241 67 1246 101
rect 1246 67 1275 101
rect 1314 67 1348 101
rect 1387 67 1416 101
rect 1416 67 1421 101
rect 1460 67 1484 101
rect 1484 67 1494 101
rect 1533 67 1552 101
rect 1552 67 1567 101
rect 1606 67 1620 101
rect 1620 67 1640 101
rect 1678 67 1688 101
rect 1688 67 1712 101
rect 1750 67 1756 101
rect 1756 67 1784 101
rect 1822 67 1824 101
rect 1824 67 1856 101
rect 1894 67 1926 101
rect 1926 67 1928 101
rect 1966 67 1994 101
rect 1994 67 2000 101
<< metal1 >>
rect 1409 3682 1415 3734
rect 1467 3682 1483 3734
rect 1535 3682 1551 3734
rect 1603 3682 1618 3734
rect 1670 3682 1685 3734
rect 1737 3682 1752 3734
rect 1804 3682 1810 3734
rect 1409 3646 1810 3682
rect 1409 3594 1415 3646
rect 1467 3594 1483 3646
rect 1535 3594 1551 3646
rect 1603 3594 1618 3646
rect 1670 3594 1685 3646
rect 1737 3594 1752 3646
rect 1804 3594 1810 3646
rect 1890 3594 2291 3734
rect 2240 3390 2246 3442
rect 2298 3390 2316 3442
rect 2368 3390 2385 3442
rect 2437 3390 2454 3442
rect 2506 3390 2523 3442
rect 2575 3390 2581 3442
rect 2240 3354 2581 3390
rect 2240 3302 2246 3354
rect 2298 3302 2316 3354
rect 2368 3302 2385 3354
rect 2437 3302 2454 3354
rect 2506 3302 2523 3354
rect 2575 3302 2581 3354
rect 2638 3370 2803 3376
rect 2690 3318 2750 3370
rect 2802 3318 2803 3370
rect 2638 3262 2803 3318
rect 1409 3188 1415 3240
rect 1467 3188 1483 3240
rect 1535 3188 1551 3240
rect 1603 3188 1618 3240
rect 1670 3188 1685 3240
rect 1737 3188 1752 3240
rect 1804 3188 1810 3240
rect 1409 3166 1810 3188
rect 1409 3114 1415 3166
rect 1467 3114 1483 3166
rect 1535 3114 1551 3166
rect 1603 3114 1618 3166
rect 1670 3114 1685 3166
rect 1737 3114 1752 3166
rect 1804 3114 1810 3166
rect 1409 3092 1810 3114
rect 1409 3040 1415 3092
rect 1467 3040 1483 3092
rect 1535 3040 1551 3092
rect 1603 3040 1618 3092
rect 1670 3040 1685 3092
rect 1737 3040 1752 3092
rect 1804 3040 1810 3092
rect 1890 3040 2291 3240
rect 2690 3210 2750 3262
rect 2802 3210 2803 3262
rect 2638 3153 2803 3210
rect 2690 3101 2750 3153
rect 2802 3101 2803 3153
rect 2638 3095 2803 3101
rect 2638 3009 2644 3061
rect 2696 3009 2745 3061
rect 2797 3009 2803 3061
rect 147 2781 831 2981
rect 1214 2975 1314 2981
rect 1214 2923 1238 2975
rect 1290 2923 1314 2975
rect 1214 2907 1314 2923
rect 2638 2965 2803 3009
rect 2638 2913 2644 2965
rect 2696 2913 2745 2965
rect 2797 2913 2803 2965
rect 1214 2855 1238 2907
rect 1290 2855 1314 2907
rect 1214 2839 1314 2855
rect 1214 2787 1238 2839
rect 1290 2787 1314 2839
rect 1214 2781 1314 2787
rect 2638 2872 2803 2878
rect 2690 2820 2750 2872
rect 2802 2820 2803 2872
rect 2638 2782 2803 2820
rect 147 2381 549 2781
tri 549 2571 759 2781 nw
rect 999 2739 1127 2745
rect 999 2687 1005 2739
rect 1057 2687 1069 2739
rect 1121 2687 1127 2739
rect 999 2625 1127 2687
rect 999 2573 1005 2625
rect 1057 2573 1069 2625
rect 1121 2573 1127 2625
rect 999 2567 1127 2573
rect 1890 2693 2246 2745
rect 2298 2693 2339 2745
rect 2391 2693 2431 2745
rect 2483 2693 2523 2745
rect 2575 2693 2581 2745
rect 1890 2619 2581 2693
rect 2690 2730 2750 2782
rect 2802 2730 2803 2782
rect 2638 2692 2803 2730
rect 2690 2640 2750 2692
rect 2802 2640 2803 2692
rect 2638 2634 2803 2640
rect 1890 2567 2246 2619
rect 2298 2567 2339 2619
rect 2391 2567 2431 2619
rect 2483 2567 2523 2619
rect 2575 2567 2581 2619
rect 1409 2363 1415 2415
rect 1467 2363 1483 2415
rect 1535 2363 1551 2415
rect 1603 2363 1618 2415
rect 1670 2363 1685 2415
rect 1737 2363 1752 2415
rect 1804 2363 1810 2415
rect 1409 2327 1810 2363
rect 1409 2275 1415 2327
rect 1467 2275 1483 2327
rect 1535 2275 1551 2327
rect 1603 2275 1618 2327
rect 1670 2275 1685 2327
rect 1737 2275 1752 2327
rect 1804 2275 1810 2327
rect 1890 2275 2291 2415
rect 2986 2257 3095 2437
rect 1005 2117 1121 2123
rect 1057 2065 1069 2117
rect 1005 2003 1121 2065
rect 1057 1951 1069 2003
rect 1005 1945 1121 1951
rect 1890 2071 2246 2123
rect 2298 2071 2339 2123
rect 2391 2071 2431 2123
rect 2483 2071 2523 2123
rect 2575 2071 2581 2123
rect 1890 1997 2581 2071
rect 1890 1945 2246 1997
rect 2298 1945 2339 1997
rect 2391 1945 2431 1997
rect 2483 1945 2523 1997
rect 2575 1945 2581 1997
rect 2638 2051 2803 2057
rect 2690 1999 2750 2051
rect 2802 1999 2803 2051
rect 2638 1961 2803 1999
rect 2690 1909 2750 1961
rect 2802 1909 2803 1961
rect 1005 1903 1121 1909
rect 1057 1851 1069 1903
rect 1005 1835 1121 1851
rect 1057 1783 1069 1835
rect 1005 1767 1121 1783
rect 1057 1715 1069 1767
rect 1005 1709 1121 1715
rect 1890 1857 2246 1909
rect 2298 1857 2388 1909
rect 2440 1857 2446 1909
rect 1890 1835 2446 1857
rect 1890 1783 2246 1835
rect 2298 1783 2388 1835
rect 2440 1783 2446 1835
rect 2638 1870 2803 1909
rect 2690 1818 2750 1870
rect 2802 1818 2803 1870
rect 2638 1812 2803 1818
rect 1890 1761 2446 1783
rect 1890 1709 2246 1761
rect 2298 1709 2388 1761
rect 2440 1709 2446 1761
rect 2638 1777 2803 1778
rect 2638 1725 2644 1777
rect 2696 1725 2745 1777
rect 2797 1725 2803 1777
rect 2638 1681 2803 1725
rect 1214 1644 1314 1650
rect 1214 1592 1238 1644
rect 1290 1592 1314 1644
rect 2638 1629 2644 1681
rect 2696 1629 2745 1681
rect 2797 1629 2803 1681
rect 1214 1576 1314 1592
rect 1214 1524 1238 1576
rect 1290 1524 1314 1576
rect 1214 1508 1314 1524
rect 1214 1456 1238 1508
rect 1290 1456 1314 1508
rect 1214 1450 1314 1456
rect 2638 1589 2803 1595
rect 2690 1537 2750 1589
rect 2802 1537 2803 1589
rect 2638 1481 2803 1537
rect 2607 1418 2622 1430
rect 2690 1429 2750 1481
rect 2802 1429 2803 1481
rect 1890 1336 2246 1388
rect 2298 1336 2339 1388
rect 2391 1336 2431 1388
rect 2483 1336 2523 1388
rect 2575 1336 2581 1388
rect 1890 1300 2581 1336
rect 2638 1372 2803 1429
rect 2690 1320 2750 1372
rect 2802 1320 2803 1372
rect 2638 1314 2803 1320
rect 1890 1248 2246 1300
rect 2298 1248 2339 1300
rect 2391 1248 2431 1300
rect 2483 1248 2523 1300
rect 2575 1248 2581 1300
rect 1409 1044 1415 1096
rect 1467 1044 1483 1096
rect 1535 1044 1551 1096
rect 1603 1044 1618 1096
rect 1670 1044 1685 1096
rect 1737 1044 1752 1096
rect 1804 1044 1810 1096
rect 1409 1008 1810 1044
rect 1409 956 1415 1008
rect 1467 956 1483 1008
rect 1535 956 1551 1008
rect 1603 956 1618 1008
rect 1670 956 1685 1008
rect 1737 956 1752 1008
rect 1804 956 1810 1008
tri 1998 922 2032 956 ne
rect 2032 823 2078 956
tri 2078 922 2112 956 nw
rect 798 754 844 766
rect 798 720 804 754
rect 838 720 844 754
rect 798 681 844 720
rect 798 647 804 681
rect 838 647 844 681
rect 798 608 844 647
rect 798 574 804 608
rect 838 574 844 608
rect 798 535 844 574
rect 798 501 804 535
rect 838 501 844 535
rect 798 462 844 501
rect 798 428 804 462
rect 838 428 844 462
rect 798 389 844 428
rect 798 355 804 389
rect 838 355 844 389
rect 798 317 844 355
rect 798 283 804 317
rect 838 283 844 317
rect 798 245 844 283
rect 999 750 1005 802
rect 1057 750 1069 802
rect 1121 796 1127 802
rect 1121 790 1877 796
rect 1131 756 1190 790
rect 1224 756 1283 790
rect 1317 756 1381 790
rect 1415 756 1457 790
rect 1491 756 1533 790
rect 1567 756 1609 790
rect 1643 756 1685 790
rect 1719 756 1761 790
rect 1795 756 1877 790
rect 1121 750 1877 756
rect 999 718 1046 750
rect 999 684 1005 718
rect 1039 717 1046 718
tri 1046 717 1079 750 nw
tri 1797 717 1830 750 ne
rect 1830 717 1877 750
rect 1039 684 1045 717
tri 1045 716 1046 717 nw
tri 1830 716 1831 717 ne
rect 999 634 1045 684
rect 1831 712 1877 717
rect 999 600 1005 634
rect 1039 600 1045 634
rect 1214 631 1220 683
rect 1272 674 1299 683
rect 1351 674 1378 683
rect 1430 674 1779 683
rect 1272 640 1298 674
rect 1351 640 1370 674
rect 1430 640 1442 674
rect 1476 640 1514 674
rect 1548 640 1586 674
rect 1620 640 1658 674
rect 1692 640 1730 674
rect 1764 640 1779 674
rect 1272 631 1299 640
rect 1351 631 1378 640
rect 1430 631 1779 640
rect 1831 678 1837 712
rect 1871 678 1877 712
rect 999 551 1045 600
rect 1831 607 1877 678
rect 999 517 1005 551
rect 1039 517 1045 551
rect 999 468 1045 517
rect 1078 591 1130 598
rect 1078 527 1130 539
rect 1078 468 1130 475
rect 1831 573 1837 607
rect 1871 573 1877 607
rect 1831 530 1877 573
rect 1831 496 1837 530
rect 1871 496 1877 530
rect 999 434 1005 468
rect 1039 434 1045 468
rect 999 385 1045 434
rect 1831 452 1877 496
rect 999 351 1005 385
rect 1039 351 1045 385
rect 1213 375 1219 427
rect 1271 375 1285 427
rect 1337 418 1351 427
rect 1403 418 1416 427
rect 1468 418 1758 427
rect 1341 384 1351 418
rect 1468 384 1469 418
rect 1503 384 1550 418
rect 1584 384 1631 418
rect 1665 384 1712 418
rect 1746 384 1758 418
rect 1337 375 1351 384
rect 1403 375 1416 384
rect 1468 375 1758 384
rect 1831 418 1837 452
rect 1871 418 1877 452
rect 999 340 1045 351
rect 1831 374 1877 418
tri 1045 340 1047 342 sw
tri 1829 340 1831 342 se
rect 1831 340 1837 374
rect 1871 340 1877 374
rect 999 319 1047 340
tri 1047 319 1068 340 sw
tri 1808 319 1829 340 se
rect 1829 319 1877 340
rect 999 308 1068 319
tri 1068 308 1079 319 sw
tri 1797 308 1808 319 se
rect 1808 308 1877 319
rect 999 302 1877 308
rect 999 268 1077 302
rect 1111 268 1153 302
rect 1187 268 1229 302
rect 1263 268 1305 302
rect 1339 268 1381 302
rect 1415 268 1457 302
rect 1491 268 1533 302
rect 1567 268 1609 302
rect 1643 268 1685 302
rect 1719 268 1761 302
rect 1795 268 1877 302
rect 999 262 1877 268
rect 2032 789 2038 823
rect 2072 789 2078 823
rect 2032 751 2078 789
rect 2032 717 2038 751
rect 2072 717 2078 751
rect 2032 679 2078 717
rect 2032 645 2038 679
rect 2072 645 2078 679
rect 2032 607 2078 645
rect 2032 573 2038 607
rect 2072 573 2078 607
rect 2032 535 2078 573
rect 2032 501 2038 535
rect 2072 501 2078 535
rect 2032 463 2078 501
rect 2032 429 2038 463
rect 2072 429 2078 463
rect 2032 391 2078 429
rect 2032 357 2038 391
rect 2072 357 2078 391
rect 2032 319 2078 357
rect 2032 285 2038 319
rect 2072 285 2078 319
rect 798 211 804 245
rect 838 211 844 245
rect 798 173 844 211
rect 220 116 443 157
rect 798 139 804 173
rect 838 139 844 173
rect 2032 246 2078 285
rect 2032 212 2038 246
rect 2072 212 2078 246
rect 2032 173 2078 212
tri 844 139 849 144 sw
tri 2027 139 2032 144 se
rect 2032 139 2038 173
rect 2072 139 2078 173
rect 798 110 849 139
tri 849 110 878 139 sw
tri 1998 110 2027 139 se
rect 2027 110 2078 139
rect 798 101 1688 110
rect 1740 101 1752 110
rect 1804 101 2078 110
rect 798 67 876 101
rect 910 67 949 101
rect 983 67 1022 101
rect 1056 67 1095 101
rect 1129 67 1168 101
rect 1202 67 1241 101
rect 1275 67 1314 101
rect 1348 67 1387 101
rect 1421 67 1460 101
rect 1494 67 1533 101
rect 1567 67 1606 101
rect 1640 67 1678 101
rect 1740 67 1750 101
rect 1804 67 1822 101
rect 1856 67 1894 101
rect 1928 67 1966 101
rect 2000 67 2078 101
rect 798 58 1688 67
rect 1740 58 1752 67
rect 1804 58 2078 67
<< via1 >>
rect 1415 3682 1467 3734
rect 1483 3682 1535 3734
rect 1551 3682 1603 3734
rect 1618 3682 1670 3734
rect 1685 3682 1737 3734
rect 1752 3682 1804 3734
rect 1415 3594 1467 3646
rect 1483 3594 1535 3646
rect 1551 3594 1603 3646
rect 1618 3594 1670 3646
rect 1685 3594 1737 3646
rect 1752 3594 1804 3646
rect 2246 3390 2298 3442
rect 2316 3390 2368 3442
rect 2385 3390 2437 3442
rect 2454 3390 2506 3442
rect 2523 3390 2575 3442
rect 2246 3302 2298 3354
rect 2316 3302 2368 3354
rect 2385 3302 2437 3354
rect 2454 3302 2506 3354
rect 2523 3302 2575 3354
rect 2638 3318 2690 3370
rect 2750 3318 2802 3370
rect 1415 3188 1467 3240
rect 1483 3188 1535 3240
rect 1551 3188 1603 3240
rect 1618 3188 1670 3240
rect 1685 3188 1737 3240
rect 1752 3188 1804 3240
rect 1415 3114 1467 3166
rect 1483 3114 1535 3166
rect 1551 3114 1603 3166
rect 1618 3114 1670 3166
rect 1685 3114 1737 3166
rect 1752 3114 1804 3166
rect 1415 3040 1467 3092
rect 1483 3040 1535 3092
rect 1551 3040 1603 3092
rect 1618 3040 1670 3092
rect 1685 3040 1737 3092
rect 1752 3040 1804 3092
rect 2638 3210 2690 3262
rect 2750 3210 2802 3262
rect 2638 3101 2690 3153
rect 2750 3101 2802 3153
rect 2644 3009 2696 3061
rect 2745 3009 2797 3061
rect 1238 2923 1290 2975
rect 2644 2913 2696 2965
rect 2745 2913 2797 2965
rect 1238 2855 1290 2907
rect 1238 2787 1290 2839
rect 2638 2820 2690 2872
rect 2750 2820 2802 2872
rect 1005 2687 1057 2739
rect 1069 2687 1121 2739
rect 1005 2573 1057 2625
rect 1069 2573 1121 2625
rect 2246 2693 2298 2745
rect 2339 2693 2391 2745
rect 2431 2693 2483 2745
rect 2523 2693 2575 2745
rect 2638 2730 2690 2782
rect 2750 2730 2802 2782
rect 2638 2640 2690 2692
rect 2750 2640 2802 2692
rect 2246 2567 2298 2619
rect 2339 2567 2391 2619
rect 2431 2567 2483 2619
rect 2523 2567 2575 2619
rect 1415 2363 1467 2415
rect 1483 2363 1535 2415
rect 1551 2363 1603 2415
rect 1618 2363 1670 2415
rect 1685 2363 1737 2415
rect 1752 2363 1804 2415
rect 1415 2275 1467 2327
rect 1483 2275 1535 2327
rect 1551 2275 1603 2327
rect 1618 2275 1670 2327
rect 1685 2275 1737 2327
rect 1752 2275 1804 2327
rect 1005 2065 1057 2117
rect 1069 2065 1121 2117
rect 1005 1951 1057 2003
rect 1069 1951 1121 2003
rect 2246 2071 2298 2123
rect 2339 2071 2391 2123
rect 2431 2071 2483 2123
rect 2523 2071 2575 2123
rect 2246 1945 2298 1997
rect 2339 1945 2391 1997
rect 2431 1945 2483 1997
rect 2523 1945 2575 1997
rect 2638 1999 2690 2051
rect 2750 1999 2802 2051
rect 2638 1909 2690 1961
rect 2750 1909 2802 1961
rect 1005 1851 1057 1903
rect 1069 1851 1121 1903
rect 1005 1783 1057 1835
rect 1069 1783 1121 1835
rect 1005 1715 1057 1767
rect 1069 1715 1121 1767
rect 2246 1857 2298 1909
rect 2388 1857 2440 1909
rect 2246 1783 2298 1835
rect 2388 1783 2440 1835
rect 2638 1818 2690 1870
rect 2750 1818 2802 1870
rect 2246 1709 2298 1761
rect 2388 1709 2440 1761
rect 2644 1725 2696 1777
rect 2745 1725 2797 1777
rect 1238 1592 1290 1644
rect 2644 1629 2696 1681
rect 2745 1629 2797 1681
rect 1238 1524 1290 1576
rect 1238 1456 1290 1508
rect 2638 1537 2690 1589
rect 2750 1537 2802 1589
rect 2638 1429 2690 1481
rect 2750 1429 2802 1481
rect 2246 1336 2298 1388
rect 2339 1336 2391 1388
rect 2431 1336 2483 1388
rect 2523 1336 2575 1388
rect 2638 1320 2690 1372
rect 2750 1320 2802 1372
rect 2246 1248 2298 1300
rect 2339 1248 2391 1300
rect 2431 1248 2483 1300
rect 2523 1248 2575 1300
rect 1415 1044 1467 1096
rect 1483 1044 1535 1096
rect 1551 1044 1603 1096
rect 1618 1044 1670 1096
rect 1685 1044 1737 1096
rect 1752 1044 1804 1096
rect 1415 956 1467 1008
rect 1483 956 1535 1008
rect 1551 956 1603 1008
rect 1618 956 1670 1008
rect 1685 956 1737 1008
rect 1752 956 1804 1008
rect 1005 750 1057 802
rect 1069 790 1121 802
rect 1069 756 1097 790
rect 1097 756 1121 790
rect 1069 750 1121 756
rect 1220 674 1272 683
rect 1299 674 1351 683
rect 1378 674 1430 683
rect 1220 640 1226 674
rect 1226 640 1260 674
rect 1260 640 1272 674
rect 1299 640 1332 674
rect 1332 640 1351 674
rect 1378 640 1404 674
rect 1404 640 1430 674
rect 1220 631 1272 640
rect 1299 631 1351 640
rect 1378 631 1430 640
rect 1078 586 1130 591
rect 1078 552 1087 586
rect 1087 552 1121 586
rect 1121 552 1130 586
rect 1078 539 1130 552
rect 1078 514 1130 527
rect 1078 480 1087 514
rect 1087 480 1121 514
rect 1121 480 1130 514
rect 1078 475 1130 480
rect 1219 418 1271 427
rect 1219 384 1225 418
rect 1225 384 1259 418
rect 1259 384 1271 418
rect 1219 375 1271 384
rect 1285 418 1337 427
rect 1351 418 1403 427
rect 1416 418 1468 427
rect 1285 384 1307 418
rect 1307 384 1337 418
rect 1351 384 1388 418
rect 1388 384 1403 418
rect 1416 384 1422 418
rect 1422 384 1468 418
rect 1285 375 1337 384
rect 1351 375 1403 384
rect 1416 375 1468 384
rect 1688 101 1740 110
rect 1752 101 1804 110
rect 1688 67 1712 101
rect 1712 67 1740 101
rect 1752 67 1784 101
rect 1784 67 1804 101
rect 1688 58 1740 67
rect 1752 58 1804 67
<< metal2 >>
rect 1409 3682 1415 3734
rect 1467 3682 1483 3734
rect 1535 3682 1551 3734
rect 1603 3682 1618 3734
rect 1670 3682 1685 3734
rect 1737 3682 1752 3734
rect 1804 3682 1810 3734
rect 1409 3646 1810 3682
rect 1409 3594 1415 3646
rect 1467 3594 1483 3646
rect 1535 3594 1551 3646
rect 1603 3594 1618 3646
rect 1670 3594 1685 3646
rect 1737 3594 1752 3646
rect 1804 3594 1810 3646
rect 1409 3240 1810 3594
rect 1409 3188 1415 3240
rect 1467 3188 1483 3240
rect 1535 3188 1551 3240
rect 1603 3188 1618 3240
rect 1670 3188 1685 3240
rect 1737 3188 1752 3240
rect 1804 3188 1810 3240
rect 1409 3166 1810 3188
rect 1409 3114 1415 3166
rect 1467 3114 1483 3166
rect 1535 3114 1551 3166
rect 1603 3114 1618 3166
rect 1670 3114 1685 3166
rect 1737 3114 1752 3166
rect 1804 3114 1810 3166
rect 1409 3092 1810 3114
rect 1409 3040 1415 3092
rect 1467 3040 1483 3092
rect 1535 3040 1551 3092
rect 1603 3040 1618 3092
rect 1670 3040 1685 3092
rect 1737 3040 1752 3092
rect 1804 3040 1810 3092
rect 1214 2975 1314 2981
rect 1214 2923 1238 2975
rect 1290 2923 1314 2975
rect 1214 2907 1314 2923
rect 1214 2855 1238 2907
rect 1290 2855 1314 2907
rect 1214 2839 1314 2855
rect 1214 2787 1238 2839
rect 1290 2787 1314 2839
rect 999 2739 1127 2745
rect 999 2687 1005 2739
rect 1057 2687 1069 2739
rect 1121 2687 1127 2739
rect 999 2625 1127 2687
rect 999 2573 1005 2625
rect 1057 2573 1069 2625
rect 1121 2573 1127 2625
rect 999 2117 1127 2573
rect 999 2065 1005 2117
rect 1057 2065 1069 2117
rect 1121 2065 1127 2117
rect 999 2003 1127 2065
rect 999 1951 1005 2003
rect 1057 1951 1069 2003
rect 1121 1951 1127 2003
rect 999 1903 1127 1951
rect 999 1851 1005 1903
rect 1057 1851 1069 1903
rect 1121 1851 1127 1903
rect 999 1835 1127 1851
rect 999 1783 1005 1835
rect 1057 1783 1069 1835
rect 1121 1783 1127 1835
rect 999 1767 1127 1783
rect 999 1715 1005 1767
rect 1057 1715 1069 1767
rect 1121 1715 1127 1767
rect 999 802 1127 1715
rect 999 750 1005 802
rect 1057 750 1069 802
rect 1121 750 1127 802
rect 1214 1644 1314 2787
rect 1214 1592 1238 1644
rect 1290 1592 1314 1644
rect 1214 1576 1314 1592
rect 1214 1524 1238 1576
rect 1290 1524 1314 1576
rect 1214 1508 1314 1524
rect 1214 1456 1238 1508
rect 1290 1456 1314 1508
tri 1180 683 1214 717 se
rect 1214 683 1314 1456
rect 1409 2415 1810 3040
rect 1409 2363 1415 2415
rect 1467 2363 1483 2415
rect 1535 2363 1551 2415
rect 1603 2363 1618 2415
rect 1670 2363 1685 2415
rect 1737 2363 1752 2415
rect 1804 2363 1810 2415
rect 1409 2327 1810 2363
rect 1409 2275 1415 2327
rect 1467 2275 1483 2327
rect 1535 2275 1551 2327
rect 1603 2275 1618 2327
rect 1670 2275 1685 2327
rect 1737 2275 1752 2327
rect 1804 2275 1810 2327
rect 1409 1096 1810 2275
rect 1409 1044 1415 1096
rect 1467 1044 1483 1096
rect 1535 1044 1551 1096
rect 1603 1044 1618 1096
rect 1670 1044 1685 1096
rect 1737 1044 1752 1096
rect 1804 1044 1810 1096
rect 1409 1008 1810 1044
rect 1409 956 1415 1008
rect 1467 956 1483 1008
rect 1535 956 1551 1008
rect 1603 956 1618 1008
rect 1670 956 1685 1008
rect 1737 956 1752 1008
rect 1804 956 1810 1008
tri 1648 922 1682 956 ne
tri 1314 683 1348 717 sw
rect 719 631 1220 683
rect 1272 631 1299 683
rect 1351 631 1378 683
rect 1430 631 1436 683
tri 1072 591 1078 597 se
rect 1078 591 1130 597
tri 1060 579 1072 591 se
rect 1072 579 1078 591
rect 639 539 1078 579
rect 639 527 1130 539
rect 639 510 1078 527
tri 1044 476 1078 510 ne
rect 1078 469 1130 475
rect 559 375 1219 427
rect 1271 375 1285 427
rect 1337 375 1351 427
rect 1403 375 1416 427
rect 1468 375 1474 427
rect 1682 110 1810 956
rect 2240 3442 2581 3734
rect 2240 3390 2246 3442
rect 2298 3390 2316 3442
rect 2368 3390 2385 3442
rect 2437 3390 2454 3442
rect 2506 3390 2523 3442
rect 2575 3390 2581 3442
rect 2240 3354 2581 3390
rect 2240 3302 2246 3354
rect 2298 3302 2316 3354
rect 2368 3302 2385 3354
rect 2437 3302 2454 3354
rect 2506 3302 2523 3354
rect 2575 3302 2581 3354
rect 2240 2745 2581 3302
rect 2240 2693 2246 2745
rect 2298 2693 2339 2745
rect 2391 2693 2431 2745
rect 2483 2693 2523 2745
rect 2575 2693 2581 2745
rect 2240 2619 2581 2693
rect 2240 2567 2246 2619
rect 2298 2567 2339 2619
rect 2391 2567 2431 2619
rect 2483 2567 2523 2619
rect 2575 2567 2581 2619
rect 2240 2123 2581 2567
rect 2240 2071 2246 2123
rect 2298 2071 2339 2123
rect 2391 2071 2431 2123
rect 2483 2071 2523 2123
rect 2575 2071 2581 2123
rect 2240 1997 2581 2071
rect 2240 1945 2246 1997
rect 2298 1945 2339 1997
rect 2391 1945 2431 1997
rect 2483 1945 2523 1997
rect 2575 1945 2581 1997
rect 2240 1909 2581 1945
rect 2240 1857 2246 1909
rect 2298 1857 2388 1909
rect 2440 1857 2581 1909
rect 2240 1835 2581 1857
rect 2240 1783 2246 1835
rect 2298 1783 2388 1835
rect 2440 1783 2581 1835
rect 2240 1761 2581 1783
rect 2240 1709 2246 1761
rect 2298 1709 2388 1761
rect 2440 1709 2581 1761
rect 2240 1388 2581 1709
rect 2240 1336 2246 1388
rect 2298 1336 2339 1388
rect 2391 1336 2431 1388
rect 2483 1336 2523 1388
rect 2575 1336 2581 1388
rect 2240 1300 2581 1336
rect 2240 1248 2246 1300
rect 2298 1248 2339 1300
rect 2391 1248 2431 1300
rect 2483 1248 2523 1300
rect 2575 1248 2581 1300
rect 2240 844 2581 1248
rect 2638 3370 2803 3735
rect 2690 3318 2750 3370
rect 2802 3318 2803 3370
rect 2638 3262 2803 3318
rect 2690 3210 2750 3262
rect 2802 3210 2803 3262
rect 2638 3153 2803 3210
rect 2690 3101 2750 3153
rect 2802 3101 2803 3153
rect 2638 3061 2803 3101
rect 2638 3009 2644 3061
rect 2696 3009 2745 3061
rect 2797 3009 2803 3061
rect 2638 2965 2803 3009
rect 2638 2913 2644 2965
rect 2696 2913 2745 2965
rect 2797 2913 2803 2965
rect 2638 2872 2803 2913
rect 2690 2820 2750 2872
rect 2802 2820 2803 2872
rect 2638 2782 2803 2820
rect 2690 2730 2750 2782
rect 2802 2730 2803 2782
rect 2638 2692 2803 2730
rect 2690 2640 2750 2692
rect 2802 2640 2803 2692
rect 2638 2051 2803 2640
rect 2690 1999 2750 2051
rect 2802 1999 2803 2051
rect 2638 1961 2803 1999
rect 2690 1909 2750 1961
rect 2802 1909 2803 1961
rect 2638 1870 2803 1909
rect 2690 1818 2750 1870
rect 2802 1818 2803 1870
rect 2638 1777 2803 1818
rect 2638 1725 2644 1777
rect 2696 1725 2745 1777
rect 2797 1725 2803 1777
rect 2638 1681 2803 1725
rect 2638 1629 2644 1681
rect 2696 1629 2745 1681
rect 2797 1629 2803 1681
rect 2638 1589 2803 1629
rect 2690 1537 2750 1589
rect 2802 1537 2803 1589
rect 2638 1481 2803 1537
rect 2690 1429 2750 1481
rect 2802 1429 2803 1481
rect 2638 1372 2803 1429
rect 2690 1320 2750 1372
rect 2802 1320 2803 1372
rect 2638 956 2803 1320
rect 1682 58 1688 110
rect 1740 58 1752 110
rect 1804 58 1810 110
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1624855509
transform 0 -1 1130 1 0 469
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_0
timestamp 1624855509
transform 1 0 1226 0 -1 674
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1624855509
transform 0 -1 1121 -1 0 586
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1624855509
transform -1 0 1137 0 -1 629
box 0 0 1 1
use sky130_fd_io__res250only_small  sky130_fd_io__res250only_small_0
timestamp 1624855509
transform 0 1 146 1 0 116
box 0 0 2270 404
use sky130_fd_pr__nfet_01v8__example_55959141808555  sky130_fd_pr__nfet_01v8__example_55959141808555_0
timestamp 1624855509
transform 0 -1 1763 1 0 429
box -28 0 228 267
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_0
timestamp 1624855509
transform 0 1 737 -1 0 2481
box 0 0 1591 2424
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_1
timestamp 1624855509
transform 0 1 737 1 0 2209
box 0 0 1591 2424
<< labels >>
flabel metal2 s 736 511 830 579 3 FreeSans 200 0 0 0 VTRIP_SEL_H
flabel metal2 s 712 384 811 421 3 FreeSans 200 0 0 0 OUT_VT
flabel metal2 s 1454 3376 1777 3567 3 FreeSans 200 0 0 0 VDDIO_Q
flabel metal2 s 2245 3422 2573 3559 3 FreeSans 200 0 0 0 VSSD
flabel metal2 s 743 637 826 674 3 FreeSans 200 0 0 0 OUT_H
flabel metal1 s 220 116 443 157 3 FreeSans 200 0 0 0 IN_H
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 6240672
string GDS_START 6212544
<< end >>
