magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 1063 391 1105 493
rect 1063 357 1180 391
rect 1146 323 1180 357
rect 1223 323 1273 493
rect 18 215 88 255
rect 205 289 549 323
rect 205 215 304 289
rect 338 215 449 255
rect 483 215 549 289
rect 601 289 955 323
rect 1146 289 1384 323
rect 601 215 721 289
rect 905 255 955 289
rect 755 215 871 255
rect 905 215 1007 255
rect 1315 181 1384 289
rect 1047 147 1384 181
rect 1047 145 1281 147
rect 1047 51 1113 145
rect 1215 51 1281 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 29 291 79 527
rect 113 391 163 493
rect 197 425 247 527
rect 281 459 499 493
rect 281 425 331 459
rect 449 425 499 459
rect 533 425 685 527
rect 719 459 937 493
rect 719 425 769 459
rect 887 425 937 459
rect 971 425 1021 527
rect 365 391 415 425
rect 803 391 853 425
rect 1139 425 1189 527
rect 113 357 1029 391
rect 113 289 169 357
rect 995 323 1029 357
rect 1307 359 1357 527
rect 17 95 69 179
rect 122 173 169 289
rect 995 289 1075 323
rect 1041 255 1075 289
rect 1041 215 1281 255
rect 103 129 169 173
rect 203 95 237 181
rect 271 145 945 181
rect 271 143 777 145
rect 271 129 507 143
rect 17 51 591 95
rect 629 17 677 109
rect 711 51 777 143
rect 811 17 845 111
rect 879 51 945 145
rect 979 17 1013 181
rect 1147 17 1181 111
rect 1315 17 1366 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 905 255 955 289 6 A1
port 1 nsew signal input
rlabel locali s 905 215 1007 255 6 A1
port 1 nsew signal input
rlabel locali s 601 289 955 323 6 A1
port 1 nsew signal input
rlabel locali s 601 215 721 289 6 A1
port 1 nsew signal input
rlabel locali s 755 215 871 255 6 A2
port 2 nsew signal input
rlabel locali s 483 215 549 289 6 B1
port 3 nsew signal input
rlabel locali s 205 289 549 323 6 B1
port 3 nsew signal input
rlabel locali s 205 215 304 289 6 B1
port 3 nsew signal input
rlabel locali s 338 215 449 255 6 B2
port 4 nsew signal input
rlabel locali s 18 215 88 255 6 C1
port 5 nsew signal input
rlabel locali s 1315 181 1384 289 6 X
port 10 nsew signal output
rlabel locali s 1223 323 1273 493 6 X
port 10 nsew signal output
rlabel locali s 1215 51 1281 145 6 X
port 10 nsew signal output
rlabel locali s 1146 323 1180 357 6 X
port 10 nsew signal output
rlabel locali s 1146 289 1384 323 6 X
port 10 nsew signal output
rlabel locali s 1063 391 1105 493 6 X
port 10 nsew signal output
rlabel locali s 1063 357 1180 391 6 X
port 10 nsew signal output
rlabel locali s 1047 147 1384 181 6 X
port 10 nsew signal output
rlabel locali s 1047 145 1281 147 6 X
port 10 nsew signal output
rlabel locali s 1047 51 1113 145 6 X
port 10 nsew signal output
rlabel metal1 s 0 -48 1472 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1510 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4105808
string GDS_START 4094998
<< end >>
