magic
tech sky130A
magscale 1 2
timestamp 1624855514
<< obsli1 >>
rect 0 37 15000 39844
<< metal1 >>
rect 4981 0 5027 1995
<< obsm1 >>
rect 0 2051 15000 39842
rect 0 0 4925 2051
rect 5083 0 15000 2051
<< metal2 >>
rect 2252 7204 2430 7256
rect 2252 6318 2304 7204
rect 2225 6296 2304 6318
rect 2225 6291 2252 6296
rect 2299 6291 2304 6296
rect 2173 6267 2225 6291
rect 2254 6267 2299 6291
rect 2173 6253 2299 6267
rect 2173 6246 2225 6253
rect 2254 6246 2299 6253
rect 2173 6217 2254 6246
rect 2173 5725 2225 6217
rect 2130 5630 2225 5725
rect 2182 5629 2225 5630
rect 2130 5587 2225 5629
rect 2130 5460 2182 5587
rect 2130 5322 2225 5460
rect 2173 2020 2225 5322
rect 2099 1946 2225 2020
rect 6073 3270 6125 4099
rect 5999 3196 6125 3270
rect 5954 3179 5999 3196
rect 6006 3179 6073 3196
rect 5954 3129 6073 3179
rect 5954 2307 6006 3129
rect 2033 1920 2099 1946
rect 2107 1920 2173 1946
rect 2033 1892 2173 1920
rect 2033 1880 2099 1892
rect 2107 1880 2173 1892
rect 5880 2233 6006 2307
rect 1993 1864 2033 1880
rect 2067 1864 2107 1880
rect 1993 1850 2107 1864
rect 1993 1840 2033 1850
rect 2067 1840 2107 1850
rect 1947 1822 1993 1840
rect 1999 1822 2067 1840
rect 1947 1772 2067 1822
rect 1947 915 1999 1772
rect 5864 2217 5880 2233
rect 5916 2217 5954 2233
rect 5864 2195 5954 2217
rect 5864 1094 5916 2195
rect 5816 1072 5916 1094
rect 5816 1046 5864 1072
rect 5890 1046 5916 1072
rect 5750 1031 5816 1046
rect 5824 1031 5890 1046
rect 5750 989 5890 1031
rect 5750 980 5816 989
rect 5824 980 5890 989
rect 5731 961 5750 980
rect 5753 961 5824 980
rect 3103 951 5824 961
rect 2009 915 2075 916
rect 1947 865 2075 915
rect 1947 850 2001 865
rect 2009 850 2075 865
rect 3103 937 3177 951
rect 4472 937 4532 951
rect 5753 937 5824 951
rect 3103 909 5824 937
rect 3103 887 3199 909
rect 2001 837 2070 850
rect 2075 837 2139 850
rect 2001 809 2139 837
rect 2001 781 2070 809
rect 2075 786 2139 809
rect 3029 813 3177 887
rect 4412 852 4589 909
rect 4412 849 4532 852
rect 2975 795 3029 813
rect 3049 795 3103 813
rect 2139 781 2186 786
rect 2070 753 2186 781
rect 2975 767 3103 795
rect 2975 759 3029 767
rect 3049 759 3103 767
rect 2070 729 2136 753
rect 2139 739 2186 753
rect 2955 739 2975 759
rect 2977 739 3049 759
rect 2164 729 3049 739
rect 2070 715 3049 729
rect 2136 687 3049 715
rect 2457 0 2509 294
rect 2911 0 3027 197
rect 4472 0 4532 849
rect 5516 0 5646 66
rect 6101 0 6231 66
rect 6552 0 6604 128
<< obsm2 >>
rect 68 7312 14983 39842
rect 68 6374 2196 7312
rect 68 6347 2169 6374
rect 68 5781 2117 6347
rect 2486 7148 14983 7312
rect 2360 6235 14983 7148
rect 68 5266 2074 5781
rect 2355 6190 14983 6235
rect 2310 6161 14983 6190
rect 2281 5531 14983 6161
rect 2238 5516 14983 5531
rect 68 2076 2117 5266
rect 68 2002 2043 2076
rect 68 1936 1977 2002
rect 2281 4155 14983 5516
rect 2281 3326 6017 4155
rect 2281 3252 5943 3326
rect 2281 2363 5898 3252
rect 6181 3140 14983 4155
rect 2281 2289 5824 2363
rect 6129 3073 14983 3140
rect 68 1896 1937 1936
rect 68 794 1891 1896
rect 2281 1890 5808 2289
rect 2229 1824 5808 1890
rect 2163 1784 5808 1824
rect 2123 1716 5808 1784
rect 2055 1150 5808 1716
rect 2055 1102 5760 1150
rect 2055 1036 5694 1102
rect 6062 2177 14983 3073
rect 6010 2139 14983 2177
rect 2055 1017 5675 1036
rect 2055 972 3047 1017
rect 5972 990 14983 2139
rect 2131 943 3047 972
rect 2131 906 2973 943
rect 2195 869 2973 906
rect 5946 924 14983 990
rect 2195 842 2919 869
rect 68 725 1945 794
rect 2242 815 2919 842
rect 2242 795 2899 815
rect 3255 831 4356 853
rect 5880 853 14983 924
rect 3233 793 4356 831
rect 3233 757 4416 793
rect 68 659 2014 725
rect 3159 703 4416 757
rect 68 631 2080 659
rect 3105 631 4416 703
rect 68 350 4416 631
rect 68 0 2401 350
rect 2565 253 4416 350
rect 2565 0 2855 253
rect 3083 0 4416 253
rect 4645 796 14983 853
rect 4588 184 14983 796
rect 4588 122 6496 184
rect 4588 0 5460 122
rect 5702 0 6045 122
rect 6287 0 6496 122
rect 6660 0 14983 184
<< metal3 >>
rect 12972 14480 13198 18929
rect 12972 14442 13236 14480
rect 12972 14416 13232 14442
rect 13236 14416 13478 14442
rect 12972 14240 13478 14416
rect 12972 14180 13208 14240
rect 13236 14200 13478 14240
rect 13478 14180 13671 14200
rect 12972 14150 13671 14180
rect 13208 14007 13671 14150
rect 13208 14000 13478 14007
rect 13671 14000 13861 14007
rect 13208 13940 13861 14000
rect 13208 13910 13478 13940
rect 13671 13910 13861 13940
rect 13208 13880 13861 13910
rect 13478 13820 13861 13880
rect 13478 13790 13651 13820
rect 13671 13817 13861 13820
rect 13861 13790 14118 13817
rect 13478 13760 14118 13790
rect 13478 13707 13651 13760
rect 13861 13730 14118 13760
rect 13658 13707 14118 13730
rect 13651 13610 14118 13707
rect 13651 13550 13838 13610
rect 13861 13560 14118 13610
rect 14118 13550 14438 13560
rect 13651 13520 14438 13550
rect 13838 13240 14438 13520
rect 14118 12920 14785 13240
rect 14438 9997 14785 12920
rect 14652 9984 14785 9997
rect 1794 6799 4455 6825
rect 1794 6769 1879 6799
rect 1794 6740 4455 6769
rect 1690 6709 1794 6740
rect 1823 6739 4455 6740
rect 1690 6679 4455 6709
rect 1690 6636 1794 6679
rect 1836 6636 1879 6679
rect 1573 6601 1690 6636
rect 1719 6601 1836 6636
rect 1573 6541 1836 6601
rect 1573 6519 1690 6541
rect 1719 6519 1836 6541
rect 1430 6481 1573 6519
rect 1576 6481 1719 6519
rect 1430 6391 1719 6481
rect 1430 6376 1573 6391
rect 1576 6376 1719 6391
rect 1355 6331 1430 6376
rect 1459 6331 1576 6376
rect 1355 6259 1576 6331
rect 1355 3524 1459 6259
rect 1355 3469 1574 3524
rect 1355 3409 1458 3469
rect 1459 3409 1574 3469
rect 1355 3379 1666 3409
rect 1458 3349 1666 3379
rect 1458 3289 1548 3349
rect 1574 3317 1666 3349
rect 1666 3289 1784 3317
rect 1548 3259 1784 3289
rect 1548 3199 1638 3259
rect 1666 3199 1784 3259
rect 1638 3157 1784 3199
rect 1680 0 1784 3157
rect 4581 1996 4810 2453
rect 4268 1899 4810 1996
rect 4268 1880 4581 1899
rect 4594 1880 4810 1899
rect 4268 1700 4810 1880
rect 4268 1683 4581 1700
rect 4594 1683 4810 1700
rect 5634 2182 5780 2954
rect 5634 2089 5933 2182
rect 5634 2029 5727 2089
rect 5780 2029 5933 2089
rect 5727 1969 5933 2029
rect 4212 1627 4268 1683
rect 4538 1627 4594 1683
rect 3449 0 3782 627
rect 4015 1580 4212 1627
rect 4245 1580 4538 1627
rect 4015 1334 4538 1580
rect 4015 0 4245 1334
rect 5787 0 5933 1969
rect 14438 9864 14785 9984
rect 14438 0 14652 9864
<< obsm3 >>
rect 193 19009 14940 40000
rect 193 14070 12892 19009
rect 13278 14560 14940 19009
rect 13316 14522 14940 14560
rect 13558 14280 14940 14522
rect 193 13800 13128 14070
rect 13751 14087 14940 14280
rect 13941 13897 14940 14087
rect 193 13627 13398 13800
rect 193 13440 13571 13627
rect 14198 13640 14940 13897
rect 193 13160 13758 13440
rect 14518 13320 14940 13640
rect 193 12840 14038 13160
rect 193 6905 14358 12840
rect 193 6820 1714 6905
rect 193 6716 1610 6820
rect 193 6599 1493 6716
rect 193 6456 1350 6599
rect 4535 6599 14358 6905
rect 1959 6556 14358 6599
rect 193 3299 1275 6456
rect 1916 6439 14358 6556
rect 1799 6296 14358 6439
rect 1656 6179 14358 6296
rect 1539 3604 14358 6179
rect 1654 3489 14358 3604
rect 1746 3397 14358 3489
rect 193 3209 1378 3299
rect 193 3119 1468 3209
rect 193 3077 1558 3119
rect 193 125 1600 3077
rect 1864 3034 14358 3397
rect 1864 2533 5554 3034
rect 1864 2076 4501 2533
rect 1864 1763 4188 2076
rect 1864 1707 4132 1763
rect 1864 707 3935 1707
rect 4890 1949 5554 2533
rect 5860 2262 14358 3034
rect 4890 1889 5647 1949
rect 1864 125 3369 707
rect 3862 125 3935 707
rect 4890 1603 5707 1889
rect 4674 1547 5707 1603
rect 4618 1254 5707 1547
rect 4325 125 5707 1254
rect 6013 125 14358 2262
rect 14865 9784 14940 13320
rect 14732 125 14940 9784
<< metal4 >>
rect 0 10625 15000 11221
rect 0 9673 15000 10269
<< obsm4 >>
rect 0 11301 15000 40000
rect 0 10349 15000 10545
rect 0 407 15000 9593
<< metal5 >>
rect 1220 20802 13760 33325
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14807 3007 15000 3657
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 0 33645 15000 40000
rect 0 20482 900 33645
rect 14080 20482 15000 33645
rect 0 19317 15000 20482
rect 0 8017 14426 19317
rect 0 7367 15000 8017
rect 0 4867 14426 7367
rect 0 3977 15000 4867
rect 0 3007 14487 3977
rect 0 427 14426 3007
<< labels >>
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal2 s 6552 0 6604 128 6 DISABLE_PULLUP_H
port 3 nsew signal input
rlabel metal2 s 2457 0 2509 294 6 ENABLE_H
port 4 nsew signal input
rlabel metal3 s 1355 3379 1458 3482 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1355 3482 1459 6280 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1355 3482 1480 3503 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1355 3503 1459 3524 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1355 3524 1459 6259 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1355 6280 1480 6301 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1355 6301 1430 6376 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1368 3469 1501 3482 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1385 6301 1501 6331 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1430 6376 1573 6519 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1458 3289 1548 3379 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1458 3379 1574 3409 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1459 3409 1574 3524 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1459 6259 1576 6376 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1475 6391 1591 6421 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1488 3349 1604 3379 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1505 6421 1621 6451 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1535 6451 1651 6481 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1548 3199 1638 3289 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1573 6519 1690 6636 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1574 3317 1666 3409 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1576 6376 1719 6519 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1578 3259 1694 3289 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1625 6541 1741 6571 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1638 3157 1680 3199 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1655 6571 1771 6601 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1666 3199 1784 3317 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1680 0 1784 3157 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1680 227 1784 3199 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1690 6636 1794 6740 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1719 6519 1836 6636 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1763 6679 4455 6709 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1794 6740 1879 6825 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1823 6739 4455 6769 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1836 6636 1879 6679 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal3 s 1879 6799 4455 6825 6 ENABLE_VDDIO
port 5 nsew signal input
rlabel metal2 s 2001 781 2070 850 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2009 850 2075 916 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2017 1850 2077 1864 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2028 823 2088 837 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2033 1880 2099 1946 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2042 809 2102 823 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2059 1892 2119 1906 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2067 1840 2107 1880 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2070 715 2136 781 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2073 1906 2133 1920 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2075 786 2139 850 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2084 767 2144 781 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2098 753 2158 767 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2099 1946 2173 2020 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2107 1880 2173 1946 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2115 1948 2175 1962 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2129 1962 2189 1976 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5322 2173 5365 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5365 2225 5417 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5417 2182 5601 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5417 2211 5431 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5431 2197 5445 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5459 2182 5460 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5460 2182 5587 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5601 2196 5615 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5615 2210 5629 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5630 2225 5682 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2130 5682 2173 5725 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2131 5364 2225 5365 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2136 687 2164 715 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2136 715 3005 729 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2139 739 2186 786 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2143 1976 2203 1990 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2144 5682 2225 5696 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2145 5350 2225 5364 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2158 5696 2225 5710 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2164 687 2977 739 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 2009 2225 2020 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 2020 2225 5322 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 5630 2225 6228 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 5724 2225 5725 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 5725 2225 6217 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 6228 2236 6239 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 6239 2225 6291 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 1946 2225 1998 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2173 1998 2225 5417 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2182 5417 2225 5460 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2182 5587 2225 5630 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2201 6253 2261 6267 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2225 6217 2254 6246 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2225 6291 2252 6318 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2252 6296 2304 7204 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2252 6307 2304 6318 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2252 7204 2430 7256 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2254 6246 2299 6291 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2299 6291 2304 6296 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2955 739 2975 759 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2975 759 3029 813 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2977 687 3049 759 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 2997 767 3057 781 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3011 781 3071 795 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3029 813 3103 887 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3049 759 3103 813 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3053 823 3113 837 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3067 837 3127 851 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3081 851 3141 865 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3103 813 3177 887 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3103 887 3177 961 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3123 893 3183 907 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3139 909 5753 923 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3153 923 5767 937 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3177 887 3199 909 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 3177 951 5795 961 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4412 849 4472 909 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4413 908 4588 909 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4427 894 4574 908 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4441 880 4560 894 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4469 852 4532 866 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4470 851 4532 852 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4472 0 4532 849 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4472 234 4532 961 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 4532 852 4589 909 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5731 961 5750 980 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5750 980 5816 1046 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5753 909 5824 980 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5773 989 5833 1003 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5787 1003 5847 1017 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5801 1017 5861 1031 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5816 1046 5864 1094 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5824 980 5890 1046 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5864 2206 5927 2217 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5864 2217 5880 2233 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5864 1072 5916 2206 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5864 1083 5916 1094 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5864 1094 5916 2195 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5880 2233 5954 2307 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5890 1046 5916 1072 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5906 2245 5966 2259 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5916 2195 5954 2233 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5920 2259 5980 2273 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5954 2233 6006 2285 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5954 2285 6006 3140 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5954 2296 6006 2307 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5954 2307 6006 3129 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5954 3140 6017 3151 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5954 3151 5999 3196 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5968 3151 6028 3165 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5982 3165 6042 3179 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 5999 3196 6073 3270 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 6006 3129 6073 3196 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 6024 3207 6084 3221 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 6038 3221 6098 3235 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 6073 3196 6125 3248 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 6073 3248 6125 3270 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 6073 3270 6125 4099 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1947 850 2001 904 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1947 904 2010 915 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1947 904 1999 1783 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1947 915 1999 926 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1947 926 1999 1772 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1947 1783 2010 1794 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1947 1794 1993 1840 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1958 893 2021 904 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1961 1794 2021 1808 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1972 879 2032 893 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1975 1808 2035 1822 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1986 865 2046 879 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1993 1840 2033 1880 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal2 s 1999 1772 2067 1840 6 EN_VDDIO_SIG_H
port 6 nsew signal input
rlabel metal3 s 4015 0 4245 1334 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4015 682 4245 1364 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4015 1364 4275 1394 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4015 1394 4305 1424 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4015 1424 4335 1430 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4015 1430 4212 1627 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4045 1430 4341 1460 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4075 1460 4371 1490 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4105 1490 4401 1520 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4135 1520 4431 1550 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4165 1550 4461 1580 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4212 1627 4268 1683 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4245 1334 4538 1627 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4268 1683 4581 1996 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4315 1700 4611 1730 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4345 1730 4641 1760 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4375 1760 4671 1790 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4405 1790 4701 1820 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4435 1820 4731 1850 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4465 1850 4761 1880 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4514 1899 4810 1929 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4538 1627 4594 1683 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4544 1929 4810 1959 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4581 1899 4810 1996 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4581 1996 4810 2453 6 FILT_IN_H
port 7 nsew signal input
rlabel metal3 s 4594 1683 4810 1899 6 FILT_IN_H
port 7 nsew signal input
rlabel metal1 s 4981 0 5027 1995 6 INP_SEL_H
port 8 nsew signal input
rlabel metal5 s 1220 20802 13760 33325 6 PAD
port 9 nsew signal bidirectional
rlabel metal3 s 3449 0 3782 627 6 PAD_A_ESD_H
port 10 nsew signal bidirectional
rlabel metal2 s 2911 0 3027 197 6 PULLUP_H
port 11 nsew signal bidirectional
rlabel metal2 s 6101 0 6231 66 6 TIE_HI_ESD
port 12 nsew signal output
rlabel metal2 s 5516 0 5646 66 6 TIE_LO_ESD
port 13 nsew signal output
rlabel metal3 s 12972 14150 13208 14386 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 12972 14386 13198 14480 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 12972 14386 13262 14416 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 12972 14416 13232 14446 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 12972 14480 13198 18929 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 12998 14360 13292 14386 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13028 14330 13318 14360 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13058 14300 13348 14330 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13088 14270 13378 14300 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13118 14240 13408 14270 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13198 14442 13236 14480 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13208 13880 13478 14150 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13208 14150 13498 14180 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13236 14200 13478 14442 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13238 14120 13528 14150 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13268 14090 13558 14120 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13298 14060 13588 14090 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13328 14030 13618 14060 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13388 13970 13678 14000 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13418 13940 13708 13970 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13478 13707 13651 13880 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13478 13880 13768 13910 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13478 14007 13671 14200 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13508 13850 13798 13880 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13538 13820 13828 13850 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13598 13760 13888 13790 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13651 13520 13838 13707 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13658 13700 13948 13730 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13671 13817 13861 14007 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13688 13670 13978 13700 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13718 13640 14008 13670 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13748 13610 14038 13640 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13838 13240 14118 13520 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13838 13520 14128 13550 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13861 13560 14118 13817 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13868 13490 14158 13520 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13898 13460 14188 13490 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13928 13430 14218 13460 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13958 13400 14248 13430 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 13988 13370 14278 13400 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14018 13340 14308 13370 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14048 13310 14338 13340 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14078 13280 14368 13310 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14118 12920 14438 13240 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14118 13240 14438 13560 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14168 13190 14458 13220 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14198 13160 14488 13190 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14228 13130 14518 13160 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14258 13100 14548 13130 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14288 13070 14578 13100 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14318 13040 14608 13070 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14348 13010 14638 13040 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14378 12980 14668 13010 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 0 14652 9864 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 145 14652 9894 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 9894 14682 9924 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 9924 14712 9954 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 9954 14742 9984 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 9997 14785 12893 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 12893 14772 12906 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 12893 14785 13240 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 12906 14759 12919 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14438 12919 14758 12920 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 14652 9864 14785 9997 6 TIE_WEAK_HI_H
port 14 nsew signal bidirectional
rlabel metal3 s 5634 2029 5727 2122 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5634 2122 5780 2182 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5634 2122 5810 2152 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5634 2182 5780 2954 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5637 2119 5840 2122 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5667 2089 5843 2119 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5727 1969 5787 2029 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5780 2029 5933 2182 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5787 0 5933 1969 6 XRES_H_N
port 15 nsew signal output
rlabel metal3 s 5787 801 5933 2029 6 XRES_H_N
port 15 nsew signal output
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 16 nsew power input
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 17 nsew power input
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 18 nsew power input
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 19 nsew power input
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 20 nsew power input
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 21 nsew ground input
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 22 nsew ground input
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 23 nsew ground input
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 24 nsew ground input
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 25 nsew power input
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 40000
string LEFsymmetry R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 13341894
string GDS_START 9248522
<< end >>
