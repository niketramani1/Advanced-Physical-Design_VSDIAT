magic
tech sky130A
magscale 1 2
timestamp 1624855598
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 125 265 191 485
rect 293 288 349 493
rect 293 265 342 288
rect 125 199 342 265
rect 125 75 175 199
rect 293 185 342 199
rect 293 70 345 185
rect 599 215 712 265
rect 1521 289 1637 323
rect 1521 199 1555 289
rect 1685 215 1767 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 57 298 91 527
rect 225 299 259 527
rect 383 443 450 527
rect 486 447 780 481
rect 921 447 987 527
rect 1054 455 1673 489
rect 1755 455 1822 527
rect 486 409 520 447
rect 1054 413 1088 455
rect 383 375 520 409
rect 588 379 1088 413
rect 383 265 417 375
rect 463 307 780 341
rect 376 199 417 265
rect 57 17 91 147
rect 225 17 259 147
rect 382 173 417 199
rect 382 139 497 173
rect 379 17 429 105
rect 463 85 497 139
rect 531 119 565 307
rect 746 265 780 307
rect 814 305 891 339
rect 835 275 891 305
rect 746 199 801 265
rect 625 159 701 181
rect 835 159 869 275
rect 925 241 959 379
rect 1005 289 1089 343
rect 625 125 869 159
rect 903 207 959 241
rect 903 91 937 207
rect 690 85 777 91
rect 463 51 777 85
rect 811 57 937 91
rect 971 17 1005 173
rect 1041 83 1089 289
rect 1125 119 1159 421
rect 1193 178 1227 455
rect 1856 421 1915 493
rect 1263 323 1346 409
rect 1453 387 1915 421
rect 1263 289 1419 323
rect 1266 199 1351 254
rect 1193 165 1235 178
rect 1193 144 1275 165
rect 1201 131 1275 144
rect 1125 97 1167 119
rect 1125 53 1207 97
rect 1241 64 1275 131
rect 1309 126 1351 199
rect 1385 85 1419 289
rect 1453 119 1487 387
rect 1818 375 1915 387
rect 1671 299 1835 341
rect 1801 265 1835 299
rect 1589 189 1651 255
rect 1801 199 1847 265
rect 1589 146 1630 189
rect 1801 181 1835 199
rect 1687 150 1835 181
rect 1679 147 1835 150
rect 1521 85 1614 93
rect 1385 51 1614 85
rect 1679 59 1737 147
rect 1881 117 1915 375
rect 1771 17 1805 113
rect 1855 51 1915 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< obsm1 >>
rect 845 320 903 329
rect 1305 320 1363 329
rect 845 292 1363 320
rect 845 283 903 292
rect 1305 283 1363 292
rect 1029 184 1087 193
rect 1305 184 1363 193
rect 1581 184 1639 193
rect 1029 156 1639 184
rect 1029 147 1087 156
rect 1305 147 1363 156
rect 1581 147 1639 156
rect 1121 116 1179 125
rect 1673 116 1731 125
rect 1121 88 1731 116
rect 1121 79 1179 88
rect 1673 79 1731 88
<< labels >>
rlabel locali s 1685 215 1767 265 6 A
port 1 nsew signal input
rlabel locali s 1521 289 1637 323 6 B
port 2 nsew signal input
rlabel locali s 1521 199 1555 289 6 B
port 2 nsew signal input
rlabel locali s 599 215 712 265 6 C
port 3 nsew signal input
rlabel locali s 293 288 349 493 6 X
port 8 nsew signal output
rlabel locali s 293 265 342 288 6 X
port 8 nsew signal output
rlabel locali s 293 185 342 199 6 X
port 8 nsew signal output
rlabel locali s 293 70 345 185 6 X
port 8 nsew signal output
rlabel locali s 125 265 191 485 6 X
port 8 nsew signal output
rlabel locali s 125 199 342 265 6 X
port 8 nsew signal output
rlabel locali s 125 75 175 199 6 X
port 8 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3275496
string GDS_START 3262310
<< end >>
