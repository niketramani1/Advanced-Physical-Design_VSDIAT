magic
tech sky130A
magscale 1 2
timestamp 1624855595
<< checkpaint >>
rect -1298 -1308 2402 1852
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 16 -26 72 30
<< scnmos >>
rect 79 47 1025 157
<< scpmoshvt >>
rect 79 323 1025 497
<< ndiff >>
rect 27 112 79 157
rect 27 78 35 112
rect 69 78 79 112
rect 27 47 79 78
rect 1025 112 1077 157
rect 1025 78 1035 112
rect 1069 78 1077 112
rect 1025 47 1077 78
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 323 79 451
rect 1025 485 1077 497
rect 1025 451 1035 485
rect 1069 451 1077 485
rect 1025 323 1077 451
<< ndiffc >>
rect 35 78 69 112
rect 1035 78 1069 112
<< pdiffc >>
rect 35 451 69 485
rect 1035 451 1069 485
<< poly >>
rect 79 497 1025 523
rect 79 297 1025 323
rect 79 275 529 297
rect 79 241 351 275
rect 385 241 529 275
rect 79 225 529 241
rect 571 239 1025 255
rect 571 205 715 239
rect 749 205 1025 239
rect 571 183 1025 205
rect 79 157 1025 183
rect 79 21 1025 47
<< polycont >>
rect 351 241 385 275
rect 715 205 749 239
<< locali >>
rect 0 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 485 1086 527
rect 17 451 35 485
rect 69 451 1035 485
rect 1069 451 1086 485
rect 17 440 1086 451
rect 334 275 402 292
rect 334 241 351 275
rect 385 241 402 275
rect 334 126 402 241
rect 698 239 768 440
rect 698 205 715 239
rect 749 205 768 239
rect 698 190 768 205
rect 17 112 1086 126
rect 17 78 35 112
rect 69 78 1035 112
rect 1069 78 1086 112
rect 17 17 1086 78
rect 0 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel metal1 s 0 -48 1104 48 0 FreeSans 250 0 0 0 VGND
port 3 nsew ground input
flabel metal1 s 0 496 1104 592 0 FreeSans 250 0 0 0 VPWR
port 1 nsew power input
flabel nwell s -38 261 1142 582 0 FreeSans 250 0 0 0 VPB
port 2 nsew default input
flabel pwell s 16 -26 72 30 0 FreeSans 250 0 0 0 VNB
port 4 nsew default input
rlabel metal1 0 0 0 0 4 decap_12
rlabel viali s 1041 -17 1075 17 1 VGND
port 3 nsew ground input
rlabel viali s 949 -17 983 17 1 VGND
port 3 nsew ground input
rlabel viali s 857 -17 891 17 1 VGND
port 3 nsew ground input
rlabel viali s 765 -17 799 17 1 VGND
port 3 nsew ground input
rlabel viali s 673 -17 707 17 1 VGND
port 3 nsew ground input
rlabel viali s 581 -17 615 17 1 VGND
port 3 nsew ground input
rlabel viali s 489 -17 523 17 1 VGND
port 3 nsew ground input
rlabel viali s 397 -17 431 17 1 VGND
port 3 nsew ground input
rlabel viali s 305 -17 339 17 1 VGND
port 3 nsew ground input
rlabel viali s 213 -17 247 17 1 VGND
port 3 nsew ground input
rlabel viali s 121 -17 155 17 1 VGND
port 3 nsew ground input
rlabel locali s 0 -17 1104 17 1 VGND
port 3 nsew ground input
rlabel locali s 17 17 1086 126 1 VGND
port 3 nsew ground input
rlabel locali s 334 126 402 292 1 VGND
port 3 nsew ground input
rlabel viali s 1041 527 1075 561 1 VPWR
port 1 nsew power input
rlabel viali s 949 527 983 561 1 VPWR
port 1 nsew power input
rlabel viali s 857 527 891 561 1 VPWR
port 1 nsew power input
rlabel viali s 765 527 799 561 1 VPWR
port 1 nsew power input
rlabel viali s 673 527 707 561 1 VPWR
port 1 nsew power input
rlabel viali s 581 527 615 561 1 VPWR
port 1 nsew power input
rlabel viali s 489 527 523 561 1 VPWR
port 1 nsew power input
rlabel viali s 397 527 431 561 1 VPWR
port 1 nsew power input
rlabel viali s 305 527 339 561 1 VPWR
port 1 nsew power input
rlabel viali s 213 527 247 561 1 VPWR
port 1 nsew power input
rlabel viali s 121 527 155 561 1 VPWR
port 1 nsew power input
rlabel locali s 698 190 768 440 1 VPWR
port 1 nsew power input
rlabel locali s 17 440 1086 527 1 VPWR
port 1 nsew power input
rlabel locali s 0 527 1104 561 1 VPWR
port 1 nsew power input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 1104 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ef_sc_hd__decap_12.gds
string GDS_END 3582
string GDS_START 142
<< end >>
